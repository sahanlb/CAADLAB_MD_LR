localparam [0:49228][125:0] P_INFO_NEW = {
  1'd1,  4'd0, 27'h00000255, 4'd3, 27'h000003bd, 4'd2, 27'h000001c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001b2, 4'd2, 27'h0000028d, 4'd6, 27'h000001a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001c3, 4'd4, 27'h0000000b, 4'd13, 27'h000002f4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000030b, 4'd6, 27'h000003ba, 4'd0, 27'h00000266, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000358, 4'd7, 27'h0000030a, 4'd8, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000144, 4'd8, 27'h0000022b, 4'd11, 27'h000002ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000b7, 4'd10, 27'h00000307, 4'd2, 27'h000001ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000294, 4'd12, 27'h00000245, 4'd8, 27'h0000004c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000163, 4'd12, 27'h00000115, 4'd11, 27'h000002e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003c0, 4'd1, 27'h0000016d, 4'd0, 27'h0000003f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000337, 4'd2, 27'h00000048, 4'd5, 27'h00000295, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000064, 4'd2, 27'h00000355, 4'd11, 27'h000002dd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002ec, 4'd6, 27'h00000101, 4'd3, 27'h00000381, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001d7, 4'd5, 27'h00000291, 4'd9, 27'h00000141, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002ef, 4'd7, 27'h00000097, 4'd11, 27'h000000e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001f1, 4'd10, 27'h0000036c, 4'd3, 27'h000002e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000286, 4'd14, 27'h00000193, 4'd5, 27'h0000002f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000010f, 4'd14, 27'h00000382, 4'd12, 27'h000002f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003e2, 4'd2, 27'h000001f7, 4'd4, 27'h00000373, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000a3, 4'd3, 27'h00000100, 4'd5, 27'h00000170, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000013f, 4'd0, 27'h000003b9, 4'd13, 27'h000003a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001ca, 4'd9, 27'h00000265, 4'd1, 27'h000003ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000238, 4'd7, 27'h000003f0, 4'd5, 27'h000003c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000fd, 4'd5, 27'h00000174, 4'd11, 27'h0000005f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000017d, 4'd13, 27'h0000031a, 4'd3, 27'h00000120, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000010c, 4'd13, 27'h000002e0, 4'd9, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000244, 4'd13, 27'h00000214, 4'd12, 27'h0000033d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000ce, 4'd2, 27'h000002a5, 4'd1, 27'h0000011b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000393, 4'd1, 27'h000000c0, 4'd8, 27'h00000339, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000167, 4'd4, 27'h000003b3, 4'd11, 27'h000002f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000374, 4'd9, 27'h00000304, 4'd1, 27'h000002c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000131, 4'd6, 27'h00000074, 4'd7, 27'h000002bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000035b, 4'd6, 27'h0000011e, 4'd10, 27'h00000321, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000ea, 4'd10, 27'h000001c2, 4'd3, 27'h0000027c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000020c, 4'd11, 27'h000001e2, 4'd7, 27'h000001a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000283, 4'd10, 27'h00000393, 4'd11, 27'h00000376, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001d5, 4'd4, 27'h00000172, 4'd4, 27'h0000025e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000010b, 4'd0, 27'h00000312, 4'd8, 27'h00000159, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000002a, 4'd4, 27'h00000344, 4'd12, 27'h00000084, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b1, 4'd7, 27'h00000183, 4'd1, 27'h000002b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000366, 4'd6, 27'h0000002f, 4'd8, 27'h0000025a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000015f, 4'd7, 27'h0000019d, 4'd13, 27'h000000f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000e3, 4'd14, 27'h00000017, 4'd0, 27'h000000f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001b5, 4'd14, 27'h0000020c, 4'd8, 27'h0000011a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002d2, 4'd14, 27'h000002db, 4'd13, 27'h00000189, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002a6, 4'd3, 27'h0000010d, 4'd2, 27'h00000086, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000007c, 4'd4, 27'h0000013d, 4'd5, 27'h000001f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000002f, 4'd1, 27'h000003e7, 4'd11, 27'h000000ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000097, 4'd7, 27'h00000243, 4'd0, 27'h00000177, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000027a, 4'd5, 27'h000003dc, 4'd9, 27'h00000109, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000036e, 4'd6, 27'h000002b8, 4'd12, 27'h000001ef, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000017, 4'd13, 27'h00000207, 4'd1, 27'h00000146, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000199, 4'd11, 27'h00000143, 4'd6, 27'h000000ee, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000018, 4'd10, 27'h000000cc, 4'd14, 27'h0000038b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000260, 4'd3, 27'h000002d2, 4'd3, 27'h00000321, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003b4, 4'd2, 27'h000000fb, 4'd5, 27'h0000002b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000c3, 4'd2, 27'h00000201, 4'd10, 27'h00000288, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000126, 4'd7, 27'h0000021e, 4'd1, 27'h00000261, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000d2, 4'd9, 27'h00000146, 4'd7, 27'h000003e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002e4, 4'd7, 27'h0000019e, 4'd12, 27'h000002e3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000044, 4'd10, 27'h0000004c, 4'd4, 27'h00000246, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001d5, 4'd11, 27'h0000019e, 4'd9, 27'h00000078, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001d6, 4'd13, 27'h0000030f, 4'd11, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b8, 4'd4, 27'h000003b4, 4'd3, 27'h00000123, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000036f, 4'd1, 27'h0000003d, 4'd9, 27'h000001bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000220, 4'd1, 27'h0000005a, 4'd13, 27'h000001ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000217, 4'd8, 27'h0000023e, 4'd4, 27'h000001b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000d6, 4'd9, 27'h000003d9, 4'd9, 27'h00000390, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000052, 4'd6, 27'h0000030d, 4'd12, 27'h000002ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000016c, 4'd14, 27'h00000184, 4'd1, 27'h00000252, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000016, 4'd13, 27'h00000112, 4'd5, 27'h000002b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000016b, 4'd14, 27'h0000026c, 4'd12, 27'h00000319, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002c7, 4'd2, 27'h0000034f, 4'd0, 27'h00000047, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003ca, 4'd4, 27'h00000153, 4'd6, 27'h000002d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000005e, 4'd1, 27'h000000e3, 4'd10, 27'h0000013e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000154, 4'd9, 27'h0000002f, 4'd4, 27'h000000cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000017d, 4'd6, 27'h0000019a, 4'd5, 27'h00000198, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003ee, 4'd9, 27'h000001c5, 4'd12, 27'h0000024e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000038e, 4'd11, 27'h00000251, 4'd1, 27'h000002c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000c8, 4'd11, 27'h00000350, 4'd5, 27'h000001cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000184, 4'd13, 27'h0000021f, 4'd13, 27'h0000012f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002d1, 4'd1, 27'h0000001d, 4'd4, 27'h00000003, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003a0, 4'd3, 27'h0000001d, 4'd8, 27'h00000304, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000329, 4'd3, 27'h0000013b, 4'd12, 27'h00000204, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003fc, 4'd9, 27'h00000202, 4'd1, 27'h00000121, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000387, 4'd7, 27'h00000033, 4'd5, 27'h000001ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000116, 4'd6, 27'h00000260, 4'd14, 27'h000003b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000030b, 4'd11, 27'h0000017c, 4'd1, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000356, 4'd14, 27'h0000003c, 4'd8, 27'h0000005a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000248, 4'd10, 27'h00000029, 4'd13, 27'h00000220, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000033b, 4'd1, 27'h0000005f, 4'd3, 27'h00000048, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000088, 4'd4, 27'h000003ad, 4'd9, 27'h00000361, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000028, 4'd2, 27'h0000031e, 4'd11, 27'h000001b4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000008c, 4'd5, 27'h0000011e, 4'd3, 27'h000002c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002f5, 4'd9, 27'h000002ec, 4'd9, 27'h0000022f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000007c, 4'd5, 27'h000002b5, 4'd11, 27'h0000009c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000db, 4'd13, 27'h00000257, 4'd1, 27'h00000179, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000031b, 4'd14, 27'h00000345, 4'd6, 27'h000003cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000306, 4'd14, 27'h00000155, 4'd12, 27'h00000112, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002a9, 4'd2, 27'h00000082, 4'd4, 27'h00000226, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002d0, 4'd3, 27'h0000005b, 4'd9, 27'h000001a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000033f, 4'd4, 27'h0000036b, 4'd14, 27'h00000363, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000332, 4'd6, 27'h00000250, 4'd3, 27'h000001d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000067, 4'd7, 27'h000003de, 4'd7, 27'h00000380, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000256, 4'd5, 27'h00000134, 4'd11, 27'h00000286, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002d2, 4'd12, 27'h0000006e, 4'd4, 27'h000001ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000246, 4'd11, 27'h0000038c, 4'd9, 27'h000000a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003af, 4'd10, 27'h000003d0, 4'd12, 27'h0000002d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000110, 4'd2, 27'h000003ae, 4'd4, 27'h000002a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000d7, 4'd4, 27'h000002f0, 4'd8, 27'h0000032a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000074, 4'd2, 27'h000002fb, 4'd11, 27'h00000321, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000354, 4'd7, 27'h000001af, 4'd1, 27'h00000028, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000002c, 4'd5, 27'h000002de, 4'd9, 27'h000003a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000ae, 4'd9, 27'h0000039d, 4'd13, 27'h000000a0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000011c, 4'd12, 27'h0000020d, 4'd1, 27'h00000284, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000121, 4'd14, 27'h00000279, 4'd7, 27'h000003aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c3, 4'd13, 27'h000003f5, 4'd13, 27'h0000016a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ce, 4'd4, 27'h00000314, 4'd0, 27'h00000002, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b2, 4'd4, 27'h0000004a, 4'd8, 27'h0000004a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002a2, 4'd3, 27'h0000036b, 4'd12, 27'h000002d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000021f, 4'd7, 27'h0000003f, 4'd1, 27'h00000165, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000048, 4'd8, 27'h0000010c, 4'd8, 27'h000001fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002fe, 4'd8, 27'h00000281, 4'd14, 27'h0000027d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003e0, 4'd11, 27'h00000284, 4'd2, 27'h000000d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002f5, 4'd10, 27'h000000b4, 4'd5, 27'h000002bb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000375, 4'd13, 27'h000003e0, 4'd13, 27'h000001e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001ff, 4'd0, 27'h000000b9, 4'd2, 27'h000003fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000001f, 4'd3, 27'h000002ef, 4'd5, 27'h000003ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000014f, 4'd0, 27'h0000012d, 4'd11, 27'h00000102, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000345, 4'd8, 27'h000002b1, 4'd4, 27'h000003e4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003bd, 4'd7, 27'h000000e8, 4'd5, 27'h000002a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000381, 4'd9, 27'h00000246, 4'd11, 27'h00000288, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000ec, 4'd11, 27'h00000275, 4'd0, 27'h00000078, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e5, 4'd13, 27'h000003f2, 4'd9, 27'h000000e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000377, 4'd12, 27'h00000146, 4'd10, 27'h0000019b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000382, 4'd0, 27'h0000012b, 4'd2, 27'h00000010, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000390, 4'd1, 27'h00000375, 4'd8, 27'h0000003b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000b8, 4'd2, 27'h0000009c, 4'd12, 27'h0000002f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000006a, 4'd9, 27'h000000fa, 4'd4, 27'h0000033f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000028d, 4'd6, 27'h000003e7, 4'd9, 27'h000001ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000021b, 4'd5, 27'h00000353, 4'd12, 27'h000001be, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001f8, 4'd12, 27'h00000305, 4'd0, 27'h000001d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000399, 4'd14, 27'h00000309, 4'd6, 27'h0000033d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000b3, 4'd11, 27'h000002ef, 4'd11, 27'h00000003, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000337, 4'd3, 27'h0000013f, 4'd1, 27'h000003b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000360, 4'd1, 27'h00000246, 4'd5, 27'h000002d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002b1, 4'd4, 27'h00000300, 4'd14, 27'h000000d7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000122, 4'd8, 27'h000002e9, 4'd4, 27'h000000f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000227, 4'd9, 27'h0000018e, 4'd6, 27'h000003cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001fb, 4'd9, 27'h000003cc, 4'd13, 27'h000002d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000026e, 4'd13, 27'h0000019d, 4'd2, 27'h000001b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000359, 4'd12, 27'h00000351, 4'd8, 27'h000001d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001e4, 4'd11, 27'h000002db, 4'd10, 27'h0000023a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002de, 4'd3, 27'h00000199, 4'd0, 27'h0000010a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000035c, 4'd3, 27'h0000011d, 4'd5, 27'h000002d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003e3, 4'd2, 27'h00000198, 4'd11, 27'h00000053, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000008e, 4'd6, 27'h0000006f, 4'd1, 27'h000002db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003e4, 4'd6, 27'h000002c1, 4'd7, 27'h000000e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001c3, 4'd6, 27'h0000021c, 4'd14, 27'h000003af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001c7, 4'd13, 27'h000003a8, 4'd3, 27'h00000266, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002a4, 4'd11, 27'h00000033, 4'd9, 27'h000002f6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003ec, 4'd10, 27'h000001d9, 4'd10, 27'h00000130, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000285, 4'd2, 27'h00000044, 4'd1, 27'h00000192, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003c2, 4'd2, 27'h00000139, 4'd8, 27'h000003aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000357, 4'd4, 27'h000003ea, 4'd11, 27'h0000021d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000fb, 4'd6, 27'h000001cb, 4'd1, 27'h00000386, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000fe, 4'd5, 27'h0000000e, 4'd5, 27'h00000184, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000261, 4'd6, 27'h00000257, 4'd10, 27'h00000016, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001b1, 4'd14, 27'h000002c0, 4'd0, 27'h000003ee, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000239, 4'd10, 27'h0000034f, 4'd8, 27'h00000397, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001eb, 4'd11, 27'h000001b7, 4'd12, 27'h000003d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001d4, 4'd4, 27'h0000010f, 4'd4, 27'h00000324, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000250, 4'd1, 27'h0000006a, 4'd5, 27'h00000124, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000016, 4'd2, 27'h000001c4, 4'd11, 27'h000001a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000346, 4'd6, 27'h00000354, 4'd1, 27'h00000271, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000385, 4'd7, 27'h000001c6, 4'd5, 27'h000001b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000292, 4'd7, 27'h000002b7, 4'd13, 27'h000000f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000263, 4'd13, 27'h00000358, 4'd0, 27'h00000247, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000140, 4'd13, 27'h00000183, 4'd9, 27'h0000008e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003a0, 4'd13, 27'h00000075, 4'd14, 27'h000000f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000ae, 4'd0, 27'h000003e5, 4'd3, 27'h000000fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000d2, 4'd3, 27'h0000008c, 4'd5, 27'h000000e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001d7, 4'd2, 27'h0000021c, 4'd11, 27'h0000015e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000036f, 4'd7, 27'h000001d7, 4'd3, 27'h0000020f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000d4, 4'd9, 27'h0000039f, 4'd9, 27'h000003ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000160, 4'd7, 27'h00000383, 4'd14, 27'h00000153, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000018c, 4'd14, 27'h000003c9, 4'd2, 27'h000002bb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000367, 4'd14, 27'h0000035a, 4'd7, 27'h00000363, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003a2, 4'd11, 27'h0000020f, 4'd10, 27'h00000324, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000019a, 4'd2, 27'h00000216, 4'd3, 27'h000001eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003bb, 4'd3, 27'h00000067, 4'd5, 27'h0000011e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000028c, 4'd3, 27'h00000256, 4'd10, 27'h0000026f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001d6, 4'd5, 27'h000001d7, 4'd3, 27'h00000134, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000315, 4'd7, 27'h000001ea, 4'd5, 27'h0000009c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003c4, 4'd7, 27'h000002b0, 4'd11, 27'h000001bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000290, 4'd12, 27'h0000036d, 4'd1, 27'h000001ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000035f, 4'd12, 27'h00000140, 4'd5, 27'h000001dd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000f4, 4'd14, 27'h00000269, 4'd10, 27'h00000177, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000277, 4'd0, 27'h000001c2, 4'd0, 27'h000002c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000025c, 4'd0, 27'h000001fb, 4'd7, 27'h000001b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000161, 4'd4, 27'h0000021c, 4'd12, 27'h00000068, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003f8, 4'd6, 27'h0000012f, 4'd2, 27'h000001b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ce, 4'd7, 27'h0000020c, 4'd9, 27'h0000028b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000220, 4'd9, 27'h00000115, 4'd11, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000002, 4'd12, 27'h00000005, 4'd0, 27'h000002db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000118, 4'd12, 27'h00000260, 4'd6, 27'h00000285, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001f1, 4'd11, 27'h000003b2, 4'd11, 27'h00000357, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000006d, 4'd4, 27'h00000187, 4'd3, 27'h00000202, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000000d, 4'd1, 27'h00000179, 4'd6, 27'h00000193, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000e0, 4'd2, 27'h0000002f, 4'd12, 27'h0000018e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000329, 4'd7, 27'h000001eb, 4'd1, 27'h0000004e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000025c, 4'd6, 27'h0000015e, 4'd5, 27'h000002b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000329, 4'd5, 27'h0000000d, 4'd11, 27'h000001e8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000129, 4'd13, 27'h00000312, 4'd0, 27'h0000017e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000027, 4'd14, 27'h00000238, 4'd9, 27'h00000123, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001ba, 4'd14, 27'h0000022e, 4'd10, 27'h00000396, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000068, 4'd4, 27'h000000e5, 4'd4, 27'h000002c0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000088, 4'd2, 27'h0000007b, 4'd7, 27'h00000384, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000148, 4'd2, 27'h0000024e, 4'd13, 27'h00000330, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000002c, 4'd9, 27'h000001bf, 4'd4, 27'h000001bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003f8, 4'd8, 27'h0000033c, 4'd7, 27'h00000260, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002ed, 4'd6, 27'h000002fa, 4'd11, 27'h00000010, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000128, 4'd14, 27'h000002f4, 4'd3, 27'h000001e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003af, 4'd10, 27'h00000179, 4'd6, 27'h00000274, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000027c, 4'd13, 27'h0000039b, 4'd14, 27'h00000281, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000011e, 4'd3, 27'h000000ee, 4'd2, 27'h00000346, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002a7, 4'd4, 27'h000002fc, 4'd5, 27'h00000085, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000142, 4'd0, 27'h00000226, 4'd11, 27'h00000259, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000350, 4'd8, 27'h00000154, 4'd3, 27'h00000161, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000024d, 4'd6, 27'h000002cf, 4'd7, 27'h00000381, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000325, 4'd7, 27'h000003c7, 4'd10, 27'h00000277, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000bf, 4'd10, 27'h0000011e, 4'd1, 27'h000001a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000100, 4'd10, 27'h00000021, 4'd7, 27'h000003bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000107, 4'd13, 27'h000002a9, 4'd14, 27'h000003dd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000dd, 4'd2, 27'h000001fe, 4'd1, 27'h00000097, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002e4, 4'd4, 27'h000000ff, 4'd7, 27'h00000384, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000013, 4'd1, 27'h00000140, 4'd13, 27'h00000099, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001e6, 4'd7, 27'h00000366, 4'd4, 27'h000001ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000175, 4'd6, 27'h000002c2, 4'd5, 27'h0000003a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003c8, 4'd9, 27'h00000207, 4'd14, 27'h00000055, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001c5, 4'd11, 27'h000002ce, 4'd4, 27'h000000ca, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000336, 4'd11, 27'h000001fd, 4'd8, 27'h00000245, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001b3, 4'd12, 27'h00000021, 4'd14, 27'h00000029, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000129, 4'd4, 27'h0000016a, 4'd3, 27'h000002d9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000f6, 4'd2, 27'h00000033, 4'd5, 27'h0000026d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000248, 4'd4, 27'h00000079, 4'd11, 27'h0000004c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000093, 4'd5, 27'h0000009d, 4'd4, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000003a, 4'd6, 27'h0000013a, 4'd5, 27'h00000399, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000013c, 4'd7, 27'h000003e4, 4'd11, 27'h000002e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001bd, 4'd14, 27'h00000156, 4'd4, 27'h00000317, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003dd, 4'd12, 27'h0000035f, 4'd8, 27'h00000099, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000341, 4'd10, 27'h00000364, 4'd14, 27'h000002fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000e5, 4'd3, 27'h00000028, 4'd3, 27'h0000026d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001b6, 4'd4, 27'h000000ab, 4'd5, 27'h000003d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000182, 4'd0, 27'h00000260, 4'd14, 27'h0000027d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000336, 4'd9, 27'h000002c9, 4'd1, 27'h00000392, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000170, 4'd6, 27'h000003c9, 4'd9, 27'h0000034e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000252, 4'd9, 27'h000001db, 4'd14, 27'h000000d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000179, 4'd13, 27'h000003bc, 4'd2, 27'h0000015c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000108, 4'd12, 27'h0000018e, 4'd6, 27'h000001b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000329, 4'd11, 27'h000000cf, 4'd11, 27'h00000137, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000319, 4'd2, 27'h00000137, 4'd0, 27'h00000299, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000074, 4'd0, 27'h00000364, 4'd6, 27'h00000151, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000025e, 4'd0, 27'h000001f2, 4'd14, 27'h000000dc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003e5, 4'd7, 27'h00000343, 4'd4, 27'h00000379, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001eb, 4'd8, 27'h00000393, 4'd8, 27'h0000024e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000000a, 4'd5, 27'h0000037c, 4'd12, 27'h00000204, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000015c, 4'd11, 27'h0000001f, 4'd1, 27'h000000cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000027e, 4'd13, 27'h000000a5, 4'd6, 27'h00000035, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000038b, 4'd11, 27'h00000158, 4'd11, 27'h00000233, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000386, 4'd0, 27'h0000035a, 4'd1, 27'h0000009b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000b6, 4'd1, 27'h0000005c, 4'd9, 27'h000001f1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000037f, 4'd3, 27'h0000008b, 4'd13, 27'h000001a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000008b, 4'd6, 27'h00000176, 4'd0, 27'h000002c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000381, 4'd6, 27'h000001ff, 4'd8, 27'h00000156, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000092, 4'd5, 27'h0000030d, 4'd12, 27'h00000224, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002cb, 4'd13, 27'h00000288, 4'd4, 27'h0000014a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000217, 4'd12, 27'h000000d0, 4'd7, 27'h000001f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000005, 4'd14, 27'h000002dd, 4'd14, 27'h00000095, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000098, 4'd1, 27'h000003e1, 4'd1, 27'h000001c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000fd, 4'd1, 27'h000001ed, 4'd8, 27'h0000019b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000036c, 4'd4, 27'h00000324, 4'd12, 27'h00000156, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000299, 4'd8, 27'h00000088, 4'd4, 27'h000000b4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000023, 4'd7, 27'h000002ed, 4'd7, 27'h000002bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000238, 4'd8, 27'h0000018b, 4'd12, 27'h0000031c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000027f, 4'd14, 27'h0000008f, 4'd3, 27'h00000395, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002a4, 4'd14, 27'h000003f0, 4'd7, 27'h000002e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000022b, 4'd11, 27'h00000270, 4'd14, 27'h000000fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000110, 4'd3, 27'h00000243, 4'd3, 27'h0000004c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003fb, 4'd2, 27'h00000259, 4'd8, 27'h000003ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001a2, 4'd3, 27'h000002d1, 4'd11, 27'h000001e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000104, 4'd7, 27'h00000213, 4'd1, 27'h000002ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a1, 4'd9, 27'h00000087, 4'd7, 27'h00000331, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001fe, 4'd8, 27'h00000283, 4'd13, 27'h0000024b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000031, 4'd13, 27'h000000be, 4'd4, 27'h0000012a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001dd, 4'd10, 27'h000002d2, 4'd7, 27'h00000278, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000fa, 4'd11, 27'h00000006, 4'd11, 27'h00000053, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003d7, 4'd4, 27'h00000375, 4'd2, 27'h00000321, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002cb, 4'd4, 27'h000000d8, 4'd5, 27'h000002d7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000000e, 4'd2, 27'h00000268, 4'd14, 27'h000000ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000193, 4'd6, 27'h0000010d, 4'd2, 27'h000003ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000000e, 4'd5, 27'h00000007, 4'd6, 27'h0000001a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001f1, 4'd7, 27'h000001e8, 4'd10, 27'h0000014b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000329, 4'd10, 27'h000002cd, 4'd3, 27'h00000080, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000255, 4'd14, 27'h00000026, 4'd6, 27'h0000011f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001f9, 4'd14, 27'h0000019b, 4'd11, 27'h00000199, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000021e, 4'd2, 27'h0000027d, 4'd3, 27'h000003d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000062, 4'd2, 27'h00000083, 4'd7, 27'h00000212, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000ac, 4'd1, 27'h0000003a, 4'd13, 27'h000000de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000017f, 4'd5, 27'h000000fa, 4'd3, 27'h00000258, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002b8, 4'd6, 27'h0000016b, 4'd9, 27'h000000d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003fc, 4'd6, 27'h0000018a, 4'd13, 27'h000000f1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000006e, 4'd11, 27'h00000248, 4'd0, 27'h00000219, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001a6, 4'd12, 27'h0000007a, 4'd6, 27'h000003c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000003, 4'd10, 27'h000001c8, 4'd12, 27'h000001ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001f9, 4'd2, 27'h00000127, 4'd0, 27'h000000fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000033c, 4'd1, 27'h00000179, 4'd6, 27'h00000028, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000197, 4'd2, 27'h0000003c, 4'd10, 27'h00000201, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001e4, 4'd5, 27'h000002cc, 4'd1, 27'h00000308, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000310, 4'd6, 27'h00000259, 4'd6, 27'h000000f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000085, 4'd7, 27'h000002d7, 4'd13, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000025f, 4'd13, 27'h00000334, 4'd0, 27'h000003c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000026f, 4'd13, 27'h00000047, 4'd6, 27'h000001d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000064, 4'd10, 27'h00000044, 4'd11, 27'h00000145, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000303, 4'd4, 27'h00000372, 4'd2, 27'h0000032f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000010a, 4'd1, 27'h000000dd, 4'd6, 27'h0000022d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003f6, 4'd4, 27'h0000011d, 4'd13, 27'h0000027f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000018b, 4'd7, 27'h0000009d, 4'd1, 27'h00000210, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000264, 4'd8, 27'h00000347, 4'd5, 27'h00000372, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000015, 4'd5, 27'h000001ae, 4'd10, 27'h00000219, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000034e, 4'd10, 27'h000002dd, 4'd0, 27'h00000339, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000032a, 4'd11, 27'h00000056, 4'd8, 27'h00000364, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003b5, 4'd10, 27'h000000ca, 4'd12, 27'h00000255, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002be, 4'd1, 27'h00000279, 4'd1, 27'h000002c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000013c, 4'd3, 27'h00000227, 4'd9, 27'h000002a7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000036a, 4'd0, 27'h000002c9, 4'd12, 27'h000002d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000038a, 4'd5, 27'h000001e4, 4'd4, 27'h000003d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000348, 4'd5, 27'h0000004f, 4'd6, 27'h000001fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000d2, 4'd9, 27'h0000004f, 4'd10, 27'h00000286, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003d9, 4'd12, 27'h000001d3, 4'd2, 27'h00000151, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000043, 4'd11, 27'h0000014e, 4'd7, 27'h0000013c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003d8, 4'd13, 27'h0000020e, 4'd10, 27'h000003d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000341, 4'd0, 27'h000002af, 4'd4, 27'h000000c0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000001b, 4'd1, 27'h00000153, 4'd6, 27'h000001f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003dd, 4'd2, 27'h000000c3, 4'd11, 27'h0000018e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000020b, 4'd6, 27'h00000277, 4'd0, 27'h000001cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000140, 4'd5, 27'h000001e4, 4'd9, 27'h000001e2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000302, 4'd7, 27'h00000391, 4'd11, 27'h0000014f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000279, 4'd11, 27'h000003b3, 4'd3, 27'h0000002e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e1, 4'd14, 27'h000001b9, 4'd8, 27'h0000036d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002c8, 4'd10, 27'h0000006a, 4'd12, 27'h000001c0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000df, 4'd1, 27'h000000b7, 4'd0, 27'h0000031e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000ad, 4'd2, 27'h00000135, 4'd6, 27'h000002f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001bc, 4'd0, 27'h000000a4, 4'd12, 27'h00000197, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000038b, 4'd6, 27'h000001b1, 4'd4, 27'h000001cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003ba, 4'd9, 27'h000002cb, 4'd9, 27'h000001a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000222, 4'd9, 27'h00000378, 4'd12, 27'h000003af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000036d, 4'd12, 27'h000001de, 4'd3, 27'h000000bc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000342, 4'd13, 27'h00000064, 4'd7, 27'h000003bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000004f, 4'd10, 27'h0000017c, 4'd14, 27'h0000005e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000253, 4'd2, 27'h00000105, 4'd2, 27'h000003b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000023a, 4'd0, 27'h00000321, 4'd8, 27'h00000055, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003d7, 4'd3, 27'h0000010a, 4'd11, 27'h0000007e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003d2, 4'd6, 27'h0000012d, 4'd4, 27'h00000086, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000cb, 4'd8, 27'h000001a6, 4'd8, 27'h00000002, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003fa, 4'd6, 27'h00000228, 4'd11, 27'h00000000, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000022d, 4'd10, 27'h00000095, 4'd2, 27'h00000235, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000032, 4'd12, 27'h000001aa, 4'd7, 27'h000000d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000211, 4'd11, 27'h00000108, 4'd13, 27'h000000a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002f8, 4'd1, 27'h000001d3, 4'd4, 27'h000000ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000260, 4'd2, 27'h00000381, 4'd8, 27'h00000208, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000380, 4'd2, 27'h00000205, 4'd14, 27'h00000098, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000032d, 4'd5, 27'h00000204, 4'd2, 27'h000003fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ee, 4'd6, 27'h000001e0, 4'd7, 27'h000000f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000015b, 4'd9, 27'h000001c9, 4'd13, 27'h000002f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000002d, 4'd10, 27'h0000029e, 4'd1, 27'h00000043, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ef, 4'd10, 27'h00000128, 4'd5, 27'h000002c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000003d, 4'd10, 27'h00000212, 4'd13, 27'h0000019b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000022a, 4'd3, 27'h00000067, 4'd1, 27'h00000199, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000385, 4'd4, 27'h00000053, 4'd5, 27'h000002aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000027b, 4'd3, 27'h00000203, 4'd10, 27'h0000016c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000024f, 4'd6, 27'h00000131, 4'd3, 27'h0000031b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000109, 4'd6, 27'h00000073, 4'd7, 27'h0000016e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003e4, 4'd6, 27'h000003ed, 4'd12, 27'h0000034d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000036c, 4'd10, 27'h000001e4, 4'd2, 27'h00000009, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000099, 4'd11, 27'h00000080, 4'd8, 27'h00000259, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001bc, 4'd11, 27'h0000033e, 4'd11, 27'h000003da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000223, 4'd4, 27'h0000005e, 4'd2, 27'h00000022, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000027d, 4'd4, 27'h00000109, 4'd9, 27'h000000d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000352, 4'd4, 27'h00000393, 4'd11, 27'h0000014b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000006c, 4'd9, 27'h0000034e, 4'd4, 27'h00000070, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003e1, 4'd9, 27'h000002a5, 4'd8, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000011f, 4'd9, 27'h0000005e, 4'd13, 27'h000002b3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000356, 4'd13, 27'h00000104, 4'd1, 27'h0000022e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001b4, 4'd10, 27'h00000392, 4'd8, 27'h00000399, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000368, 4'd12, 27'h0000011f, 4'd13, 27'h00000018, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000259, 4'd3, 27'h000000da, 4'd3, 27'h00000090, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002d8, 4'd0, 27'h00000343, 4'd5, 27'h00000162, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000004, 4'd4, 27'h00000010, 4'd14, 27'h000002af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000378, 4'd9, 27'h00000053, 4'd4, 27'h000001ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000348, 4'd5, 27'h00000003, 4'd8, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000dd, 4'd5, 27'h000001a2, 4'd14, 27'h00000015, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000037f, 4'd13, 27'h00000133, 4'd0, 27'h000002f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000f2, 4'd13, 27'h00000396, 4'd8, 27'h00000041, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000010e, 4'd13, 27'h000002a5, 4'd10, 27'h00000143, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000033f, 4'd3, 27'h00000365, 4'd1, 27'h0000025e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002d6, 4'd4, 27'h00000109, 4'd5, 27'h000003f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000dd, 4'd1, 27'h00000036, 4'd12, 27'h000001d4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002c1, 4'd7, 27'h00000371, 4'd1, 27'h000003d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001ee, 4'd8, 27'h000002af, 4'd9, 27'h00000105, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000054, 4'd7, 27'h000003c6, 4'd13, 27'h00000112, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000020e, 4'd12, 27'h0000012f, 4'd0, 27'h000000a7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002ae, 4'd13, 27'h0000026e, 4'd6, 27'h0000028e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000033b, 4'd14, 27'h00000309, 4'd12, 27'h00000327, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000027f, 4'd3, 27'h0000001a, 4'd0, 27'h0000035f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000267, 4'd1, 27'h00000163, 4'd6, 27'h000003ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000f9, 4'd1, 27'h000001a9, 4'd12, 27'h0000034e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000037, 4'd5, 27'h000003a2, 4'd4, 27'h00000259, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003ba, 4'd7, 27'h000002ad, 4'd9, 27'h000002bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001ab, 4'd7, 27'h000001db, 4'd14, 27'h000001b0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000281, 4'd11, 27'h000003f1, 4'd4, 27'h000001c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000cd, 4'd10, 27'h00000116, 4'd7, 27'h00000101, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000011c, 4'd12, 27'h0000029d, 4'd13, 27'h000001d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000032a, 4'd0, 27'h00000069, 4'd0, 27'h00000182, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000b2, 4'd3, 27'h00000336, 4'd7, 27'h00000159, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000035b, 4'd2, 27'h00000200, 4'd13, 27'h000003d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000001b, 4'd6, 27'h0000024b, 4'd3, 27'h000002a7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001f1, 4'd8, 27'h000000a6, 4'd6, 27'h00000107, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003bf, 4'd9, 27'h0000018e, 4'd11, 27'h00000087, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000323, 4'd12, 27'h0000007c, 4'd2, 27'h000003a2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002b1, 4'd14, 27'h000001cf, 4'd8, 27'h000002d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000023f, 4'd11, 27'h0000028b, 4'd13, 27'h000001f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000ae, 4'd1, 27'h000003c1, 4'd1, 27'h00000327, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001a1, 4'd0, 27'h00000276, 4'd6, 27'h0000003e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001f8, 4'd1, 27'h0000011f, 4'd12, 27'h00000119, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000008f, 4'd8, 27'h00000258, 4'd0, 27'h00000200, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000281, 4'd6, 27'h000003f7, 4'd7, 27'h00000183, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000086, 4'd8, 27'h00000360, 4'd12, 27'h000001cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000367, 4'd14, 27'h00000228, 4'd1, 27'h00000199, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000211, 4'd10, 27'h0000020d, 4'd9, 27'h00000326, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001fd, 4'd12, 27'h0000022e, 4'd12, 27'h0000020a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003a0, 4'd3, 27'h00000090, 4'd2, 27'h000002e0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000274, 4'd1, 27'h0000003c, 4'd8, 27'h000002e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000045, 4'd3, 27'h000000a0, 4'd10, 27'h00000038, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000012, 4'd6, 27'h000002f3, 4'd3, 27'h00000166, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000015, 4'd9, 27'h00000320, 4'd9, 27'h000000d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000277, 4'd7, 27'h00000318, 4'd14, 27'h000002b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000c8, 4'd10, 27'h000003cc, 4'd1, 27'h00000065, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000133, 4'd13, 27'h000000be, 4'd8, 27'h00000384, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002ff, 4'd13, 27'h00000215, 4'd12, 27'h0000024b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000016f, 4'd4, 27'h0000024f, 4'd1, 27'h000001cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e0, 4'd1, 27'h0000029a, 4'd6, 27'h000003ad, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001a5, 4'd1, 27'h000003ee, 4'd12, 27'h000000f6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000383, 4'd8, 27'h000000dc, 4'd4, 27'h000001fc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000283, 4'd7, 27'h0000001d, 4'd7, 27'h000000e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002d4, 4'd5, 27'h000001a0, 4'd12, 27'h0000004a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000196, 4'd13, 27'h00000151, 4'd1, 27'h0000030e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002a4, 4'd10, 27'h00000221, 4'd6, 27'h00000186, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000086, 4'd11, 27'h000002f3, 4'd10, 27'h0000034c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000106, 4'd1, 27'h00000336, 4'd0, 27'h00000215, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001fc, 4'd2, 27'h00000033, 4'd6, 27'h00000224, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000dc, 4'd0, 27'h000000f6, 4'd12, 27'h000000db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c9, 4'd6, 27'h00000277, 4'd0, 27'h00000208, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000184, 4'd8, 27'h0000037d, 4'd9, 27'h0000002b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000082, 4'd8, 27'h0000014f, 4'd10, 27'h0000017b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000a8, 4'd14, 27'h00000036, 4'd3, 27'h0000012c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000204, 4'd12, 27'h000001fb, 4'd5, 27'h00000010, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002a4, 4'd13, 27'h000002bc, 4'd11, 27'h0000023d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001ef, 4'd1, 27'h0000020d, 4'd4, 27'h000000a7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000093, 4'd4, 27'h000001ee, 4'd8, 27'h0000031a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000334, 4'd3, 27'h00000182, 4'd12, 27'h00000160, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000137, 4'd7, 27'h00000291, 4'd1, 27'h000000be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002f9, 4'd9, 27'h000003c9, 4'd5, 27'h0000009c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000093, 4'd7, 27'h000001d2, 4'd10, 27'h00000242, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001d3, 4'd11, 27'h00000365, 4'd3, 27'h000003dd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b7, 4'd10, 27'h00000070, 4'd6, 27'h000003b3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000319, 4'd13, 27'h000001dc, 4'd11, 27'h0000021f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000151, 4'd2, 27'h00000212, 4'd0, 27'h0000009f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000395, 4'd2, 27'h000002bb, 4'd8, 27'h0000013b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002bb, 4'd0, 27'h000002ec, 4'd14, 27'h00000042, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001b5, 4'd8, 27'h000003c5, 4'd4, 27'h000000c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000141, 4'd6, 27'h00000215, 4'd5, 27'h000001cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000f2, 4'd6, 27'h00000108, 4'd14, 27'h00000065, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000125, 4'd12, 27'h00000087, 4'd2, 27'h000002dc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001ab, 4'd10, 27'h00000354, 4'd7, 27'h0000024c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000030, 4'd12, 27'h0000002c, 4'd11, 27'h00000168, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000031b, 4'd1, 27'h00000014, 4'd2, 27'h0000009d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003a2, 4'd1, 27'h00000246, 4'd5, 27'h000003d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000b9, 4'd1, 27'h0000022a, 4'd13, 27'h0000018e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000037b, 4'd5, 27'h00000134, 4'd2, 27'h000001ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001a0, 4'd7, 27'h0000015b, 4'd9, 27'h000002da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000035a, 4'd9, 27'h00000106, 4'd13, 27'h000002df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000b1, 4'd10, 27'h000000de, 4'd1, 27'h00000336, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000001e, 4'd11, 27'h00000355, 4'd6, 27'h00000325, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003db, 4'd13, 27'h00000077, 4'd10, 27'h0000008f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001f7, 4'd1, 27'h000001bc, 4'd3, 27'h00000050, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b5, 4'd2, 27'h00000379, 4'd5, 27'h000000aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000000e, 4'd1, 27'h00000273, 4'd14, 27'h0000037e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000197, 4'd7, 27'h000003c5, 4'd4, 27'h0000011b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000264, 4'd8, 27'h00000372, 4'd5, 27'h000003d1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000011e, 4'd8, 27'h000001a9, 4'd10, 27'h000003a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000146, 4'd10, 27'h0000013c, 4'd0, 27'h00000146, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003fc, 4'd13, 27'h00000079, 4'd5, 27'h000001c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003f0, 4'd13, 27'h00000119, 4'd10, 27'h000001db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000fc, 4'd4, 27'h0000026b, 4'd0, 27'h000003c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000212, 4'd1, 27'h000001b8, 4'd6, 27'h000003fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000030b, 4'd0, 27'h00000045, 4'd11, 27'h00000053, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000019f, 4'd9, 27'h00000236, 4'd0, 27'h00000339, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000123, 4'd9, 27'h00000376, 4'd8, 27'h0000020c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002ce, 4'd9, 27'h00000221, 4'd13, 27'h000002c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000036a, 4'd14, 27'h00000391, 4'd4, 27'h00000310, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000107, 4'd12, 27'h00000335, 4'd7, 27'h0000027f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000001, 4'd13, 27'h00000363, 4'd12, 27'h0000003a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003be, 4'd4, 27'h0000016a, 4'd1, 27'h00000351, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000021e, 4'd3, 27'h000001de, 4'd8, 27'h00000367, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001c9, 4'd0, 27'h00000312, 4'd11, 27'h00000373, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000dc, 4'd7, 27'h000003aa, 4'd2, 27'h000003c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001f4, 4'd7, 27'h00000135, 4'd6, 27'h000002cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000023f, 4'd5, 27'h0000022e, 4'd14, 27'h00000344, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001b6, 4'd10, 27'h00000328, 4'd1, 27'h0000033b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002ba, 4'd11, 27'h00000032, 4'd7, 27'h00000222, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002ed, 4'd11, 27'h0000016e, 4'd10, 27'h00000073, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000380, 4'd1, 27'h000000a4, 4'd4, 27'h000003f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000069, 4'd4, 27'h00000192, 4'd7, 27'h0000003a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000015b, 4'd0, 27'h0000009a, 4'd11, 27'h00000029, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002ef, 4'd7, 27'h000003ea, 4'd3, 27'h000002e4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000350, 4'd5, 27'h00000022, 4'd7, 27'h00000225, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001e1, 4'd6, 27'h000001e9, 4'd13, 27'h000000ad, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000054, 4'd13, 27'h000002cf, 4'd4, 27'h00000054, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000095, 4'd14, 27'h00000104, 4'd9, 27'h0000023d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002c1, 4'd14, 27'h00000146, 4'd11, 27'h000001ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000184, 4'd3, 27'h000002c1, 4'd2, 27'h0000008c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003bd, 4'd2, 27'h000002da, 4'd6, 27'h000000d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000fd, 4'd3, 27'h000003df, 4'd13, 27'h00000250, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000179, 4'd8, 27'h0000014f, 4'd4, 27'h00000359, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000351, 4'd9, 27'h000002a2, 4'd9, 27'h00000012, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000234, 4'd7, 27'h0000000a, 4'd12, 27'h00000333, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000358, 4'd10, 27'h00000285, 4'd1, 27'h000001df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000189, 4'd10, 27'h00000279, 4'd8, 27'h00000366, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001d9, 4'd13, 27'h0000006e, 4'd11, 27'h000000af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001d2, 4'd2, 27'h00000165, 4'd2, 27'h000001c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000351, 4'd4, 27'h00000154, 4'd9, 27'h000002fc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000166, 4'd4, 27'h00000074, 4'd13, 27'h0000036a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003b3, 4'd8, 27'h000002fc, 4'd2, 27'h00000067, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ad, 4'd7, 27'h00000314, 4'd5, 27'h000002ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000022d, 4'd8, 27'h0000016f, 4'd11, 27'h000002ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000271, 4'd11, 27'h0000016e, 4'd1, 27'h00000005, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002ad, 4'd12, 27'h000001ac, 4'd9, 27'h00000272, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003ea, 4'd10, 27'h0000028c, 4'd13, 27'h00000219, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000023a, 4'd1, 27'h0000022f, 4'd4, 27'h0000039d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002ad, 4'd4, 27'h00000115, 4'd9, 27'h00000360, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000018c, 4'd1, 27'h0000032a, 4'd14, 27'h0000019d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000105, 4'd6, 27'h00000210, 4'd4, 27'h000000a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000096, 4'd9, 27'h00000123, 4'd8, 27'h0000014d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000de, 4'd5, 27'h0000014e, 4'd12, 27'h00000078, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000110, 4'd14, 27'h000001f8, 4'd3, 27'h000000d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000038b, 4'd13, 27'h00000083, 4'd7, 27'h000003f1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000266, 4'd13, 27'h00000290, 4'd11, 27'h00000117, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000e3, 4'd1, 27'h000001c6, 4'd0, 27'h0000024d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000313, 4'd3, 27'h0000024c, 4'd5, 27'h00000090, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002e7, 4'd4, 27'h00000204, 4'd13, 27'h000001a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000141, 4'd5, 27'h00000181, 4'd3, 27'h0000037d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000032d, 4'd8, 27'h00000069, 4'd8, 27'h00000094, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000216, 4'd6, 27'h00000249, 4'd10, 27'h0000024c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003a9, 4'd13, 27'h000001d2, 4'd4, 27'h000001f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001bc, 4'd10, 27'h0000016a, 4'd8, 27'h00000245, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000211, 4'd11, 27'h00000079, 4'd14, 27'h00000092, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000e7, 4'd0, 27'h00000322, 4'd2, 27'h00000135, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002f4, 4'd2, 27'h00000306, 4'd6, 27'h0000028c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000004b, 4'd0, 27'h000000b8, 4'd10, 27'h000001fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003a6, 4'd5, 27'h00000069, 4'd3, 27'h0000006b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000011, 4'd8, 27'h000001a6, 4'd8, 27'h000002f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001c0, 4'd6, 27'h00000237, 4'd14, 27'h00000038, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002c5, 4'd12, 27'h00000142, 4'd0, 27'h00000384, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000304, 4'd12, 27'h000003e3, 4'd5, 27'h00000271, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000024a, 4'd10, 27'h00000157, 4'd12, 27'h000003fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000b8, 4'd3, 27'h0000018f, 4'd2, 27'h000002ff, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003e3, 4'd1, 27'h000000ef, 4'd8, 27'h000000ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001b2, 4'd4, 27'h00000230, 4'd14, 27'h0000009f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000220, 4'd8, 27'h000002d0, 4'd3, 27'h000003d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000c1, 4'd6, 27'h00000135, 4'd9, 27'h0000028b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000332, 4'd5, 27'h0000025c, 4'd11, 27'h00000053, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000110, 4'd12, 27'h0000002d, 4'd0, 27'h000003d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000056, 4'd12, 27'h0000005b, 4'd5, 27'h0000017e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000029d, 4'd13, 27'h00000190, 4'd14, 27'h0000002a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000012f, 4'd0, 27'h000000f1, 4'd1, 27'h000003a3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000ba, 4'd4, 27'h0000010f, 4'd6, 27'h00000265, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001ad, 4'd3, 27'h0000026c, 4'd11, 27'h00000212, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002c2, 4'd6, 27'h000000ad, 4'd1, 27'h000000da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001e9, 4'd9, 27'h00000148, 4'd5, 27'h00000380, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000230, 4'd8, 27'h00000155, 4'd14, 27'h00000243, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000222, 4'd14, 27'h000000f7, 4'd4, 27'h00000032, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001d7, 4'd13, 27'h000002c8, 4'd6, 27'h0000019f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000000, 4'd11, 27'h000003b3, 4'd14, 27'h0000033a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000009c, 4'd0, 27'h000001e1, 4'd1, 27'h000001d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002ca, 4'd4, 27'h00000244, 4'd6, 27'h00000232, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003c3, 4'd2, 27'h00000128, 4'd10, 27'h00000015, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000ab, 4'd7, 27'h0000029b, 4'd0, 27'h00000031, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000039a, 4'd6, 27'h00000277, 4'd6, 27'h000002a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000012b, 4'd6, 27'h000002d1, 4'd14, 27'h000003c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000273, 4'd13, 27'h00000033, 4'd2, 27'h000003bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000021a, 4'd14, 27'h000002cf, 4'd9, 27'h000002ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000ff, 4'd12, 27'h00000164, 4'd12, 27'h0000032b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002e7, 4'd1, 27'h000003df, 4'd1, 27'h00000237, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000253, 4'd2, 27'h000001d0, 4'd6, 27'h00000289, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000261, 4'd1, 27'h000003e5, 4'd10, 27'h000000b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000014, 4'd5, 27'h00000114, 4'd0, 27'h00000126, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000217, 4'd7, 27'h000003e8, 4'd6, 27'h000002ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000396, 4'd8, 27'h000003a7, 4'd14, 27'h0000000b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000146, 4'd11, 27'h000000cd, 4'd4, 27'h00000066, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002e5, 4'd13, 27'h0000011e, 4'd7, 27'h00000339, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000033, 4'd11, 27'h0000031a, 4'd10, 27'h0000008f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003f6, 4'd0, 27'h00000070, 4'd4, 27'h00000188, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001b5, 4'd2, 27'h0000013b, 4'd7, 27'h00000029, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000103, 4'd3, 27'h000000fa, 4'd13, 27'h0000017a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002f5, 4'd7, 27'h000002cc, 4'd1, 27'h0000039a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000fc, 4'd9, 27'h0000004f, 4'd7, 27'h0000029b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001b2, 4'd8, 27'h00000339, 4'd12, 27'h00000164, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000187, 4'd10, 27'h000001ac, 4'd0, 27'h000001ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000298, 4'd10, 27'h00000309, 4'd8, 27'h00000253, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ed, 4'd14, 27'h00000321, 4'd11, 27'h0000000f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003a3, 4'd3, 27'h00000250, 4'd0, 27'h000002fb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000063, 4'd4, 27'h0000015a, 4'd5, 27'h00000348, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000195, 4'd3, 27'h00000064, 4'd14, 27'h0000017c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000039c, 4'd9, 27'h00000341, 4'd3, 27'h0000012f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000002, 4'd8, 27'h00000182, 4'd8, 27'h0000011f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000022, 4'd6, 27'h000002e1, 4'd13, 27'h00000208, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000029a, 4'd13, 27'h0000039c, 4'd0, 27'h0000020f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000024f, 4'd13, 27'h00000257, 4'd6, 27'h000000e9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000069, 4'd11, 27'h00000214, 4'd13, 27'h000001ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000004c, 4'd2, 27'h000002b5, 4'd0, 27'h000003c0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000012d, 4'd3, 27'h0000025c, 4'd5, 27'h0000036d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000048, 4'd4, 27'h0000020d, 4'd10, 27'h000003e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000225, 4'd6, 27'h00000113, 4'd2, 27'h000001ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003b2, 4'd5, 27'h0000016e, 4'd8, 27'h00000095, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000018, 4'd9, 27'h000001dc, 4'd10, 27'h000003f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000087, 4'd13, 27'h000001fe, 4'd4, 27'h0000034a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000369, 4'd10, 27'h000002ba, 4'd5, 27'h000002c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000034b, 4'd14, 27'h000002dc, 4'd10, 27'h000003d7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000026c, 4'd3, 27'h00000387, 4'd4, 27'h000003f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003c4, 4'd2, 27'h000003cf, 4'd8, 27'h000003ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000d9, 4'd0, 27'h0000023d, 4'd12, 27'h0000030a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003c9, 4'd5, 27'h0000004e, 4'd4, 27'h0000015f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000310, 4'd9, 27'h00000060, 4'd7, 27'h00000160, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000208, 4'd6, 27'h000002d1, 4'd13, 27'h000003d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001da, 4'd13, 27'h00000010, 4'd3, 27'h00000161, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003ee, 4'd14, 27'h00000120, 4'd5, 27'h000001b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003e7, 4'd13, 27'h00000077, 4'd12, 27'h00000163, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000052, 4'd3, 27'h00000229, 4'd1, 27'h000002ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003d7, 4'd4, 27'h00000145, 4'd8, 27'h000002d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002e9, 4'd3, 27'h000000af, 4'd11, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002b2, 4'd8, 27'h0000001e, 4'd3, 27'h00000202, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000290, 4'd6, 27'h00000171, 4'd7, 27'h000000ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000030b, 4'd9, 27'h000000dd, 4'd12, 27'h0000035a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000e1, 4'd12, 27'h00000234, 4'd4, 27'h0000028b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001a9, 4'd13, 27'h00000271, 4'd6, 27'h00000102, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000284, 4'd11, 27'h000002e6, 4'd13, 27'h00000346, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001f3, 4'd3, 27'h0000000f, 4'd0, 27'h000002f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000aa, 4'd0, 27'h000001c2, 4'd9, 27'h000003e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003e2, 4'd4, 27'h000000c7, 4'd14, 27'h00000264, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002bd, 4'd7, 27'h000002d5, 4'd0, 27'h000002bb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000000b, 4'd5, 27'h00000325, 4'd7, 27'h00000090, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000287, 4'd9, 27'h000001ce, 4'd11, 27'h00000339, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000113, 4'd13, 27'h000000f0, 4'd2, 27'h0000029f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000052, 4'd14, 27'h00000048, 4'd7, 27'h00000238, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000313, 4'd13, 27'h0000028b, 4'd11, 27'h000000b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002a7, 4'd0, 27'h000003ba, 4'd1, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000028c, 4'd4, 27'h000000a5, 4'd9, 27'h00000365, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000181, 4'd1, 27'h0000003d, 4'd13, 27'h00000216, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000381, 4'd9, 27'h00000322, 4'd1, 27'h00000245, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000140, 4'd6, 27'h000002ae, 4'd7, 27'h0000015c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002b9, 4'd7, 27'h00000353, 4'd14, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000000b, 4'd10, 27'h000000de, 4'd4, 27'h00000297, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000029e, 4'd12, 27'h000002cc, 4'd7, 27'h00000341, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000a4, 4'd10, 27'h000001b8, 4'd11, 27'h000000ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000145, 4'd4, 27'h000002da, 4'd1, 27'h000003fb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003b5, 4'd4, 27'h00000316, 4'd5, 27'h00000342, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000bd, 4'd0, 27'h0000006a, 4'd10, 27'h00000081, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000154, 4'd5, 27'h00000251, 4'd1, 27'h00000211, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000019b, 4'd6, 27'h00000320, 4'd5, 27'h0000034c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000d0, 4'd8, 27'h00000294, 4'd14, 27'h00000036, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000062, 4'd11, 27'h00000138, 4'd4, 27'h00000249, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000262, 4'd11, 27'h00000181, 4'd9, 27'h0000039e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000142, 4'd11, 27'h00000078, 4'd11, 27'h000002af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000ec, 4'd0, 27'h0000001e, 4'd3, 27'h00000292, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000013e, 4'd3, 27'h00000397, 4'd8, 27'h00000059, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003db, 4'd2, 27'h0000039c, 4'd11, 27'h0000033b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b3, 4'd8, 27'h00000289, 4'd1, 27'h000002b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000011c, 4'd6, 27'h00000362, 4'd9, 27'h00000396, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002f6, 4'd7, 27'h00000063, 4'd10, 27'h00000024, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000004f, 4'd14, 27'h000003f8, 4'd0, 27'h000001c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000274, 4'd11, 27'h000000b4, 4'd8, 27'h00000353, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003be, 4'd14, 27'h0000010b, 4'd13, 27'h000001a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000045, 4'd1, 27'h000001f0, 4'd4, 27'h000003a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000098, 4'd0, 27'h0000033b, 4'd8, 27'h00000105, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000214, 4'd3, 27'h00000050, 4'd10, 27'h000000cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000005d, 4'd7, 27'h00000157, 4'd3, 27'h00000240, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000187, 4'd5, 27'h000003c7, 4'd5, 27'h000003bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000196, 4'd8, 27'h00000025, 4'd14, 27'h000000d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000121, 4'd10, 27'h00000066, 4'd3, 27'h00000168, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000101, 4'd11, 27'h000002a7, 4'd6, 27'h000003a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000207, 4'd14, 27'h00000065, 4'd14, 27'h00000176, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000358, 4'd0, 27'h00000034, 4'd0, 27'h000003d8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000395, 4'd0, 27'h00000341, 4'd6, 27'h000000e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000394, 4'd2, 27'h000000c3, 4'd11, 27'h00000191, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000017c, 4'd9, 27'h00000174, 4'd2, 27'h000002ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000163, 4'd6, 27'h00000024, 4'd5, 27'h000001ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000015a, 4'd9, 27'h000003df, 4'd11, 27'h00000091, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000067, 4'd11, 27'h00000245, 4'd3, 27'h00000249, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001ef, 4'd13, 27'h00000285, 4'd5, 27'h0000003e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002d4, 4'd10, 27'h00000054, 4'd13, 27'h00000304, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000035a, 4'd2, 27'h000001e6, 4'd4, 27'h0000014d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b6, 4'd4, 27'h0000012b, 4'd7, 27'h000000df, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000232, 4'd2, 27'h000002d3, 4'd14, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000078, 4'd7, 27'h00000382, 4'd1, 27'h000002fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000038b, 4'd7, 27'h000003a0, 4'd9, 27'h0000016c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003de, 4'd5, 27'h000001e1, 4'd14, 27'h0000022d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001a8, 4'd12, 27'h00000166, 4'd3, 27'h00000019, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000297, 4'd12, 27'h0000003f, 4'd7, 27'h0000028d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000020d, 4'd10, 27'h0000031d, 4'd12, 27'h000000cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000137, 4'd0, 27'h00000186, 4'd4, 27'h000002e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000054, 4'd4, 27'h000002bd, 4'd8, 27'h00000307, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000275, 4'd2, 27'h00000165, 4'd10, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000039, 4'd8, 27'h000002c2, 4'd1, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000147, 4'd8, 27'h00000379, 4'd9, 27'h000000e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000045, 4'd8, 27'h0000000a, 4'd14, 27'h00000070, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001e6, 4'd11, 27'h00000195, 4'd3, 27'h0000030d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002e1, 4'd11, 27'h0000010d, 4'd9, 27'h00000074, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000025d, 4'd10, 27'h00000095, 4'd14, 27'h000001b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000336, 4'd4, 27'h00000272, 4'd0, 27'h000002f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000273, 4'd3, 27'h0000012c, 4'd5, 27'h000003d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001ad, 4'd4, 27'h00000080, 4'd10, 27'h000000fc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000353, 4'd6, 27'h00000129, 4'd0, 27'h0000011a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001a2, 4'd7, 27'h000000ea, 4'd9, 27'h000001bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003b2, 4'd9, 27'h00000165, 4'd12, 27'h000000e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003ba, 4'd11, 27'h0000010a, 4'd0, 27'h000000eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000006c, 4'd11, 27'h000003d1, 4'd7, 27'h00000393, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000102, 4'd13, 27'h0000031e, 4'd14, 27'h000002ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000f0, 4'd1, 27'h00000137, 4'd1, 27'h000003bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000039a, 4'd4, 27'h00000335, 4'd5, 27'h0000030f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001ff, 4'd0, 27'h000001b1, 4'd10, 27'h000000ed, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000033c, 4'd8, 27'h000003a0, 4'd3, 27'h00000309, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000031a, 4'd8, 27'h000000a4, 4'd9, 27'h0000009e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000004f, 4'd6, 27'h00000197, 4'd14, 27'h00000026, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000014d, 4'd13, 27'h0000019b, 4'd3, 27'h0000010c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000bd, 4'd10, 27'h00000275, 4'd5, 27'h00000252, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002cb, 4'd11, 27'h0000011a, 4'd14, 27'h00000319, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000108, 4'd3, 27'h000003e0, 4'd2, 27'h0000021b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000004, 4'd1, 27'h0000016b, 4'd6, 27'h00000243, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000192, 4'd3, 27'h00000262, 4'd10, 27'h00000221, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e7, 4'd9, 27'h00000006, 4'd4, 27'h000002a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002c5, 4'd6, 27'h00000315, 4'd9, 27'h00000021, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000ef, 4'd8, 27'h000003f2, 4'd14, 27'h000000d8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000028a, 4'd14, 27'h000002bd, 4'd3, 27'h0000019c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003a8, 4'd10, 27'h00000229, 4'd9, 27'h00000256, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000016, 4'd14, 27'h0000005d, 4'd11, 27'h000000f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000005b, 4'd4, 27'h000001ec, 4'd4, 27'h00000099, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002bf, 4'd0, 27'h0000027c, 4'd7, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002f6, 4'd0, 27'h000001e2, 4'd13, 27'h0000012c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000024f, 4'd9, 27'h000003a5, 4'd2, 27'h0000003d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000032f, 4'd6, 27'h0000024a, 4'd7, 27'h0000011f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000219, 4'd5, 27'h000002d0, 4'd13, 27'h000002d1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000ce, 4'd10, 27'h000001cc, 4'd1, 27'h000003b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002a0, 4'd14, 27'h00000168, 4'd5, 27'h00000139, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000e3, 4'd13, 27'h00000226, 4'd14, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003cc, 4'd2, 27'h00000230, 4'd0, 27'h00000001, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003f4, 4'd2, 27'h0000002b, 4'd5, 27'h0000009a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000153, 4'd0, 27'h00000290, 4'd13, 27'h000000d4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b1, 4'd9, 27'h000001e5, 4'd1, 27'h0000017f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000151, 4'd7, 27'h000002ee, 4'd8, 27'h00000288, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003ee, 4'd5, 27'h000002b2, 4'd12, 27'h0000010e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000364, 4'd14, 27'h00000009, 4'd3, 27'h000003f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000022, 4'd14, 27'h00000001, 4'd7, 27'h000003ca, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000047, 4'd12, 27'h000003c3, 4'd10, 27'h00000301, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000397, 4'd3, 27'h000003ec, 4'd3, 27'h000000a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000174, 4'd3, 27'h00000262, 4'd6, 27'h00000181, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000173, 4'd3, 27'h00000087, 4'd10, 27'h000001c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000146, 4'd9, 27'h000003c4, 4'd1, 27'h0000026b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000b9, 4'd9, 27'h0000035e, 4'd8, 27'h00000144, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001d6, 4'd6, 27'h000002e3, 4'd12, 27'h000000b0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000022d, 4'd11, 27'h000003f2, 4'd1, 27'h0000023b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000a9, 4'd13, 27'h000000d8, 4'd5, 27'h000001a4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000035b, 4'd11, 27'h0000015e, 4'd14, 27'h00000273, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000293, 4'd1, 27'h000000b1, 4'd0, 27'h00000042, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000156, 4'd0, 27'h0000017c, 4'd7, 27'h0000034b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000002c, 4'd0, 27'h0000021e, 4'd11, 27'h000001af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001ad, 4'd5, 27'h0000030f, 4'd1, 27'h0000033c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000029a, 4'd9, 27'h000002cb, 4'd6, 27'h0000021d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000e5, 4'd9, 27'h000003b2, 4'd14, 27'h00000077, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000005d, 4'd13, 27'h00000332, 4'd4, 27'h0000013f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000357, 4'd12, 27'h00000126, 4'd9, 27'h000001aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003df, 4'd14, 27'h00000295, 4'd13, 27'h000003e3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000ed, 4'd4, 27'h000002d9, 4'd1, 27'h0000024f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000025c, 4'd0, 27'h000001c5, 4'd7, 27'h0000018d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000004a, 4'd0, 27'h0000039c, 4'd13, 27'h000000a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003fb, 4'd8, 27'h00000272, 4'd1, 27'h00000375, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000262, 4'd5, 27'h00000163, 4'd5, 27'h0000006a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000250, 4'd5, 27'h00000393, 4'd10, 27'h0000021e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001f4, 4'd12, 27'h000003df, 4'd0, 27'h000001eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b6, 4'd12, 27'h00000148, 4'd9, 27'h00000299, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003aa, 4'd11, 27'h000002c0, 4'd13, 27'h000000bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a1, 4'd0, 27'h000003f8, 4'd3, 27'h0000030e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000242, 4'd2, 27'h00000092, 4'd8, 27'h00000181, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001c9, 4'd0, 27'h0000005f, 4'd13, 27'h000000aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000008f, 4'd5, 27'h000000e4, 4'd4, 27'h00000190, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000218, 4'd9, 27'h0000021f, 4'd6, 27'h00000221, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003c0, 4'd6, 27'h000002a2, 4'd11, 27'h0000036f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003bd, 4'd10, 27'h0000012b, 4'd1, 27'h0000016a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000275, 4'd14, 27'h000003b8, 4'd7, 27'h0000030b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000285, 4'd14, 27'h0000032a, 4'd13, 27'h00000373, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000017d, 4'd2, 27'h0000039c, 4'd0, 27'h0000006e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000295, 4'd4, 27'h00000121, 4'd5, 27'h000003b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000263, 4'd0, 27'h00000178, 4'd11, 27'h000003b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002df, 4'd7, 27'h0000036a, 4'd0, 27'h000003d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000029a, 4'd7, 27'h00000096, 4'd9, 27'h000001d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000004f, 4'd5, 27'h00000076, 4'd13, 27'h00000111, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000251, 4'd12, 27'h0000032f, 4'd2, 27'h000000eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000036b, 4'd13, 27'h0000026c, 4'd7, 27'h00000237, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000c8, 4'd12, 27'h0000007e, 4'd10, 27'h000000ee, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000018c, 4'd2, 27'h000001c4, 4'd3, 27'h0000035f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003a3, 4'd2, 27'h000003e7, 4'd8, 27'h000001be, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000da, 4'd0, 27'h0000027e, 4'd12, 27'h000003ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000002a, 4'd5, 27'h00000046, 4'd1, 27'h0000006b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000321, 4'd6, 27'h00000147, 4'd8, 27'h000000e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003ee, 4'd8, 27'h000001da, 4'd13, 27'h000003e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000245, 4'd12, 27'h00000099, 4'd1, 27'h00000206, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000017f, 4'd10, 27'h000003fe, 4'd6, 27'h00000372, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000030c, 4'd14, 27'h000000bf, 4'd13, 27'h0000019a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000357, 4'd0, 27'h00000074, 4'd0, 27'h00000166, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000238, 4'd1, 27'h00000336, 4'd8, 27'h00000212, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000275, 4'd2, 27'h00000143, 4'd10, 27'h00000105, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002a4, 4'd7, 27'h00000023, 4'd1, 27'h00000214, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000325, 4'd9, 27'h0000019c, 4'd6, 27'h00000094, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002af, 4'd5, 27'h0000036a, 4'd11, 27'h000000e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000005a, 4'd12, 27'h000001be, 4'd2, 27'h0000012f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000047, 4'd14, 27'h0000034f, 4'd7, 27'h000001c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000023d, 4'd10, 27'h00000190, 4'd13, 27'h0000031a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000211, 4'd0, 27'h0000006b, 4'd0, 27'h00000014, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000017b, 4'd4, 27'h000000b6, 4'd7, 27'h000000db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000009, 4'd2, 27'h00000090, 4'd13, 27'h0000004c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000002f, 4'd7, 27'h000003a6, 4'd2, 27'h000001d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001a4, 4'd6, 27'h0000025a, 4'd8, 27'h00000269, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002b5, 4'd5, 27'h000003ff, 4'd11, 27'h00000374, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002ce, 4'd10, 27'h000003cc, 4'd3, 27'h0000005e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000299, 4'd11, 27'h00000155, 4'd7, 27'h00000280, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000132, 4'd10, 27'h00000013, 4'd12, 27'h0000005f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000011b, 4'd4, 27'h00000034, 4'd3, 27'h00000179, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002ee, 4'd0, 27'h000002a1, 4'd8, 27'h00000118, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000028b, 4'd2, 27'h0000013e, 4'd10, 27'h0000038a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000122, 4'd7, 27'h000002ee, 4'd2, 27'h00000107, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000020, 4'd8, 27'h00000251, 4'd9, 27'h0000036e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003d9, 4'd7, 27'h00000337, 4'd13, 27'h000003b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000331, 4'd10, 27'h000000a0, 4'd3, 27'h00000398, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001e0, 4'd14, 27'h000000d2, 4'd9, 27'h00000016, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001a4, 4'd12, 27'h00000334, 4'd12, 27'h00000365, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002a3, 4'd3, 27'h000003c7, 4'd3, 27'h0000030b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003d5, 4'd1, 27'h000000fb, 4'd5, 27'h0000024b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000014c, 4'd2, 27'h000001d8, 4'd11, 27'h000001cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000019f, 4'd8, 27'h0000020e, 4'd4, 27'h0000039d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000054, 4'd9, 27'h000000ad, 4'd8, 27'h0000015e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000210, 4'd8, 27'h0000015e, 4'd11, 27'h0000001d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002f3, 4'd13, 27'h00000332, 4'd3, 27'h0000029a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000012e, 4'd10, 27'h0000039b, 4'd5, 27'h00000117, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000c0, 4'd13, 27'h000002d2, 4'd12, 27'h000001e4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000087, 4'd2, 27'h00000391, 4'd4, 27'h000002af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000296, 4'd1, 27'h00000259, 4'd6, 27'h00000184, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000af, 4'd0, 27'h000003bd, 4'd12, 27'h00000266, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001cd, 4'd8, 27'h00000259, 4'd0, 27'h000001bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000181, 4'd8, 27'h00000355, 4'd6, 27'h000001a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000203, 4'd6, 27'h00000190, 4'd12, 27'h000000ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002ea, 4'd12, 27'h0000005c, 4'd3, 27'h0000013d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000037b, 4'd12, 27'h000001e8, 4'd9, 27'h000003e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000005e, 4'd10, 27'h0000006b, 4'd12, 27'h000001d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000155, 4'd2, 27'h0000014c, 4'd4, 27'h00000254, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000cf, 4'd3, 27'h000002be, 4'd6, 27'h00000135, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000018f, 4'd0, 27'h000002e1, 4'd12, 27'h0000021d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000269, 4'd6, 27'h000003b0, 4'd1, 27'h000003d8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000345, 4'd8, 27'h000001fa, 4'd5, 27'h0000008a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000338, 4'd9, 27'h0000003c, 4'd10, 27'h00000150, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000f0, 4'd10, 27'h000003c3, 4'd2, 27'h000000ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002bd, 4'd13, 27'h000002df, 4'd8, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000122, 4'd13, 27'h000001c5, 4'd11, 27'h000001a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000038c, 4'd2, 27'h00000226, 4'd3, 27'h000000c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002a3, 4'd0, 27'h000000a8, 4'd9, 27'h00000254, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000004a, 4'd4, 27'h000002e4, 4'd10, 27'h000001f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002e1, 4'd8, 27'h0000014a, 4'd1, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003bd, 4'd5, 27'h0000023b, 4'd8, 27'h0000039f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a7, 4'd5, 27'h00000329, 4'd13, 27'h00000199, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000024, 4'd13, 27'h0000026a, 4'd3, 27'h000001a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000397, 4'd13, 27'h0000017c, 4'd7, 27'h00000229, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000b8, 4'd12, 27'h00000324, 4'd10, 27'h00000023, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000033a, 4'd2, 27'h0000008f, 4'd0, 27'h00000139, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002fe, 4'd2, 27'h000002d2, 4'd9, 27'h000002c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000204, 4'd3, 27'h000000d8, 4'd13, 27'h0000017d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003bb, 4'd7, 27'h0000011d, 4'd4, 27'h000002a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000035e, 4'd9, 27'h000000fd, 4'd7, 27'h00000179, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000357, 4'd6, 27'h000000a2, 4'd11, 27'h00000228, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000138, 4'd13, 27'h00000217, 4'd1, 27'h000003d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000032e, 4'd14, 27'h0000016a, 4'd9, 27'h0000028d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002cc, 4'd10, 27'h0000022f, 4'd11, 27'h00000130, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000178, 4'd0, 27'h00000299, 4'd1, 27'h000000d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000036e, 4'd4, 27'h000000b6, 4'd7, 27'h000000d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000024a, 4'd0, 27'h00000177, 4'd12, 27'h00000041, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001b7, 4'd6, 27'h00000285, 4'd4, 27'h0000033f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003c7, 4'd8, 27'h0000013c, 4'd6, 27'h00000003, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002d7, 4'd5, 27'h00000147, 4'd11, 27'h00000018, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000388, 4'd10, 27'h0000028c, 4'd3, 27'h000002a7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000191, 4'd12, 27'h00000291, 4'd6, 27'h00000200, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003e2, 4'd11, 27'h0000007f, 4'd13, 27'h000001c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000024c, 4'd0, 27'h00000090, 4'd2, 27'h00000346, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002fe, 4'd1, 27'h0000029c, 4'd7, 27'h0000011f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001da, 4'd2, 27'h00000281, 4'd12, 27'h00000322, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000021e, 4'd9, 27'h00000322, 4'd2, 27'h000001fc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003ab, 4'd7, 27'h0000014a, 4'd6, 27'h00000297, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000e7, 4'd5, 27'h0000035c, 4'd14, 27'h000003a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002ca, 4'd12, 27'h00000392, 4'd1, 27'h000002b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000150, 4'd10, 27'h00000128, 4'd8, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001b1, 4'd13, 27'h000001ec, 4'd14, 27'h0000004b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002e8, 4'd1, 27'h00000158, 4'd1, 27'h00000285, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000390, 4'd3, 27'h00000248, 4'd7, 27'h00000275, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003c0, 4'd1, 27'h00000000, 4'd12, 27'h00000086, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002ff, 4'd5, 27'h00000002, 4'd0, 27'h000003f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000382, 4'd7, 27'h000001f4, 4'd6, 27'h0000036c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000380, 4'd8, 27'h000003bf, 4'd12, 27'h00000041, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003cc, 4'd14, 27'h000001ff, 4'd4, 27'h0000025d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002cf, 4'd11, 27'h00000280, 4'd9, 27'h00000141, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000235, 4'd14, 27'h00000092, 4'd12, 27'h0000036b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000012c, 4'd1, 27'h000001fb, 4'd3, 27'h00000118, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000020b, 4'd4, 27'h00000358, 4'd6, 27'h00000104, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000213, 4'd1, 27'h0000028c, 4'd13, 27'h000001f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001da, 4'd9, 27'h00000274, 4'd1, 27'h000003ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000078, 4'd8, 27'h000001c4, 4'd9, 27'h000001c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000191, 4'd8, 27'h000002d5, 4'd13, 27'h0000000f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000013c, 4'd11, 27'h000002cb, 4'd4, 27'h0000024b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000ce, 4'd10, 27'h0000034d, 4'd8, 27'h000001bb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000023b, 4'd13, 27'h000002ac, 4'd10, 27'h000000fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002e5, 4'd1, 27'h000003c7, 4'd1, 27'h0000005f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000094, 4'd0, 27'h000003d5, 4'd9, 27'h000001c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002c4, 4'd3, 27'h000001e0, 4'd14, 27'h000002a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003fe, 4'd5, 27'h00000188, 4'd1, 27'h0000010b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002a2, 4'd5, 27'h000002f6, 4'd7, 27'h00000230, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000211, 4'd9, 27'h00000095, 4'd13, 27'h000000ba, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000038c, 4'd14, 27'h000000ac, 4'd0, 27'h00000023, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000039, 4'd12, 27'h0000000e, 4'd8, 27'h0000014e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000a4, 4'd14, 27'h00000054, 4'd11, 27'h0000018d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000018c, 4'd3, 27'h0000027c, 4'd1, 27'h000000ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000272, 4'd1, 27'h0000010f, 4'd7, 27'h000003d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000086, 4'd2, 27'h0000032d, 4'd12, 27'h000002f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000035a, 4'd6, 27'h00000121, 4'd4, 27'h000001f1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003a0, 4'd8, 27'h000000ce, 4'd5, 27'h000000ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002f7, 4'd9, 27'h0000003a, 4'd11, 27'h00000283, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000027e, 4'd11, 27'h00000009, 4'd2, 27'h000003ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000027a, 4'd11, 27'h000001fb, 4'd8, 27'h00000324, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000385, 4'd14, 27'h00000023, 4'd11, 27'h0000007f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000020, 4'd0, 27'h00000194, 4'd2, 27'h0000039a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000181, 4'd4, 27'h000001d3, 4'd6, 27'h00000335, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000380, 4'd1, 27'h00000390, 4'd11, 27'h00000342, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000028d, 4'd9, 27'h0000037c, 4'd0, 27'h0000035d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002f5, 4'd7, 27'h000000e8, 4'd9, 27'h00000322, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001fb, 4'd5, 27'h000002b9, 4'd12, 27'h0000032f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000331, 4'd11, 27'h0000012e, 4'd3, 27'h00000113, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000036b, 4'd12, 27'h00000297, 4'd9, 27'h000000b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000039b, 4'd12, 27'h0000017a, 4'd11, 27'h00000089, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000019c, 4'd3, 27'h000000e1, 4'd1, 27'h0000039d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001f5, 4'd1, 27'h00000004, 4'd5, 27'h00000191, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000d0, 4'd1, 27'h0000035c, 4'd13, 27'h000000bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000014e, 4'd7, 27'h000002df, 4'd4, 27'h0000005a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000268, 4'd7, 27'h0000014a, 4'd6, 27'h000003ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000147, 4'd7, 27'h000003c7, 4'd11, 27'h000003ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000237, 4'd14, 27'h00000120, 4'd2, 27'h00000373, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000138, 4'd11, 27'h00000078, 4'd8, 27'h00000280, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000202, 4'd13, 27'h000001e6, 4'd11, 27'h00000202, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000085, 4'd3, 27'h0000023d, 4'd3, 27'h00000123, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000273, 4'd1, 27'h0000012e, 4'd9, 27'h00000217, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000014, 4'd0, 27'h00000343, 4'd13, 27'h00000365, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000000c, 4'd5, 27'h00000065, 4'd2, 27'h00000216, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000034f, 4'd6, 27'h0000018b, 4'd8, 27'h000003db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003ea, 4'd9, 27'h00000318, 4'd10, 27'h00000241, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000020d, 4'd14, 27'h000000cc, 4'd2, 27'h000002e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000017, 4'd14, 27'h0000007d, 4'd5, 27'h0000020a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003ee, 4'd10, 27'h0000019f, 4'd11, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000d5, 4'd2, 27'h00000277, 4'd3, 27'h000000a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001f5, 4'd3, 27'h0000037c, 4'd5, 27'h000001a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003bd, 4'd3, 27'h0000015f, 4'd14, 27'h000001a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000014c, 4'd9, 27'h0000016e, 4'd1, 27'h00000278, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000009c, 4'd8, 27'h00000091, 4'd6, 27'h000001e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000232, 4'd8, 27'h000002d4, 4'd11, 27'h000002bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002c7, 4'd10, 27'h0000031b, 4'd1, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000035e, 4'd11, 27'h0000018c, 4'd5, 27'h00000145, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000010a, 4'd11, 27'h0000036a, 4'd14, 27'h00000314, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003ab, 4'd2, 27'h0000021b, 4'd3, 27'h0000028b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000033f, 4'd1, 27'h0000004f, 4'd7, 27'h00000122, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000391, 4'd0, 27'h00000207, 4'd14, 27'h00000350, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000015d, 4'd8, 27'h000002e7, 4'd4, 27'h000002e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ba, 4'd6, 27'h00000350, 4'd6, 27'h0000017f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000029d, 4'd7, 27'h000001ac, 4'd13, 27'h000002dd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000276, 4'd14, 27'h00000111, 4'd4, 27'h00000065, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000077, 4'd13, 27'h00000068, 4'd5, 27'h000003f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000017e, 4'd10, 27'h000003e7, 4'd10, 27'h000003fc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003a1, 4'd1, 27'h00000268, 4'd4, 27'h0000004c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003c2, 4'd3, 27'h0000032f, 4'd7, 27'h000001c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003fd, 4'd4, 27'h0000036d, 4'd11, 27'h00000118, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000039b, 4'd7, 27'h00000385, 4'd2, 27'h000003f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001c2, 4'd6, 27'h0000019f, 4'd6, 27'h000001f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000039c, 4'd8, 27'h00000220, 4'd13, 27'h00000292, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000130, 4'd13, 27'h00000111, 4'd2, 27'h00000082, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000085, 4'd14, 27'h000001d2, 4'd7, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002cb, 4'd11, 27'h0000037b, 4'd11, 27'h000001ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000025a, 4'd0, 27'h00000292, 4'd3, 27'h00000010, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003f1, 4'd2, 27'h000001da, 4'd9, 27'h0000006a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002ed, 4'd3, 27'h00000075, 4'd13, 27'h0000028c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002a9, 4'd9, 27'h0000039e, 4'd1, 27'h0000018f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000024, 4'd9, 27'h00000329, 4'd7, 27'h0000034b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000020b, 4'd5, 27'h000003f7, 4'd11, 27'h00000191, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000073, 4'd11, 27'h00000350, 4'd0, 27'h0000010c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001f3, 4'd13, 27'h0000021d, 4'd6, 27'h00000220, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000037a, 4'd14, 27'h00000229, 4'd13, 27'h00000205, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000389, 4'd0, 27'h0000013e, 4'd2, 27'h000003e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000017a, 4'd3, 27'h000002a8, 4'd9, 27'h00000336, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001b1, 4'd2, 27'h00000367, 4'd11, 27'h0000032a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000295, 4'd9, 27'h0000006c, 4'd2, 27'h000003f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000008b, 4'd6, 27'h00000278, 4'd7, 27'h000000e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002b7, 4'd6, 27'h000002c8, 4'd11, 27'h00000311, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000023, 4'd10, 27'h0000003a, 4'd2, 27'h000002fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000034c, 4'd13, 27'h000000b1, 4'd8, 27'h000000f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002ce, 4'd10, 27'h0000030a, 4'd14, 27'h0000036c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000259, 4'd1, 27'h000003e0, 4'd3, 27'h00000165, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000175, 4'd3, 27'h00000356, 4'd9, 27'h00000384, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000284, 4'd3, 27'h00000246, 4'd14, 27'h00000270, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000202, 4'd9, 27'h00000078, 4'd1, 27'h00000099, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000024d, 4'd8, 27'h000003b9, 4'd5, 27'h00000301, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000315, 4'd5, 27'h00000327, 4'd11, 27'h00000384, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001a0, 4'd12, 27'h0000013d, 4'd1, 27'h000001ef, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000395, 4'd10, 27'h00000323, 4'd5, 27'h000002ba, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000245, 4'd11, 27'h00000092, 4'd11, 27'h00000358, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000003, 4'd4, 27'h00000382, 4'd4, 27'h00000399, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003e7, 4'd2, 27'h0000015c, 4'd9, 27'h00000135, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000090, 4'd3, 27'h00000294, 4'd10, 27'h00000163, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b9, 4'd9, 27'h00000071, 4'd4, 27'h000002ca, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000248, 4'd5, 27'h0000021f, 4'd8, 27'h000001df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000275, 4'd6, 27'h000000bd, 4'd11, 27'h0000009f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002b5, 4'd13, 27'h00000107, 4'd1, 27'h00000260, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001c1, 4'd14, 27'h00000358, 4'd9, 27'h0000007e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000308, 4'd11, 27'h000000e8, 4'd12, 27'h00000241, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003a9, 4'd3, 27'h0000022e, 4'd1, 27'h000000d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000314, 4'd3, 27'h000001a5, 4'd8, 27'h0000032a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003c0, 4'd4, 27'h000001e2, 4'd14, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003ba, 4'd5, 27'h000000c9, 4'd4, 27'h000003b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000006b, 4'd9, 27'h000000c8, 4'd8, 27'h00000211, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000328, 4'd8, 27'h000000d0, 4'd10, 27'h00000107, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000006e, 4'd13, 27'h000000a9, 4'd4, 27'h000000d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000034, 4'd10, 27'h000003a0, 4'd6, 27'h00000178, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000383, 4'd12, 27'h00000370, 4'd10, 27'h000003a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000041, 4'd2, 27'h00000332, 4'd0, 27'h000001da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000065, 4'd1, 27'h0000033f, 4'd7, 27'h00000166, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002dd, 4'd3, 27'h000000cb, 4'd13, 27'h000000a4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000147, 4'd5, 27'h00000392, 4'd2, 27'h0000032f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000329, 4'd5, 27'h00000382, 4'd9, 27'h0000033a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000064, 4'd6, 27'h0000010b, 4'd10, 27'h00000384, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000056, 4'd13, 27'h00000387, 4'd1, 27'h00000398, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000ec, 4'd12, 27'h00000299, 4'd7, 27'h000003d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003ee, 4'd12, 27'h000002f0, 4'd10, 27'h0000002a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003af, 4'd3, 27'h0000027a, 4'd2, 27'h000002ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000299, 4'd1, 27'h000000c0, 4'd8, 27'h000003c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000e7, 4'd0, 27'h000001f5, 4'd12, 27'h000000b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b1, 4'd8, 27'h00000170, 4'd4, 27'h00000299, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000e0, 4'd5, 27'h000001fe, 4'd9, 27'h00000337, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001f8, 4'd5, 27'h00000009, 4'd11, 27'h00000108, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003e9, 4'd13, 27'h00000324, 4'd3, 27'h000000c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000365, 4'd13, 27'h000000ab, 4'd7, 27'h0000009a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000026b, 4'd11, 27'h0000034a, 4'd11, 27'h00000283, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001b2, 4'd1, 27'h00000213, 4'd3, 27'h00000198, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000236, 4'd4, 27'h0000017c, 4'd5, 27'h000000b5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000154, 4'd1, 27'h00000278, 4'd11, 27'h000003e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000024f, 4'd9, 27'h00000126, 4'd3, 27'h0000035e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000317, 4'd8, 27'h00000237, 4'd7, 27'h00000221, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003bf, 4'd9, 27'h00000029, 4'd13, 27'h0000016f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a8, 4'd14, 27'h000003f0, 4'd1, 27'h00000132, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001e9, 4'd11, 27'h000002a3, 4'd9, 27'h0000020c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002f9, 4'd10, 27'h00000040, 4'd12, 27'h0000001b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000058, 4'd1, 27'h000000c3, 4'd1, 27'h000000cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000020e, 4'd0, 27'h000000b9, 4'd6, 27'h000002cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001d7, 4'd3, 27'h000002bf, 4'd13, 27'h00000107, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002a0, 4'd5, 27'h00000065, 4'd1, 27'h0000000f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000002c, 4'd7, 27'h00000026, 4'd5, 27'h00000006, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000163, 4'd9, 27'h00000138, 4'd10, 27'h000002fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000372, 4'd12, 27'h000003b7, 4'd4, 27'h00000229, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000137, 4'd14, 27'h00000054, 4'd9, 27'h00000189, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000144, 4'd14, 27'h000000ae, 4'd10, 27'h00000319, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000fb, 4'd4, 27'h000002bb, 4'd4, 27'h000001cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000a0, 4'd1, 27'h0000000e, 4'd8, 27'h000000ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000fd, 4'd3, 27'h0000014b, 4'd11, 27'h00000117, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000117, 4'd8, 27'h00000052, 4'd4, 27'h00000012, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000036, 4'd6, 27'h0000024d, 4'd8, 27'h0000017b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000168, 4'd9, 27'h000002d5, 4'd10, 27'h00000176, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000017f, 4'd13, 27'h0000031a, 4'd1, 27'h000001ad, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000356, 4'd11, 27'h00000147, 4'd5, 27'h00000271, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003da, 4'd10, 27'h0000015d, 4'd10, 27'h000000fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000064, 4'd0, 27'h000003d6, 4'd0, 27'h000003cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000071, 4'd1, 27'h0000037e, 4'd9, 27'h000003d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e4, 4'd1, 27'h000000ed, 4'd13, 27'h0000016b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000023c, 4'd7, 27'h00000149, 4'd4, 27'h0000011c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000b4, 4'd9, 27'h000002ef, 4'd9, 27'h00000275, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000035b, 4'd9, 27'h0000000a, 4'd11, 27'h000001dc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002cc, 4'd10, 27'h00000393, 4'd3, 27'h0000036a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000014f, 4'd10, 27'h000003ce, 4'd6, 27'h0000001e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000204, 4'd11, 27'h000003ac, 4'd12, 27'h000002cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002dd, 4'd4, 27'h0000004b, 4'd1, 27'h000002e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003bf, 4'd4, 27'h00000070, 4'd8, 27'h00000216, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000130, 4'd3, 27'h0000007e, 4'd13, 27'h000003cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c6, 4'd7, 27'h0000009d, 4'd4, 27'h0000019a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000ee, 4'd5, 27'h000001f3, 4'd6, 27'h00000151, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002cf, 4'd7, 27'h00000171, 4'd13, 27'h00000163, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002f5, 4'd12, 27'h000000ff, 4'd1, 27'h000002a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001a3, 4'd11, 27'h000003e8, 4'd9, 27'h00000034, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000370, 4'd12, 27'h000000ed, 4'd12, 27'h00000206, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000c3, 4'd4, 27'h00000018, 4'd0, 27'h00000342, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002e3, 4'd4, 27'h0000024d, 4'd5, 27'h00000049, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000184, 4'd2, 27'h00000205, 4'd13, 27'h0000016d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000155, 4'd8, 27'h00000347, 4'd1, 27'h0000032e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002cb, 4'd5, 27'h0000015e, 4'd5, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000372, 4'd7, 27'h000001a1, 4'd12, 27'h000001b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001c8, 4'd13, 27'h00000395, 4'd4, 27'h00000141, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000007d, 4'd10, 27'h00000368, 4'd8, 27'h000003c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003f4, 4'd13, 27'h0000013d, 4'd11, 27'h0000000f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000009c, 4'd4, 27'h0000015e, 4'd1, 27'h000000e4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000395, 4'd1, 27'h00000202, 4'd5, 27'h0000011f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000029, 4'd1, 27'h00000306, 4'd14, 27'h000002b0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003c4, 4'd8, 27'h00000120, 4'd3, 27'h000000f6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003b4, 4'd7, 27'h00000126, 4'd7, 27'h0000026f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000172, 4'd6, 27'h00000197, 4'd13, 27'h0000013e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003d9, 4'd13, 27'h00000156, 4'd0, 27'h00000071, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000a2, 4'd14, 27'h00000287, 4'd7, 27'h000003b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003d5, 4'd13, 27'h00000196, 4'd13, 27'h00000345, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000214, 4'd3, 27'h00000170, 4'd0, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001e7, 4'd2, 27'h0000013e, 4'd5, 27'h000001e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000013, 4'd2, 27'h000001c5, 4'd13, 27'h00000142, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000060, 4'd7, 27'h000000b3, 4'd4, 27'h00000202, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003f1, 4'd7, 27'h00000222, 4'd7, 27'h0000037a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000025a, 4'd8, 27'h00000339, 4'd10, 27'h00000285, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000009e, 4'd13, 27'h00000111, 4'd0, 27'h000000fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002b0, 4'd12, 27'h00000322, 4'd8, 27'h000003f1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000027a, 4'd11, 27'h00000035, 4'd10, 27'h000003be, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000253, 4'd2, 27'h000003eb, 4'd0, 27'h00000044, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000b1, 4'd2, 27'h00000082, 4'd5, 27'h000000d7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001b1, 4'd0, 27'h000001a1, 4'd14, 27'h00000062, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002a8, 4'd8, 27'h00000382, 4'd4, 27'h000002b5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000399, 4'd8, 27'h0000027b, 4'd5, 27'h00000153, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000044, 4'd5, 27'h00000216, 4'd13, 27'h000001d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000331, 4'd14, 27'h000002ca, 4'd1, 27'h000001a4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001b3, 4'd14, 27'h0000008d, 4'd6, 27'h000003a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001fd, 4'd13, 27'h00000075, 4'd13, 27'h00000182, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000166, 4'd2, 27'h00000356, 4'd2, 27'h0000003b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000d4, 4'd4, 27'h0000028d, 4'd8, 27'h00000210, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000cc, 4'd0, 27'h00000001, 4'd13, 27'h00000031, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000017, 4'd7, 27'h000003d8, 4'd0, 27'h00000177, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000002e, 4'd6, 27'h0000035d, 4'd9, 27'h000003f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000188, 4'd6, 27'h000003d5, 4'd10, 27'h0000033f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000290, 4'd14, 27'h00000390, 4'd1, 27'h00000069, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000aa, 4'd10, 27'h000001c3, 4'd5, 27'h00000219, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000004f, 4'd12, 27'h00000383, 4'd10, 27'h000000d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002bb, 4'd4, 27'h00000180, 4'd4, 27'h00000189, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000281, 4'd3, 27'h00000067, 4'd9, 27'h00000186, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000016e, 4'd4, 27'h00000373, 4'd13, 27'h000002be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000307, 4'd9, 27'h00000315, 4'd0, 27'h00000030, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000023d, 4'd5, 27'h00000005, 4'd8, 27'h0000002e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000229, 4'd8, 27'h00000072, 4'd11, 27'h000001f1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002ee, 4'd13, 27'h00000118, 4'd3, 27'h00000128, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000013, 4'd13, 27'h00000263, 4'd8, 27'h00000156, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000344, 4'd12, 27'h00000231, 4'd11, 27'h000002ce, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000073, 4'd2, 27'h00000130, 4'd0, 27'h0000002d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000030d, 4'd3, 27'h00000235, 4'd5, 27'h00000049, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001b4, 4'd3, 27'h000001ba, 4'd12, 27'h000002ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000149, 4'd5, 27'h00000079, 4'd0, 27'h0000017b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b1, 4'd5, 27'h00000316, 4'd5, 27'h000000af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000009f, 4'd9, 27'h00000366, 4'd11, 27'h0000037b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000300, 4'd14, 27'h000000a5, 4'd4, 27'h00000044, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001cd, 4'd11, 27'h00000299, 4'd9, 27'h00000298, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000241, 4'd13, 27'h0000039c, 4'd12, 27'h00000159, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000205, 4'd3, 27'h000000f5, 4'd4, 27'h00000019, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000254, 4'd3, 27'h00000154, 4'd8, 27'h00000083, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000b9, 4'd1, 27'h00000201, 4'd14, 27'h00000100, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000009c, 4'd5, 27'h00000267, 4'd2, 27'h00000135, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000201, 4'd6, 27'h00000347, 4'd7, 27'h0000034f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002f9, 4'd7, 27'h000000a1, 4'd13, 27'h000002e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000037f, 4'd11, 27'h000003d1, 4'd3, 27'h00000174, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000003a, 4'd11, 27'h00000189, 4'd5, 27'h000002b4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001b5, 4'd14, 27'h00000233, 4'd11, 27'h000000de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000019b, 4'd2, 27'h0000030f, 4'd0, 27'h00000123, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000b7, 4'd1, 27'h0000034c, 4'd8, 27'h0000031c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003ca, 4'd1, 27'h00000111, 4'd14, 27'h0000036f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001a7, 4'd7, 27'h00000061, 4'd4, 27'h0000000a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000c7, 4'd5, 27'h00000282, 4'd5, 27'h00000026, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000349, 4'd6, 27'h00000018, 4'd12, 27'h00000062, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000071, 4'd14, 27'h000000e6, 4'd4, 27'h0000034e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000de, 4'd11, 27'h00000273, 4'd7, 27'h00000179, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000e3, 4'd13, 27'h0000023f, 4'd13, 27'h000002c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003b9, 4'd3, 27'h00000383, 4'd2, 27'h000000f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ce, 4'd1, 27'h000000af, 4'd7, 27'h00000152, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000268, 4'd3, 27'h000000a7, 4'd12, 27'h000003d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003c3, 4'd7, 27'h000003bb, 4'd2, 27'h000001a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000012c, 4'd9, 27'h00000076, 4'd9, 27'h000003f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003c1, 4'd7, 27'h000001e7, 4'd13, 27'h0000024e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000039e, 4'd10, 27'h00000193, 4'd2, 27'h00000088, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002c8, 4'd12, 27'h00000388, 4'd7, 27'h000003db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000032c, 4'd11, 27'h0000018f, 4'd10, 27'h00000093, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000281, 4'd1, 27'h00000381, 4'd0, 27'h0000004c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001e7, 4'd0, 27'h000002de, 4'd9, 27'h00000230, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000199, 4'd0, 27'h000002b0, 4'd12, 27'h00000000, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000084, 4'd6, 27'h00000244, 4'd2, 27'h0000004d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002c2, 4'd9, 27'h000002ee, 4'd5, 27'h00000174, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000312, 4'd6, 27'h00000049, 4'd11, 27'h00000229, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000147, 4'd14, 27'h000001f9, 4'd0, 27'h00000264, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000241, 4'd10, 27'h000002b1, 4'd6, 27'h000000e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000126, 4'd10, 27'h00000381, 4'd10, 27'h00000095, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000020a, 4'd0, 27'h00000083, 4'd3, 27'h00000110, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000022f, 4'd2, 27'h00000340, 4'd6, 27'h000001c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000378, 4'd4, 27'h00000262, 4'd12, 27'h0000027b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000106, 4'd8, 27'h000003e4, 4'd3, 27'h0000000c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000118, 4'd6, 27'h0000023e, 4'd5, 27'h000003b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000093, 4'd8, 27'h00000048, 4'd12, 27'h00000294, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000025, 4'd14, 27'h000000ef, 4'd3, 27'h00000243, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000007f, 4'd10, 27'h000001f2, 4'd9, 27'h00000150, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000d5, 4'd13, 27'h000002af, 4'd12, 27'h00000156, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ee, 4'd1, 27'h00000019, 4'd2, 27'h000000a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000066, 4'd4, 27'h00000249, 4'd9, 27'h00000064, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000164, 4'd3, 27'h0000031a, 4'd13, 27'h00000097, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002b5, 4'd5, 27'h00000123, 4'd2, 27'h00000124, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000f5, 4'd9, 27'h0000006f, 4'd7, 27'h000001d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000008d, 4'd7, 27'h000001ba, 4'd13, 27'h00000394, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002be, 4'd11, 27'h0000005d, 4'd1, 27'h0000039b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000091, 4'd14, 27'h000002c4, 4'd5, 27'h000003ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000036, 4'd14, 27'h00000170, 4'd14, 27'h0000036b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002da, 4'd1, 27'h00000097, 4'd4, 27'h00000299, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000004b, 4'd3, 27'h000001cf, 4'd9, 27'h000003f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000229, 4'd1, 27'h00000302, 4'd11, 27'h0000009b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001b7, 4'd6, 27'h00000223, 4'd3, 27'h000002a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002b7, 4'd5, 27'h00000340, 4'd7, 27'h000002d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000254, 4'd5, 27'h000000dd, 4'd11, 27'h00000343, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002e6, 4'd10, 27'h00000035, 4'd3, 27'h000001b8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000006, 4'd11, 27'h000001b1, 4'd7, 27'h000001b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000226, 4'd10, 27'h00000195, 4'd14, 27'h00000307, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000000a, 4'd1, 27'h000002f5, 4'd3, 27'h0000018a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000245, 4'd3, 27'h0000010f, 4'd5, 27'h000000d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000159, 4'd2, 27'h00000221, 4'd11, 27'h000002c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000200, 4'd5, 27'h000000c7, 4'd3, 27'h000002e4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002de, 4'd6, 27'h000003bb, 4'd6, 27'h0000014a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000339, 4'd6, 27'h000003b8, 4'd13, 27'h000000eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002df, 4'd12, 27'h00000134, 4'd2, 27'h00000275, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000017f, 4'd14, 27'h000002f8, 4'd9, 27'h000001d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000001c, 4'd11, 27'h00000372, 4'd13, 27'h0000028f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000039c, 4'd3, 27'h0000023b, 4'd4, 27'h000001cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000026b, 4'd1, 27'h0000005d, 4'd5, 27'h000002d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000167, 4'd0, 27'h00000367, 4'd13, 27'h00000264, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000231, 4'd7, 27'h000002ca, 4'd0, 27'h00000001, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000298, 4'd5, 27'h00000260, 4'd6, 27'h0000000a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000345, 4'd7, 27'h000002d0, 4'd14, 27'h000003ea, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000b9, 4'd12, 27'h0000024e, 4'd2, 27'h000000fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000244, 4'd12, 27'h00000001, 4'd5, 27'h000000a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000140, 4'd12, 27'h00000271, 4'd10, 27'h00000065, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000207, 4'd4, 27'h0000028d, 4'd0, 27'h00000267, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000034c, 4'd3, 27'h0000008f, 4'd7, 27'h000001d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000019f, 4'd4, 27'h00000036, 4'd14, 27'h0000011c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003a0, 4'd5, 27'h000002b3, 4'd3, 27'h00000358, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003a0, 4'd6, 27'h000001c4, 4'd5, 27'h00000040, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000199, 4'd5, 27'h00000062, 4'd14, 27'h00000165, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000097, 4'd12, 27'h000001a1, 4'd4, 27'h000002e2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002c3, 4'd13, 27'h00000191, 4'd7, 27'h0000023a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003fd, 4'd14, 27'h00000069, 4'd14, 27'h0000024c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000c6, 4'd0, 27'h000002a5, 4'd0, 27'h0000037e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000171, 4'd1, 27'h00000081, 4'd7, 27'h000000e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000387, 4'd1, 27'h0000012c, 4'd12, 27'h000000cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000039b, 4'd9, 27'h00000343, 4'd3, 27'h00000327, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000192, 4'd5, 27'h00000339, 4'd5, 27'h0000008a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000f4, 4'd9, 27'h000000d9, 4'd13, 27'h00000249, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000023d, 4'd14, 27'h000002e4, 4'd3, 27'h0000017a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000240, 4'd13, 27'h000001f9, 4'd5, 27'h00000075, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000305, 4'd14, 27'h00000257, 4'd13, 27'h0000003d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000209, 4'd4, 27'h00000021, 4'd2, 27'h00000150, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000121, 4'd3, 27'h0000004c, 4'd9, 27'h00000015, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000006a, 4'd0, 27'h00000047, 4'd10, 27'h000001ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000193, 4'd7, 27'h00000195, 4'd2, 27'h00000355, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003cd, 4'd9, 27'h0000026d, 4'd8, 27'h00000128, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000010f, 4'd5, 27'h000002ae, 4'd13, 27'h000003e3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000070, 4'd11, 27'h000002b2, 4'd3, 27'h00000003, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000031d, 4'd14, 27'h000002ed, 4'd8, 27'h0000029b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001e1, 4'd12, 27'h000000a6, 4'd11, 27'h000002b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003c6, 4'd2, 27'h000003d6, 4'd4, 27'h00000380, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000160, 4'd0, 27'h00000368, 4'd5, 27'h00000343, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000020b, 4'd4, 27'h0000007b, 4'd11, 27'h000002da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000386, 4'd8, 27'h00000133, 4'd4, 27'h000002d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000295, 4'd7, 27'h0000025e, 4'd8, 27'h000003b8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000032a, 4'd8, 27'h000002f8, 4'd12, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000204, 4'd10, 27'h000001b8, 4'd3, 27'h00000170, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000342, 4'd10, 27'h000002a7, 4'd7, 27'h00000190, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000014e, 4'd12, 27'h000000ce, 4'd12, 27'h000001b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003aa, 4'd3, 27'h00000244, 4'd1, 27'h000003fc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000d6, 4'd3, 27'h0000022b, 4'd5, 27'h000003a0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000310, 4'd3, 27'h00000115, 4'd13, 27'h000000d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003e4, 4'd9, 27'h0000002d, 4'd2, 27'h00000397, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000cb, 4'd8, 27'h000001a8, 4'd9, 27'h000000f4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000e0, 4'd9, 27'h00000107, 4'd10, 27'h00000004, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001e1, 4'd11, 27'h000000bd, 4'd2, 27'h00000240, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000039a, 4'd12, 27'h00000392, 4'd5, 27'h0000012e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003ce, 4'd10, 27'h000000dc, 4'd12, 27'h0000012c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002b9, 4'd2, 27'h00000316, 4'd2, 27'h000000e4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000a1, 4'd1, 27'h0000029b, 4'd8, 27'h000003bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000106, 4'd0, 27'h000000e4, 4'd12, 27'h000002ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003cb, 4'd8, 27'h00000330, 4'd4, 27'h00000078, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001d8, 4'd9, 27'h0000005d, 4'd6, 27'h0000038f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002b5, 4'd6, 27'h00000336, 4'd13, 27'h00000195, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000064, 4'd12, 27'h00000205, 4'd0, 27'h0000013a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002fc, 4'd14, 27'h000000e6, 4'd9, 27'h00000194, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000004f, 4'd10, 27'h00000221, 4'd11, 27'h0000012d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000338, 4'd2, 27'h000003bf, 4'd2, 27'h00000028, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001b4, 4'd0, 27'h00000092, 4'd8, 27'h000000e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000164, 4'd2, 27'h0000015c, 4'd11, 27'h0000009b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003d9, 4'd8, 27'h00000146, 4'd1, 27'h00000180, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001af, 4'd7, 27'h000002a1, 4'd5, 27'h0000013f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000067, 4'd7, 27'h000002ea, 4'd13, 27'h000003b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002f7, 4'd14, 27'h00000089, 4'd2, 27'h00000213, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000353, 4'd14, 27'h00000189, 4'd8, 27'h00000119, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003f6, 4'd14, 27'h000000a2, 4'd11, 27'h00000083, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000236, 4'd0, 27'h0000018d, 4'd3, 27'h0000006e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000011b, 4'd4, 27'h00000286, 4'd9, 27'h00000100, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000028, 4'd0, 27'h0000008a, 4'd12, 27'h0000034b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000218, 4'd9, 27'h000000f1, 4'd4, 27'h0000006d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000125, 4'd8, 27'h00000339, 4'd9, 27'h000003a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002a3, 4'd6, 27'h0000000c, 4'd10, 27'h000003a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001c3, 4'd10, 27'h000001a1, 4'd1, 27'h000001df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000015, 4'd13, 27'h00000052, 4'd5, 27'h00000086, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000240, 4'd13, 27'h000000da, 4'd11, 27'h0000019b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000373, 4'd2, 27'h00000217, 4'd0, 27'h000001ed, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000036b, 4'd0, 27'h000003ec, 4'd7, 27'h00000150, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000039f, 4'd4, 27'h00000052, 4'd14, 27'h00000167, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001b9, 4'd9, 27'h0000027d, 4'd4, 27'h000002dd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003b7, 4'd7, 27'h0000008d, 4'd8, 27'h000002eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000316, 4'd8, 27'h000001ed, 4'd10, 27'h0000021d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003b9, 4'd11, 27'h00000214, 4'd1, 27'h00000223, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000290, 4'd12, 27'h0000035b, 4'd8, 27'h000000ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000141, 4'd14, 27'h0000035d, 4'd11, 27'h000002c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000ac, 4'd1, 27'h00000341, 4'd1, 27'h00000030, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000011a, 4'd3, 27'h000001c6, 4'd6, 27'h000000dd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000008, 4'd1, 27'h00000088, 4'd14, 27'h000001ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000341, 4'd8, 27'h00000306, 4'd0, 27'h0000012b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000028b, 4'd6, 27'h0000020b, 4'd7, 27'h0000022b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003b0, 4'd7, 27'h00000111, 4'd14, 27'h0000001a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001db, 4'd12, 27'h000001d7, 4'd0, 27'h0000019a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000238, 4'd13, 27'h000003a7, 4'd7, 27'h000001d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000291, 4'd11, 27'h0000037d, 4'd11, 27'h00000280, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000013e, 4'd2, 27'h00000061, 4'd3, 27'h0000023e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000038c, 4'd0, 27'h0000008e, 4'd5, 27'h0000009d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000037b, 4'd1, 27'h00000263, 4'd14, 27'h000000f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000283, 4'd6, 27'h000001b0, 4'd2, 27'h000001c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000036e, 4'd7, 27'h0000005b, 4'd8, 27'h00000006, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000230, 4'd8, 27'h00000371, 4'd13, 27'h0000009c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000038a, 4'd14, 27'h00000211, 4'd4, 27'h00000233, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000211, 4'd10, 27'h00000165, 4'd9, 27'h00000104, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000137, 4'd14, 27'h00000299, 4'd10, 27'h00000036, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000277, 4'd1, 27'h000002ec, 4'd1, 27'h000003ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000029b, 4'd0, 27'h000003d9, 4'd5, 27'h00000247, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000030e, 4'd0, 27'h00000397, 4'd10, 27'h0000002e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000197, 4'd8, 27'h00000190, 4'd2, 27'h000002f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000252, 4'd9, 27'h00000398, 4'd7, 27'h0000017b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000306, 4'd9, 27'h00000099, 4'd14, 27'h00000201, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000004e, 4'd10, 27'h000002b0, 4'd0, 27'h000001c4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000019d, 4'd11, 27'h0000016e, 4'd5, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000007c, 4'd10, 27'h0000007d, 4'd12, 27'h0000036b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000245, 4'd1, 27'h00000050, 4'd1, 27'h00000214, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000f4, 4'd3, 27'h000003bd, 4'd8, 27'h000000b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003fa, 4'd2, 27'h000000e1, 4'd12, 27'h0000019f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003d1, 4'd7, 27'h000003cf, 4'd2, 27'h00000085, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000084, 4'd6, 27'h000001d7, 4'd6, 27'h000001eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000002e, 4'd8, 27'h000000ef, 4'd10, 27'h000002a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000393, 4'd13, 27'h00000340, 4'd3, 27'h000002ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002e3, 4'd11, 27'h00000304, 4'd8, 27'h000002ba, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001f2, 4'd14, 27'h000001a3, 4'd12, 27'h00000019, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000206, 4'd4, 27'h00000222, 4'd1, 27'h000000b8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000003b, 4'd1, 27'h00000276, 4'd8, 27'h000000b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000350, 4'd3, 27'h000000d8, 4'd10, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000394, 4'd7, 27'h0000020c, 4'd2, 27'h0000031a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000011a, 4'd9, 27'h0000038f, 4'd6, 27'h000001d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000114, 4'd9, 27'h0000008d, 4'd11, 27'h00000287, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003c8, 4'd14, 27'h0000014f, 4'd3, 27'h000001a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000006a, 4'd13, 27'h0000004d, 4'd8, 27'h000002e2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002fb, 4'd13, 27'h00000148, 4'd14, 27'h0000020c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000112, 4'd3, 27'h0000027f, 4'd1, 27'h0000006e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000ce, 4'd0, 27'h00000203, 4'd5, 27'h0000032f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002a0, 4'd3, 27'h00000027, 4'd10, 27'h0000030c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002f1, 4'd8, 27'h0000034c, 4'd1, 27'h00000215, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000288, 4'd8, 27'h00000218, 4'd7, 27'h00000247, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000349, 4'd8, 27'h000003d3, 4'd12, 27'h00000397, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003cf, 4'd11, 27'h0000016e, 4'd0, 27'h00000351, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002db, 4'd12, 27'h0000007f, 4'd7, 27'h00000357, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000324, 4'd10, 27'h00000075, 4'd14, 27'h00000091, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003fb, 4'd4, 27'h00000368, 4'd0, 27'h00000325, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000383, 4'd1, 27'h000001a1, 4'd7, 27'h00000018, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003e8, 4'd2, 27'h000002ea, 4'd14, 27'h00000184, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000024a, 4'd9, 27'h00000289, 4'd0, 27'h000001cf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000023, 4'd9, 27'h00000269, 4'd7, 27'h00000302, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000e5, 4'd7, 27'h0000018c, 4'd14, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000da, 4'd10, 27'h000000e7, 4'd0, 27'h0000010f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000385, 4'd14, 27'h000002f9, 4'd5, 27'h000000ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000013a, 4'd13, 27'h000003c5, 4'd10, 27'h0000025d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003d7, 4'd2, 27'h000003b6, 4'd0, 27'h0000024c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000038c, 4'd1, 27'h00000198, 4'd5, 27'h000002c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000015a, 4'd2, 27'h00000199, 4'd13, 27'h000000d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000076, 4'd8, 27'h000001f3, 4'd1, 27'h00000294, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000016f, 4'd9, 27'h0000001c, 4'd5, 27'h0000039e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000ff, 4'd6, 27'h000000aa, 4'd14, 27'h0000013e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003cd, 4'd11, 27'h00000002, 4'd1, 27'h000001bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000332, 4'd14, 27'h00000038, 4'd9, 27'h0000019d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000280, 4'd14, 27'h0000016b, 4'd14, 27'h00000077, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000072, 4'd1, 27'h00000180, 4'd0, 27'h0000009c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002cc, 4'd2, 27'h00000102, 4'd7, 27'h00000336, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003aa, 4'd3, 27'h0000002c, 4'd12, 27'h000001b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000248, 4'd8, 27'h0000038a, 4'd4, 27'h00000182, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000362, 4'd5, 27'h00000077, 4'd5, 27'h0000022b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000063, 4'd9, 27'h000002e1, 4'd14, 27'h00000393, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002e9, 4'd10, 27'h00000094, 4'd3, 27'h000002eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000378, 4'd10, 27'h00000161, 4'd8, 27'h000003ef, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000202, 4'd11, 27'h0000031f, 4'd12, 27'h000003c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000363, 4'd1, 27'h00000306, 4'd3, 27'h000001cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000022c, 4'd4, 27'h000001b1, 4'd8, 27'h00000027, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003a4, 4'd0, 27'h0000036c, 4'd13, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000037b, 4'd9, 27'h0000022f, 4'd4, 27'h000003d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000dc, 4'd7, 27'h00000217, 4'd5, 27'h000001a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000040, 4'd6, 27'h00000131, 4'd11, 27'h000000e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000086, 4'd13, 27'h000000e6, 4'd3, 27'h00000113, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001d7, 4'd13, 27'h00000077, 4'd9, 27'h000002b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003e1, 4'd13, 27'h00000103, 4'd10, 27'h0000037e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000085, 4'd4, 27'h00000055, 4'd3, 27'h00000224, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000299, 4'd0, 27'h000000e4, 4'd9, 27'h000001bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003f1, 4'd4, 27'h0000002d, 4'd14, 27'h000001cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000ca, 4'd5, 27'h00000299, 4'd4, 27'h00000149, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003f1, 4'd5, 27'h00000035, 4'd7, 27'h00000369, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000033c, 4'd6, 27'h00000159, 4'd14, 27'h00000243, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000084, 4'd14, 27'h0000018f, 4'd0, 27'h00000100, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000032b, 4'd13, 27'h00000209, 4'd9, 27'h000000d7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000123, 4'd10, 27'h000003b1, 4'd10, 27'h00000018, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000071, 4'd1, 27'h00000350, 4'd4, 27'h00000005, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002c2, 4'd0, 27'h00000248, 4'd8, 27'h000000ba, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000254, 4'd0, 27'h00000004, 4'd14, 27'h00000061, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001c7, 4'd6, 27'h0000033d, 4'd0, 27'h00000222, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000095, 4'd6, 27'h000000b5, 4'd9, 27'h0000034b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000012d, 4'd5, 27'h00000021, 4'd11, 27'h000002c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002d5, 4'd10, 27'h000002d3, 4'd1, 27'h0000033e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000363, 4'd12, 27'h000002bb, 4'd6, 27'h00000292, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000cf, 4'd14, 27'h000003a5, 4'd14, 27'h00000253, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000c2, 4'd4, 27'h000002a7, 4'd1, 27'h000001aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000012a, 4'd2, 27'h0000003d, 4'd5, 27'h000003e5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000364, 4'd1, 27'h000002aa, 4'd13, 27'h00000273, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003d6, 4'd9, 27'h0000007c, 4'd2, 27'h0000007e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002c9, 4'd9, 27'h00000063, 4'd5, 27'h0000026a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000306, 4'd6, 27'h000002b0, 4'd11, 27'h00000062, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000389, 4'd11, 27'h00000192, 4'd0, 27'h00000331, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000269, 4'd13, 27'h00000153, 4'd8, 27'h00000165, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000033d, 4'd12, 27'h00000225, 4'd11, 27'h000000a3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000275, 4'd1, 27'h00000189, 4'd3, 27'h000001c0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002de, 4'd0, 27'h00000215, 4'd7, 27'h00000121, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000de, 4'd1, 27'h00000210, 4'd11, 27'h000002f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000138, 4'd5, 27'h0000003d, 4'd4, 27'h0000000c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000383, 4'd9, 27'h000002cb, 4'd9, 27'h000001c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000023c, 4'd6, 27'h000003a5, 4'd10, 27'h000001fc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001cf, 4'd13, 27'h00000009, 4'd4, 27'h0000010c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000016e, 4'd13, 27'h00000161, 4'd7, 27'h00000099, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000017b, 4'd11, 27'h0000039c, 4'd11, 27'h00000143, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000030, 4'd3, 27'h0000009a, 4'd0, 27'h000000ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000071, 4'd1, 27'h000002aa, 4'd9, 27'h00000213, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000150, 4'd1, 27'h000002f9, 4'd12, 27'h00000100, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000145, 4'd6, 27'h00000106, 4'd2, 27'h00000154, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002d0, 4'd5, 27'h0000031c, 4'd8, 27'h0000017f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000143, 4'd6, 27'h0000013a, 4'd13, 27'h00000092, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001ca, 4'd10, 27'h00000174, 4'd3, 27'h0000036d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000030c, 4'd13, 27'h000003b9, 4'd7, 27'h00000290, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000036a, 4'd10, 27'h00000279, 4'd10, 27'h0000015e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000135, 4'd4, 27'h000000e0, 4'd4, 27'h00000302, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000012b, 4'd0, 27'h00000353, 4'd5, 27'h000000df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002fe, 4'd4, 27'h00000298, 4'd11, 27'h000000d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000011d, 4'd7, 27'h0000034f, 4'd4, 27'h0000037e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000032e, 4'd8, 27'h000003be, 4'd6, 27'h00000010, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000080, 4'd8, 27'h0000004e, 4'd11, 27'h0000034c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002a7, 4'd12, 27'h0000033a, 4'd1, 27'h00000282, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002d4, 4'd12, 27'h000003fd, 4'd7, 27'h000002d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000287, 4'd11, 27'h00000288, 4'd13, 27'h000001b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000006c, 4'd1, 27'h00000118, 4'd2, 27'h0000031d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000011e, 4'd0, 27'h00000185, 4'd5, 27'h00000182, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000033b, 4'd4, 27'h000002e1, 4'd11, 27'h000000ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000010, 4'd5, 27'h00000183, 4'd3, 27'h000001cf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000357, 4'd8, 27'h000003c3, 4'd6, 27'h0000014f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001cc, 4'd5, 27'h000003ab, 4'd12, 27'h000001e9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002b0, 4'd14, 27'h000000c3, 4'd0, 27'h000003e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000089, 4'd12, 27'h00000399, 4'd6, 27'h0000023e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000078, 4'd11, 27'h00000367, 4'd13, 27'h0000014d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000219, 4'd0, 27'h0000035b, 4'd1, 27'h000000b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000b8, 4'd3, 27'h00000136, 4'd5, 27'h00000014, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000370, 4'd1, 27'h00000310, 4'd12, 27'h0000031e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001a4, 4'd7, 27'h000003cf, 4'd2, 27'h000003fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000061, 4'd7, 27'h000003e5, 4'd7, 27'h00000231, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000007b, 4'd9, 27'h000002ea, 4'd10, 27'h000003c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000376, 4'd11, 27'h00000070, 4'd1, 27'h000003b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000dd, 4'd14, 27'h000001e9, 4'd6, 27'h00000026, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002d9, 4'd13, 27'h00000397, 4'd12, 27'h00000129, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000329, 4'd3, 27'h00000007, 4'd2, 27'h000002d1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003be, 4'd4, 27'h0000032d, 4'd5, 27'h00000235, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000019b, 4'd3, 27'h000000e2, 4'd13, 27'h000002ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003b8, 4'd7, 27'h0000000f, 4'd1, 27'h000000de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000005a, 4'd9, 27'h000003b4, 4'd8, 27'h00000189, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001cd, 4'd6, 27'h00000063, 4'd12, 27'h00000019, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000097, 4'd11, 27'h0000017a, 4'd2, 27'h0000012a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000342, 4'd10, 27'h000000a6, 4'd9, 27'h0000005e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001df, 4'd12, 27'h0000015d, 4'd10, 27'h00000345, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000081, 4'd0, 27'h0000005d, 4'd1, 27'h0000025d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002fb, 4'd4, 27'h00000142, 4'd7, 27'h000001c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000181, 4'd1, 27'h000000e3, 4'd10, 27'h00000011, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000008d, 4'd5, 27'h00000203, 4'd1, 27'h0000021b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000139, 4'd6, 27'h00000303, 4'd8, 27'h0000025f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000253, 4'd6, 27'h0000021f, 4'd12, 27'h000003ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000032c, 4'd12, 27'h000000a7, 4'd2, 27'h00000064, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000011e, 4'd11, 27'h0000026f, 4'd5, 27'h000000d9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000389, 4'd11, 27'h000001fb, 4'd12, 27'h0000023b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003b2, 4'd0, 27'h0000039a, 4'd1, 27'h0000003b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000012a, 4'd1, 27'h000002a0, 4'd6, 27'h0000010f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000ad, 4'd2, 27'h000003cb, 4'd12, 27'h0000001b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000022e, 4'd9, 27'h00000326, 4'd0, 27'h00000042, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000c7, 4'd5, 27'h000003ce, 4'd6, 27'h00000130, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000292, 4'd8, 27'h00000383, 4'd11, 27'h00000284, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000193, 4'd13, 27'h0000026d, 4'd4, 27'h000001b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000005, 4'd13, 27'h00000100, 4'd5, 27'h00000033, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000a7, 4'd10, 27'h00000378, 4'd10, 27'h000002d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001ca, 4'd0, 27'h000000e0, 4'd3, 27'h00000005, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000007, 4'd2, 27'h000002e7, 4'd7, 27'h000001ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000c6, 4'd0, 27'h00000212, 4'd14, 27'h00000051, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000155, 4'd7, 27'h000000c7, 4'd2, 27'h00000120, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001b2, 4'd5, 27'h000003af, 4'd6, 27'h0000032f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000025c, 4'd8, 27'h00000015, 4'd14, 27'h0000031a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000111, 4'd14, 27'h00000377, 4'd3, 27'h00000133, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000fc, 4'd10, 27'h0000013e, 4'd7, 27'h0000001b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000e1, 4'd11, 27'h0000016c, 4'd11, 27'h00000047, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000035a, 4'd0, 27'h000002d5, 4'd0, 27'h00000339, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001db, 4'd1, 27'h000000bb, 4'd5, 27'h0000026a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000089, 4'd0, 27'h000000e5, 4'd11, 27'h00000101, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001e4, 4'd6, 27'h00000193, 4'd2, 27'h000002e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000321, 4'd7, 27'h0000026d, 4'd6, 27'h00000244, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000d2, 4'd5, 27'h00000327, 4'd12, 27'h00000225, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003ad, 4'd10, 27'h00000092, 4'd3, 27'h000002bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000398, 4'd13, 27'h000003a3, 4'd8, 27'h00000186, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000029d, 4'd13, 27'h000003eb, 4'd11, 27'h00000263, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000318, 4'd3, 27'h0000012d, 4'd4, 27'h00000399, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001d6, 4'd4, 27'h000000f0, 4'd6, 27'h00000087, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002e1, 4'd2, 27'h000003a0, 4'd13, 27'h0000028e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000164, 4'd6, 27'h000003a0, 4'd3, 27'h000003f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000029e, 4'd5, 27'h000003fb, 4'd5, 27'h00000322, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003f4, 4'd9, 27'h00000025, 4'd11, 27'h0000031f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000c3, 4'd11, 27'h0000036f, 4'd4, 27'h0000038c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000348, 4'd10, 27'h00000074, 4'd8, 27'h00000359, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001f2, 4'd13, 27'h000003d0, 4'd14, 27'h0000018d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000012, 4'd2, 27'h00000347, 4'd1, 27'h000001ad, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000108, 4'd3, 27'h0000019b, 4'd8, 27'h0000037d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000109, 4'd0, 27'h000000f2, 4'd10, 27'h00000217, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e7, 4'd8, 27'h000000b4, 4'd4, 27'h000001a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000017e, 4'd6, 27'h0000028f, 4'd8, 27'h000000c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000013c, 4'd7, 27'h000000e1, 4'd10, 27'h00000239, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000e2, 4'd10, 27'h000001c6, 4'd4, 27'h00000092, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003de, 4'd14, 27'h000000e4, 4'd7, 27'h000001ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000013a, 4'd11, 27'h0000008b, 4'd14, 27'h00000118, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000248, 4'd4, 27'h000002e6, 4'd2, 27'h000000d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000083, 4'd3, 27'h0000034d, 4'd8, 27'h00000151, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000164, 4'd2, 27'h0000032a, 4'd10, 27'h00000047, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000082, 4'd9, 27'h00000151, 4'd3, 27'h000001ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000013a, 4'd7, 27'h00000165, 4'd9, 27'h00000145, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000261, 4'd7, 27'h0000002f, 4'd13, 27'h000003f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000129, 4'd14, 27'h0000025a, 4'd2, 27'h00000214, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c0, 4'd14, 27'h000003fb, 4'd9, 27'h00000002, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000e5, 4'd10, 27'h000002b5, 4'd12, 27'h0000022a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003cd, 4'd0, 27'h0000023e, 4'd3, 27'h00000069, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000122, 4'd1, 27'h000003c9, 4'd8, 27'h0000009a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000c5, 4'd3, 27'h0000010a, 4'd13, 27'h00000227, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000144, 4'd5, 27'h000003e8, 4'd0, 27'h0000007e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000022, 4'd9, 27'h00000071, 4'd9, 27'h00000019, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001db, 4'd6, 27'h000003a7, 4'd10, 27'h0000023f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000009a, 4'd10, 27'h000003a4, 4'd3, 27'h000002fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001c7, 4'd14, 27'h000003a0, 4'd8, 27'h0000025b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000025a, 4'd14, 27'h00000268, 4'd14, 27'h0000001a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000a0, 4'd2, 27'h000000b0, 4'd3, 27'h000001da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000379, 4'd3, 27'h0000006b, 4'd5, 27'h00000382, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000054, 4'd1, 27'h00000199, 4'd13, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000008e, 4'd6, 27'h000003dd, 4'd1, 27'h000003ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000111, 4'd6, 27'h00000385, 4'd5, 27'h00000104, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000040, 4'd7, 27'h000003ae, 4'd13, 27'h00000338, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001fe, 4'd13, 27'h0000018c, 4'd0, 27'h0000006c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003ca, 4'd11, 27'h000001e5, 4'd6, 27'h000001dc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003e1, 4'd12, 27'h000003cc, 4'd11, 27'h000003e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000241, 4'd3, 27'h000003fb, 4'd1, 27'h0000003b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000314, 4'd0, 27'h0000000b, 4'd8, 27'h0000019c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000376, 4'd4, 27'h00000156, 4'd11, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000006a, 4'd6, 27'h00000169, 4'd3, 27'h000001ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000123, 4'd6, 27'h00000162, 4'd6, 27'h000001b3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000017d, 4'd8, 27'h000001ab, 4'd12, 27'h0000001c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003db, 4'd13, 27'h000003b5, 4'd3, 27'h000003eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000042, 4'd12, 27'h00000364, 4'd9, 27'h0000035b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001bc, 4'd11, 27'h00000310, 4'd11, 27'h0000021b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000f0, 4'd0, 27'h00000076, 4'd4, 27'h000002a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003d3, 4'd4, 27'h00000210, 4'd7, 27'h00000188, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001f4, 4'd2, 27'h00000058, 4'd10, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000b3, 4'd8, 27'h0000024e, 4'd4, 27'h000002c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000dd, 4'd6, 27'h00000184, 4'd5, 27'h000003c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003be, 4'd6, 27'h00000017, 4'd10, 27'h000002f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001a1, 4'd12, 27'h0000016a, 4'd1, 27'h0000022f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003d6, 4'd14, 27'h00000048, 4'd8, 27'h00000218, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001c3, 4'd11, 27'h0000020a, 4'd13, 27'h00000248, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000018f, 4'd0, 27'h0000027f, 4'd1, 27'h00000198, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000024c, 4'd2, 27'h00000109, 4'd9, 27'h000000f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000008, 4'd3, 27'h0000033a, 4'd12, 27'h0000005f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003f6, 4'd6, 27'h0000016f, 4'd4, 27'h00000010, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000192, 4'd8, 27'h00000297, 4'd6, 27'h000000ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000d0, 4'd7, 27'h0000006c, 4'd14, 27'h0000034c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000004a, 4'd12, 27'h00000022, 4'd0, 27'h00000279, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000022c, 4'd11, 27'h0000038b, 4'd9, 27'h00000060, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000018a, 4'd10, 27'h000002c5, 4'd14, 27'h000002d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000022f, 4'd3, 27'h000000d2, 4'd1, 27'h000002ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000029b, 4'd0, 27'h0000009f, 4'd6, 27'h000000a2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000398, 4'd3, 27'h000003e8, 4'd10, 27'h000001a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000038d, 4'd8, 27'h00000242, 4'd1, 27'h000001f1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000022c, 4'd6, 27'h00000206, 4'd9, 27'h000002c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000176, 4'd6, 27'h00000395, 4'd10, 27'h000001e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000048, 4'd13, 27'h000003a5, 4'd1, 27'h000000be, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000039a, 4'd10, 27'h0000021a, 4'd6, 27'h0000027f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003e3, 4'd14, 27'h00000078, 4'd11, 27'h00000235, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000280, 4'd1, 27'h000001b7, 4'd4, 27'h000003a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000af, 4'd4, 27'h000000bf, 4'd9, 27'h00000144, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000e2, 4'd0, 27'h000002e8, 4'd12, 27'h000000a7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b8, 4'd9, 27'h00000073, 4'd4, 27'h0000021a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000009d, 4'd9, 27'h000001b0, 4'd6, 27'h000000c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000328, 4'd6, 27'h000002ee, 4'd12, 27'h000003b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000304, 4'd14, 27'h000003a5, 4'd2, 27'h00000150, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002d6, 4'd11, 27'h0000034c, 4'd5, 27'h0000025e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001dc, 4'd11, 27'h00000200, 4'd12, 27'h000003e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000026b, 4'd3, 27'h00000212, 4'd0, 27'h000000ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000251, 4'd0, 27'h000001a3, 4'd5, 27'h000000af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000bf, 4'd0, 27'h000000d5, 4'd11, 27'h00000053, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002dd, 4'd9, 27'h00000354, 4'd0, 27'h000002bc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001be, 4'd9, 27'h000003ae, 4'd5, 27'h00000229, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000eb, 4'd6, 27'h00000305, 4'd13, 27'h0000028c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000225, 4'd10, 27'h000000a0, 4'd2, 27'h0000023a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001bb, 4'd14, 27'h00000056, 4'd8, 27'h0000035b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a3, 4'd12, 27'h0000023a, 4'd10, 27'h00000238, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000192, 4'd3, 27'h000000e4, 4'd1, 27'h000003bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002bb, 4'd3, 27'h00000122, 4'd8, 27'h000000fb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000e9, 4'd3, 27'h000002cc, 4'd10, 27'h000003e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000271, 4'd9, 27'h00000146, 4'd3, 27'h0000004c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002ee, 4'd5, 27'h000000af, 4'd6, 27'h00000234, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000002f, 4'd6, 27'h0000039c, 4'd13, 27'h0000007e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000114, 4'd13, 27'h00000332, 4'd0, 27'h00000062, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001fb, 4'd10, 27'h0000011c, 4'd8, 27'h00000128, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000024, 4'd12, 27'h00000051, 4'd11, 27'h000000ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001a3, 4'd2, 27'h000001fe, 4'd2, 27'h00000053, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000380, 4'd3, 27'h00000394, 4'd7, 27'h000001cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000332, 4'd1, 27'h0000012f, 4'd13, 27'h000002b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000042, 4'd6, 27'h000002ba, 4'd2, 27'h0000014a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000345, 4'd9, 27'h00000244, 4'd6, 27'h00000278, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000037c, 4'd5, 27'h00000396, 4'd13, 27'h0000008b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000391, 4'd12, 27'h0000005a, 4'd1, 27'h000001fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001b8, 4'd14, 27'h000003b0, 4'd7, 27'h0000020e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000003, 4'd14, 27'h000000dc, 4'd11, 27'h000001d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000009c, 4'd3, 27'h00000226, 4'd3, 27'h00000135, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000c8, 4'd2, 27'h00000100, 4'd5, 27'h000001f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000249, 4'd1, 27'h00000232, 4'd11, 27'h00000055, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000013f, 4'd7, 27'h000003b7, 4'd1, 27'h00000386, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000040, 4'd9, 27'h000000c2, 4'd6, 27'h0000023d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000012d, 4'd9, 27'h00000350, 4'd14, 27'h00000042, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001aa, 4'd13, 27'h00000001, 4'd0, 27'h000001c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000048, 4'd10, 27'h00000213, 4'd8, 27'h000002db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000015c, 4'd11, 27'h0000027a, 4'd10, 27'h00000243, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002f9, 4'd2, 27'h00000182, 4'd1, 27'h00000045, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000009d, 4'd3, 27'h0000010b, 4'd9, 27'h00000292, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000203, 4'd4, 27'h00000083, 4'd14, 27'h000003c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001d5, 4'd6, 27'h000003d8, 4'd1, 27'h000000e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000019f, 4'd8, 27'h000003f8, 4'd9, 27'h00000394, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000000c, 4'd8, 27'h0000037d, 4'd14, 27'h00000069, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001e9, 4'd13, 27'h00000376, 4'd4, 27'h00000142, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000271, 4'd12, 27'h000002c5, 4'd8, 27'h000000aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000081, 4'd11, 27'h00000174, 4'd14, 27'h00000398, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000024a, 4'd2, 27'h000001d2, 4'd0, 27'h0000026a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000392, 4'd4, 27'h0000009e, 4'd8, 27'h000003a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000024b, 4'd4, 27'h000001cf, 4'd10, 27'h00000148, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000119, 4'd5, 27'h0000003e, 4'd3, 27'h000001cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003c9, 4'd6, 27'h0000013d, 4'd9, 27'h000002f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000000, 4'd8, 27'h0000018b, 4'd10, 27'h00000313, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003aa, 4'd14, 27'h000003ea, 4'd0, 27'h000003ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000002c, 4'd11, 27'h000001fb, 4'd7, 27'h00000332, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000396, 4'd10, 27'h000002df, 4'd10, 27'h000000e0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000052, 4'd2, 27'h000002dd, 4'd3, 27'h000001b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000175, 4'd0, 27'h00000296, 4'd8, 27'h00000192, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000c6, 4'd2, 27'h000000fc, 4'd12, 27'h000001f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000025, 4'd9, 27'h0000021c, 4'd2, 27'h000000a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000137, 4'd7, 27'h00000169, 4'd5, 27'h00000360, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001e0, 4'd9, 27'h00000201, 4'd10, 27'h000001ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000305, 4'd14, 27'h000001b0, 4'd4, 27'h00000224, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000266, 4'd14, 27'h00000204, 4'd9, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001bb, 4'd13, 27'h000003cf, 4'd10, 27'h000000d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000153, 4'd4, 27'h00000351, 4'd4, 27'h0000013b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000007f, 4'd1, 27'h0000016d, 4'd5, 27'h00000183, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000305, 4'd2, 27'h00000377, 4'd13, 27'h00000390, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000039a, 4'd6, 27'h000002d9, 4'd2, 27'h000002fe, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000130, 4'd7, 27'h0000002e, 4'd9, 27'h000003af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000028f, 4'd5, 27'h00000394, 4'd13, 27'h000000b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001e2, 4'd12, 27'h00000286, 4'd0, 27'h000002b3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000027b, 4'd12, 27'h00000238, 4'd5, 27'h0000019a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002cd, 4'd11, 27'h00000195, 4'd14, 27'h000001ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002ab, 4'd2, 27'h000001ef, 4'd0, 27'h00000297, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000002d, 4'd4, 27'h00000284, 4'd6, 27'h000002b8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000209, 4'd2, 27'h00000355, 4'd10, 27'h00000315, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000015, 4'd8, 27'h000002dc, 4'd3, 27'h00000183, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000017d, 4'd7, 27'h0000023f, 4'd9, 27'h0000024b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000150, 4'd7, 27'h00000213, 4'd11, 27'h0000035b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000ef, 4'd10, 27'h00000059, 4'd0, 27'h000003e5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001bf, 4'd12, 27'h0000032f, 4'd6, 27'h000000a0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000343, 4'd13, 27'h000003aa, 4'd14, 27'h0000001f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003a8, 4'd2, 27'h00000291, 4'd0, 27'h00000165, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001ae, 4'd0, 27'h000003d5, 4'd5, 27'h0000006c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000026d, 4'd1, 27'h000002d7, 4'd12, 27'h00000238, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000022d, 4'd5, 27'h000000bf, 4'd3, 27'h00000391, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000ab, 4'd6, 27'h000002ce, 4'd9, 27'h000001aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000191, 4'd5, 27'h000003c3, 4'd13, 27'h00000218, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000067, 4'd12, 27'h000002f8, 4'd4, 27'h000000c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000013e, 4'd12, 27'h0000019c, 4'd5, 27'h00000368, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000105, 4'd11, 27'h00000160, 4'd14, 27'h000001ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000132, 4'd1, 27'h0000020a, 4'd2, 27'h0000034b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000080, 4'd4, 27'h00000269, 4'd6, 27'h0000025d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000026, 4'd1, 27'h0000020f, 4'd13, 27'h000002f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000305, 4'd7, 27'h0000009b, 4'd0, 27'h0000008e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001a0, 4'd8, 27'h00000105, 4'd8, 27'h00000139, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001d5, 4'd8, 27'h0000039f, 4'd12, 27'h00000005, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001bf, 4'd13, 27'h000002d3, 4'd4, 27'h0000010d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003d7, 4'd14, 27'h00000173, 4'd9, 27'h0000006d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000279, 4'd14, 27'h00000158, 4'd10, 27'h00000130, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000158, 4'd0, 27'h000003c5, 4'd3, 27'h00000045, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003f1, 4'd1, 27'h0000039f, 4'd9, 27'h0000004d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000ff, 4'd0, 27'h00000006, 4'd13, 27'h00000213, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003b4, 4'd6, 27'h0000016a, 4'd4, 27'h000001d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000007d, 4'd6, 27'h0000001c, 4'd6, 27'h0000020a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000224, 4'd6, 27'h00000296, 4'd10, 27'h00000115, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001a1, 4'd10, 27'h000002d2, 4'd4, 27'h000001ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b8, 4'd12, 27'h00000155, 4'd5, 27'h00000333, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000003f, 4'd13, 27'h00000232, 4'd14, 27'h000000a7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000ab, 4'd4, 27'h00000237, 4'd2, 27'h00000249, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002dd, 4'd2, 27'h00000377, 4'd5, 27'h000001a3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001ee, 4'd4, 27'h0000032b, 4'd10, 27'h0000011d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001e8, 4'd8, 27'h00000254, 4'd1, 27'h000000c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003df, 4'd9, 27'h000001de, 4'd5, 27'h0000014f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000ab, 4'd7, 27'h0000004c, 4'd10, 27'h0000002e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000036, 4'd11, 27'h00000384, 4'd3, 27'h000003ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000050, 4'd12, 27'h00000172, 4'd6, 27'h000003e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000041, 4'd10, 27'h000000ef, 4'd14, 27'h000002f6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000115, 4'd4, 27'h00000255, 4'd4, 27'h000003b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000369, 4'd4, 27'h000002cf, 4'd7, 27'h000001ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000288, 4'd1, 27'h000003fb, 4'd13, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000011e, 4'd9, 27'h000003aa, 4'd0, 27'h000003af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000023a, 4'd9, 27'h000000f9, 4'd5, 27'h00000068, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000350, 4'd9, 27'h00000180, 4'd12, 27'h0000026c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002d4, 4'd12, 27'h00000086, 4'd0, 27'h000001d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000090, 4'd10, 27'h000000cc, 4'd9, 27'h00000376, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000304, 4'd12, 27'h00000049, 4'd11, 27'h000003c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000020f, 4'd3, 27'h00000241, 4'd2, 27'h0000024f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000c0, 4'd0, 27'h000003ce, 4'd5, 27'h00000097, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002e8, 4'd3, 27'h0000018e, 4'd11, 27'h0000015a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000203, 4'd8, 27'h000001de, 4'd0, 27'h000002b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000216, 4'd9, 27'h00000341, 4'd8, 27'h0000020d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003ac, 4'd6, 27'h000000da, 4'd13, 27'h0000002a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001ee, 4'd12, 27'h00000092, 4'd4, 27'h000002f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000330, 4'd13, 27'h0000024c, 4'd6, 27'h000003b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000050, 4'd11, 27'h0000016d, 4'd11, 27'h000002ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000009f, 4'd1, 27'h00000165, 4'd4, 27'h0000038a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002b2, 4'd1, 27'h0000016a, 4'd8, 27'h000003f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003d2, 4'd2, 27'h00000262, 4'd12, 27'h00000177, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000021f, 4'd6, 27'h000002f5, 4'd2, 27'h00000371, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000373, 4'd8, 27'h00000025, 4'd5, 27'h0000014a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000317, 4'd5, 27'h00000284, 4'd14, 27'h00000230, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003c5, 4'd14, 27'h000000e1, 4'd0, 27'h000001b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000160, 4'd14, 27'h000001ad, 4'd6, 27'h0000025e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002a9, 4'd13, 27'h000000b6, 4'd10, 27'h00000225, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001a6, 4'd0, 27'h000000e5, 4'd4, 27'h0000011c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000326, 4'd3, 27'h00000119, 4'd9, 27'h00000341, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002e2, 4'd3, 27'h00000398, 4'd10, 27'h000002c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000386, 4'd9, 27'h000001a9, 4'd1, 27'h00000197, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001be, 4'd6, 27'h00000348, 4'd6, 27'h00000318, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000006b, 4'd9, 27'h0000017b, 4'd14, 27'h00000100, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003fa, 4'd14, 27'h000000f4, 4'd2, 27'h000002b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003d7, 4'd13, 27'h00000355, 4'd9, 27'h000002f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000008d, 4'd13, 27'h0000014f, 4'd11, 27'h000003aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000f8, 4'd2, 27'h0000007f, 4'd0, 27'h000000a1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000092, 4'd1, 27'h000000e3, 4'd9, 27'h00000104, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000191, 4'd0, 27'h000003ce, 4'd10, 27'h000003dc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000034b, 4'd6, 27'h0000017f, 4'd0, 27'h000002a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000013a, 4'd6, 27'h00000390, 4'd9, 27'h0000023f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002a5, 4'd8, 27'h000001fa, 4'd11, 27'h00000364, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002e9, 4'd14, 27'h0000029a, 4'd3, 27'h000000f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000287, 4'd14, 27'h0000022c, 4'd8, 27'h000000f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000002f, 4'd11, 27'h000000be, 4'd13, 27'h000001c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000016d, 4'd4, 27'h0000001a, 4'd2, 27'h00000189, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000154, 4'd3, 27'h00000300, 4'd6, 27'h00000314, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003b3, 4'd0, 27'h0000011e, 4'd12, 27'h00000380, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000344, 4'd7, 27'h00000296, 4'd3, 27'h00000162, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002c0, 4'd8, 27'h0000019e, 4'd9, 27'h0000002e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000052, 4'd8, 27'h0000032b, 4'd13, 27'h0000017f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000007e, 4'd10, 27'h00000310, 4'd2, 27'h000001a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000163, 4'd14, 27'h0000032b, 4'd8, 27'h00000108, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000017d, 4'd10, 27'h00000131, 4'd12, 27'h0000032d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000005d, 4'd0, 27'h00000236, 4'd2, 27'h000001c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000090, 4'd1, 27'h00000033, 4'd9, 27'h00000117, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000312, 4'd1, 27'h0000035c, 4'd12, 27'h000001d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000372, 4'd9, 27'h000002cf, 4'd1, 27'h0000000b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c4, 4'd6, 27'h000003c5, 4'd9, 27'h000001a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000005d, 4'd8, 27'h00000146, 4'd10, 27'h00000115, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000262, 4'd10, 27'h000003fb, 4'd2, 27'h0000011c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000f3, 4'd11, 27'h00000222, 4'd5, 27'h000002bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000029a, 4'd10, 27'h00000251, 4'd13, 27'h00000283, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001d8, 4'd1, 27'h00000366, 4'd0, 27'h00000382, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000298, 4'd3, 27'h00000350, 4'd7, 27'h0000021d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000000a, 4'd1, 27'h0000018d, 4'd14, 27'h0000006e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000005, 4'd5, 27'h000000a4, 4'd0, 27'h000000dd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000006f, 4'd7, 27'h00000209, 4'd6, 27'h00000331, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000332, 4'd5, 27'h00000349, 4'd11, 27'h00000220, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000023b, 4'd12, 27'h000001f2, 4'd4, 27'h0000018e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003fd, 4'd11, 27'h00000400, 4'd5, 27'h0000035f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000ea, 4'd12, 27'h000003fb, 4'd14, 27'h000003e8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002cf, 4'd4, 27'h0000001e, 4'd0, 27'h00000181, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000a3, 4'd3, 27'h00000211, 4'd8, 27'h000002b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000ca, 4'd2, 27'h00000282, 4'd12, 27'h000001f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000013d, 4'd6, 27'h000000e6, 4'd2, 27'h00000171, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000018c, 4'd7, 27'h000003b3, 4'd9, 27'h0000036e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000032, 4'd7, 27'h00000226, 4'd13, 27'h00000372, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000233, 4'd12, 27'h00000266, 4'd3, 27'h000002cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003c5, 4'd12, 27'h0000020c, 4'd6, 27'h000003b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000017f, 4'd13, 27'h00000070, 4'd10, 27'h00000067, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003d7, 4'd1, 27'h000003f1, 4'd1, 27'h000002c7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001ed, 4'd0, 27'h000002cb, 4'd9, 27'h0000021e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000268, 4'd1, 27'h000001a9, 4'd11, 27'h00000125, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000034f, 4'd8, 27'h000000bd, 4'd2, 27'h0000033d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001c6, 4'd5, 27'h00000259, 4'd9, 27'h00000264, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000069, 4'd9, 27'h0000011f, 4'd10, 27'h0000005d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000014, 4'd11, 27'h00000386, 4'd3, 27'h000003e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003ae, 4'd13, 27'h000002a1, 4'd7, 27'h00000044, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000323, 4'd11, 27'h000001be, 4'd14, 27'h00000347, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002a7, 4'd2, 27'h00000351, 4'd0, 27'h0000022e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000023a, 4'd1, 27'h000003b6, 4'd5, 27'h000000a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000031a, 4'd1, 27'h00000289, 4'd13, 27'h000003e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000239, 4'd6, 27'h000003a5, 4'd1, 27'h00000079, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000018b, 4'd7, 27'h000001a7, 4'd6, 27'h00000369, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000235, 4'd7, 27'h0000016f, 4'd14, 27'h000003b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000239, 4'd11, 27'h00000343, 4'd4, 27'h000001fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000111, 4'd10, 27'h00000075, 4'd6, 27'h00000029, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000257, 4'd11, 27'h00000029, 4'd12, 27'h0000007b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001e5, 4'd3, 27'h00000229, 4'd4, 27'h00000211, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002c3, 4'd3, 27'h0000027e, 4'd8, 27'h000001b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001da, 4'd3, 27'h00000087, 4'd13, 27'h000001c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000133, 4'd5, 27'h0000002b, 4'd4, 27'h000003e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000021c, 4'd8, 27'h0000032e, 4'd8, 27'h000003ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001e5, 4'd5, 27'h00000262, 4'd13, 27'h0000038a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000039e, 4'd10, 27'h00000290, 4'd4, 27'h000003c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002c2, 4'd13, 27'h000000f4, 4'd7, 27'h000000c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000ff, 4'd12, 27'h00000276, 4'd13, 27'h000001a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000014, 4'd3, 27'h00000198, 4'd3, 27'h000003f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002d4, 4'd1, 27'h0000008a, 4'd6, 27'h0000016e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000006e, 4'd3, 27'h000001ec, 4'd10, 27'h00000333, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000bc, 4'd9, 27'h00000072, 4'd4, 27'h00000235, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000067, 4'd7, 27'h0000035e, 4'd5, 27'h0000000b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000007a, 4'd7, 27'h00000247, 4'd12, 27'h000002df, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000239, 4'd11, 27'h0000030c, 4'd4, 27'h00000101, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003a1, 4'd14, 27'h000002ef, 4'd9, 27'h0000030d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000005a, 4'd11, 27'h000003bc, 4'd10, 27'h00000033, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000349, 4'd1, 27'h000003ef, 4'd0, 27'h000000c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000101, 4'd0, 27'h00000174, 4'd7, 27'h00000271, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000030b, 4'd0, 27'h00000355, 4'd13, 27'h0000037c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001ca, 4'd5, 27'h00000189, 4'd3, 27'h000001c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001ee, 4'd8, 27'h000001ea, 4'd9, 27'h00000203, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000008b, 4'd8, 27'h000000dd, 4'd10, 27'h00000025, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002c3, 4'd11, 27'h000001a8, 4'd1, 27'h00000353, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000010b, 4'd13, 27'h0000029c, 4'd8, 27'h0000004a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000006c, 4'd13, 27'h0000023a, 4'd12, 27'h000000c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000097, 4'd2, 27'h0000033c, 4'd4, 27'h0000018a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001f7, 4'd0, 27'h00000161, 4'd8, 27'h000003e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000c6, 4'd4, 27'h0000028d, 4'd14, 27'h00000263, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000048, 4'd9, 27'h000003f8, 4'd3, 27'h0000018b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000187, 4'd7, 27'h00000363, 4'd5, 27'h0000030d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000002b, 4'd5, 27'h000000d8, 4'd10, 27'h00000033, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000391, 4'd13, 27'h00000269, 4'd2, 27'h00000117, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000149, 4'd14, 27'h00000271, 4'd5, 27'h0000004c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001be, 4'd14, 27'h0000014d, 4'd10, 27'h000003c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ed, 4'd1, 27'h0000031c, 4'd3, 27'h000001e2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000013d, 4'd4, 27'h00000398, 4'd6, 27'h000002ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000012e, 4'd3, 27'h00000336, 4'd13, 27'h0000017a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000340, 4'd6, 27'h00000241, 4'd1, 27'h0000000a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003e7, 4'd7, 27'h00000332, 4'd9, 27'h000003a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000110, 4'd8, 27'h000001e5, 4'd14, 27'h00000233, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001bc, 4'd13, 27'h00000125, 4'd4, 27'h000002e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000322, 4'd10, 27'h00000087, 4'd5, 27'h0000039e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000019, 4'd11, 27'h000001fa, 4'd13, 27'h00000009, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000016d, 4'd3, 27'h000001ab, 4'd3, 27'h00000270, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002dd, 4'd3, 27'h000001e4, 4'd9, 27'h000001c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002be, 4'd0, 27'h0000010c, 4'd10, 27'h00000177, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000023, 4'd9, 27'h000003cd, 4'd4, 27'h00000117, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000201, 4'd9, 27'h00000390, 4'd6, 27'h00000149, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000031b, 4'd5, 27'h000001ec, 4'd11, 27'h0000037c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001c8, 4'd13, 27'h00000312, 4'd1, 27'h0000015e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000032c, 4'd11, 27'h0000013f, 4'd8, 27'h000001fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ff, 4'd13, 27'h000002d0, 4'd11, 27'h00000364, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000019a, 4'd3, 27'h000003ae, 4'd1, 27'h0000030e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000002c, 4'd3, 27'h00000029, 4'd6, 27'h000003c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002ff, 4'd3, 27'h00000068, 4'd14, 27'h000002d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001e2, 4'd5, 27'h000003ea, 4'd1, 27'h00000306, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000039f, 4'd8, 27'h000001e0, 4'd7, 27'h000002a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001bf, 4'd7, 27'h000001d1, 4'd12, 27'h0000028b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000278, 4'd14, 27'h0000004b, 4'd1, 27'h000000ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000280, 4'd11, 27'h000002cb, 4'd5, 27'h000000d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000032f, 4'd14, 27'h000000ac, 4'd11, 27'h000000d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000035f, 4'd0, 27'h000003d2, 4'd0, 27'h00000230, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000186, 4'd4, 27'h000002e2, 4'd9, 27'h000001ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000002d, 4'd2, 27'h00000177, 4'd14, 27'h00000351, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000327, 4'd5, 27'h00000396, 4'd0, 27'h0000014f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001b0, 4'd9, 27'h00000043, 4'd6, 27'h0000005b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000163, 4'd6, 27'h000001fe, 4'd13, 27'h000002e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000014b, 4'd10, 27'h000003ab, 4'd3, 27'h000002c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000024b, 4'd14, 27'h0000013b, 4'd8, 27'h0000025e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000106, 4'd14, 27'h000003b8, 4'd10, 27'h0000031c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002b2, 4'd4, 27'h000000ba, 4'd2, 27'h00000191, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002b7, 4'd2, 27'h0000037a, 4'd7, 27'h00000382, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000007f, 4'd2, 27'h0000029e, 4'd14, 27'h0000013b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003f2, 4'd5, 27'h000001e3, 4'd3, 27'h000002fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001c5, 4'd6, 27'h00000260, 4'd9, 27'h000003aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000335, 4'd7, 27'h000000a1, 4'd11, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000002f, 4'd13, 27'h00000334, 4'd0, 27'h000001e5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000293, 4'd13, 27'h000002ae, 4'd8, 27'h000002ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000004, 4'd12, 27'h000003df, 4'd11, 27'h0000029e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000026c, 4'd0, 27'h000000f1, 4'd1, 27'h0000004a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000199, 4'd3, 27'h00000000, 4'd9, 27'h000003b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000330, 4'd2, 27'h0000000e, 4'd10, 27'h0000035a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000184, 4'd7, 27'h0000034b, 4'd1, 27'h0000015a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003d3, 4'd6, 27'h000003ab, 4'd9, 27'h0000032e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000006d, 4'd7, 27'h00000123, 4'd12, 27'h0000032d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000126, 4'd11, 27'h0000023f, 4'd0, 27'h00000119, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000378, 4'd10, 27'h0000026b, 4'd7, 27'h00000294, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000142, 4'd13, 27'h000002d7, 4'd10, 27'h0000007b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000035c, 4'd0, 27'h0000038d, 4'd0, 27'h00000099, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003e2, 4'd0, 27'h0000022e, 4'd8, 27'h0000023a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001ae, 4'd1, 27'h00000288, 4'd10, 27'h00000392, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000070, 4'd8, 27'h0000016a, 4'd1, 27'h00000093, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003b6, 4'd7, 27'h00000310, 4'd6, 27'h00000000, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000a8, 4'd6, 27'h00000379, 4'd13, 27'h00000008, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000339, 4'd14, 27'h000002b7, 4'd2, 27'h00000359, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000230, 4'd11, 27'h00000145, 4'd7, 27'h00000377, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000269, 4'd12, 27'h00000345, 4'd14, 27'h000000c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000029a, 4'd1, 27'h0000009c, 4'd0, 27'h00000142, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000001d, 4'd0, 27'h00000367, 4'd8, 27'h0000000c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000039e, 4'd0, 27'h000001ea, 4'd14, 27'h00000037, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000ae, 4'd9, 27'h0000019e, 4'd1, 27'h000000c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003e0, 4'd6, 27'h00000002, 4'd5, 27'h0000012b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000016d, 4'd7, 27'h00000357, 4'd11, 27'h00000115, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002c5, 4'd14, 27'h0000009d, 4'd3, 27'h00000056, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000036a, 4'd10, 27'h00000329, 4'd5, 27'h00000194, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000013, 4'd12, 27'h00000339, 4'd10, 27'h00000168, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000014, 4'd3, 27'h000002c1, 4'd1, 27'h000001b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000170, 4'd4, 27'h00000222, 4'd6, 27'h00000044, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000132, 4'd2, 27'h0000022e, 4'd12, 27'h00000206, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000318, 4'd5, 27'h000001f5, 4'd2, 27'h000001f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000310, 4'd5, 27'h000000dc, 4'd9, 27'h00000071, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000028c, 4'd8, 27'h000002b7, 4'd13, 27'h00000295, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001c9, 4'd13, 27'h000003ea, 4'd4, 27'h0000002f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002ff, 4'd10, 27'h00000190, 4'd5, 27'h000000b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000e9, 4'd11, 27'h000003a2, 4'd10, 27'h000000a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000002, 4'd3, 27'h00000319, 4'd1, 27'h00000091, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000130, 4'd4, 27'h00000391, 4'd9, 27'h00000391, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000008c, 4'd3, 27'h00000277, 4'd14, 27'h0000002f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000281, 4'd9, 27'h000002c6, 4'd1, 27'h000002fb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000007e, 4'd8, 27'h000002ac, 4'd6, 27'h00000308, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001d7, 4'd5, 27'h000000cd, 4'd14, 27'h00000119, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002f2, 4'd10, 27'h00000135, 4'd3, 27'h000001d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001a7, 4'd10, 27'h00000241, 4'd5, 27'h000000b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000200, 4'd11, 27'h00000125, 4'd11, 27'h00000016, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000172, 4'd3, 27'h0000003d, 4'd3, 27'h0000014b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000060, 4'd1, 27'h00000091, 4'd7, 27'h00000339, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002bc, 4'd1, 27'h0000038a, 4'd12, 27'h000003b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b4, 4'd7, 27'h00000025, 4'd3, 27'h00000021, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002f8, 4'd6, 27'h0000027b, 4'd5, 27'h00000291, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000353, 4'd7, 27'h000002e6, 4'd10, 27'h000000cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000189, 4'd10, 27'h000001a3, 4'd2, 27'h000000c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000325, 4'd13, 27'h000001ab, 4'd7, 27'h00000248, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000039b, 4'd13, 27'h00000323, 4'd10, 27'h00000238, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000347, 4'd2, 27'h00000251, 4'd1, 27'h000000b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000010e, 4'd2, 27'h0000007a, 4'd7, 27'h00000070, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000160, 4'd4, 27'h00000063, 4'd11, 27'h0000039d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000202, 4'd6, 27'h000002a4, 4'd2, 27'h000001bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000023, 4'd8, 27'h0000007a, 4'd9, 27'h000003e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000010d, 4'd8, 27'h00000041, 4'd12, 27'h00000179, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003e3, 4'd11, 27'h000000ef, 4'd4, 27'h0000033d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000295, 4'd14, 27'h00000126, 4'd7, 27'h000002e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000034c, 4'd14, 27'h00000343, 4'd11, 27'h000002e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000087, 4'd3, 27'h0000021a, 4'd2, 27'h00000238, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002ab, 4'd4, 27'h0000039d, 4'd9, 27'h0000018f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000379, 4'd4, 27'h000002d4, 4'd11, 27'h00000242, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000037d, 4'd7, 27'h000001bc, 4'd4, 27'h00000212, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000052, 4'd7, 27'h000002f1, 4'd6, 27'h0000039f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000026b, 4'd9, 27'h0000032f, 4'd13, 27'h0000019b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002b2, 4'd10, 27'h00000086, 4'd0, 27'h000001bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000083, 4'd11, 27'h000003fc, 4'd9, 27'h00000206, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003ff, 4'd11, 27'h000000c1, 4'd14, 27'h00000256, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000001d, 4'd0, 27'h0000035e, 4'd0, 27'h0000030e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000314, 4'd3, 27'h000002e1, 4'd9, 27'h0000009f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000d2, 4'd3, 27'h00000094, 4'd13, 27'h0000011b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000ca, 4'd8, 27'h000001b8, 4'd0, 27'h00000017, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000039a, 4'd8, 27'h00000000, 4'd6, 27'h00000324, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001a4, 4'd8, 27'h00000107, 4'd13, 27'h00000200, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003a0, 4'd10, 27'h000000d3, 4'd4, 27'h000001b8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000020, 4'd10, 27'h00000193, 4'd5, 27'h000002f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000032e, 4'd14, 27'h000000e0, 4'd14, 27'h0000009e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000012d, 4'd3, 27'h000001c0, 4'd4, 27'h00000093, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000071, 4'd0, 27'h000003a4, 4'd9, 27'h000001c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001e3, 4'd1, 27'h000001c2, 4'd14, 27'h00000235, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002a6, 4'd8, 27'h00000344, 4'd0, 27'h0000004a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001f9, 4'd8, 27'h000002aa, 4'd6, 27'h0000019f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000392, 4'd9, 27'h000003fa, 4'd14, 27'h000001df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000039a, 4'd13, 27'h00000056, 4'd0, 27'h000002f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000144, 4'd13, 27'h000001be, 4'd5, 27'h00000343, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000071, 4'd11, 27'h000002e8, 4'd10, 27'h000000da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002cd, 4'd3, 27'h00000200, 4'd2, 27'h000000c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000227, 4'd3, 27'h0000030b, 4'd9, 27'h00000116, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000170, 4'd2, 27'h000003f2, 4'd10, 27'h00000377, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000de, 4'd6, 27'h000001b8, 4'd2, 27'h00000374, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000023, 4'd8, 27'h00000075, 4'd8, 27'h000001de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003e0, 4'd7, 27'h00000384, 4'd11, 27'h00000317, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000314, 4'd10, 27'h00000309, 4'd4, 27'h00000109, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000205, 4'd13, 27'h00000068, 4'd5, 27'h00000320, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000006e, 4'd10, 27'h000000f9, 4'd13, 27'h0000022e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000fb, 4'd2, 27'h0000028c, 4'd0, 27'h000003a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000002f, 4'd4, 27'h0000007d, 4'd9, 27'h00000108, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000266, 4'd4, 27'h000001b6, 4'd11, 27'h0000014f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000204, 4'd5, 27'h00000003, 4'd4, 27'h000000cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003f4, 4'd8, 27'h000003a7, 4'd9, 27'h00000111, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000031b, 4'd8, 27'h00000211, 4'd10, 27'h000000c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003ae, 4'd12, 27'h0000029e, 4'd0, 27'h00000331, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000026b, 4'd13, 27'h000000c9, 4'd9, 27'h0000026c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000335, 4'd14, 27'h00000230, 4'd11, 27'h0000022c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000025d, 4'd1, 27'h00000038, 4'd1, 27'h000003fb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000245, 4'd1, 27'h000002b3, 4'd8, 27'h000000c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000008e, 4'd4, 27'h000002de, 4'd14, 27'h000003c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000262, 4'd7, 27'h000002a0, 4'd4, 27'h0000031a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000387, 4'd9, 27'h000003de, 4'd9, 27'h000001d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000197, 4'd9, 27'h00000256, 4'd11, 27'h00000225, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ef, 4'd14, 27'h0000024f, 4'd3, 27'h0000022b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003e6, 4'd13, 27'h0000008c, 4'd6, 27'h00000274, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000016e, 4'd13, 27'h00000089, 4'd10, 27'h00000091, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000000f, 4'd3, 27'h0000020b, 4'd4, 27'h00000186, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003cc, 4'd3, 27'h0000026b, 4'd6, 27'h000002ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002ee, 4'd3, 27'h00000311, 4'd14, 27'h0000034e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000023c, 4'd6, 27'h000001c9, 4'd0, 27'h000001f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000001c, 4'd5, 27'h000001c7, 4'd5, 27'h00000155, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000394, 4'd5, 27'h00000105, 4'd14, 27'h000000a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000e9, 4'd13, 27'h0000039c, 4'd1, 27'h00000132, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000d4, 4'd13, 27'h000003eb, 4'd7, 27'h00000350, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000376, 4'd11, 27'h00000342, 4'd12, 27'h000000ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000034e, 4'd4, 27'h0000020f, 4'd0, 27'h00000371, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000368, 4'd2, 27'h000003e9, 4'd9, 27'h0000001d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002ac, 4'd3, 27'h000002ca, 4'd14, 27'h0000000d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000f1, 4'd5, 27'h000001f8, 4'd4, 27'h000001ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000203, 4'd9, 27'h00000352, 4'd5, 27'h000003f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000002f, 4'd8, 27'h000003b5, 4'd12, 27'h0000011b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000029a, 4'd13, 27'h000002d2, 4'd4, 27'h000003d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001d5, 4'd13, 27'h00000253, 4'd9, 27'h000001ff, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000367, 4'd12, 27'h0000038f, 4'd12, 27'h00000233, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000169, 4'd4, 27'h00000003, 4'd4, 27'h00000146, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000313, 4'd3, 27'h00000078, 4'd8, 27'h000000e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000001d, 4'd3, 27'h000000cc, 4'd12, 27'h00000270, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001e0, 4'd6, 27'h00000172, 4'd2, 27'h00000041, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000257, 4'd9, 27'h0000007c, 4'd8, 27'h0000039a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003f1, 4'd6, 27'h000000a4, 4'd13, 27'h00000325, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000229, 4'd13, 27'h00000249, 4'd4, 27'h000000e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001d1, 4'd12, 27'h00000365, 4'd9, 27'h00000251, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003f5, 4'd14, 27'h00000356, 4'd13, 27'h00000328, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000216, 4'd4, 27'h0000019f, 4'd1, 27'h0000007b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ae, 4'd0, 27'h000000ef, 4'd8, 27'h000000ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000332, 4'd2, 27'h00000015, 4'd13, 27'h00000167, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002d3, 4'd5, 27'h00000298, 4'd4, 27'h00000163, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000001a, 4'd8, 27'h000003b0, 4'd5, 27'h000002d2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000293, 4'd8, 27'h000003a7, 4'd11, 27'h0000037b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000277, 4'd11, 27'h00000340, 4'd1, 27'h000000e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000023d, 4'd12, 27'h00000046, 4'd9, 27'h00000159, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000012c, 4'd11, 27'h00000122, 4'd13, 27'h0000026f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003d4, 4'd4, 27'h0000035a, 4'd0, 27'h0000019e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000255, 4'd4, 27'h00000194, 4'd8, 27'h000002d6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000073, 4'd1, 27'h00000304, 4'd13, 27'h00000393, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000033, 4'd7, 27'h00000285, 4'd2, 27'h00000179, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000f0, 4'd9, 27'h00000375, 4'd8, 27'h00000393, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000122, 4'd8, 27'h0000014c, 4'd12, 27'h0000000f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000007b, 4'd13, 27'h000001c1, 4'd3, 27'h000003e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000029b, 4'd12, 27'h00000283, 4'd9, 27'h000001a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000029f, 4'd14, 27'h000000b4, 4'd12, 27'h000002e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000028d, 4'd3, 27'h000001da, 4'd4, 27'h00000289, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000020d, 4'd1, 27'h000002cc, 4'd6, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000151, 4'd1, 27'h00000326, 4'd12, 27'h000003f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000003c, 4'd8, 27'h0000004d, 4'd0, 27'h00000234, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000d0, 4'd5, 27'h00000150, 4'd8, 27'h000001e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002ec, 4'd6, 27'h000002ac, 4'd12, 27'h0000018b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000284, 4'd11, 27'h000001d6, 4'd1, 27'h000003b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000176, 4'd12, 27'h000001d5, 4'd8, 27'h000001c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000d5, 4'd11, 27'h00000266, 4'd10, 27'h0000019c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000297, 4'd4, 27'h00000307, 4'd2, 27'h000001ff, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000013f, 4'd2, 27'h0000030a, 4'd9, 27'h0000002f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000376, 4'd1, 27'h00000167, 4'd13, 27'h00000329, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002fb, 4'd6, 27'h00000054, 4'd0, 27'h0000021a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000031b, 4'd7, 27'h000003ae, 4'd8, 27'h000000af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000dd, 4'd6, 27'h00000013, 4'd10, 27'h00000270, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000bc, 4'd11, 27'h000002ff, 4'd4, 27'h00000341, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000019f, 4'd12, 27'h000002e9, 4'd5, 27'h000000c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000122, 4'd12, 27'h00000210, 4'd10, 27'h00000383, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000066, 4'd0, 27'h000003bb, 4'd2, 27'h00000272, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000018b, 4'd3, 27'h00000020, 4'd8, 27'h0000019e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000369, 4'd4, 27'h00000126, 4'd13, 27'h0000005c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000dc, 4'd6, 27'h000000ce, 4'd4, 27'h000003fb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000232, 4'd5, 27'h000001e3, 4'd9, 27'h000001b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000197, 4'd7, 27'h000003c3, 4'd13, 27'h000003cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001bf, 4'd13, 27'h00000148, 4'd1, 27'h00000088, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000010a, 4'd13, 27'h00000255, 4'd6, 27'h00000175, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000088, 4'd14, 27'h0000023b, 4'd10, 27'h000003ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000221, 4'd0, 27'h00000294, 4'd4, 27'h00000232, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000205, 4'd4, 27'h0000024c, 4'd9, 27'h000000f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003d3, 4'd4, 27'h000002d3, 4'd14, 27'h000001bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000251, 4'd7, 27'h000002c1, 4'd2, 27'h0000008f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000c5, 4'd7, 27'h0000012e, 4'd5, 27'h000000e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000265, 4'd8, 27'h0000016a, 4'd12, 27'h00000288, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000032c, 4'd11, 27'h000003e0, 4'd0, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000067, 4'd13, 27'h00000185, 4'd9, 27'h000001db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000023, 4'd11, 27'h000002e4, 4'd14, 27'h00000292, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001b3, 4'd1, 27'h000003fe, 4'd4, 27'h000001e3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003da, 4'd2, 27'h0000030e, 4'd9, 27'h00000028, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002e2, 4'd3, 27'h000003e0, 4'd11, 27'h000002f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000094, 4'd6, 27'h000000a7, 4'd1, 27'h00000096, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000001c, 4'd8, 27'h00000392, 4'd5, 27'h000002c4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000a6, 4'd9, 27'h0000010a, 4'd11, 27'h000002d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003e2, 4'd11, 27'h0000028d, 4'd4, 27'h00000059, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000184, 4'd13, 27'h000002d9, 4'd7, 27'h000002ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000dd, 4'd11, 27'h000002ae, 4'd10, 27'h0000031a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000245, 4'd2, 27'h00000234, 4'd1, 27'h000001e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000033c, 4'd2, 27'h00000285, 4'd8, 27'h00000126, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000384, 4'd1, 27'h00000346, 4'd13, 27'h00000328, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000a4, 4'd8, 27'h000000a2, 4'd3, 27'h000000d2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000a8, 4'd8, 27'h0000033a, 4'd6, 27'h000003b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000b7, 4'd7, 27'h00000021, 4'd12, 27'h00000270, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000038, 4'd11, 27'h000002cf, 4'd4, 27'h00000231, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000229, 4'd13, 27'h00000299, 4'd8, 27'h000002cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000258, 4'd13, 27'h0000024a, 4'd10, 27'h0000004c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002ef, 4'd0, 27'h0000020c, 4'd2, 27'h000000f4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003a6, 4'd4, 27'h000003b8, 4'd5, 27'h000000b3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000328, 4'd3, 27'h00000338, 4'd11, 27'h00000059, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002da, 4'd8, 27'h00000093, 4'd3, 27'h000002cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000102, 4'd6, 27'h0000003b, 4'd8, 27'h0000011d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000010d, 4'd8, 27'h000001c2, 4'd12, 27'h0000003f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000391, 4'd12, 27'h000001ad, 4'd4, 27'h00000081, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003a6, 4'd10, 27'h000001ac, 4'd8, 27'h0000010d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003fd, 4'd10, 27'h000001bf, 4'd10, 27'h0000011e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000024, 4'd3, 27'h00000001, 4'd3, 27'h00000325, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000004d, 4'd0, 27'h000000d8, 4'd6, 27'h0000039f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000324, 4'd1, 27'h00000196, 4'd13, 27'h0000021c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000017b, 4'd9, 27'h0000018c, 4'd1, 27'h00000042, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001bf, 4'd9, 27'h00000171, 4'd9, 27'h00000179, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000358, 4'd6, 27'h000000d1, 4'd11, 27'h000000de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003db, 4'd12, 27'h000001a8, 4'd0, 27'h000001df, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000262, 4'd10, 27'h000002d6, 4'd9, 27'h000001a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003b1, 4'd14, 27'h00000381, 4'd11, 27'h0000006a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000392, 4'd4, 27'h000003f2, 4'd1, 27'h00000144, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001e4, 4'd0, 27'h00000264, 4'd7, 27'h000001ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000d5, 4'd4, 27'h000000e7, 4'd13, 27'h0000024c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003fa, 4'd5, 27'h000000b3, 4'd4, 27'h000002ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003a1, 4'd5, 27'h0000029f, 4'd8, 27'h00000375, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001a8, 4'd7, 27'h00000251, 4'd13, 27'h00000382, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000036, 4'd12, 27'h00000374, 4'd0, 27'h000001d6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000239, 4'd12, 27'h00000152, 4'd7, 27'h00000323, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003fc, 4'd14, 27'h000001ac, 4'd11, 27'h0000017f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000004b, 4'd2, 27'h000000c6, 4'd1, 27'h00000220, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000356, 4'd4, 27'h00000384, 4'd8, 27'h00000386, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002bc, 4'd3, 27'h00000340, 4'd11, 27'h0000006b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000035a, 4'd7, 27'h00000196, 4'd3, 27'h000003a7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000185, 4'd7, 27'h00000078, 4'd5, 27'h00000367, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000219, 4'd6, 27'h0000023f, 4'd13, 27'h000000f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002de, 4'd10, 27'h0000017f, 4'd2, 27'h000002cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000116, 4'd12, 27'h000003bc, 4'd5, 27'h0000023b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000167, 4'd11, 27'h000000f1, 4'd14, 27'h00000120, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002b6, 4'd4, 27'h000002fd, 4'd0, 27'h000000db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000227, 4'd0, 27'h00000391, 4'd9, 27'h0000023a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000033, 4'd0, 27'h0000023b, 4'd10, 27'h00000029, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001ff, 4'd5, 27'h00000364, 4'd0, 27'h000003a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003af, 4'd5, 27'h00000316, 4'd7, 27'h0000013b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000022c, 4'd5, 27'h00000206, 4'd13, 27'h0000005a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000026b, 4'd12, 27'h0000010c, 4'd4, 27'h000003a2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000037e, 4'd11, 27'h000000f5, 4'd8, 27'h000000ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000018d, 4'd13, 27'h00000194, 4'd11, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ad, 4'd0, 27'h00000286, 4'd4, 27'h0000020a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000be, 4'd1, 27'h0000020d, 4'd8, 27'h00000351, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003f2, 4'd1, 27'h000001c9, 4'd13, 27'h000003fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002c3, 4'd8, 27'h00000377, 4'd1, 27'h0000007a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000017f, 4'd9, 27'h0000010b, 4'd7, 27'h00000359, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000006a, 4'd8, 27'h000002da, 4'd10, 27'h00000374, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000019a, 4'd11, 27'h000002ae, 4'd0, 27'h0000031d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000092, 4'd14, 27'h0000020f, 4'd7, 27'h0000018d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000158, 4'd12, 27'h000001ce, 4'd12, 27'h00000100, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000259, 4'd3, 27'h0000014a, 4'd2, 27'h000003a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000aa, 4'd1, 27'h0000016c, 4'd6, 27'h000002a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000039a, 4'd0, 27'h00000252, 4'd11, 27'h000003b0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000da, 4'd6, 27'h00000086, 4'd3, 27'h0000035d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001c0, 4'd5, 27'h00000057, 4'd5, 27'h00000148, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000112, 4'd9, 27'h00000372, 4'd13, 27'h00000138, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000238, 4'd12, 27'h0000029e, 4'd0, 27'h000001f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000049, 4'd11, 27'h00000131, 4'd9, 27'h00000394, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003fa, 4'd14, 27'h00000131, 4'd14, 27'h000000f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003d2, 4'd3, 27'h000001be, 4'd0, 27'h000000c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003e6, 4'd4, 27'h00000299, 4'd9, 27'h00000363, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002ca, 4'd1, 27'h000001c9, 4'd14, 27'h00000395, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003c4, 4'd9, 27'h000003a5, 4'd3, 27'h000002ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002d8, 4'd5, 27'h0000018f, 4'd9, 27'h0000020b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000301, 4'd5, 27'h000000eb, 4'd11, 27'h0000038b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000105, 4'd14, 27'h00000336, 4'd2, 27'h000002ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003e8, 4'd13, 27'h00000165, 4'd7, 27'h000000a4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002cc, 4'd12, 27'h000003b8, 4'd12, 27'h00000377, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002cb, 4'd0, 27'h000001f1, 4'd3, 27'h00000204, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002e9, 4'd0, 27'h00000394, 4'd7, 27'h000001e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000010d, 4'd4, 27'h00000152, 4'd13, 27'h0000032d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001b4, 4'd5, 27'h0000031f, 4'd0, 27'h000002e2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003db, 4'd7, 27'h0000023c, 4'd9, 27'h00000310, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002f4, 4'd5, 27'h00000346, 4'd13, 27'h00000106, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000018d, 4'd12, 27'h00000267, 4'd4, 27'h0000039e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000198, 4'd12, 27'h000001ef, 4'd6, 27'h00000214, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000003b, 4'd11, 27'h000000b7, 4'd12, 27'h00000096, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001ed, 4'd4, 27'h00000273, 4'd0, 27'h00000316, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000264, 4'd4, 27'h000000b1, 4'd9, 27'h000001ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000016d, 4'd3, 27'h000002a5, 4'd14, 27'h0000007a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000039d, 4'd5, 27'h00000289, 4'd2, 27'h00000088, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000004, 4'd9, 27'h0000013f, 4'd7, 27'h00000291, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000132, 4'd6, 27'h000003e7, 4'd10, 27'h000000b8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000365, 4'd12, 27'h000000a2, 4'd2, 27'h0000033e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002f9, 4'd10, 27'h00000313, 4'd6, 27'h000001e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000080, 4'd11, 27'h00000236, 4'd14, 27'h00000193, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003a5, 4'd0, 27'h000001bd, 4'd2, 27'h0000035d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003fe, 4'd1, 27'h000002a9, 4'd8, 27'h00000375, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000156, 4'd2, 27'h000003e2, 4'd12, 27'h00000371, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002d5, 4'd8, 27'h00000104, 4'd4, 27'h00000017, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000038a, 4'd5, 27'h000003ae, 4'd9, 27'h000003a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003a9, 4'd7, 27'h00000239, 4'd11, 27'h00000319, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003bd, 4'd12, 27'h00000170, 4'd3, 27'h000003c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000026a, 4'd13, 27'h000003ef, 4'd8, 27'h000002a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000013d, 4'd13, 27'h000001ad, 4'd10, 27'h0000001c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000038e, 4'd1, 27'h000000e1, 4'd1, 27'h000003b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000288, 4'd1, 27'h00000137, 4'd9, 27'h00000122, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003cb, 4'd0, 27'h00000377, 4'd14, 27'h00000309, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000210, 4'd7, 27'h00000224, 4'd2, 27'h00000154, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000014, 4'd9, 27'h000001a7, 4'd6, 27'h000002ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000377, 4'd9, 27'h0000033c, 4'd11, 27'h00000270, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000b9, 4'd12, 27'h000000c7, 4'd0, 27'h000002a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000179, 4'd13, 27'h000000c2, 4'd8, 27'h00000149, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002e6, 4'd13, 27'h0000012f, 4'd14, 27'h000000c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003a0, 4'd1, 27'h00000003, 4'd0, 27'h000001ae, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000018c, 4'd4, 27'h000002fc, 4'd9, 27'h000001dc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000258, 4'd0, 27'h00000201, 4'd13, 27'h0000016b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002a3, 4'd9, 27'h00000221, 4'd2, 27'h000001af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000082, 4'd8, 27'h0000008e, 4'd7, 27'h000002f1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000a0, 4'd6, 27'h0000015b, 4'd11, 27'h00000338, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000210, 4'd14, 27'h000003e0, 4'd4, 27'h00000072, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000d8, 4'd10, 27'h00000267, 4'd5, 27'h0000026e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000008d, 4'd11, 27'h000001b5, 4'd12, 27'h000003aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000158, 4'd3, 27'h0000022a, 4'd1, 27'h000002e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001ff, 4'd1, 27'h000001fd, 4'd8, 27'h000002e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000033c, 4'd0, 27'h000001df, 4'd12, 27'h0000028f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003b6, 4'd8, 27'h000002cc, 4'd1, 27'h00000362, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000012a, 4'd8, 27'h0000029b, 4'd5, 27'h000003cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000016f, 4'd9, 27'h0000024a, 4'd14, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000068, 4'd14, 27'h000003ad, 4'd0, 27'h000002da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000028e, 4'd10, 27'h0000020f, 4'd5, 27'h00000171, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000298, 4'd10, 27'h00000281, 4'd12, 27'h00000112, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002ca, 4'd2, 27'h0000032d, 4'd1, 27'h0000036f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000a5, 4'd3, 27'h0000023e, 4'd9, 27'h0000030c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000fa, 4'd0, 27'h00000257, 4'd10, 27'h0000025d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000007a, 4'd8, 27'h000000d3, 4'd3, 27'h00000391, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000002e, 4'd9, 27'h000000e1, 4'd9, 27'h000002e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000018, 4'd6, 27'h00000265, 4'd14, 27'h0000016e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000027b, 4'd10, 27'h0000028e, 4'd0, 27'h00000263, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000012f, 4'd11, 27'h00000385, 4'd8, 27'h00000256, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003e9, 4'd13, 27'h000001ac, 4'd13, 27'h0000028b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000217, 4'd0, 27'h0000011c, 4'd4, 27'h0000015f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000316, 4'd0, 27'h000000c8, 4'd9, 27'h00000392, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000029f, 4'd4, 27'h000000e1, 4'd14, 27'h000003d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003b1, 4'd5, 27'h0000020f, 4'd4, 27'h00000382, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000031d, 4'd7, 27'h0000008a, 4'd6, 27'h000001df, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000025b, 4'd5, 27'h000002a7, 4'd12, 27'h00000108, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000207, 4'd14, 27'h0000027d, 4'd2, 27'h000000b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001fd, 4'd12, 27'h0000036c, 4'd9, 27'h000001ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000005d, 4'd13, 27'h000003bc, 4'd12, 27'h000000a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000369, 4'd0, 27'h0000018a, 4'd2, 27'h0000036d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000f0, 4'd4, 27'h00000038, 4'd5, 27'h000002bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000003b, 4'd4, 27'h00000395, 4'd14, 27'h0000039b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000029c, 4'd7, 27'h000002a9, 4'd1, 27'h000001f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000376, 4'd7, 27'h00000269, 4'd6, 27'h00000127, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000099, 4'd7, 27'h0000021d, 4'd11, 27'h0000039f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001d7, 4'd14, 27'h000001ca, 4'd4, 27'h0000012e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000013a, 4'd11, 27'h000003e2, 4'd9, 27'h000002eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000119, 4'd14, 27'h0000024c, 4'd12, 27'h000001ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000290, 4'd0, 27'h000002e8, 4'd4, 27'h000001b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001a9, 4'd3, 27'h00000052, 4'd5, 27'h00000008, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000029c, 4'd0, 27'h00000361, 4'd13, 27'h0000020f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000038d, 4'd8, 27'h000003d7, 4'd0, 27'h00000066, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000107, 4'd6, 27'h000001b5, 4'd8, 27'h00000057, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000020, 4'd8, 27'h00000240, 4'd13, 27'h0000028d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000020b, 4'd11, 27'h000002ca, 4'd0, 27'h000001c0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000028b, 4'd11, 27'h000001c5, 4'd9, 27'h000002f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000180, 4'd13, 27'h00000380, 4'd13, 27'h000003c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000001e, 4'd1, 27'h000003b3, 4'd2, 27'h00000006, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001a2, 4'd4, 27'h000002c0, 4'd6, 27'h00000058, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003d1, 4'd3, 27'h0000018b, 4'd12, 27'h0000030a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000033c, 4'd5, 27'h000003ed, 4'd2, 27'h000001f1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003ae, 4'd5, 27'h0000004b, 4'd9, 27'h00000052, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000f0, 4'd5, 27'h000002d7, 4'd12, 27'h000003ca, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000024f, 4'd10, 27'h00000292, 4'd0, 27'h000001b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000026b, 4'd10, 27'h000003d7, 4'd8, 27'h00000148, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000013f, 4'd11, 27'h000003c5, 4'd11, 27'h000003f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000057, 4'd0, 27'h00000150, 4'd3, 27'h000001cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002b1, 4'd2, 27'h000000b1, 4'd5, 27'h00000029, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000d3, 4'd2, 27'h000001dc, 4'd10, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001e4, 4'd8, 27'h00000022, 4'd1, 27'h00000238, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000019c, 4'd5, 27'h00000245, 4'd6, 27'h00000098, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000005c, 4'd5, 27'h0000005e, 4'd10, 27'h0000038d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000229, 4'd10, 27'h00000298, 4'd0, 27'h0000020e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000089, 4'd14, 27'h0000013b, 4'd8, 27'h0000006a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002f3, 4'd12, 27'h000000d1, 4'd10, 27'h0000026c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002ad, 4'd1, 27'h00000093, 4'd4, 27'h000000d1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000006, 4'd2, 27'h00000106, 4'd5, 27'h00000362, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000032f, 4'd2, 27'h00000216, 4'd11, 27'h00000201, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000027, 4'd9, 27'h000003d7, 4'd2, 27'h00000237, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003ea, 4'd5, 27'h000001ea, 4'd9, 27'h00000038, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000007, 4'd9, 27'h0000020f, 4'd14, 27'h00000321, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002f7, 4'd10, 27'h00000319, 4'd0, 27'h0000008a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000027, 4'd13, 27'h00000254, 4'd7, 27'h0000033b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000063, 4'd11, 27'h0000000c, 4'd13, 27'h000000e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000011, 4'd4, 27'h0000036c, 4'd2, 27'h0000025e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000ab, 4'd4, 27'h0000027d, 4'd7, 27'h000000bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000148, 4'd1, 27'h000003e9, 4'd14, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000358, 4'd5, 27'h000002dd, 4'd0, 27'h0000038b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000003a, 4'd5, 27'h000003e8, 4'd8, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000014, 4'd5, 27'h00000373, 4'd14, 27'h000000b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000309, 4'd14, 27'h000003a4, 4'd4, 27'h000002f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000017c, 4'd12, 27'h0000005e, 4'd6, 27'h00000382, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000341, 4'd13, 27'h0000002d, 4'd11, 27'h00000349, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000271, 4'd1, 27'h0000030d, 4'd2, 27'h00000270, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000260, 4'd0, 27'h0000037b, 4'd6, 27'h0000032d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000032a, 4'd4, 27'h0000024b, 4'd12, 27'h0000014c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000337, 4'd9, 27'h00000326, 4'd3, 27'h000002f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001fd, 4'd8, 27'h00000173, 4'd5, 27'h000000ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001ee, 4'd5, 27'h000000e5, 4'd12, 27'h00000158, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000087, 4'd14, 27'h00000204, 4'd4, 27'h0000027a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000033, 4'd11, 27'h00000341, 4'd9, 27'h00000268, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000007a, 4'd12, 27'h000002fe, 4'd14, 27'h000001c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000359, 4'd3, 27'h0000039a, 4'd0, 27'h00000343, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000235, 4'd2, 27'h00000372, 4'd8, 27'h00000327, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000286, 4'd1, 27'h000001b2, 4'd13, 27'h00000399, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000143, 4'd5, 27'h00000339, 4'd3, 27'h000002fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000254, 4'd8, 27'h00000179, 4'd6, 27'h00000219, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000006f, 4'd6, 27'h00000178, 4'd13, 27'h00000104, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000020a, 4'd14, 27'h00000206, 4'd3, 27'h00000118, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001f2, 4'd10, 27'h000000b5, 4'd7, 27'h000002b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001e8, 4'd12, 27'h0000035e, 4'd10, 27'h00000057, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000297, 4'd2, 27'h00000038, 4'd2, 27'h00000128, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000034, 4'd3, 27'h000002a5, 4'd6, 27'h000002e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000303, 4'd2, 27'h0000025e, 4'd13, 27'h00000046, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000b5, 4'd7, 27'h00000057, 4'd0, 27'h000001c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000054, 4'd9, 27'h000003e0, 4'd9, 27'h0000030f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000294, 4'd7, 27'h00000357, 4'd14, 27'h0000028c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000396, 4'd12, 27'h00000043, 4'd0, 27'h00000263, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000159, 4'd14, 27'h00000225, 4'd8, 27'h00000162, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000120, 4'd12, 27'h000000ef, 4'd11, 27'h00000395, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000088, 4'd3, 27'h00000270, 4'd0, 27'h000002b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000245, 4'd3, 27'h0000018d, 4'd8, 27'h00000188, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000292, 4'd4, 27'h0000000b, 4'd12, 27'h000001bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000000c, 4'd8, 27'h0000017f, 4'd4, 27'h000001c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002cf, 4'd7, 27'h0000028c, 4'd8, 27'h000000b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001b9, 4'd5, 27'h00000018, 4'd12, 27'h00000084, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000017, 4'd14, 27'h0000011b, 4'd1, 27'h000001f5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002d7, 4'd13, 27'h0000012e, 4'd7, 27'h00000039, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000fa, 4'd11, 27'h00000369, 4'd12, 27'h00000066, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000340, 4'd0, 27'h000000ef, 4'd4, 27'h00000259, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000016d, 4'd1, 27'h000002d3, 4'd7, 27'h00000270, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000215, 4'd2, 27'h000000f7, 4'd13, 27'h0000012b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001ec, 4'd9, 27'h00000316, 4'd2, 27'h0000026d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001e5, 4'd6, 27'h000000e4, 4'd9, 27'h000003e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000023c, 4'd6, 27'h000003d6, 4'd12, 27'h000003ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000030f, 4'd12, 27'h00000349, 4'd0, 27'h00000360, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000031d, 4'd14, 27'h000002fb, 4'd9, 27'h000001d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001fa, 4'd12, 27'h0000006c, 4'd11, 27'h000001c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002f6, 4'd4, 27'h00000374, 4'd2, 27'h0000034c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000012f, 4'd1, 27'h000003e0, 4'd6, 27'h000003e3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003a5, 4'd2, 27'h0000004a, 4'd13, 27'h0000020d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000003a, 4'd8, 27'h00000066, 4'd2, 27'h0000013e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e2, 4'd5, 27'h000001bb, 4'd6, 27'h000000bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000099, 4'd7, 27'h000001f8, 4'd11, 27'h0000000f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000293, 4'd12, 27'h000000ea, 4'd2, 27'h00000111, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000034d, 4'd14, 27'h000000a8, 4'd7, 27'h0000037c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001ff, 4'd14, 27'h000000d1, 4'd14, 27'h0000013c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001cb, 4'd0, 27'h0000025f, 4'd4, 27'h00000009, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000c2, 4'd2, 27'h0000007b, 4'd9, 27'h0000020d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000096, 4'd4, 27'h000002c8, 4'd14, 27'h000001ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000004, 4'd9, 27'h00000310, 4'd3, 27'h000003bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000076, 4'd5, 27'h0000039a, 4'd9, 27'h00000184, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001fd, 4'd6, 27'h0000019e, 4'd14, 27'h0000009e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000090, 4'd12, 27'h000003bf, 4'd2, 27'h0000008c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000031c, 4'd13, 27'h00000211, 4'd8, 27'h000000b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000331, 4'd14, 27'h00000279, 4'd13, 27'h00000278, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000018d, 4'd2, 27'h00000249, 4'd2, 27'h00000093, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003e3, 4'd4, 27'h000000d1, 4'd6, 27'h00000102, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b1, 4'd1, 27'h00000063, 4'd10, 27'h00000345, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000141, 4'd6, 27'h0000000c, 4'd4, 27'h00000036, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000020f, 4'd7, 27'h00000355, 4'd7, 27'h000003e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002fe, 4'd5, 27'h00000236, 4'd12, 27'h000002c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000016c, 4'd12, 27'h0000029c, 4'd3, 27'h00000004, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000013c, 4'd13, 27'h00000135, 4'd5, 27'h000002e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000009, 4'd12, 27'h00000322, 4'd12, 27'h00000170, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000005b, 4'd2, 27'h00000013, 4'd2, 27'h0000000b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001de, 4'd0, 27'h000003fe, 4'd7, 27'h000000d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003d6, 4'd2, 27'h000002d4, 4'd14, 27'h0000022a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002e2, 4'd9, 27'h000003bd, 4'd3, 27'h00000041, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001ac, 4'd8, 27'h0000020e, 4'd9, 27'h00000180, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000186, 4'd9, 27'h0000016f, 4'd11, 27'h00000301, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000157, 4'd11, 27'h00000064, 4'd3, 27'h000001ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001fa, 4'd12, 27'h0000010b, 4'd9, 27'h0000030c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000021e, 4'd12, 27'h000002c5, 4'd11, 27'h000001f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000006c, 4'd1, 27'h00000104, 4'd3, 27'h00000155, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002b1, 4'd4, 27'h000000ec, 4'd8, 27'h00000086, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000222, 4'd4, 27'h000000eb, 4'd13, 27'h000003cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000031e, 4'd9, 27'h000000ae, 4'd2, 27'h0000033b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000013c, 4'd7, 27'h00000023, 4'd8, 27'h0000030f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003af, 4'd7, 27'h00000268, 4'd10, 27'h00000300, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000045, 4'd10, 27'h000000ed, 4'd3, 27'h0000029f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000d8, 4'd10, 27'h000002f4, 4'd9, 27'h00000157, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000185, 4'd13, 27'h00000249, 4'd12, 27'h00000379, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000382, 4'd0, 27'h000001aa, 4'd3, 27'h00000227, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000152, 4'd4, 27'h000001ba, 4'd9, 27'h000001ea, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000038b, 4'd4, 27'h0000022a, 4'd10, 27'h0000032e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000354, 4'd8, 27'h000000fe, 4'd4, 27'h00000396, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000307, 4'd6, 27'h000000fc, 4'd8, 27'h00000073, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000c7, 4'd9, 27'h00000010, 4'd10, 27'h00000083, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000282, 4'd10, 27'h0000036b, 4'd3, 27'h00000050, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001e4, 4'd10, 27'h000003b2, 4'd9, 27'h00000179, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000364, 4'd12, 27'h0000021c, 4'd10, 27'h00000079, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000200, 4'd0, 27'h0000006a, 4'd3, 27'h000001c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000326, 4'd0, 27'h00000192, 4'd9, 27'h00000348, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000344, 4'd2, 27'h000001c7, 4'd10, 27'h000003f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000010d, 4'd9, 27'h000003ea, 4'd2, 27'h0000018b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000202, 4'd9, 27'h000001e6, 4'd6, 27'h0000019c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000059, 4'd7, 27'h00000171, 4'd13, 27'h00000171, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000286, 4'd13, 27'h000001f9, 4'd3, 27'h000001e5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000e0, 4'd12, 27'h000000bc, 4'd8, 27'h000003df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000006d, 4'd12, 27'h00000110, 4'd11, 27'h0000022c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001e7, 4'd2, 27'h000002f2, 4'd1, 27'h0000007c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000257, 4'd2, 27'h000003eb, 4'd7, 27'h000000c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001c0, 4'd1, 27'h000002b2, 4'd10, 27'h00000218, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000125, 4'd7, 27'h0000002f, 4'd1, 27'h00000241, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001b0, 4'd9, 27'h00000393, 4'd6, 27'h0000028d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000113, 4'd6, 27'h000001f3, 4'd14, 27'h000001e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000031e, 4'd11, 27'h000001ee, 4'd2, 27'h00000020, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000034d, 4'd13, 27'h00000111, 4'd5, 27'h000002ff, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000368, 4'd12, 27'h0000030b, 4'd13, 27'h000001e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b3, 4'd4, 27'h0000017d, 4'd2, 27'h00000327, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000f6, 4'd0, 27'h00000149, 4'd8, 27'h0000016c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000144, 4'd3, 27'h000002e0, 4'd11, 27'h00000302, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001fb, 4'd6, 27'h00000291, 4'd2, 27'h00000204, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000254, 4'd6, 27'h00000057, 4'd5, 27'h00000257, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000311, 4'd5, 27'h000003ad, 4'd14, 27'h0000010c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003fb, 4'd13, 27'h000003e8, 4'd4, 27'h000000ca, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000134, 4'd11, 27'h0000030b, 4'd5, 27'h00000028, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000012a, 4'd11, 27'h00000112, 4'd13, 27'h0000001c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ac, 4'd2, 27'h0000002c, 4'd0, 27'h000001bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000292, 4'd3, 27'h000001a3, 4'd7, 27'h000003d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000136, 4'd1, 27'h00000189, 4'd13, 27'h000003ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000315, 4'd8, 27'h000000d3, 4'd3, 27'h000000db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000263, 4'd5, 27'h00000147, 4'd7, 27'h000003f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000018f, 4'd5, 27'h00000002, 4'd11, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001e1, 4'd14, 27'h0000026e, 4'd4, 27'h00000177, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000038f, 4'd10, 27'h00000291, 4'd9, 27'h00000247, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000020f, 4'd13, 27'h000002e8, 4'd11, 27'h000001a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000018, 4'd1, 27'h00000213, 4'd2, 27'h000002f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000018f, 4'd4, 27'h000002e6, 4'd8, 27'h0000007f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001ff, 4'd2, 27'h00000307, 4'd14, 27'h0000022b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000101, 4'd7, 27'h00000029, 4'd0, 27'h00000260, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000d9, 4'd9, 27'h00000207, 4'd7, 27'h000003e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000333, 4'd7, 27'h000003f2, 4'd11, 27'h000002f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001c9, 4'd10, 27'h00000008, 4'd1, 27'h000001b5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000018b, 4'd10, 27'h00000116, 4'd8, 27'h000001c0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000000a, 4'd10, 27'h00000128, 4'd12, 27'h000001b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000028b, 4'd2, 27'h000002e5, 4'd1, 27'h00000009, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000108, 4'd1, 27'h0000037e, 4'd5, 27'h00000196, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000005f, 4'd4, 27'h0000014b, 4'd11, 27'h0000015d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000305, 4'd9, 27'h0000028c, 4'd0, 27'h000000b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003fd, 4'd6, 27'h0000036a, 4'd6, 27'h000002a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000cb, 4'd9, 27'h00000087, 4'd12, 27'h00000090, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000005c, 4'd14, 27'h0000031c, 4'd0, 27'h000001a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000091, 4'd11, 27'h000001f6, 4'd5, 27'h00000082, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000150, 4'd11, 27'h0000013b, 4'd12, 27'h000001ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000108, 4'd4, 27'h0000036d, 4'd2, 27'h00000016, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002d4, 4'd2, 27'h00000018, 4'd5, 27'h000001b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c3, 4'd1, 27'h00000301, 4'd10, 27'h000003f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000384, 4'd6, 27'h000003c4, 4'd4, 27'h000001c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000071, 4'd8, 27'h00000296, 4'd9, 27'h00000052, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001e6, 4'd5, 27'h000003f1, 4'd11, 27'h000002a7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000026c, 4'd10, 27'h000002dc, 4'd2, 27'h000001f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a9, 4'd11, 27'h000002af, 4'd8, 27'h00000330, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000191, 4'd11, 27'h0000006e, 4'd12, 27'h000002a4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000138, 4'd1, 27'h0000009d, 4'd2, 27'h00000300, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000312, 4'd3, 27'h00000394, 4'd7, 27'h00000389, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000067, 4'd4, 27'h00000201, 4'd13, 27'h00000334, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000212, 4'd5, 27'h000002a1, 4'd0, 27'h000000c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000022c, 4'd9, 27'h00000313, 4'd6, 27'h000002e0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000016a, 4'd5, 27'h000000c3, 4'd14, 27'h00000116, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000b6, 4'd13, 27'h00000042, 4'd3, 27'h0000011d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000277, 4'd14, 27'h0000003f, 4'd9, 27'h00000007, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000069, 4'd10, 27'h000001a8, 4'd14, 27'h00000106, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000240, 4'd0, 27'h0000034c, 4'd1, 27'h00000019, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000020b, 4'd3, 27'h0000004d, 4'd8, 27'h0000003d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000228, 4'd2, 27'h000000a6, 4'd10, 27'h0000037f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000007c, 4'd9, 27'h000000a8, 4'd0, 27'h00000075, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000153, 4'd8, 27'h00000243, 4'd7, 27'h00000397, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000032c, 4'd8, 27'h000002f8, 4'd12, 27'h000002de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000e7, 4'd13, 27'h000002f6, 4'd3, 27'h000003d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000360, 4'd13, 27'h00000323, 4'd5, 27'h00000069, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000262, 4'd11, 27'h00000399, 4'd13, 27'h0000021b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000265, 4'd0, 27'h0000000f, 4'd3, 27'h000000f4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003b9, 4'd2, 27'h0000024a, 4'd5, 27'h000001dd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003ba, 4'd1, 27'h00000119, 4'd11, 27'h0000020b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000150, 4'd7, 27'h000003df, 4'd1, 27'h00000127, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003ba, 4'd6, 27'h000000f9, 4'd6, 27'h000001d4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002dd, 4'd9, 27'h000003fd, 4'd13, 27'h00000102, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c8, 4'd11, 27'h000000c3, 4'd4, 27'h000003a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000004, 4'd13, 27'h00000323, 4'd9, 27'h0000008b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000283, 4'd13, 27'h000001b2, 4'd11, 27'h00000124, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000268, 4'd1, 27'h00000263, 4'd0, 27'h00000071, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002be, 4'd1, 27'h000001e1, 4'd9, 27'h000001d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000019d, 4'd4, 27'h000001a3, 4'd12, 27'h00000297, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000221, 4'd7, 27'h0000028b, 4'd1, 27'h0000030d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000182, 4'd8, 27'h000001c7, 4'd9, 27'h0000037a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000227, 4'd5, 27'h000003be, 4'd12, 27'h000002cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000166, 4'd11, 27'h00000027, 4'd1, 27'h00000365, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000324, 4'd10, 27'h00000044, 4'd5, 27'h00000049, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000387, 4'd14, 27'h0000029c, 4'd10, 27'h000000c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001a6, 4'd0, 27'h00000315, 4'd1, 27'h000003d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000153, 4'd4, 27'h00000386, 4'd5, 27'h000003fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000308, 4'd4, 27'h0000020f, 4'd12, 27'h0000019d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000122, 4'd7, 27'h00000106, 4'd1, 27'h0000022a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000208, 4'd8, 27'h000001c2, 4'd5, 27'h00000316, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000010e, 4'd7, 27'h00000146, 4'd10, 27'h000002b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001f1, 4'd12, 27'h0000014f, 4'd4, 27'h00000238, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001fc, 4'd12, 27'h0000028a, 4'd8, 27'h0000028b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001a8, 4'd14, 27'h0000024c, 4'd13, 27'h000003fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000261, 4'd3, 27'h00000216, 4'd3, 27'h000003d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000192, 4'd2, 27'h000001ec, 4'd9, 27'h00000126, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000123, 4'd3, 27'h00000367, 4'd13, 27'h0000030c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001f0, 4'd9, 27'h00000183, 4'd2, 27'h0000016d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000259, 4'd5, 27'h00000079, 4'd6, 27'h000002ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002f5, 4'd8, 27'h00000279, 4'd11, 27'h000001eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003fb, 4'd11, 27'h000000c9, 4'd0, 27'h0000006a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001f2, 4'd13, 27'h0000038b, 4'd7, 27'h000003f4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000d0, 4'd14, 27'h00000058, 4'd12, 27'h000003a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003bb, 4'd2, 27'h0000017e, 4'd1, 27'h000003ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000006, 4'd3, 27'h00000394, 4'd6, 27'h000001f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002c1, 4'd3, 27'h0000038a, 4'd12, 27'h0000019f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001d0, 4'd8, 27'h00000266, 4'd2, 27'h000002d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003a6, 4'd9, 27'h00000277, 4'd9, 27'h00000040, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002e0, 4'd9, 27'h00000196, 4'd14, 27'h000002f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001c7, 4'd10, 27'h00000025, 4'd4, 27'h00000373, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000d7, 4'd13, 27'h000000da, 4'd7, 27'h000000db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000ae, 4'd13, 27'h00000290, 4'd12, 27'h000002c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000062, 4'd0, 27'h0000037d, 4'd2, 27'h00000167, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002fa, 4'd0, 27'h00000268, 4'd5, 27'h00000315, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000062, 4'd3, 27'h000002e7, 4'd14, 27'h00000303, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000010, 4'd6, 27'h0000015a, 4'd0, 27'h000002cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003e5, 4'd5, 27'h000003b5, 4'd8, 27'h000000dc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000066, 4'd7, 27'h000000f0, 4'd14, 27'h0000005b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000024a, 4'd14, 27'h00000090, 4'd4, 27'h00000065, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000260, 4'd10, 27'h0000014e, 4'd9, 27'h000001f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003e3, 4'd12, 27'h00000334, 4'd12, 27'h00000084, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000d6, 4'd0, 27'h0000003b, 4'd3, 27'h000000da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003ce, 4'd2, 27'h000001c2, 4'd5, 27'h00000317, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001ca, 4'd2, 27'h000003b2, 4'd12, 27'h00000209, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000225, 4'd6, 27'h000000a9, 4'd0, 27'h000003ff, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000039f, 4'd7, 27'h000000c7, 4'd8, 27'h0000000a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000019c, 4'd9, 27'h000003ea, 4'd12, 27'h00000282, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000238, 4'd13, 27'h00000132, 4'd1, 27'h0000032e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000a0, 4'd11, 27'h00000304, 4'd7, 27'h000001f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e3, 4'd12, 27'h000001a0, 4'd11, 27'h00000122, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000201, 4'd1, 27'h00000038, 4'd3, 27'h0000026a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000115, 4'd1, 27'h0000001d, 4'd8, 27'h000003be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003da, 4'd3, 27'h0000009a, 4'd13, 27'h00000134, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000379, 4'd5, 27'h000001a9, 4'd3, 27'h00000190, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000176, 4'd6, 27'h0000021c, 4'd8, 27'h00000011, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000072, 4'd7, 27'h000003d4, 4'd14, 27'h00000182, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002e5, 4'd12, 27'h00000281, 4'd0, 27'h000002b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000338, 4'd10, 27'h000000b6, 4'd9, 27'h00000301, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001cc, 4'd14, 27'h00000094, 4'd13, 27'h0000005b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000251, 4'd4, 27'h000000f9, 4'd0, 27'h00000037, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000208, 4'd3, 27'h00000188, 4'd7, 27'h0000033b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000179, 4'd0, 27'h0000026e, 4'd10, 27'h000003e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000364, 4'd6, 27'h000003d3, 4'd1, 27'h000001d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000031c, 4'd9, 27'h00000305, 4'd7, 27'h0000036c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002e0, 4'd7, 27'h00000268, 4'd10, 27'h0000022a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000012b, 4'd11, 27'h0000028a, 4'd4, 27'h000001fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000192, 4'd14, 27'h00000299, 4'd8, 27'h00000237, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000019e, 4'd12, 27'h00000397, 4'd10, 27'h000003c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000375, 4'd2, 27'h0000038e, 4'd2, 27'h00000122, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000383, 4'd3, 27'h00000111, 4'd6, 27'h000000cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000038e, 4'd1, 27'h00000241, 4'd11, 27'h0000000d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003a4, 4'd6, 27'h000000b4, 4'd4, 27'h000003da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000242, 4'd6, 27'h000001f7, 4'd7, 27'h00000206, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000153, 4'd6, 27'h000001a0, 4'd14, 27'h0000037a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000215, 4'd11, 27'h000002cc, 4'd4, 27'h00000121, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000224, 4'd13, 27'h000000b2, 4'd9, 27'h0000034c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000236, 4'd12, 27'h00000299, 4'd11, 27'h00000165, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000138, 4'd2, 27'h00000359, 4'd1, 27'h000003da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000117, 4'd3, 27'h000003a2, 4'd8, 27'h000002ff, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000020b, 4'd0, 27'h00000357, 4'd10, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002bd, 4'd7, 27'h00000312, 4'd4, 27'h000000bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002a3, 4'd5, 27'h0000031d, 4'd7, 27'h000002a3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000345, 4'd9, 27'h00000013, 4'd13, 27'h00000058, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003be, 4'd10, 27'h000001cc, 4'd2, 27'h000000fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000c4, 4'd11, 27'h00000051, 4'd7, 27'h000001ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000339, 4'd12, 27'h00000229, 4'd11, 27'h00000136, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000009f, 4'd0, 27'h000003ed, 4'd2, 27'h000002ee, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000075, 4'd2, 27'h0000000b, 4'd8, 27'h00000045, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000026c, 4'd0, 27'h00000005, 4'd14, 27'h0000004a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000200, 4'd8, 27'h000001ae, 4'd4, 27'h0000016f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000a6, 4'd5, 27'h000003e8, 4'd7, 27'h00000178, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002d5, 4'd6, 27'h0000032e, 4'd12, 27'h0000017b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002d6, 4'd12, 27'h00000038, 4'd2, 27'h000002cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000018, 4'd10, 27'h000002e1, 4'd9, 27'h00000064, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000320, 4'd14, 27'h00000270, 4'd13, 27'h000002d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000020f, 4'd4, 27'h000000c1, 4'd1, 27'h0000029b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000036c, 4'd0, 27'h000001aa, 4'd7, 27'h000002aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003dd, 4'd1, 27'h00000158, 4'd14, 27'h00000194, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003d7, 4'd9, 27'h00000347, 4'd1, 27'h000003a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000021b, 4'd7, 27'h00000199, 4'd5, 27'h00000090, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000b2, 4'd9, 27'h00000045, 4'd14, 27'h000003a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003e4, 4'd13, 27'h000000cd, 4'd0, 27'h00000147, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002b8, 4'd14, 27'h0000011c, 4'd6, 27'h00000063, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001f0, 4'd10, 27'h000003be, 4'd11, 27'h000002d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000174, 4'd2, 27'h000003a0, 4'd3, 27'h000002bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000027a, 4'd1, 27'h0000003e, 4'd6, 27'h00000322, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000373, 4'd2, 27'h00000375, 4'd12, 27'h000002fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000139, 4'd8, 27'h000002d5, 4'd1, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000009c, 4'd6, 27'h0000032e, 4'd9, 27'h00000121, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003ec, 4'd9, 27'h000001b2, 4'd14, 27'h000001ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000161, 4'd13, 27'h00000220, 4'd2, 27'h00000021, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000d8, 4'd10, 27'h00000154, 4'd8, 27'h000000b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000048, 4'd13, 27'h000003d1, 4'd11, 27'h000003ef, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002db, 4'd3, 27'h0000030d, 4'd1, 27'h00000152, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002fb, 4'd4, 27'h00000255, 4'd7, 27'h000000a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000102, 4'd1, 27'h00000130, 4'd10, 27'h0000021c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000020a, 4'd9, 27'h0000037d, 4'd2, 27'h000000eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000212, 4'd6, 27'h000003c2, 4'd5, 27'h00000098, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000290, 4'd7, 27'h000000f3, 4'd13, 27'h000001bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000084, 4'd12, 27'h00000029, 4'd2, 27'h00000187, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003a6, 4'd12, 27'h000003a9, 4'd6, 27'h0000038a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000300, 4'd12, 27'h00000288, 4'd11, 27'h000000ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003fc, 4'd1, 27'h000000b9, 4'd3, 27'h000000f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000286, 4'd0, 27'h00000342, 4'd5, 27'h00000111, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000098, 4'd1, 27'h000002bf, 4'd14, 27'h00000249, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001c7, 4'd9, 27'h00000211, 4'd2, 27'h000002bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000b8, 4'd6, 27'h00000340, 4'd6, 27'h0000028d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000020a, 4'd7, 27'h0000018a, 4'd13, 27'h0000035b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000255, 4'd11, 27'h000001c7, 4'd4, 27'h0000002b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001e6, 4'd14, 27'h00000118, 4'd6, 27'h000003fb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003f1, 4'd13, 27'h000001c7, 4'd14, 27'h00000301, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000f9, 4'd0, 27'h000000bf, 4'd1, 27'h000002e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003b4, 4'd3, 27'h00000230, 4'd6, 27'h000000ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001e7, 4'd0, 27'h0000034e, 4'd13, 27'h00000145, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000012f, 4'd8, 27'h000002ee, 4'd1, 27'h00000114, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000200, 4'd5, 27'h000002e4, 4'd9, 27'h0000032d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000252, 4'd9, 27'h00000285, 4'd13, 27'h0000032c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000003f, 4'd12, 27'h00000269, 4'd4, 27'h0000007a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000346, 4'd13, 27'h00000064, 4'd7, 27'h000003e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000e1, 4'd10, 27'h00000396, 4'd14, 27'h00000276, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003c9, 4'd0, 27'h0000008c, 4'd0, 27'h000001bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000c4, 4'd3, 27'h000000e8, 4'd7, 27'h000002af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000145, 4'd1, 27'h0000009a, 4'd12, 27'h000000d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000024e, 4'd6, 27'h000001f1, 4'd2, 27'h000001a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003e5, 4'd5, 27'h000002a6, 4'd9, 27'h0000002c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001a7, 4'd6, 27'h000003f3, 4'd13, 27'h0000019c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000308, 4'd12, 27'h00000101, 4'd4, 27'h00000141, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000029b, 4'd12, 27'h000000ae, 4'd8, 27'h000001ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000c7, 4'd14, 27'h000001a8, 4'd10, 27'h000001b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000209, 4'd1, 27'h000000a5, 4'd4, 27'h00000131, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000362, 4'd4, 27'h00000030, 4'd7, 27'h00000161, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003ef, 4'd2, 27'h00000077, 4'd12, 27'h0000024b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000031, 4'd9, 27'h0000026a, 4'd0, 27'h00000024, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001f1, 4'd5, 27'h00000319, 4'd9, 27'h00000250, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002b2, 4'd5, 27'h00000309, 4'd11, 27'h000002a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000023b, 4'd10, 27'h000003e0, 4'd1, 27'h0000015e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000347, 4'd11, 27'h000001d8, 4'd9, 27'h000002fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000030a, 4'd13, 27'h00000348, 4'd10, 27'h000002fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000012b, 4'd0, 27'h000003aa, 4'd4, 27'h0000026c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001d9, 4'd2, 27'h00000124, 4'd7, 27'h000001bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000186, 4'd4, 27'h000000fb, 4'd11, 27'h0000021a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000016, 4'd7, 27'h000003de, 4'd4, 27'h000001f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000155, 4'd5, 27'h0000018f, 4'd5, 27'h000003a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000032e, 4'd6, 27'h00000293, 4'd11, 27'h000000a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000fb, 4'd14, 27'h00000106, 4'd1, 27'h000000f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000185, 4'd12, 27'h000003cf, 4'd5, 27'h0000028c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000012c, 4'd13, 27'h00000364, 4'd10, 27'h000000d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000308, 4'd2, 27'h00000015, 4'd4, 27'h00000384, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000022f, 4'd2, 27'h0000011c, 4'd8, 27'h000003ea, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000357, 4'd2, 27'h000002d5, 4'd10, 27'h00000253, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000043, 4'd6, 27'h00000187, 4'd0, 27'h000003d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001d6, 4'd5, 27'h00000202, 4'd8, 27'h0000000c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001eb, 4'd5, 27'h000002bb, 4'd10, 27'h000000d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000cd, 4'd11, 27'h00000170, 4'd3, 27'h0000007f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003e7, 4'd12, 27'h00000107, 4'd5, 27'h00000087, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000104, 4'd10, 27'h000000d0, 4'd12, 27'h0000025a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000223, 4'd0, 27'h000001c1, 4'd3, 27'h0000025a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000004c, 4'd0, 27'h000002df, 4'd6, 27'h00000362, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000374, 4'd4, 27'h00000338, 4'd13, 27'h0000035d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000023a, 4'd6, 27'h0000021e, 4'd4, 27'h0000010f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000de, 4'd7, 27'h000002d0, 4'd9, 27'h000002ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000221, 4'd9, 27'h00000027, 4'd13, 27'h00000323, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000011a, 4'd12, 27'h000001d5, 4'd4, 27'h00000112, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000a9, 4'd10, 27'h00000294, 4'd6, 27'h000002df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001b4, 4'd10, 27'h00000091, 4'd13, 27'h000001cf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000126, 4'd0, 27'h000002e4, 4'd4, 27'h00000108, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000150, 4'd0, 27'h00000193, 4'd8, 27'h000003f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000c8, 4'd3, 27'h00000390, 4'd12, 27'h000001f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003c6, 4'd5, 27'h000002a7, 4'd1, 27'h00000239, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000093, 4'd6, 27'h00000197, 4'd8, 27'h00000212, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000317, 4'd5, 27'h0000031b, 4'd11, 27'h0000009f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000003b, 4'd13, 27'h000000d9, 4'd1, 27'h00000190, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000039f, 4'd11, 27'h00000247, 4'd7, 27'h000001d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000342, 4'd10, 27'h00000152, 4'd10, 27'h000002a0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000274, 4'd3, 27'h000002b1, 4'd3, 27'h0000021b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003cd, 4'd1, 27'h0000007c, 4'd6, 27'h00000332, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003c4, 4'd1, 27'h000002ae, 4'd14, 27'h000002b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002b4, 4'd7, 27'h00000054, 4'd0, 27'h00000235, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002f7, 4'd9, 27'h00000018, 4'd8, 27'h000003f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000190, 4'd6, 27'h0000035a, 4'd14, 27'h0000038e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000236, 4'd14, 27'h000002e0, 4'd0, 27'h00000014, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000036d, 4'd12, 27'h000002f4, 4'd6, 27'h00000321, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002fb, 4'd10, 27'h0000036a, 4'd13, 27'h00000247, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000d9, 4'd2, 27'h00000202, 4'd1, 27'h00000023, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003bb, 4'd0, 27'h0000033b, 4'd7, 27'h00000332, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000017a, 4'd0, 27'h0000007f, 4'd13, 27'h0000039d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000093, 4'd5, 27'h000001de, 4'd1, 27'h00000385, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000379, 4'd5, 27'h000002fb, 4'd9, 27'h00000119, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001ba, 4'd7, 27'h00000062, 4'd11, 27'h00000354, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000258, 4'd11, 27'h00000301, 4'd4, 27'h000002fb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000028c, 4'd12, 27'h000003ae, 4'd8, 27'h0000008e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000ce, 4'd10, 27'h000000f3, 4'd13, 27'h000002ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003ca, 4'd0, 27'h000003d9, 4'd3, 27'h000002b5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000238, 4'd3, 27'h0000037c, 4'd7, 27'h00000186, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000202, 4'd1, 27'h00000391, 4'd12, 27'h0000016e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000014d, 4'd7, 27'h00000193, 4'd4, 27'h00000337, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000c1, 4'd5, 27'h00000296, 4'd8, 27'h00000203, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000142, 4'd6, 27'h000003a4, 4'd14, 27'h00000109, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000028, 4'd10, 27'h0000005c, 4'd2, 27'h00000002, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000211, 4'd13, 27'h000002bb, 4'd8, 27'h00000372, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000101, 4'd14, 27'h0000033f, 4'd14, 27'h000003e8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002d8, 4'd3, 27'h000002da, 4'd2, 27'h00000125, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000398, 4'd4, 27'h00000317, 4'd5, 27'h000000d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001df, 4'd4, 27'h00000159, 4'd11, 27'h0000032f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000204, 4'd5, 27'h00000313, 4'd1, 27'h000001c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003a2, 4'd8, 27'h000000ec, 4'd5, 27'h00000080, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001e3, 4'd8, 27'h000001db, 4'd13, 27'h0000035d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001ea, 4'd11, 27'h00000183, 4'd1, 27'h000003f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003d7, 4'd13, 27'h000002ca, 4'd9, 27'h0000019f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000055, 4'd13, 27'h0000012e, 4'd11, 27'h0000016d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000370, 4'd0, 27'h000003e8, 4'd0, 27'h0000015c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001dc, 4'd1, 27'h00000011, 4'd7, 27'h000001ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002f3, 4'd0, 27'h0000004d, 4'd10, 27'h00000254, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001bc, 4'd5, 27'h00000281, 4'd1, 27'h000002ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000254, 4'd5, 27'h000002f3, 4'd7, 27'h00000298, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002fa, 4'd9, 27'h000000d2, 4'd10, 27'h00000373, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000d1, 4'd14, 27'h00000152, 4'd0, 27'h000001b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000028b, 4'd14, 27'h00000079, 4'd9, 27'h000003a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000237, 4'd10, 27'h000002a1, 4'd12, 27'h000000aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000006e, 4'd2, 27'h000000f8, 4'd0, 27'h00000004, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000012d, 4'd4, 27'h00000017, 4'd5, 27'h000002ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002b9, 4'd2, 27'h00000231, 4'd12, 27'h000003d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000022b, 4'd5, 27'h00000043, 4'd1, 27'h00000107, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003ee, 4'd8, 27'h0000001b, 4'd7, 27'h000001a2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000213, 4'd6, 27'h00000043, 4'd13, 27'h00000107, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000131, 4'd13, 27'h000000f2, 4'd3, 27'h00000126, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000379, 4'd13, 27'h00000291, 4'd7, 27'h00000212, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000b7, 4'd12, 27'h0000027a, 4'd14, 27'h0000023e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000027f, 4'd4, 27'h000002d4, 4'd0, 27'h000002ed, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002d2, 4'd2, 27'h00000089, 4'd8, 27'h0000012d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000022f, 4'd3, 27'h000003ba, 4'd14, 27'h00000036, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000360, 4'd9, 27'h00000160, 4'd3, 27'h0000027a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000006e, 4'd9, 27'h0000002b, 4'd9, 27'h000003b4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001b9, 4'd8, 27'h00000248, 4'd10, 27'h000001f4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000127, 4'd10, 27'h000001fb, 4'd1, 27'h000003ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000ca, 4'd13, 27'h0000035c, 4'd5, 27'h00000272, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000369, 4'd10, 27'h0000010f, 4'd13, 27'h000001b5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000011a, 4'd0, 27'h000002bd, 4'd2, 27'h00000311, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000032a, 4'd4, 27'h00000325, 4'd5, 27'h000002c7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000376, 4'd3, 27'h000000e0, 4'd12, 27'h000001bc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000267, 4'd9, 27'h000003f3, 4'd3, 27'h00000083, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000043, 4'd7, 27'h00000089, 4'd5, 27'h00000160, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003e8, 4'd7, 27'h000001ce, 4'd11, 27'h0000012c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000105, 4'd12, 27'h0000018a, 4'd4, 27'h00000245, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000041, 4'd10, 27'h000003c0, 4'd7, 27'h000000db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c5, 4'd13, 27'h000000bb, 4'd12, 27'h000002b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000322, 4'd3, 27'h000001e0, 4'd2, 27'h000001fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000038f, 4'd2, 27'h000001f6, 4'd7, 27'h000001ba, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000181, 4'd4, 27'h000001e4, 4'd14, 27'h00000127, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000016, 4'd5, 27'h000003ef, 4'd3, 27'h00000218, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001eb, 4'd8, 27'h000000e9, 4'd7, 27'h000002d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000099, 4'd8, 27'h00000281, 4'd13, 27'h0000038d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000307, 4'd10, 27'h0000015e, 4'd2, 27'h00000398, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000117, 4'd13, 27'h0000022f, 4'd7, 27'h00000309, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000302, 4'd14, 27'h000002ca, 4'd14, 27'h00000309, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000309, 4'd1, 27'h000003c7, 4'd0, 27'h000003b9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000038c, 4'd3, 27'h000003f9, 4'd6, 27'h000002c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002db, 4'd3, 27'h000003bf, 4'd12, 27'h0000025c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002d7, 4'd9, 27'h000002bd, 4'd3, 27'h000000d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001eb, 4'd8, 27'h000003a7, 4'd9, 27'h00000250, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001f8, 4'd7, 27'h00000272, 4'd12, 27'h000001b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000003b, 4'd13, 27'h00000307, 4'd4, 27'h000001e3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002a9, 4'd14, 27'h000003db, 4'd8, 27'h000000ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003f2, 4'd14, 27'h0000001b, 4'd12, 27'h000001bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000a9, 4'd3, 27'h00000100, 4'd1, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000357, 4'd1, 27'h0000011a, 4'd9, 27'h00000005, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003fd, 4'd3, 27'h00000155, 4'd12, 27'h00000061, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000f7, 4'd8, 27'h00000253, 4'd1, 27'h00000337, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000025c, 4'd6, 27'h00000247, 4'd7, 27'h0000016d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000f9, 4'd9, 27'h000003c7, 4'd12, 27'h0000028b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002af, 4'd11, 27'h000003e0, 4'd1, 27'h00000199, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000137, 4'd14, 27'h000001b4, 4'd5, 27'h000000e0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001b3, 4'd13, 27'h00000291, 4'd12, 27'h0000037f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001fb, 4'd2, 27'h000002ef, 4'd3, 27'h000001c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001b2, 4'd2, 27'h000000f2, 4'd6, 27'h00000257, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002d5, 4'd2, 27'h00000335, 4'd12, 27'h00000098, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000125, 4'd7, 27'h00000340, 4'd3, 27'h0000025f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000029a, 4'd8, 27'h000001c6, 4'd8, 27'h0000023c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000292, 4'd7, 27'h00000025, 4'd11, 27'h000003a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000034c, 4'd13, 27'h000000af, 4'd3, 27'h00000397, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000132, 4'd14, 27'h00000349, 4'd9, 27'h000000d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000019d, 4'd11, 27'h000003c4, 4'd11, 27'h00000166, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000231, 4'd0, 27'h0000020b, 4'd3, 27'h000000f7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000023d, 4'd3, 27'h000002dc, 4'd7, 27'h000003ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000027f, 4'd0, 27'h0000016f, 4'd10, 27'h00000328, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000012a, 4'd6, 27'h000003e2, 4'd3, 27'h0000020f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000bf, 4'd5, 27'h000003d7, 4'd7, 27'h00000357, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b9, 4'd6, 27'h0000007c, 4'd12, 27'h000002c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000089, 4'd11, 27'h000000d0, 4'd2, 27'h000003ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000ea, 4'd13, 27'h00000081, 4'd8, 27'h00000226, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000259, 4'd14, 27'h0000017c, 4'd10, 27'h00000284, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000cb, 4'd2, 27'h000002bc, 4'd1, 27'h0000027a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000031d, 4'd4, 27'h000000d0, 4'd6, 27'h00000244, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000202, 4'd3, 27'h00000364, 4'd13, 27'h00000146, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000003e, 4'd6, 27'h00000332, 4'd4, 27'h000003e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000052, 4'd7, 27'h00000084, 4'd8, 27'h000002d6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000383, 4'd7, 27'h0000029b, 4'd14, 27'h000000d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002b6, 4'd14, 27'h00000186, 4'd3, 27'h0000003b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000380, 4'd10, 27'h0000037d, 4'd5, 27'h000001b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000010d, 4'd13, 27'h0000033b, 4'd12, 27'h00000385, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002ee, 4'd3, 27'h000000de, 4'd1, 27'h00000118, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000007a, 4'd1, 27'h00000014, 4'd9, 27'h000002a7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002d0, 4'd2, 27'h000001c0, 4'd14, 27'h00000393, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000020e, 4'd5, 27'h00000184, 4'd0, 27'h000003e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000314, 4'd8, 27'h000000ca, 4'd9, 27'h00000357, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000083, 4'd5, 27'h00000046, 4'd12, 27'h00000309, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000018b, 4'd14, 27'h00000173, 4'd0, 27'h000000f4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000006e, 4'd14, 27'h0000032a, 4'd9, 27'h00000202, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000019e, 4'd14, 27'h000002ab, 4'd13, 27'h000003d9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000000d, 4'd2, 27'h0000012d, 4'd0, 27'h0000002b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002ca, 4'd2, 27'h00000364, 4'd5, 27'h00000273, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002e6, 4'd1, 27'h000002c3, 4'd14, 27'h00000096, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000005c, 4'd8, 27'h000001cb, 4'd1, 27'h0000010e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001e7, 4'd8, 27'h00000256, 4'd6, 27'h00000235, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000023f, 4'd7, 27'h00000025, 4'd13, 27'h000000a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003d2, 4'd14, 27'h0000023a, 4'd2, 27'h000001c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000133, 4'd12, 27'h000003e1, 4'd5, 27'h000002c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000005b, 4'd10, 27'h000002c3, 4'd11, 27'h0000036a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000014c, 4'd3, 27'h0000002a, 4'd2, 27'h000000fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000011e, 4'd2, 27'h00000063, 4'd6, 27'h00000201, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000b5, 4'd1, 27'h0000024f, 4'd13, 27'h00000230, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000330, 4'd8, 27'h0000016d, 4'd0, 27'h000001f1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000085, 4'd9, 27'h00000387, 4'd9, 27'h0000026f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000084, 4'd8, 27'h000003c3, 4'd14, 27'h00000198, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000216, 4'd13, 27'h000001b6, 4'd4, 27'h000002b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000045, 4'd14, 27'h000001db, 4'd9, 27'h000003eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002dd, 4'd12, 27'h00000390, 4'd10, 27'h0000027d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000228, 4'd0, 27'h000002eb, 4'd3, 27'h000001a4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000025b, 4'd1, 27'h0000021a, 4'd8, 27'h0000006a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000fa, 4'd3, 27'h00000028, 4'd10, 27'h000003be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003cb, 4'd5, 27'h00000283, 4'd1, 27'h000002a7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000ff, 4'd8, 27'h00000303, 4'd7, 27'h00000166, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000244, 4'd8, 27'h00000398, 4'd14, 27'h00000294, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002c1, 4'd12, 27'h0000007f, 4'd0, 27'h00000151, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003a9, 4'd14, 27'h000003b3, 4'd6, 27'h0000000e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001a9, 4'd14, 27'h000003d4, 4'd11, 27'h0000020a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000010c, 4'd2, 27'h000000fa, 4'd2, 27'h00000115, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000c5, 4'd3, 27'h00000260, 4'd5, 27'h00000207, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000a0, 4'd1, 27'h00000317, 4'd12, 27'h00000263, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000273, 4'd5, 27'h00000051, 4'd3, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000008c, 4'd7, 27'h000000d3, 4'd5, 27'h00000285, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000306, 4'd9, 27'h000001ad, 4'd10, 27'h000001be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000018a, 4'd14, 27'h000003d0, 4'd1, 27'h0000022d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000057, 4'd10, 27'h00000355, 4'd6, 27'h00000377, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002fc, 4'd14, 27'h000003b9, 4'd12, 27'h000001f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000021a, 4'd4, 27'h000001e3, 4'd3, 27'h000000d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000023d, 4'd4, 27'h000001ee, 4'd7, 27'h0000036a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000285, 4'd1, 27'h00000094, 4'd14, 27'h0000011d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000085, 4'd7, 27'h000001ce, 4'd2, 27'h00000115, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003a0, 4'd8, 27'h00000241, 4'd9, 27'h00000232, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000031c, 4'd7, 27'h000000e6, 4'd13, 27'h000002c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000055, 4'd11, 27'h000001d5, 4'd4, 27'h00000017, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000013d, 4'd10, 27'h000003b9, 4'd5, 27'h00000300, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000022, 4'd12, 27'h000000a3, 4'd12, 27'h0000016c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000039c, 4'd1, 27'h000001c2, 4'd3, 27'h00000143, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000017d, 4'd3, 27'h000003f9, 4'd5, 27'h0000013f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000032e, 4'd0, 27'h00000113, 4'd10, 27'h00000003, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000d4, 4'd6, 27'h00000311, 4'd0, 27'h00000214, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000339, 4'd5, 27'h000000d5, 4'd5, 27'h0000013c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000274, 4'd7, 27'h000002cd, 4'd14, 27'h0000003f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003f3, 4'd11, 27'h0000011b, 4'd3, 27'h0000029c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000000, 4'd14, 27'h0000015b, 4'd7, 27'h000003e0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000022b, 4'd13, 27'h000003ae, 4'd12, 27'h000001de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000023f, 4'd0, 27'h00000318, 4'd4, 27'h00000199, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000025a, 4'd1, 27'h000003f9, 4'd6, 27'h0000026f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000155, 4'd0, 27'h00000212, 4'd10, 27'h00000177, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003c1, 4'd5, 27'h0000015b, 4'd1, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001d1, 4'd6, 27'h000003e1, 4'd8, 27'h00000190, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000188, 4'd7, 27'h0000021d, 4'd11, 27'h0000029f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002b2, 4'd11, 27'h00000336, 4'd3, 27'h00000399, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000002a, 4'd12, 27'h0000021a, 4'd7, 27'h00000074, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000275, 4'd13, 27'h0000004a, 4'd14, 27'h000000a4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000017c, 4'd2, 27'h000002e5, 4'd2, 27'h000001ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000306, 4'd3, 27'h0000032f, 4'd8, 27'h0000000f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000003f, 4'd4, 27'h0000039f, 4'd13, 27'h00000357, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000143, 4'd5, 27'h000002d7, 4'd2, 27'h0000011d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000281, 4'd5, 27'h00000147, 4'd7, 27'h0000018f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000ae, 4'd6, 27'h00000139, 4'd11, 27'h000000dc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000036a, 4'd13, 27'h000000ea, 4'd2, 27'h00000052, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001e1, 4'd10, 27'h00000022, 4'd6, 27'h00000344, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000032d, 4'd14, 27'h0000014a, 4'd11, 27'h000002c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000160, 4'd2, 27'h00000155, 4'd2, 27'h00000127, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000321, 4'd0, 27'h00000194, 4'd9, 27'h00000164, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000ba, 4'd1, 27'h00000029, 4'd11, 27'h000002b4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000a3, 4'd5, 27'h00000168, 4'd2, 27'h00000136, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000026c, 4'd6, 27'h0000002e, 4'd8, 27'h000000d2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000b2, 4'd5, 27'h00000248, 4'd10, 27'h000000d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000021a, 4'd13, 27'h00000282, 4'd1, 27'h000001d6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003ea, 4'd12, 27'h000003d6, 4'd8, 27'h0000027a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000043, 4'd14, 27'h000003d3, 4'd12, 27'h000002fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000011d, 4'd2, 27'h00000332, 4'd0, 27'h000000c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002b7, 4'd4, 27'h000002a1, 4'd7, 27'h000001c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000159, 4'd2, 27'h000000ba, 4'd11, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000014d, 4'd7, 27'h000003e7, 4'd2, 27'h0000033e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001d6, 4'd8, 27'h00000136, 4'd8, 27'h000000d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000269, 4'd5, 27'h000003f1, 4'd14, 27'h000002c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002dc, 4'd10, 27'h0000024a, 4'd2, 27'h000000e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000154, 4'd14, 27'h0000028d, 4'd5, 27'h00000001, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b8, 4'd10, 27'h0000025d, 4'd12, 27'h000001c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000000d, 4'd4, 27'h00000078, 4'd1, 27'h000000e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003b7, 4'd2, 27'h00000273, 4'd8, 27'h00000325, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002a5, 4'd0, 27'h00000146, 4'd13, 27'h00000122, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000037e, 4'd5, 27'h000002ec, 4'd4, 27'h000002e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001cf, 4'd7, 27'h00000242, 4'd5, 27'h0000029a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001bf, 4'd7, 27'h000003c9, 4'd10, 27'h00000399, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000038b, 4'd11, 27'h00000196, 4'd1, 27'h000003e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000025b, 4'd11, 27'h0000007f, 4'd5, 27'h000001ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000005a, 4'd10, 27'h000000aa, 4'd12, 27'h00000395, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000074, 4'd0, 27'h0000033b, 4'd0, 27'h00000158, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002a2, 4'd3, 27'h000000e9, 4'd9, 27'h0000030a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000009e, 4'd3, 27'h00000112, 4'd13, 27'h000001fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000284, 4'd5, 27'h00000146, 4'd1, 27'h000002cc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000e3, 4'd6, 27'h000000c5, 4'd8, 27'h00000274, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000037, 4'd9, 27'h0000009b, 4'd13, 27'h00000092, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000091, 4'd11, 27'h000003cf, 4'd4, 27'h00000123, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000337, 4'd11, 27'h00000275, 4'd7, 27'h00000344, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000357, 4'd13, 27'h000001c9, 4'd12, 27'h000003be, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001a1, 4'd1, 27'h000000d1, 4'd1, 27'h000002ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000005c, 4'd0, 27'h00000203, 4'd5, 27'h00000378, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000028a, 4'd0, 27'h000001e7, 4'd11, 27'h0000018d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000106, 4'd6, 27'h00000246, 4'd2, 27'h00000080, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000058, 4'd8, 27'h000002f0, 4'd6, 27'h00000389, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002ca, 4'd6, 27'h0000023b, 4'd11, 27'h00000007, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000005a, 4'd12, 27'h0000010e, 4'd3, 27'h00000242, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002e2, 4'd10, 27'h00000010, 4'd8, 27'h0000031c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000070, 4'd11, 27'h000000fe, 4'd10, 27'h000003ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001fd, 4'd4, 27'h000003cc, 4'd2, 27'h00000248, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000360, 4'd2, 27'h000002e9, 4'd6, 27'h00000024, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000282, 4'd1, 27'h0000017e, 4'd14, 27'h000000c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001f9, 4'd7, 27'h000002c3, 4'd1, 27'h00000104, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000018c, 4'd6, 27'h000000ae, 4'd6, 27'h0000014e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000086, 4'd9, 27'h000003be, 4'd13, 27'h000000aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000007d, 4'd13, 27'h00000013, 4'd4, 27'h0000004a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003bb, 4'd10, 27'h00000348, 4'd7, 27'h000002ba, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003b8, 4'd14, 27'h000002df, 4'd12, 27'h00000110, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000000f, 4'd2, 27'h00000227, 4'd1, 27'h000003a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000036d, 4'd1, 27'h0000035c, 4'd9, 27'h000000eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000167, 4'd0, 27'h000000e4, 4'd13, 27'h000002b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001a3, 4'd6, 27'h00000259, 4'd3, 27'h00000050, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000020c, 4'd9, 27'h000000c3, 4'd8, 27'h0000019f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000f8, 4'd9, 27'h0000013a, 4'd14, 27'h0000004b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000019e, 4'd14, 27'h0000039a, 4'd3, 27'h0000003a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002f0, 4'd14, 27'h00000112, 4'd7, 27'h0000006c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000c4, 4'd10, 27'h000000ba, 4'd10, 27'h00000337, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000275, 4'd3, 27'h000002ad, 4'd2, 27'h00000272, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000206, 4'd0, 27'h0000019c, 4'd5, 27'h00000193, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000381, 4'd4, 27'h000001db, 4'd14, 27'h00000244, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000c4, 4'd8, 27'h000003dc, 4'd3, 27'h00000265, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003d4, 4'd7, 27'h00000287, 4'd6, 27'h000002bf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000ac, 4'd7, 27'h000002ec, 4'd13, 27'h000001c2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000024e, 4'd12, 27'h000000ea, 4'd0, 27'h00000037, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000072, 4'd10, 27'h00000380, 4'd7, 27'h000003a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000366, 4'd14, 27'h00000296, 4'd11, 27'h0000004d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000010a, 4'd3, 27'h0000032d, 4'd1, 27'h000003b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000008, 4'd1, 27'h00000114, 4'd5, 27'h000002f9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000b0, 4'd3, 27'h00000045, 4'd11, 27'h00000370, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000330, 4'd5, 27'h000003f4, 4'd2, 27'h0000023d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000023a, 4'd9, 27'h000000a4, 4'd7, 27'h00000246, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000018, 4'd6, 27'h00000364, 4'd11, 27'h0000006e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001fa, 4'd14, 27'h00000111, 4'd0, 27'h00000021, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000035f, 4'd13, 27'h00000041, 4'd8, 27'h00000045, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000142, 4'd13, 27'h000003f0, 4'd10, 27'h0000023d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000098, 4'd2, 27'h0000008a, 4'd0, 27'h00000284, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000367, 4'd3, 27'h0000006e, 4'd6, 27'h000001cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000fe, 4'd0, 27'h000002f9, 4'd11, 27'h000003f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000322, 4'd7, 27'h0000039f, 4'd0, 27'h00000337, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000073, 4'd7, 27'h000002fc, 4'd9, 27'h00000042, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000006e, 4'd9, 27'h0000023d, 4'd11, 27'h00000013, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000022f, 4'd11, 27'h00000363, 4'd4, 27'h0000024e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000027c, 4'd12, 27'h0000019f, 4'd9, 27'h00000322, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000287, 4'd10, 27'h00000294, 4'd14, 27'h000002fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000159, 4'd1, 27'h00000047, 4'd0, 27'h000002f8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000029, 4'd0, 27'h00000078, 4'd5, 27'h0000021b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000050, 4'd1, 27'h000000a4, 4'd13, 27'h0000025d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000039b, 4'd5, 27'h00000127, 4'd1, 27'h000001b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000021f, 4'd6, 27'h00000075, 4'd5, 27'h000001cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000030c, 4'd7, 27'h0000021a, 4'd11, 27'h000003e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000fd, 4'd14, 27'h00000364, 4'd3, 27'h00000362, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000ef, 4'd13, 27'h000001c9, 4'd9, 27'h000002b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000309, 4'd14, 27'h000002a3, 4'd11, 27'h000000cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003c9, 4'd2, 27'h0000004b, 4'd0, 27'h0000035a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000139, 4'd4, 27'h00000008, 4'd6, 27'h000001ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000f3, 4'd4, 27'h00000102, 4'd12, 27'h000002fb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000017c, 4'd9, 27'h00000307, 4'd4, 27'h000001da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002a2, 4'd7, 27'h00000234, 4'd7, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000db, 4'd7, 27'h00000085, 4'd11, 27'h00000255, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000140, 4'd10, 27'h0000022e, 4'd3, 27'h00000199, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000209, 4'd13, 27'h0000010e, 4'd6, 27'h00000024, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000232, 4'd14, 27'h00000336, 4'd10, 27'h00000141, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000001a, 4'd1, 27'h00000119, 4'd1, 27'h0000001a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000026f, 4'd4, 27'h000003eb, 4'd7, 27'h0000020e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000089, 4'd3, 27'h000002d1, 4'd13, 27'h0000012d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000015e, 4'd8, 27'h00000017, 4'd3, 27'h00000199, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002f7, 4'd9, 27'h000000e5, 4'd7, 27'h00000299, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001eb, 4'd6, 27'h000000ca, 4'd10, 27'h00000317, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000012d, 4'd14, 27'h0000018c, 4'd1, 27'h00000225, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000029a, 4'd11, 27'h0000012c, 4'd5, 27'h00000167, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000203, 4'd14, 27'h000002dc, 4'd11, 27'h00000104, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002f7, 4'd0, 27'h0000015f, 4'd2, 27'h0000034e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000018, 4'd4, 27'h0000033b, 4'd7, 27'h000000b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000f6, 4'd2, 27'h00000055, 4'd11, 27'h00000114, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000341, 4'd6, 27'h000002d2, 4'd4, 27'h000000ca, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000213, 4'd5, 27'h000002da, 4'd8, 27'h0000021a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000eb, 4'd7, 27'h000001fb, 4'd13, 27'h000001d9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000001d, 4'd10, 27'h0000025f, 4'd4, 27'h00000136, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000030f, 4'd12, 27'h00000366, 4'd7, 27'h00000278, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002b0, 4'd10, 27'h000002c2, 4'd13, 27'h00000111, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000208, 4'd3, 27'h00000041, 4'd4, 27'h000003c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003c6, 4'd1, 27'h000002d8, 4'd8, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000341, 4'd1, 27'h00000037, 4'd13, 27'h00000069, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000dc, 4'd8, 27'h00000245, 4'd0, 27'h00000322, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000013f, 4'd6, 27'h000003cc, 4'd8, 27'h0000004c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000e1, 4'd9, 27'h00000077, 4'd11, 27'h00000285, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000fe, 4'd12, 27'h000002b1, 4'd3, 27'h00000235, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000010f, 4'd11, 27'h00000067, 4'd5, 27'h0000035a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000042, 4'd11, 27'h00000073, 4'd13, 27'h0000038d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000000b, 4'd1, 27'h00000122, 4'd3, 27'h000001c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000174, 4'd4, 27'h00000242, 4'd6, 27'h00000237, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000223, 4'd1, 27'h000001ba, 4'd14, 27'h0000017a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000043, 4'd5, 27'h00000028, 4'd0, 27'h000003ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000c0, 4'd8, 27'h0000033f, 4'd7, 27'h000000b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000039e, 4'd6, 27'h000003f9, 4'd10, 27'h00000124, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000001, 4'd13, 27'h000000da, 4'd4, 27'h00000392, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003e1, 4'd10, 27'h000001cb, 4'd5, 27'h000003e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003be, 4'd11, 27'h0000024a, 4'd12, 27'h0000012c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000009f, 4'd1, 27'h00000348, 4'd2, 27'h000003c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000269, 4'd0, 27'h000003d0, 4'd9, 27'h0000015d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003ed, 4'd1, 27'h000000f6, 4'd13, 27'h00000065, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000095, 4'd9, 27'h00000071, 4'd2, 27'h000003fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000014, 4'd5, 27'h000000cd, 4'd9, 27'h00000187, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000053, 4'd9, 27'h00000198, 4'd12, 27'h000001be, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000356, 4'd11, 27'h000003e1, 4'd1, 27'h00000145, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000165, 4'd14, 27'h0000035a, 4'd7, 27'h00000332, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001bd, 4'd12, 27'h000000d1, 4'd12, 27'h0000020e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000013a, 4'd0, 27'h00000352, 4'd4, 27'h000002b5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001a1, 4'd0, 27'h000001ed, 4'd7, 27'h000003ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000019f, 4'd3, 27'h000000e9, 4'd14, 27'h00000235, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000280, 4'd5, 27'h00000281, 4'd0, 27'h00000337, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001da, 4'd6, 27'h000001e3, 4'd5, 27'h0000032f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000361, 4'd9, 27'h00000015, 4'd12, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000d4, 4'd10, 27'h00000181, 4'd4, 27'h000001e2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002fc, 4'd13, 27'h000003e6, 4'd8, 27'h000001f4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002de, 4'd11, 27'h000003bd, 4'd11, 27'h000003e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000015e, 4'd3, 27'h000003a5, 4'd1, 27'h00000140, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000328, 4'd3, 27'h000002ed, 4'd8, 27'h00000228, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000002f, 4'd0, 27'h00000015, 4'd12, 27'h000000ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000b2, 4'd7, 27'h00000178, 4'd0, 27'h00000171, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000198, 4'd7, 27'h0000014f, 4'd6, 27'h00000117, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001c7, 4'd9, 27'h00000269, 4'd13, 27'h00000252, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000b1, 4'd14, 27'h00000292, 4'd4, 27'h00000359, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000198, 4'd14, 27'h0000036e, 4'd7, 27'h0000030a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000002, 4'd10, 27'h0000030c, 4'd10, 27'h000003c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001ab, 4'd3, 27'h00000201, 4'd0, 27'h00000269, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000175, 4'd1, 27'h000002b7, 4'd6, 27'h00000004, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000f6, 4'd1, 27'h000000e0, 4'd13, 27'h00000379, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000201, 4'd7, 27'h00000355, 4'd3, 27'h00000124, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001e6, 4'd7, 27'h000000c4, 4'd5, 27'h000003d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000388, 4'd6, 27'h00000024, 4'd14, 27'h00000388, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003c0, 4'd10, 27'h00000203, 4'd1, 27'h00000245, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000297, 4'd13, 27'h0000030a, 4'd9, 27'h00000327, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002d0, 4'd14, 27'h000002eb, 4'd14, 27'h0000010d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000209, 4'd3, 27'h0000032c, 4'd3, 27'h000002ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000028f, 4'd4, 27'h000000ef, 4'd8, 27'h00000050, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000045, 4'd4, 27'h0000027b, 4'd10, 27'h000002db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000165, 4'd7, 27'h000001cb, 4'd4, 27'h000001e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000010f, 4'd8, 27'h00000282, 4'd9, 27'h0000018a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003a6, 4'd7, 27'h00000013, 4'd11, 27'h000000c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000214, 4'd10, 27'h0000038e, 4'd0, 27'h000002ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000054, 4'd12, 27'h0000000a, 4'd7, 27'h000003e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000006a, 4'd14, 27'h000000c3, 4'd10, 27'h00000156, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002d8, 4'd4, 27'h00000390, 4'd2, 27'h00000169, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000322, 4'd2, 27'h00000091, 4'd8, 27'h00000345, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002a4, 4'd3, 27'h000002d2, 4'd13, 27'h000001ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001de, 4'd9, 27'h0000015f, 4'd0, 27'h000000d8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000cc, 4'd8, 27'h0000011e, 4'd7, 27'h000002b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000012e, 4'd9, 27'h00000083, 4'd10, 27'h00000100, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ed, 4'd14, 27'h0000021d, 4'd1, 27'h00000015, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002a5, 4'd12, 27'h000000c5, 4'd5, 27'h000002cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000203, 4'd12, 27'h00000283, 4'd11, 27'h000000f4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000057, 4'd2, 27'h000003e0, 4'd3, 27'h00000382, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000022, 4'd4, 27'h0000039b, 4'd7, 27'h000003fb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003f2, 4'd3, 27'h00000098, 4'd12, 27'h000003ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000203, 4'd7, 27'h000002ab, 4'd1, 27'h00000100, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000203, 4'd8, 27'h000000e1, 4'd6, 27'h00000293, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000258, 4'd7, 27'h0000010b, 4'd10, 27'h00000338, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000286, 4'd13, 27'h0000037d, 4'd1, 27'h0000003f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000336, 4'd14, 27'h000000cf, 4'd5, 27'h000000b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000020c, 4'd11, 27'h00000057, 4'd13, 27'h00000387, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001f7, 4'd2, 27'h00000398, 4'd3, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000011a, 4'd2, 27'h0000021f, 4'd6, 27'h000001a2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000362, 4'd1, 27'h00000343, 4'd13, 27'h0000007f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002a2, 4'd9, 27'h0000008a, 4'd0, 27'h00000340, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003d8, 4'd6, 27'h000001d6, 4'd8, 27'h000003d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000021b, 4'd8, 27'h00000184, 4'd12, 27'h0000030a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000012c, 4'd14, 27'h00000350, 4'd0, 27'h00000263, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000238, 4'd12, 27'h000001ab, 4'd8, 27'h000000b3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003ad, 4'd13, 27'h0000011d, 4'd13, 27'h000002a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000104, 4'd0, 27'h0000000a, 4'd2, 27'h00000150, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000017, 4'd2, 27'h0000007b, 4'd7, 27'h0000000d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c5, 4'd2, 27'h00000297, 4'd12, 27'h000001b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000f7, 4'd8, 27'h000003a1, 4'd1, 27'h00000255, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000028a, 4'd7, 27'h000001cb, 4'd7, 27'h0000006f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000307, 4'd5, 27'h0000035b, 4'd14, 27'h00000029, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000078, 4'd10, 27'h0000013a, 4'd4, 27'h00000130, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000010a, 4'd14, 27'h00000337, 4'd5, 27'h0000017d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003f3, 4'd13, 27'h0000021c, 4'd10, 27'h00000059, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000dc, 4'd3, 27'h0000037c, 4'd4, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000109, 4'd3, 27'h000000d8, 4'd9, 27'h00000293, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000ec, 4'd4, 27'h00000109, 4'd12, 27'h000003a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000013f, 4'd5, 27'h000003c9, 4'd4, 27'h000001d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000356, 4'd5, 27'h00000219, 4'd7, 27'h0000008e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001ea, 4'd6, 27'h0000001d, 4'd12, 27'h0000039b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000039d, 4'd13, 27'h00000398, 4'd1, 27'h00000323, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000153, 4'd14, 27'h000003f6, 4'd7, 27'h00000222, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000370, 4'd14, 27'h00000379, 4'd12, 27'h00000194, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000018f, 4'd1, 27'h00000160, 4'd4, 27'h0000021e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000248, 4'd1, 27'h00000169, 4'd7, 27'h0000034c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000393, 4'd1, 27'h000001e6, 4'd12, 27'h000000f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002ee, 4'd8, 27'h000002b7, 4'd3, 27'h00000316, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003da, 4'd9, 27'h00000158, 4'd5, 27'h0000023b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000045, 4'd7, 27'h0000037c, 4'd11, 27'h0000005e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001df, 4'd11, 27'h00000113, 4'd1, 27'h0000005f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000003f, 4'd12, 27'h00000359, 4'd9, 27'h000000ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001fc, 4'd11, 27'h00000098, 4'd10, 27'h00000289, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000024a, 4'd3, 27'h0000029e, 4'd3, 27'h00000246, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003f5, 4'd3, 27'h0000033a, 4'd9, 27'h00000087, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000036c, 4'd2, 27'h0000035e, 4'd12, 27'h00000104, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000067, 4'd8, 27'h0000031a, 4'd2, 27'h000000be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000387, 4'd7, 27'h0000022a, 4'd6, 27'h000000d4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000336, 4'd5, 27'h00000138, 4'd13, 27'h000001f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000017e, 4'd14, 27'h00000101, 4'd1, 27'h00000033, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000293, 4'd12, 27'h000003c3, 4'd7, 27'h000001a2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000d5, 4'd13, 27'h00000128, 4'd14, 27'h00000312, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000015a, 4'd2, 27'h00000188, 4'd1, 27'h000002d4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000269, 4'd2, 27'h000003df, 4'd5, 27'h00000062, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000175, 4'd0, 27'h00000206, 4'd14, 27'h0000036c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000367, 4'd7, 27'h0000000b, 4'd1, 27'h0000036e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000152, 4'd9, 27'h000001cb, 4'd6, 27'h00000060, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001c2, 4'd5, 27'h00000359, 4'd11, 27'h00000179, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003b7, 4'd13, 27'h00000020, 4'd3, 27'h0000029e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000e3, 4'd13, 27'h0000010b, 4'd6, 27'h00000073, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000092, 4'd14, 27'h0000016d, 4'd11, 27'h00000178, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000333, 4'd4, 27'h0000001f, 4'd0, 27'h00000394, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000002b, 4'd3, 27'h000001c7, 4'd5, 27'h00000005, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000cb, 4'd2, 27'h0000006e, 4'd12, 27'h000000e5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002e7, 4'd8, 27'h00000249, 4'd3, 27'h00000299, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000009f, 4'd9, 27'h00000315, 4'd7, 27'h000001bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002ff, 4'd9, 27'h00000033, 4'd11, 27'h0000015b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000010, 4'd10, 27'h000002b5, 4'd0, 27'h0000001c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000352, 4'd11, 27'h000001a0, 4'd9, 27'h00000063, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000113, 4'd14, 27'h00000015, 4'd13, 27'h000001ea, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000374, 4'd1, 27'h00000369, 4'd1, 27'h000003e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000241, 4'd4, 27'h0000013e, 4'd5, 27'h00000063, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002ac, 4'd2, 27'h000003d6, 4'd14, 27'h00000274, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000038a, 4'd6, 27'h000003f9, 4'd0, 27'h0000030a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000395, 4'd8, 27'h00000094, 4'd7, 27'h0000004b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001f0, 4'd8, 27'h00000212, 4'd11, 27'h000000e9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000327, 4'd13, 27'h000002bc, 4'd2, 27'h000001eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000d2, 4'd10, 27'h0000033e, 4'd5, 27'h00000045, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000367, 4'd13, 27'h000001c2, 4'd14, 27'h00000210, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000034d, 4'd1, 27'h00000380, 4'd4, 27'h000001de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000169, 4'd0, 27'h00000323, 4'd9, 27'h0000039c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000007d, 4'd3, 27'h0000007f, 4'd10, 27'h00000118, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000030e, 4'd6, 27'h00000398, 4'd1, 27'h0000027c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000029a, 4'd6, 27'h0000002d, 4'd8, 27'h0000030c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001ce, 4'd5, 27'h00000145, 4'd12, 27'h00000277, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000021c, 4'd13, 27'h0000008b, 4'd1, 27'h000002fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000395, 4'd13, 27'h0000010e, 4'd6, 27'h000001ff, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000069, 4'd10, 27'h000003b5, 4'd13, 27'h000001e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000024a, 4'd0, 27'h00000057, 4'd2, 27'h000001bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000016a, 4'd0, 27'h00000316, 4'd7, 27'h000003b7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003b2, 4'd3, 27'h000001fd, 4'd13, 27'h0000014e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000244, 4'd5, 27'h000002c9, 4'd0, 27'h00000022, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002e8, 4'd7, 27'h000003dd, 4'd9, 27'h00000325, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000004, 4'd8, 27'h00000192, 4'd14, 27'h0000031d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000039d, 4'd14, 27'h00000033, 4'd3, 27'h0000028d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000179, 4'd11, 27'h000003c5, 4'd9, 27'h000001c4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000194, 4'd12, 27'h00000178, 4'd14, 27'h00000220, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001b5, 4'd4, 27'h000002a8, 4'd1, 27'h000002d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002ab, 4'd1, 27'h00000336, 4'd7, 27'h00000372, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001f7, 4'd1, 27'h0000001d, 4'd13, 27'h000003a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003a3, 4'd9, 27'h00000130, 4'd2, 27'h000000e8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000cc, 4'd5, 27'h000002cf, 4'd6, 27'h00000104, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000004a, 4'd5, 27'h0000006e, 4'd12, 27'h00000392, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001f5, 4'd12, 27'h000003b3, 4'd2, 27'h00000305, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002c3, 4'd11, 27'h00000285, 4'd5, 27'h00000360, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001db, 4'd14, 27'h0000028d, 4'd14, 27'h00000121, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003e4, 4'd0, 27'h00000257, 4'd1, 27'h00000319, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000db, 4'd4, 27'h000000e6, 4'd8, 27'h0000007e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003d3, 4'd4, 27'h0000031a, 4'd13, 27'h00000217, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000077, 4'd7, 27'h000002d4, 4'd0, 27'h00000220, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001df, 4'd7, 27'h00000148, 4'd7, 27'h0000024a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000c9, 4'd5, 27'h00000164, 4'd13, 27'h00000192, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000097, 4'd12, 27'h000000a8, 4'd2, 27'h00000189, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000db, 4'd11, 27'h000001ba, 4'd8, 27'h00000035, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000027f, 4'd11, 27'h000003c7, 4'd10, 27'h000001f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000e4, 4'd0, 27'h0000013d, 4'd0, 27'h0000033d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001e9, 4'd4, 27'h00000385, 4'd7, 27'h00000362, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000381, 4'd2, 27'h00000033, 4'd10, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000b0, 4'd8, 27'h00000195, 4'd4, 27'h00000024, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001a7, 4'd7, 27'h0000039e, 4'd6, 27'h00000013, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002e7, 4'd6, 27'h00000257, 4'd13, 27'h00000110, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000039a, 4'd11, 27'h0000018a, 4'd3, 27'h00000399, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000163, 4'd10, 27'h00000227, 4'd8, 27'h00000099, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000190, 4'd10, 27'h000000c1, 4'd10, 27'h000002de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ad, 4'd2, 27'h00000349, 4'd2, 27'h00000203, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000264, 4'd4, 27'h000001b6, 4'd6, 27'h00000020, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000301, 4'd4, 27'h00000011, 4'd14, 27'h00000149, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000013a, 4'd5, 27'h00000100, 4'd3, 27'h00000181, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000186, 4'd6, 27'h00000143, 4'd8, 27'h000002f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000369, 4'd6, 27'h00000144, 4'd11, 27'h000001e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000175, 4'd11, 27'h00000197, 4'd3, 27'h00000283, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000294, 4'd13, 27'h00000161, 4'd9, 27'h0000037b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000236, 4'd12, 27'h000003db, 4'd14, 27'h000003fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000014e, 4'd3, 27'h00000305, 4'd4, 27'h00000149, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002c7, 4'd3, 27'h000003bc, 4'd7, 27'h00000137, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000276, 4'd0, 27'h00000060, 4'd10, 27'h0000020e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000045, 4'd7, 27'h000000ff, 4'd4, 27'h0000023b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000098, 4'd5, 27'h000002c6, 4'd9, 27'h000002c8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000004a, 4'd8, 27'h00000099, 4'd11, 27'h000000e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000ef, 4'd11, 27'h00000218, 4'd3, 27'h0000005d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000233, 4'd11, 27'h000002d4, 4'd5, 27'h0000013f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000331, 4'd14, 27'h000003b9, 4'd13, 27'h00000215, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000261, 4'd4, 27'h00000393, 4'd0, 27'h0000022f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c5, 4'd0, 27'h0000022f, 4'd6, 27'h00000077, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002d7, 4'd1, 27'h0000003a, 4'd11, 27'h0000007a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000371, 4'd9, 27'h00000307, 4'd3, 27'h00000282, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000025f, 4'd7, 27'h00000161, 4'd9, 27'h00000335, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002fc, 4'd8, 27'h00000261, 4'd14, 27'h00000161, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000008b, 4'd14, 27'h00000141, 4'd0, 27'h00000248, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000367, 4'd14, 27'h00000183, 4'd6, 27'h00000394, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000048, 4'd13, 27'h0000005e, 4'd10, 27'h000002b4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002eb, 4'd1, 27'h00000046, 4'd4, 27'h000002ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000de, 4'd1, 27'h0000030e, 4'd9, 27'h000003b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003ed, 4'd2, 27'h00000021, 4'd13, 27'h000002f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002a6, 4'd9, 27'h00000072, 4'd0, 27'h0000016b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000fd, 4'd5, 27'h00000095, 4'd9, 27'h0000024b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000f8, 4'd9, 27'h00000246, 4'd12, 27'h00000143, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000ac, 4'd12, 27'h00000309, 4'd1, 27'h000000a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000038, 4'd10, 27'h000001dc, 4'd5, 27'h000003f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000bb, 4'd10, 27'h00000363, 4'd11, 27'h0000032c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000027c, 4'd0, 27'h0000005e, 4'd4, 27'h000000a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000000a, 4'd4, 27'h0000009f, 4'd7, 27'h00000216, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000033e, 4'd3, 27'h000001fc, 4'd11, 27'h00000215, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000034d, 4'd9, 27'h00000157, 4'd4, 27'h00000095, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001ff, 4'd6, 27'h00000295, 4'd9, 27'h000003fb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002f7, 4'd8, 27'h000002f3, 4'd13, 27'h000001ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000ae, 4'd11, 27'h00000025, 4'd4, 27'h00000111, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000006f, 4'd13, 27'h00000213, 4'd7, 27'h000003dc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000029f, 4'd14, 27'h00000257, 4'd14, 27'h0000026c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002e0, 4'd2, 27'h0000011c, 4'd4, 27'h000001bb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001aa, 4'd4, 27'h0000011b, 4'd8, 27'h00000314, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000134, 4'd0, 27'h000002a5, 4'd13, 27'h000000cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002d5, 4'd5, 27'h000003a2, 4'd2, 27'h00000062, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000146, 4'd8, 27'h00000210, 4'd5, 27'h000002e6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000b1, 4'd5, 27'h0000020a, 4'd11, 27'h000002e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000b7, 4'd12, 27'h00000012, 4'd0, 27'h00000326, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000020d, 4'd12, 27'h00000053, 4'd8, 27'h00000112, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000057, 4'd13, 27'h000001ee, 4'd12, 27'h00000294, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000039c, 4'd2, 27'h000003b4, 4'd2, 27'h000003e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000028, 4'd1, 27'h00000036, 4'd9, 27'h00000112, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001ab, 4'd4, 27'h00000040, 4'd11, 27'h00000317, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000277, 4'd8, 27'h000003a4, 4'd1, 27'h00000177, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002a6, 4'd6, 27'h00000202, 4'd8, 27'h0000034d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000216, 4'd6, 27'h000000af, 4'd10, 27'h000001b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000111, 4'd12, 27'h000000ae, 4'd3, 27'h00000305, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000034a, 4'd14, 27'h00000097, 4'd8, 27'h000000c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000217, 4'd12, 27'h000001e2, 4'd10, 27'h0000025e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000030f, 4'd1, 27'h000001b0, 4'd3, 27'h000003ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000032b, 4'd1, 27'h000003ec, 4'd9, 27'h00000268, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000274, 4'd0, 27'h000003a8, 4'd13, 27'h000000b3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000171, 4'd9, 27'h00000200, 4'd2, 27'h000002bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000013f, 4'd7, 27'h000001e3, 4'd6, 27'h000003fe, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000068, 4'd8, 27'h00000092, 4'd14, 27'h0000013f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000e5, 4'd14, 27'h00000311, 4'd4, 27'h00000311, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000183, 4'd10, 27'h0000024e, 4'd5, 27'h000003c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000268, 4'd12, 27'h00000196, 4'd11, 27'h000001cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000da, 4'd1, 27'h000001c2, 4'd4, 27'h0000038c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000239, 4'd3, 27'h00000147, 4'd9, 27'h0000028a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000206, 4'd1, 27'h000003dc, 4'd13, 27'h00000249, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000227, 4'd6, 27'h000001e0, 4'd3, 27'h0000033e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000168, 4'd9, 27'h0000034b, 4'd7, 27'h0000018f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000174, 4'd8, 27'h00000128, 4'd12, 27'h000001f1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000005e, 4'd13, 27'h000000a6, 4'd3, 27'h0000039d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c4, 4'd14, 27'h000001b8, 4'd8, 27'h00000207, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000006, 4'd10, 27'h000001e4, 4'd12, 27'h00000380, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000351, 4'd1, 27'h0000016c, 4'd2, 27'h0000025b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000341, 4'd4, 27'h0000028d, 4'd5, 27'h000001e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000006c, 4'd1, 27'h0000006a, 4'd14, 27'h0000013b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000008f, 4'd6, 27'h000003cf, 4'd1, 27'h00000194, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000014d, 4'd5, 27'h0000026a, 4'd8, 27'h0000030d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000a8, 4'd7, 27'h000001e5, 4'd13, 27'h0000033f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000037d, 4'd12, 27'h000003e3, 4'd3, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000103, 4'd14, 27'h000000fb, 4'd7, 27'h0000006b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002fe, 4'd12, 27'h00000225, 4'd12, 27'h00000220, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003a7, 4'd4, 27'h00000025, 4'd4, 27'h00000150, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001db, 4'd1, 27'h00000175, 4'd6, 27'h000003ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000108, 4'd2, 27'h000002bb, 4'd10, 27'h00000016, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000039b, 4'd6, 27'h0000028d, 4'd2, 27'h00000376, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000007b, 4'd5, 27'h00000077, 4'd6, 27'h00000172, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000299, 4'd9, 27'h000000eb, 4'd12, 27'h000002ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000039b, 4'd12, 27'h000000d4, 4'd3, 27'h00000036, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000164, 4'd12, 27'h0000008a, 4'd7, 27'h000001e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000247, 4'd14, 27'h000001ba, 4'd10, 27'h000000fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003a0, 4'd0, 27'h00000085, 4'd1, 27'h000003a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000c6, 4'd4, 27'h000000c3, 4'd7, 27'h000003f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000161, 4'd3, 27'h000003a1, 4'd11, 27'h000000d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000245, 4'd7, 27'h000002f2, 4'd1, 27'h000002bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003cc, 4'd9, 27'h0000015e, 4'd5, 27'h000000cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000050, 4'd9, 27'h0000017f, 4'd12, 27'h00000124, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000095, 4'd13, 27'h0000024f, 4'd1, 27'h00000290, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000008c, 4'd10, 27'h0000020d, 4'd8, 27'h00000256, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000038d, 4'd10, 27'h00000360, 4'd12, 27'h00000157, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000027e, 4'd4, 27'h00000016, 4'd2, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000371, 4'd1, 27'h00000120, 4'd6, 27'h000002ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001a8, 4'd0, 27'h000000dd, 4'd13, 27'h000000a8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000017e, 4'd6, 27'h0000021a, 4'd1, 27'h000003de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000de, 4'd9, 27'h00000060, 4'd8, 27'h00000283, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003ff, 4'd7, 27'h00000268, 4'd11, 27'h00000074, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001e3, 4'd14, 27'h00000253, 4'd1, 27'h00000110, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000009e, 4'd10, 27'h0000027b, 4'd6, 27'h00000088, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000021, 4'd13, 27'h00000139, 4'd11, 27'h0000017e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000fc, 4'd2, 27'h00000398, 4'd2, 27'h00000284, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000295, 4'd1, 27'h00000367, 4'd6, 27'h00000097, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000030d, 4'd2, 27'h000002bb, 4'd13, 27'h0000038c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000027c, 4'd5, 27'h000003d4, 4'd2, 27'h0000011e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000157, 4'd5, 27'h0000017d, 4'd6, 27'h0000012c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000003d, 4'd7, 27'h00000044, 4'd13, 27'h000000d2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001d8, 4'd12, 27'h0000001d, 4'd0, 27'h0000005c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000121, 4'd13, 27'h0000027c, 4'd7, 27'h00000091, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000a7, 4'd13, 27'h00000291, 4'd10, 27'h0000011e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000004e, 4'd0, 27'h0000033b, 4'd0, 27'h000001fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000032f, 4'd4, 27'h000003f4, 4'd8, 27'h0000037f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000103, 4'd0, 27'h0000035b, 4'd12, 27'h000003e1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003b9, 4'd6, 27'h00000027, 4'd4, 27'h0000016e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000381, 4'd8, 27'h00000051, 4'd5, 27'h00000313, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000019, 4'd5, 27'h000002a6, 4'd10, 27'h00000220, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000025b, 4'd10, 27'h00000118, 4'd3, 27'h0000026d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000034c, 4'd12, 27'h0000036e, 4'd9, 27'h0000001e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000283, 4'd13, 27'h00000238, 4'd10, 27'h00000086, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000035a, 4'd0, 27'h00000014, 4'd3, 27'h0000013e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000087, 4'd0, 27'h000003f8, 4'd9, 27'h0000031f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000012e, 4'd0, 27'h00000322, 4'd13, 27'h00000056, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000354, 4'd5, 27'h0000019f, 4'd2, 27'h0000028c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000026a, 4'd6, 27'h0000004c, 4'd7, 27'h00000249, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000038b, 4'd7, 27'h0000032f, 4'd10, 27'h000001c7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000183, 4'd10, 27'h000001a1, 4'd4, 27'h000002b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000289, 4'd13, 27'h00000041, 4'd8, 27'h0000010c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000003d, 4'd13, 27'h00000313, 4'd12, 27'h00000007, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000116, 4'd0, 27'h0000022b, 4'd1, 27'h00000282, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000057, 4'd0, 27'h000001c8, 4'd5, 27'h000002fa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000aa, 4'd3, 27'h00000039, 4'd12, 27'h00000200, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002f3, 4'd6, 27'h00000305, 4'd0, 27'h0000036a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000313, 4'd9, 27'h0000023b, 4'd8, 27'h000002de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000004, 4'd9, 27'h00000137, 4'd14, 27'h00000171, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000099, 4'd14, 27'h00000122, 4'd2, 27'h00000227, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000208, 4'd10, 27'h000000ce, 4'd8, 27'h0000013c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001c1, 4'd13, 27'h000001e8, 4'd12, 27'h000000d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000004a, 4'd2, 27'h00000007, 4'd4, 27'h00000316, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000258, 4'd3, 27'h00000116, 4'd8, 27'h00000123, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000149, 4'd1, 27'h0000024e, 4'd12, 27'h00000008, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001cb, 4'd8, 27'h00000312, 4'd4, 27'h000002be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000030a, 4'd9, 27'h0000025c, 4'd6, 27'h000003ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003bb, 4'd6, 27'h00000174, 4'd12, 27'h00000023, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001ff, 4'd13, 27'h000001f3, 4'd0, 27'h000001a8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000021b, 4'd13, 27'h000003ee, 4'd9, 27'h00000116, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002f4, 4'd13, 27'h000002da, 4'd11, 27'h00000280, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000135, 4'd3, 27'h0000039c, 4'd2, 27'h0000006a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000128, 4'd3, 27'h00000077, 4'd8, 27'h00000074, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001c8, 4'd4, 27'h000003d0, 4'd13, 27'h00000167, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000026e, 4'd6, 27'h0000022e, 4'd1, 27'h0000001a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000395, 4'd7, 27'h000002fa, 4'd9, 27'h00000308, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001d1, 4'd8, 27'h0000006a, 4'd14, 27'h000001b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000018b, 4'd11, 27'h00000355, 4'd2, 27'h00000029, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002de, 4'd14, 27'h00000043, 4'd8, 27'h000002e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000018b, 4'd14, 27'h00000340, 4'd11, 27'h000003e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003df, 4'd3, 27'h000000d2, 4'd0, 27'h000002d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000087, 4'd0, 27'h0000009c, 4'd6, 27'h000001bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000049, 4'd4, 27'h000001e9, 4'd13, 27'h00000392, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000305, 4'd9, 27'h000003b2, 4'd1, 27'h000000fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002e8, 4'd8, 27'h000003fe, 4'd9, 27'h00000030, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002e5, 4'd5, 27'h0000026e, 4'd10, 27'h0000039d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002a9, 4'd11, 27'h000000ed, 4'd4, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003f5, 4'd12, 27'h00000262, 4'd6, 27'h0000031e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003e6, 4'd11, 27'h00000317, 4'd13, 27'h000000a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000024c, 4'd1, 27'h00000152, 4'd3, 27'h00000352, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000200, 4'd0, 27'h00000046, 4'd8, 27'h00000190, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003f3, 4'd3, 27'h000001fb, 4'd12, 27'h00000011, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003e2, 4'd6, 27'h000000de, 4'd0, 27'h00000182, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000021f, 4'd8, 27'h000003cc, 4'd5, 27'h0000000f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000034e, 4'd6, 27'h0000003b, 4'd12, 27'h000000a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ce, 4'd11, 27'h00000039, 4'd2, 27'h00000303, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000008b, 4'd11, 27'h0000014f, 4'd7, 27'h000001db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000172, 4'd10, 27'h00000192, 4'd11, 27'h0000006c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000374, 4'd2, 27'h000001d5, 4'd1, 27'h0000010e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000193, 4'd3, 27'h00000138, 4'd7, 27'h00000156, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000168, 4'd4, 27'h000003be, 4'd11, 27'h0000038e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000034, 4'd5, 27'h000003a2, 4'd1, 27'h00000072, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000be, 4'd6, 27'h000003f1, 4'd6, 27'h000002c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000005, 4'd6, 27'h00000092, 4'd13, 27'h000003c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000017, 4'd13, 27'h00000394, 4'd2, 27'h000002cb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002c4, 4'd12, 27'h000002cd, 4'd5, 27'h00000066, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002f0, 4'd10, 27'h0000008d, 4'd12, 27'h000001a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000001c, 4'd4, 27'h00000373, 4'd3, 27'h00000345, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000227, 4'd3, 27'h00000033, 4'd8, 27'h0000037f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003b4, 4'd1, 27'h000000fd, 4'd13, 27'h00000048, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001ad, 4'd6, 27'h0000033c, 4'd3, 27'h00000020, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003f7, 4'd5, 27'h000003f2, 4'd7, 27'h0000008c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000335, 4'd9, 27'h0000010b, 4'd12, 27'h000001ef, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001cf, 4'd14, 27'h000002e5, 4'd1, 27'h0000033b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000035b, 4'd14, 27'h00000084, 4'd6, 27'h00000270, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000036, 4'd10, 27'h000000bd, 4'd14, 27'h000001bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002c9, 4'd0, 27'h00000376, 4'd1, 27'h000002f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000045, 4'd1, 27'h00000355, 4'd8, 27'h0000024c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000158, 4'd1, 27'h00000388, 4'd11, 27'h000000c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000f3, 4'd6, 27'h000001f1, 4'd2, 27'h000003a0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002bf, 4'd8, 27'h0000008f, 4'd6, 27'h000001eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000dc, 4'd8, 27'h00000290, 4'd11, 27'h000001bf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000201, 4'd11, 27'h00000131, 4'd0, 27'h000001d3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000034b, 4'd14, 27'h000003a8, 4'd7, 27'h00000312, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001d1, 4'd12, 27'h0000036f, 4'd12, 27'h0000027b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002c6, 4'd4, 27'h00000238, 4'd0, 27'h0000034a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002fa, 4'd0, 27'h000002f4, 4'd6, 27'h00000231, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003c7, 4'd3, 27'h0000028e, 4'd13, 27'h00000189, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000097, 4'd7, 27'h00000305, 4'd1, 27'h0000027b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000129, 4'd8, 27'h0000024f, 4'd8, 27'h0000023e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003c7, 4'd8, 27'h0000016b, 4'd12, 27'h0000009e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000020e, 4'd12, 27'h0000024e, 4'd2, 27'h000001c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001c3, 4'd10, 27'h000001e5, 4'd8, 27'h000002fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000216, 4'd14, 27'h000002d4, 4'd11, 27'h00000150, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000005c, 4'd2, 27'h000000a2, 4'd2, 27'h0000014a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002cb, 4'd3, 27'h000001d1, 4'd9, 27'h000001d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000000d, 4'd3, 27'h00000201, 4'd11, 27'h000003c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000182, 4'd6, 27'h000001cd, 4'd4, 27'h000003d7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000097, 4'd5, 27'h0000032c, 4'd6, 27'h00000062, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000341, 4'd5, 27'h0000019a, 4'd10, 27'h000003e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002f2, 4'd10, 27'h0000039b, 4'd4, 27'h000002e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ea, 4'd12, 27'h0000012a, 4'd9, 27'h000000c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000025b, 4'd13, 27'h000002b3, 4'd12, 27'h00000305, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001fa, 4'd4, 27'h000002fc, 4'd0, 27'h00000012, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000300, 4'd4, 27'h00000084, 4'd6, 27'h00000070, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000120, 4'd0, 27'h00000218, 4'd12, 27'h0000034c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000029c, 4'd8, 27'h00000376, 4'd1, 27'h00000065, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002b3, 4'd7, 27'h000003f1, 4'd5, 27'h000001db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000022d, 4'd6, 27'h00000196, 4'd10, 27'h000001b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000239, 4'd14, 27'h000001dc, 4'd0, 27'h00000130, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000387, 4'd12, 27'h000001cd, 4'd7, 27'h000003c3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001bf, 4'd14, 27'h000003bb, 4'd11, 27'h00000166, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000379, 4'd4, 27'h0000001b, 4'd1, 27'h00000352, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000ba, 4'd2, 27'h0000022d, 4'd9, 27'h000003b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000290, 4'd4, 27'h0000019a, 4'd12, 27'h000001ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000347, 4'd5, 27'h00000374, 4'd1, 27'h00000218, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000038c, 4'd5, 27'h00000001, 4'd6, 27'h0000031d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000016, 4'd9, 27'h00000291, 4'd13, 27'h000002e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000020c, 4'd11, 27'h0000022d, 4'd4, 27'h00000364, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000bf, 4'd10, 27'h000001a9, 4'd7, 27'h000003bc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000332, 4'd14, 27'h000003b7, 4'd11, 27'h00000187, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000034c, 4'd3, 27'h00000082, 4'd0, 27'h000001d3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000275, 4'd3, 27'h00000080, 4'd5, 27'h00000224, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003fd, 4'd3, 27'h00000353, 4'd14, 27'h0000004d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000028b, 4'd5, 27'h00000090, 4'd3, 27'h000002c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000258, 4'd8, 27'h00000095, 4'd9, 27'h00000184, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000305, 4'd5, 27'h000000d0, 4'd10, 27'h00000336, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000137, 4'd10, 27'h0000011e, 4'd0, 27'h000002fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003ac, 4'd12, 27'h00000199, 4'd6, 27'h0000022c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000025c, 4'd12, 27'h000002c8, 4'd14, 27'h00000244, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000163, 4'd2, 27'h00000140, 4'd3, 27'h00000297, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001fb, 4'd3, 27'h00000057, 4'd6, 27'h00000306, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000010c, 4'd1, 27'h00000009, 4'd12, 27'h0000004f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000025c, 4'd7, 27'h0000037a, 4'd4, 27'h00000031, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000361, 4'd5, 27'h000002f5, 4'd6, 27'h00000315, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001b9, 4'd9, 27'h00000134, 4'd14, 27'h000001f7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000155, 4'd12, 27'h000001c6, 4'd4, 27'h00000343, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000028c, 4'd13, 27'h0000029d, 4'd9, 27'h00000085, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001fa, 4'd13, 27'h000002aa, 4'd12, 27'h00000384, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000026b, 4'd0, 27'h00000282, 4'd2, 27'h000002ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003d4, 4'd4, 27'h0000028c, 4'd6, 27'h000000d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000007, 4'd4, 27'h000000ff, 4'd14, 27'h000002bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000009c, 4'd5, 27'h00000056, 4'd2, 27'h000002bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000398, 4'd7, 27'h00000366, 4'd9, 27'h000003c0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001e8, 4'd7, 27'h000000c5, 4'd14, 27'h00000019, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000008d, 4'd12, 27'h0000000e, 4'd0, 27'h00000100, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ab, 4'd10, 27'h00000399, 4'd9, 27'h00000308, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000075, 4'd10, 27'h0000009d, 4'd12, 27'h00000198, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002d0, 4'd4, 27'h00000243, 4'd0, 27'h00000316, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000225, 4'd3, 27'h00000369, 4'd7, 27'h000000b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003b9, 4'd2, 27'h000003ed, 4'd13, 27'h00000142, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002c7, 4'd6, 27'h000002cb, 4'd0, 27'h0000018d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001a0, 4'd5, 27'h00000369, 4'd6, 27'h00000038, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000023b, 4'd8, 27'h0000039a, 4'd13, 27'h000001df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000002d, 4'd13, 27'h0000003b, 4'd1, 27'h000003f0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000029b, 4'd10, 27'h000003b4, 4'd8, 27'h000000f3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000301, 4'd10, 27'h0000032a, 4'd10, 27'h00000133, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000020d, 4'd3, 27'h000001b9, 4'd0, 27'h00000305, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001fc, 4'd2, 27'h000000ef, 4'd8, 27'h000003ef, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000144, 4'd2, 27'h0000039b, 4'd13, 27'h00000200, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001bb, 4'd8, 27'h000003b3, 4'd4, 27'h00000117, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001c6, 4'd8, 27'h00000323, 4'd7, 27'h00000279, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000024f, 4'd6, 27'h00000106, 4'd11, 27'h00000168, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002ea, 4'd14, 27'h000002b7, 4'd1, 27'h000002d6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000b6, 4'd10, 27'h000001a0, 4'd6, 27'h000001d1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000024a, 4'd12, 27'h0000023b, 4'd10, 27'h00000049, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000169, 4'd0, 27'h00000177, 4'd1, 27'h0000037e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000dc, 4'd2, 27'h00000230, 4'd8, 27'h00000242, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001ef, 4'd1, 27'h0000039f, 4'd14, 27'h000002dc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000398, 4'd7, 27'h00000163, 4'd1, 27'h000001f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000158, 4'd6, 27'h0000011e, 4'd5, 27'h000000c7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000065, 4'd5, 27'h00000371, 4'd13, 27'h000003f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000237, 4'd11, 27'h000000cc, 4'd4, 27'h000000bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000108, 4'd14, 27'h00000082, 4'd5, 27'h0000021a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000071, 4'd11, 27'h000001bf, 4'd14, 27'h000001b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002af, 4'd4, 27'h00000342, 4'd1, 27'h00000166, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001e0, 4'd2, 27'h00000308, 4'd8, 27'h00000187, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000208, 4'd1, 27'h00000127, 4'd14, 27'h000001cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001bf, 4'd7, 27'h00000089, 4'd2, 27'h00000053, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000390, 4'd8, 27'h00000374, 4'd5, 27'h00000365, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002ed, 4'd8, 27'h00000136, 4'd14, 27'h000003d0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002cf, 4'd13, 27'h00000132, 4'd3, 27'h0000035e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000000d6, 4'd11, 27'h00000164, 4'd5, 27'h000001a3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002b5, 4'd10, 27'h0000025b, 4'd10, 27'h000000cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000027d, 4'd1, 27'h00000108, 4'd0, 27'h00000128, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000311, 4'd3, 27'h000002cd, 4'd6, 27'h00000349, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000017f, 4'd0, 27'h0000029a, 4'd12, 27'h0000036a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001b1, 4'd7, 27'h00000219, 4'd4, 27'h0000013f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001b0, 4'd7, 27'h000001e0, 4'd5, 27'h00000367, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000082, 4'd8, 27'h00000330, 4'd10, 27'h00000007, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003f8, 4'd12, 27'h0000002e, 4'd4, 27'h000003ad, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000000e, 4'd11, 27'h00000289, 4'd5, 27'h0000032f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003b2, 4'd12, 27'h0000011f, 4'd14, 27'h00000024, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000a4, 4'd3, 27'h000000b9, 4'd2, 27'h00000311, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000df, 4'd1, 27'h00000187, 4'd5, 27'h000000d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000017d, 4'd4, 27'h000002b6, 4'd10, 27'h000002a0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001aa, 4'd6, 27'h00000319, 4'd3, 27'h000002eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002ed, 4'd8, 27'h000000ea, 4'd6, 27'h0000003b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000017e, 4'd5, 27'h00000390, 4'd13, 27'h00000263, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000af, 4'd12, 27'h000003d3, 4'd0, 27'h000000f0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003c6, 4'd12, 27'h000002a4, 4'd6, 27'h000002bd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000028f, 4'd10, 27'h00000256, 4'd11, 27'h0000030e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000080, 4'd2, 27'h00000395, 4'd2, 27'h00000326, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001c7, 4'd0, 27'h000003af, 4'd8, 27'h00000229, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000009e, 4'd0, 27'h0000005a, 4'd14, 27'h0000006c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000112, 4'd9, 27'h00000284, 4'd3, 27'h000001bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000374, 4'd7, 27'h000002ec, 4'd5, 27'h000003e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000245, 4'd6, 27'h0000024f, 4'd10, 27'h0000007d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000001, 4'd13, 27'h000003c0, 4'd3, 27'h0000035c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001bc, 4'd13, 27'h00000262, 4'd7, 27'h0000029c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000240, 4'd14, 27'h00000274, 4'd12, 27'h0000038f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000062, 4'd4, 27'h00000025, 4'd3, 27'h00000175, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000f1, 4'd4, 27'h00000025, 4'd8, 27'h000001a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000038b, 4'd2, 27'h000003bf, 4'd11, 27'h000002de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000175, 4'd5, 27'h00000240, 4'd3, 27'h000001af, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000003a, 4'd5, 27'h00000257, 4'd7, 27'h00000346, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001fd, 4'd9, 27'h000002ca, 4'd10, 27'h000003d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000001d2, 4'd14, 27'h000000c8, 4'd0, 27'h0000025a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000012d, 4'd12, 27'h0000011e, 4'd9, 27'h000000cf, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000338, 4'd13, 27'h00000302, 4'd12, 27'h000002ec, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000310, 4'd3, 27'h0000010e, 4'd4, 27'h000002fc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000027d, 4'd4, 27'h0000007d, 4'd8, 27'h0000012a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000296, 4'd1, 27'h00000297, 4'd11, 27'h00000122, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000140, 4'd5, 27'h0000026a, 4'd3, 27'h0000016d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003e4, 4'd7, 27'h0000036d, 4'd5, 27'h00000290, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000315, 4'd6, 27'h00000025, 4'd12, 27'h00000362, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003e1, 4'd13, 27'h00000144, 4'd1, 27'h00000043, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000039, 4'd14, 27'h00000379, 4'd9, 27'h000000e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000011e, 4'd10, 27'h00000340, 4'd13, 27'h00000110, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000021c, 4'd0, 27'h0000012d, 4'd2, 27'h00000126, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000265, 4'd0, 27'h000000a9, 4'd9, 27'h000000e1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000038f, 4'd0, 27'h00000314, 4'd13, 27'h000003a6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000011b, 4'd5, 27'h0000034c, 4'd3, 27'h00000057, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003c0, 4'd8, 27'h000001b7, 4'd8, 27'h000000cb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000027c, 4'd9, 27'h00000094, 4'd12, 27'h00000210, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000170, 4'd10, 27'h000000cb, 4'd3, 27'h000000df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000348, 4'd13, 27'h00000131, 4'd5, 27'h000000c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000001, 4'd10, 27'h00000357, 4'd14, 27'h0000010e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000020a, 4'd0, 27'h000003da, 4'd3, 27'h000001b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002e7, 4'd3, 27'h00000274, 4'd6, 27'h00000315, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000031b, 4'd3, 27'h0000029d, 4'd10, 27'h00000262, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000210, 4'd8, 27'h000003ef, 4'd2, 27'h00000052, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000ab, 4'd9, 27'h00000137, 4'd5, 27'h000001a9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001ab, 4'd7, 27'h00000124, 4'd12, 27'h000000b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000198, 4'd13, 27'h000001c6, 4'd4, 27'h00000101, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000003, 4'd13, 27'h0000005a, 4'd8, 27'h00000397, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000001c, 4'd11, 27'h000002d1, 4'd11, 27'h00000349, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000030c, 4'd2, 27'h000003c6, 4'd2, 27'h00000218, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000351, 4'd2, 27'h00000343, 4'd5, 27'h00000031, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000096, 4'd3, 27'h00000368, 4'd10, 27'h000001aa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000030c, 4'd6, 27'h00000144, 4'd0, 27'h00000182, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000277, 4'd9, 27'h000002cf, 4'd7, 27'h0000023c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000114, 4'd7, 27'h00000203, 4'd10, 27'h00000024, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000037e, 4'd12, 27'h000000e2, 4'd1, 27'h00000306, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002f0, 4'd14, 27'h000001d5, 4'd8, 27'h0000001b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000119, 4'd13, 27'h000000f3, 4'd11, 27'h000001c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001de, 4'd2, 27'h000000ca, 4'd1, 27'h000001b9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000244, 4'd1, 27'h00000365, 4'd9, 27'h000002bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000363, 4'd3, 27'h00000205, 4'd10, 27'h000000d5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000011d, 4'd8, 27'h000000f9, 4'd1, 27'h000003ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000304, 4'd8, 27'h0000011c, 4'd8, 27'h00000303, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000003d, 4'd6, 27'h000001ff, 4'd12, 27'h00000257, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000024e, 4'd12, 27'h00000263, 4'd4, 27'h000003eb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000144, 4'd14, 27'h00000061, 4'd9, 27'h000000fd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000017f, 4'd13, 27'h000002d3, 4'd13, 27'h000000f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000036c, 4'd0, 27'h0000013b, 4'd3, 27'h00000353, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000032d, 4'd1, 27'h000000f5, 4'd7, 27'h000002b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000027c, 4'd1, 27'h000001dd, 4'd12, 27'h000003d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000200, 4'd6, 27'h00000015, 4'd4, 27'h00000203, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000001d0, 4'd6, 27'h000002f7, 4'd5, 27'h00000130, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000247, 4'd5, 27'h00000146, 4'd14, 27'h000003c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001c4, 4'd12, 27'h0000000d, 4'd4, 27'h00000132, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000a0, 4'd13, 27'h0000010a, 4'd8, 27'h000003da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000203, 4'd14, 27'h0000034c, 4'd10, 27'h00000099, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000086, 4'd1, 27'h000001ea, 4'd2, 27'h0000000f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001da, 4'd3, 27'h00000370, 4'd6, 27'h000001c4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000384, 4'd2, 27'h00000372, 4'd13, 27'h000003de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000397, 4'd9, 27'h000001e8, 4'd1, 27'h00000287, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000230, 4'd9, 27'h0000016c, 4'd7, 27'h000000a6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000035e, 4'd9, 27'h000003db, 4'd10, 27'h00000065, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001a8, 4'd13, 27'h0000010d, 4'd1, 27'h0000034d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003a9, 4'd14, 27'h000000e3, 4'd8, 27'h00000315, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000128, 4'd12, 27'h00000006, 4'd13, 27'h0000035d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000065, 4'd0, 27'h000000b3, 4'd4, 27'h0000021b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001b4, 4'd1, 27'h00000327, 4'd6, 27'h0000017e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000370, 4'd2, 27'h00000164, 4'd12, 27'h000001de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003e4, 4'd6, 27'h000000df, 4'd4, 27'h00000145, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000180, 4'd5, 27'h00000194, 4'd6, 27'h0000015c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000370, 4'd9, 27'h00000179, 4'd10, 27'h000002ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000ca, 4'd12, 27'h00000016, 4'd4, 27'h00000192, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002fe, 4'd13, 27'h000001aa, 4'd9, 27'h000003f6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000355, 4'd12, 27'h000003d9, 4'd14, 27'h00000347, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000025d, 4'd4, 27'h000002f3, 4'd0, 27'h00000390, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000020, 4'd1, 27'h0000013a, 4'd8, 27'h00000024, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003dd, 4'd4, 27'h000000e4, 4'd12, 27'h0000035f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000003, 4'd8, 27'h000002bc, 4'd3, 27'h0000025c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000009f, 4'd7, 27'h00000160, 4'd7, 27'h0000023a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000027e, 4'd5, 27'h00000239, 4'd10, 27'h0000038c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002db, 4'd14, 27'h0000005d, 4'd4, 27'h0000020d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002f1, 4'd14, 27'h00000316, 4'd8, 27'h0000009f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c0, 4'd12, 27'h00000009, 4'd13, 27'h000002a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000150, 4'd1, 27'h00000060, 4'd0, 27'h00000314, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000020c, 4'd4, 27'h00000049, 4'd7, 27'h0000024f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003a1, 4'd2, 27'h0000000f, 4'd12, 27'h000001ea, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000024a, 4'd6, 27'h00000052, 4'd1, 27'h0000017d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000002a6, 4'd9, 27'h000003be, 4'd5, 27'h00000034, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000003e, 4'd8, 27'h000002f2, 4'd13, 27'h000000ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000035a, 4'd14, 27'h00000261, 4'd0, 27'h0000028a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002c2, 4'd10, 27'h000002fd, 4'd7, 27'h000003f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000028f, 4'd11, 27'h00000242, 4'd13, 27'h00000357, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000197, 4'd0, 27'h0000014b, 4'd2, 27'h00000003, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002a1, 4'd1, 27'h000002c2, 4'd6, 27'h00000068, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000003f, 4'd1, 27'h00000371, 4'd14, 27'h0000015f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000001bf, 4'd9, 27'h000000e2, 4'd0, 27'h000001eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000097, 4'd6, 27'h0000031b, 4'd6, 27'h000001c6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000109, 4'd5, 27'h00000300, 4'd12, 27'h000000c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000017d, 4'd11, 27'h00000146, 4'd4, 27'h00000169, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003d9, 4'd12, 27'h000001f2, 4'd7, 27'h000003d6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000113, 4'd12, 27'h000000a8, 4'd14, 27'h00000006, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000066, 4'd0, 27'h0000023c, 4'd4, 27'h00000060, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000011e, 4'd3, 27'h00000375, 4'd6, 27'h00000267, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000298, 4'd0, 27'h00000097, 4'd10, 27'h000001a1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002d4, 4'd6, 27'h00000363, 4'd4, 27'h00000390, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000068, 4'd5, 27'h000001f8, 4'd8, 27'h0000034b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000033f, 4'd8, 27'h0000018b, 4'd12, 27'h00000288, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000034e, 4'd10, 27'h00000336, 4'd2, 27'h000003bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000019e, 4'd10, 27'h0000012c, 4'd8, 27'h000000b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000070, 4'd11, 27'h0000018f, 4'd11, 27'h000001d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000003b9, 4'd4, 27'h000001d7, 4'd4, 27'h000003ed, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000361, 4'd0, 27'h0000035c, 4'd8, 27'h000003fa, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002a6, 4'd1, 27'h000001f2, 4'd13, 27'h000001c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003bb, 4'd9, 27'h00000271, 4'd1, 27'h0000030d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000081, 4'd7, 27'h000003ce, 4'd8, 27'h00000288, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002d8, 4'd5, 27'h000003f1, 4'd13, 27'h000003cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000051, 4'd12, 27'h00000234, 4'd2, 27'h00000044, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001fe, 4'd13, 27'h00000243, 4'd6, 27'h0000028b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001cd, 4'd14, 27'h0000032b, 4'd12, 27'h00000044, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000e1, 4'd2, 27'h00000122, 4'd4, 27'h000003e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001b9, 4'd2, 27'h00000164, 4'd8, 27'h00000167, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000339, 4'd1, 27'h0000008f, 4'd14, 27'h0000027d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001cb, 4'd8, 27'h00000123, 4'd3, 27'h00000090, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000106, 4'd9, 27'h0000026b, 4'd8, 27'h000001e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003a3, 4'd5, 27'h000000d9, 4'd10, 27'h00000364, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002a9, 4'd13, 27'h000000ce, 4'd4, 27'h000000e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000022, 4'd14, 27'h000002f8, 4'd6, 27'h00000025, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000025a, 4'd12, 27'h000002f2, 4'd12, 27'h000001c6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003df, 4'd3, 27'h000003f9, 4'd2, 27'h0000033f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000010c, 4'd1, 27'h00000071, 4'd5, 27'h000003cf, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000005d, 4'd1, 27'h00000004, 4'd14, 27'h00000359, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000004, 4'd6, 27'h00000067, 4'd1, 27'h00000053, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003db, 4'd6, 27'h000001e7, 4'd7, 27'h00000214, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002b1, 4'd7, 27'h0000010f, 4'd12, 27'h000003c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000058, 4'd12, 27'h00000245, 4'd4, 27'h000003aa, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003ae, 4'd11, 27'h00000028, 4'd5, 27'h0000008b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000106, 4'd14, 27'h00000095, 4'd11, 27'h000003e7, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000271, 4'd1, 27'h0000019a, 4'd2, 27'h000003cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001d3, 4'd4, 27'h000000e4, 4'd9, 27'h000003c2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002ef, 4'd1, 27'h00000279, 4'd14, 27'h00000012, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001ff, 4'd8, 27'h000003d5, 4'd2, 27'h0000030d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000014d, 4'd9, 27'h000001a4, 4'd5, 27'h00000308, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000029c, 4'd8, 27'h00000243, 4'd11, 27'h0000000e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000017f, 4'd11, 27'h00000311, 4'd1, 27'h000002bd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000037d, 4'd14, 27'h00000029, 4'd5, 27'h00000099, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000336, 4'd11, 27'h000000eb, 4'd12, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000015a, 4'd2, 27'h000001f9, 4'd4, 27'h000002ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000036, 4'd3, 27'h000001e0, 4'd9, 27'h00000315, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000302, 4'd4, 27'h000003b9, 4'd13, 27'h0000004a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003a8, 4'd9, 27'h0000018f, 4'd1, 27'h00000102, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002b6, 4'd8, 27'h00000026, 4'd7, 27'h000001f2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000014e, 4'd9, 27'h000001df, 4'd13, 27'h00000001, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000287, 4'd10, 27'h00000222, 4'd3, 27'h00000236, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003df, 4'd10, 27'h00000360, 4'd9, 27'h00000356, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000011a, 4'd10, 27'h000002d0, 4'd13, 27'h0000030d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000251, 4'd1, 27'h00000133, 4'd3, 27'h0000005d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000007, 4'd1, 27'h00000296, 4'd9, 27'h00000354, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000037a, 4'd3, 27'h000003eb, 4'd14, 27'h00000171, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002bf, 4'd8, 27'h00000123, 4'd4, 27'h00000359, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000108, 4'd9, 27'h00000029, 4'd6, 27'h000000b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003b3, 4'd8, 27'h000002e3, 4'd11, 27'h00000224, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000204, 4'd12, 27'h000001c7, 4'd2, 27'h000002a1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000025d, 4'd10, 27'h000001af, 4'd7, 27'h0000018a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000000f, 4'd11, 27'h000003f0, 4'd13, 27'h0000016e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000033a, 4'd3, 27'h0000028d, 4'd1, 27'h0000004a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000038a, 4'd3, 27'h00000110, 4'd6, 27'h000000ce, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001d0, 4'd2, 27'h00000280, 4'd12, 27'h0000016a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000367, 4'd5, 27'h00000194, 4'd2, 27'h000002b0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000088, 4'd5, 27'h0000033c, 4'd9, 27'h0000004d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000039a, 4'd6, 27'h000002a3, 4'd14, 27'h0000010e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000209, 4'd11, 27'h000002ea, 4'd2, 27'h0000011c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000002b7, 4'd11, 27'h0000025a, 4'd8, 27'h00000170, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000012d, 4'd13, 27'h00000004, 4'd14, 27'h0000023c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000163, 4'd0, 27'h00000078, 4'd1, 27'h0000018b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000000ed, 4'd0, 27'h000002da, 4'd9, 27'h000003a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000322, 4'd4, 27'h00000312, 4'd11, 27'h00000357, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003d2, 4'd7, 27'h00000386, 4'd1, 27'h000001a1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000a2, 4'd9, 27'h000002d7, 4'd8, 27'h000000af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000224, 4'd7, 27'h00000257, 4'd12, 27'h00000323, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002aa, 4'd10, 27'h000002f0, 4'd2, 27'h000001b2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003c3, 4'd11, 27'h00000223, 4'd7, 27'h00000142, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000286, 4'd10, 27'h000002ea, 4'd10, 27'h00000046, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000013, 4'd0, 27'h000002e8, 4'd0, 27'h0000009f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000c7, 4'd4, 27'h000001a3, 4'd5, 27'h00000049, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000135, 4'd2, 27'h00000137, 4'd10, 27'h0000022a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003a4, 4'd5, 27'h00000366, 4'd2, 27'h00000041, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000f8, 4'd5, 27'h00000372, 4'd6, 27'h00000125, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000366, 4'd9, 27'h000000c1, 4'd12, 27'h000003ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002f9, 4'd10, 27'h00000391, 4'd4, 27'h00000289, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000021d, 4'd11, 27'h000000fd, 4'd5, 27'h000003e6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000322, 4'd12, 27'h00000389, 4'd14, 27'h00000310, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003fa, 4'd4, 27'h000001bb, 4'd4, 27'h00000214, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000111, 4'd2, 27'h00000046, 4'd9, 27'h0000018e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000378, 4'd2, 27'h0000023a, 4'd14, 27'h00000347, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003da, 4'd9, 27'h000003c5, 4'd2, 27'h000002a0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002d8, 4'd6, 27'h000000e8, 4'd5, 27'h000003ef, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000026e, 4'd6, 27'h00000379, 4'd14, 27'h00000025, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000029f, 4'd10, 27'h0000035d, 4'd1, 27'h000003ed, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001d0, 4'd13, 27'h000003f5, 4'd9, 27'h00000339, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000147, 4'd11, 27'h000002e2, 4'd10, 27'h0000026f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003da, 4'd3, 27'h0000023e, 4'd4, 27'h000001a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000012b, 4'd4, 27'h000003d3, 4'd8, 27'h000000f5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000290, 4'd3, 27'h000001cb, 4'd10, 27'h00000383, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002e7, 4'd6, 27'h00000046, 4'd0, 27'h000003d1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000025c, 4'd7, 27'h000000c5, 4'd9, 27'h000002bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001c3, 4'd6, 27'h00000176, 4'd11, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000073, 4'd14, 27'h00000223, 4'd2, 27'h000002c1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001f3, 4'd14, 27'h000001de, 4'd9, 27'h00000036, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002a5, 4'd11, 27'h000003ae, 4'd13, 27'h00000344, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001b2, 4'd3, 27'h000000c2, 4'd2, 27'h0000000c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000018c, 4'd1, 27'h0000028d, 4'd8, 27'h00000007, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000000e5, 4'd1, 27'h0000025b, 4'd11, 27'h0000009f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000016b, 4'd9, 27'h00000339, 4'd4, 27'h0000030d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000011a, 4'd5, 27'h00000227, 4'd5, 27'h000001fc, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000000ed, 4'd8, 27'h000002f8, 4'd10, 27'h000001cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000306, 4'd10, 27'h00000108, 4'd0, 27'h00000117, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003c5, 4'd10, 27'h00000243, 4'd5, 27'h000002b1, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000045, 4'd10, 27'h000003b8, 4'd13, 27'h000003df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001fd, 4'd2, 27'h00000086, 4'd1, 27'h00000258, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000002b4, 4'd2, 27'h000002d6, 4'd9, 27'h00000268, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003cf, 4'd1, 27'h00000385, 4'd10, 27'h000001c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000038d, 4'd7, 27'h00000160, 4'd0, 27'h000002f9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000028a, 4'd5, 27'h00000027, 4'd7, 27'h00000350, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000165, 4'd9, 27'h000001dd, 4'd11, 27'h000001b0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000000ed, 4'd14, 27'h000000e0, 4'd3, 27'h0000005c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000232, 4'd10, 27'h000000c9, 4'd8, 27'h00000074, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000203, 4'd12, 27'h00000118, 4'd11, 27'h000001d6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000253, 4'd0, 27'h000002c8, 4'd4, 27'h000001e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000c9, 4'd4, 27'h0000038d, 4'd7, 27'h00000381, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002e2, 4'd3, 27'h0000021f, 4'd11, 27'h00000362, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002ef, 4'd9, 27'h000000cf, 4'd3, 27'h00000363, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003b7, 4'd6, 27'h00000386, 4'd6, 27'h00000302, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003cb, 4'd8, 27'h00000166, 4'd10, 27'h0000018d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000165, 4'd10, 27'h0000038b, 4'd0, 27'h000003a3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000020f, 4'd11, 27'h0000035d, 4'd8, 27'h000003e0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000178, 4'd10, 27'h00000267, 4'd13, 27'h000002d4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000059, 4'd0, 27'h000001da, 4'd2, 27'h00000009, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003b9, 4'd1, 27'h0000021a, 4'd6, 27'h0000035d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000019, 4'd3, 27'h00000217, 4'd11, 27'h00000067, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000032e, 4'd7, 27'h0000016c, 4'd1, 27'h00000370, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003c8, 4'd7, 27'h00000391, 4'd9, 27'h00000035, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003c7, 4'd8, 27'h000001a2, 4'd12, 27'h0000030b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000358, 4'd12, 27'h000000df, 4'd4, 27'h0000030c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000000bc, 4'd14, 27'h00000310, 4'd6, 27'h000000a3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002f0, 4'd13, 27'h00000172, 4'd10, 27'h000003c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000ca, 4'd3, 27'h00000054, 4'd1, 27'h00000363, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001e9, 4'd3, 27'h000000bb, 4'd6, 27'h000003cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000082, 4'd4, 27'h00000038, 4'd13, 27'h00000070, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001a7, 4'd6, 27'h00000160, 4'd2, 27'h000002ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000341, 4'd6, 27'h000002c3, 4'd5, 27'h000000df, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000362, 4'd7, 27'h000001b6, 4'd10, 27'h000000b8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000025, 4'd13, 27'h0000030c, 4'd3, 27'h00000292, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001a6, 4'd10, 27'h00000122, 4'd5, 27'h0000010c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000008, 4'd14, 27'h00000356, 4'd13, 27'h000000be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000021d, 4'd0, 27'h0000028f, 4'd2, 27'h00000358, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000328, 4'd4, 27'h000001f4, 4'd5, 27'h0000001e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000f6, 4'd3, 27'h00000145, 4'd14, 27'h0000005d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000335, 4'd9, 27'h00000021, 4'd0, 27'h00000067, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002ab, 4'd6, 27'h0000018b, 4'd8, 27'h000000cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000039b, 4'd7, 27'h00000117, 4'd12, 27'h000003ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001e4, 4'd10, 27'h00000056, 4'd2, 27'h000003e4, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002fe, 4'd11, 27'h000000f3, 4'd9, 27'h0000033b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000158, 4'd10, 27'h00000232, 4'd13, 27'h00000193, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000014e, 4'd2, 27'h000003d3, 4'd4, 27'h00000037, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001d5, 4'd0, 27'h000000cc, 4'd6, 27'h00000281, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000034e, 4'd1, 27'h00000317, 4'd13, 27'h000001e9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001b6, 4'd8, 27'h00000051, 4'd4, 27'h000000e9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000015, 4'd7, 27'h000000c5, 4'd7, 27'h000003a9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000010f, 4'd7, 27'h000002de, 4'd14, 27'h00000364, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000044, 4'd11, 27'h0000017d, 4'd2, 27'h000001ab, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000001f1, 4'd13, 27'h0000011f, 4'd8, 27'h0000000c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000025d, 4'd13, 27'h000003f9, 4'd11, 27'h00000252, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h0000002d, 4'd1, 27'h000002b4, 4'd1, 27'h00000166, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000340, 4'd0, 27'h00000105, 4'd8, 27'h000002ce, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000140, 4'd2, 27'h00000352, 4'd11, 27'h000001ee, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000015a, 4'd8, 27'h000003a9, 4'd3, 27'h000003a5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000184, 4'd9, 27'h000002e4, 4'd7, 27'h00000006, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000000f6, 4'd5, 27'h000002a5, 4'd11, 27'h0000014e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000244, 4'd14, 27'h000003f2, 4'd1, 27'h000003ae, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000024a, 4'd11, 27'h0000007a, 4'd9, 27'h00000079, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000003a7, 4'd14, 27'h000000f5, 4'd11, 27'h0000036d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000175, 4'd4, 27'h000003da, 4'd0, 27'h0000012d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002e1, 4'd2, 27'h00000143, 4'd9, 27'h0000013e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000033b, 4'd3, 27'h00000068, 4'd10, 27'h0000001c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000000ec, 4'd6, 27'h000001b2, 4'd2, 27'h00000375, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000372, 4'd7, 27'h000003a1, 4'd6, 27'h00000268, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003b8, 4'd5, 27'h00000103, 4'd11, 27'h00000238, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001d6, 4'd14, 27'h00000148, 4'd0, 27'h00000191, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000379, 4'd13, 27'h00000144, 4'd6, 27'h000001cc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000001f5, 4'd11, 27'h0000017c, 4'd10, 27'h000001af, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000014c, 4'd0, 27'h000002ab, 4'd3, 27'h000003bb, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000004e, 4'd2, 27'h00000381, 4'd9, 27'h00000071, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000003b8, 4'd2, 27'h00000209, 4'd11, 27'h00000222, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000020d, 4'd7, 27'h000001e3, 4'd3, 27'h000001ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000236, 4'd6, 27'h000003a8, 4'd6, 27'h00000176, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000203, 4'd6, 27'h00000252, 4'd10, 27'h00000047, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000024f, 4'd11, 27'h000002a2, 4'd1, 27'h000000da, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000003f8, 4'd10, 27'h0000026a, 4'd8, 27'h00000066, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000111, 4'd13, 27'h000000c7, 4'd13, 27'h00000261, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000295, 4'd1, 27'h00000259, 4'd3, 27'h0000011f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000034c, 4'd2, 27'h000000db, 4'd7, 27'h000001b3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000034a, 4'd1, 27'h00000014, 4'd10, 27'h000001b5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003eb, 4'd9, 27'h00000107, 4'd4, 27'h0000016d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000320, 4'd8, 27'h0000026c, 4'd9, 27'h00000142, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000173, 4'd6, 27'h00000168, 4'd11, 27'h000002ba, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000026, 4'd11, 27'h00000046, 4'd0, 27'h00000329, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000023e, 4'd13, 27'h000002ba, 4'd7, 27'h0000001c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000003cb, 4'd14, 27'h0000000a, 4'd11, 27'h000002c0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000070, 4'd1, 27'h0000032a, 4'd3, 27'h0000022d, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003ea, 4'd2, 27'h000002a8, 4'd7, 27'h000002cd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000016a, 4'd0, 27'h000001ea, 4'd14, 27'h00000140, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000039d, 4'd5, 27'h000003f5, 4'd0, 27'h000003a1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001ae, 4'd9, 27'h00000369, 4'd6, 27'h00000102, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000294, 4'd9, 27'h000002b0, 4'd12, 27'h00000355, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000036e, 4'd14, 27'h00000050, 4'd2, 27'h00000243, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003af, 4'd11, 27'h0000002e, 4'd5, 27'h0000018e, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000001b6, 4'd11, 27'h0000002d, 4'd11, 27'h000000bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001c7, 4'd2, 27'h00000055, 4'd2, 27'h00000386, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h000002b9, 4'd2, 27'h00000213, 4'd7, 27'h00000165, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000028f, 4'd3, 27'h00000089, 4'd14, 27'h000000b6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000145, 4'd6, 27'h0000028b, 4'd3, 27'h00000291, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000133, 4'd6, 27'h00000075, 4'd9, 27'h00000344, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000083, 4'd5, 27'h000003cf, 4'd11, 27'h00000226, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000086, 4'd13, 27'h0000024f, 4'd3, 27'h00000089, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000052, 4'd12, 27'h000002b6, 4'd8, 27'h0000027b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003d1, 4'd14, 27'h000002f6, 4'd12, 27'h00000176, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000000dc, 4'd2, 27'h00000138, 4'd3, 27'h000003fd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003fe, 4'd2, 27'h00000149, 4'd8, 27'h00000348, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000025f, 4'd2, 27'h00000208, 4'd14, 27'h0000030b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000192, 4'd8, 27'h0000035f, 4'd1, 27'h0000033d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h00000277, 4'd8, 27'h0000030b, 4'd5, 27'h000000a2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000204, 4'd9, 27'h00000250, 4'd10, 27'h000001fe, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h0000028c, 4'd10, 27'h000000eb, 4'd0, 27'h00000394, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000003e3, 4'd13, 27'h00000032, 4'd8, 27'h00000072, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000090, 4'd11, 27'h00000148, 4'd10, 27'h00000290, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000000a8, 4'd1, 27'h00000256, 4'd4, 27'h00000382, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000003fc, 4'd3, 27'h000002ce, 4'd8, 27'h00000329, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000326, 4'd3, 27'h00000173, 4'd14, 27'h000003d2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000031e, 4'd9, 27'h00000394, 4'd2, 27'h000000fe, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000339, 4'd9, 27'h00000159, 4'd8, 27'h00000102, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000059, 4'd9, 27'h000003fb, 4'd10, 27'h00000211, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003ac, 4'd10, 27'h000000d0, 4'd4, 27'h000001bb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000001ac, 4'd11, 27'h000001cf, 4'd5, 27'h000001f3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000028a, 4'd10, 27'h0000023e, 4'd10, 27'h00000101, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000064, 4'd1, 27'h00000327, 4'd4, 27'h00000316, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000024b, 4'd2, 27'h00000317, 4'd6, 27'h000001d0, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000004f, 4'd4, 27'h00000158, 4'd10, 27'h00000091, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000100, 4'd8, 27'h00000293, 4'd1, 27'h00000178, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001c2, 4'd7, 27'h00000041, 4'd8, 27'h000003e9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000039f, 4'd7, 27'h0000035a, 4'd10, 27'h00000343, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000010, 4'd12, 27'h000003a0, 4'd0, 27'h000003ce, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000189, 4'd11, 27'h000000ec, 4'd6, 27'h0000006b, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000359, 4'd12, 27'h0000010e, 4'd12, 27'h00000117, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000267, 4'd1, 27'h000003fe, 4'd1, 27'h00000102, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001b0, 4'd4, 27'h000002c3, 4'd6, 27'h00000184, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h0000009e, 4'd0, 27'h000001e9, 4'd10, 27'h0000025d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000ee, 4'd6, 27'h000001e6, 4'd4, 27'h00000185, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000031c, 4'd8, 27'h000002fb, 4'd5, 27'h00000314, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002b0, 4'd9, 27'h000003fe, 4'd10, 27'h000001e3, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000001b8, 4'd13, 27'h00000131, 4'd3, 27'h00000265, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000271, 4'd14, 27'h00000176, 4'd9, 27'h00000243, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000336, 4'd11, 27'h000003b6, 4'd11, 27'h000001ee, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003da, 4'd4, 27'h0000032d, 4'd1, 27'h00000021, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000032a, 4'd2, 27'h00000100, 4'd5, 27'h000000dd, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000000b, 4'd4, 27'h0000031d, 4'd11, 27'h00000366, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000001a7, 4'd9, 27'h0000033a, 4'd1, 27'h00000268, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000002cf, 4'd6, 27'h00000227, 4'd7, 27'h00000135, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000044, 4'd7, 27'h00000207, 4'd10, 27'h000002c3, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000041, 4'd11, 27'h000002cf, 4'd0, 27'h000003b2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000226, 4'd10, 27'h000000be, 4'd9, 27'h000002db, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000334, 4'd11, 27'h0000007a, 4'd10, 27'h00000049, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h0000034e, 4'd2, 27'h0000028d, 4'd0, 27'h00000225, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000367, 4'd4, 27'h000002ab, 4'd6, 27'h00000224, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000346, 4'd2, 27'h00000031, 4'd10, 27'h000000c9, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000000e9, 4'd8, 27'h000001ac, 4'd0, 27'h000001f5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000090, 4'd8, 27'h000000df, 4'd6, 27'h0000015f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000009e, 4'd7, 27'h00000315, 4'd13, 27'h00000086, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000002aa, 4'd10, 27'h00000012, 4'd3, 27'h00000171, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h000001fa, 4'd12, 27'h00000284, 4'd6, 27'h000000f8, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000239, 4'd10, 27'h000002e7, 4'd11, 27'h000002be, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h000001cd, 4'd1, 27'h0000030c, 4'd3, 27'h0000014e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000216, 4'd0, 27'h00000396, 4'd8, 27'h00000283, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ce, 4'd7, 27'h0000034d, 4'd1, 27'h00000049, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000023d, 4'd8, 27'h000002b6, 4'd7, 27'h00000151, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000002fa, 4'd8, 27'h0000029a, 4'd12, 27'h00000054, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000003b0, 4'd12, 27'h000002a9, 4'd3, 27'h000001d4, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000162, 4'd14, 27'h000002e6, 4'd6, 27'h000003a5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h0000039f, 4'd13, 27'h00000259, 4'd12, 27'h000000e2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h0000001f, 4'd3, 27'h000003b6, 4'd1, 27'h000001ec, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000078, 4'd2, 27'h0000012a, 4'd7, 27'h00000069, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h000003bf, 4'd0, 27'h00000012, 4'd13, 27'h000002f6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000279, 4'd6, 27'h00000173, 4'd4, 27'h00000320, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002cc, 4'd5, 27'h0000010f, 4'd9, 27'h00000153, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h0000030e, 4'd9, 27'h000002dd, 4'd10, 27'h000003e7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000048, 4'd11, 27'h00000316, 4'd4, 27'h00000359, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000003bb, 4'd10, 27'h000000c0, 4'd9, 27'h00000172, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003e1, 4'd14, 27'h0000021e, 4'd10, 27'h0000031a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000a5, 4'd0, 27'h000001d5, 4'd2, 27'h000003de, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000000ae, 4'd4, 27'h000001c7, 4'd8, 27'h000000d2, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000016f, 4'd4, 27'h00000126, 4'd13, 27'h00000308, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000002ac, 4'd9, 27'h0000002c, 4'd3, 27'h000003bc, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000185, 4'd6, 27'h000001f2, 4'd6, 27'h0000033a, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000005, 4'd9, 27'h000002f1, 4'd14, 27'h00000261, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000003d2, 4'd13, 27'h000003bb, 4'd0, 27'h000001c1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h00000085, 4'd11, 27'h000002d5, 4'd5, 27'h000000ab, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003c5, 4'd13, 27'h000002cc, 4'd13, 27'h0000011c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h000001a9, 4'd2, 27'h0000023e, 4'd3, 27'h0000018e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000265, 4'd1, 27'h0000008f, 4'd6, 27'h0000001c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001ca, 4'd6, 27'h0000003c, 4'd3, 27'h00000280, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000b7, 4'd7, 27'h0000002a, 4'd8, 27'h00000221, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000002ab, 4'd6, 27'h00000255, 4'd14, 27'h000002c9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000303, 4'd10, 27'h00000135, 4'd2, 27'h00000356, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd4, 27'h00000216, 4'd14, 27'h000002fc, 4'd6, 27'h00000111, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000041, 4'd4, 27'h00000213, 4'd3, 27'h00000077, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000162, 4'd2, 27'h000003e3, 4'd5, 27'h00000258, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000223, 4'd2, 27'h0000036d, 4'd10, 27'h00000027, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000003b2, 4'd6, 27'h00000086, 4'd3, 27'h0000037c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000119, 4'd7, 27'h00000066, 4'd9, 27'h000000f6, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000015b, 4'd7, 27'h00000174, 4'd14, 27'h000000b0, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000362, 4'd11, 27'h000002d1, 4'd1, 27'h000002ac, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000cf, 4'd14, 27'h000001c9, 4'd6, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002a9, 4'd11, 27'h000003b1, 4'd12, 27'h0000010f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000010, 4'd3, 27'h000003c0, 4'd1, 27'h00000122, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000022a, 4'd0, 27'h000002fb, 4'd6, 27'h00000109, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000003c1, 4'd3, 27'h0000029d, 4'd12, 27'h000000db, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000196, 4'd7, 27'h000001e7, 4'd1, 27'h00000324, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000391, 4'd9, 27'h0000010f, 4'd9, 27'h00000098, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd10, 27'h000001ed, 4'd5, 27'h0000000d, 4'd13, 27'h00000175, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h0000028b, 4'd13, 27'h000003c3, 4'd1, 27'h000000de, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000338, 4'd14, 27'h00000119, 4'd5, 27'h0000005f, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000001f, 4'd12, 27'h0000010a, 4'd11, 27'h0000027f, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000266, 4'd2, 27'h00000309, 4'd1, 27'h00000366, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000311, 4'd2, 27'h000003cc, 4'd5, 27'h00000100, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000398, 4'd5, 27'h000003fd, 4'd1, 27'h00000111, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h0000016e, 4'd8, 27'h0000031e, 4'd5, 27'h0000006c, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001c2, 4'd9, 27'h0000034e, 4'd10, 27'h000000c8, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000047, 4'd14, 27'h000001b7, 4'd1, 27'h00000266, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h00000244, 4'd14, 27'h00000347, 4'd5, 27'h0000020c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002f2, 4'd2, 27'h00000224, 4'd0, 27'h00000295, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h00000155, 4'd3, 27'h000001e5, 4'd7, 27'h00000345, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000290, 4'd1, 27'h000000b1, 4'd14, 27'h000003c5, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000002a5, 4'd7, 27'h00000283, 4'd4, 27'h00000262, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h000002c7, 4'd6, 27'h000002bc, 4'd7, 27'h00000163, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h00000212, 4'd5, 27'h000002d4, 4'd11, 27'h00000139, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000002c8, 4'd13, 27'h00000028, 4'd2, 27'h0000002a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003f8, 4'd12, 27'h000000b2, 4'd5, 27'h000002b7, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd6, 27'h00000308, 4'd11, 27'h000000e4, 4'd10, 27'h0000015a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002cd, 4'd3, 27'h000001bd, 4'd1, 27'h00000107, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h0000032f, 4'd2, 27'h000000b3, 4'd8, 27'h000000fe, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000103, 4'd4, 27'h00000307, 4'd10, 27'h000001b1, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002f2, 4'd6, 27'h0000014e, 4'd2, 27'h00000083, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h00000249, 4'd7, 27'h000000cc, 4'd7, 27'h00000200, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h000002a4, 4'd6, 27'h000001e3, 4'd12, 27'h00000001, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000015e, 4'd14, 27'h00000086, 4'd1, 27'h000003eb, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000034, 4'd12, 27'h000001e2, 4'd5, 27'h00000375, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000018f, 4'd13, 27'h00000174, 4'd10, 27'h000001f2, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000bb, 4'd3, 27'h000003d4, 4'd2, 27'h000002e9, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000000f5, 4'd2, 27'h00000051, 4'd8, 27'h000000d5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h000001f0, 4'd7, 27'h000003b6, 4'd4, 27'h000002ac, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd2, 27'h00000245, 4'd9, 27'h00000354, 4'd5, 27'h00000389, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd1, 27'h000001da, 4'd9, 27'h000001f1, 4'd13, 27'h000002cd, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd3, 27'h00000342, 4'd12, 27'h00000271, 4'd3, 27'h00000373, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd0, 27'h000000ed, 4'd12, 27'h00000146, 4'd5, 27'h00000131, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h000003d9, 4'd0, 27'h0000033d, 4'd1, 27'h0000008d, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h0000033f, 4'd3, 27'h000003c7, 4'd9, 27'h0000001e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd7, 27'h0000025c, 4'd3, 27'h0000034e, 4'd11, 27'h00000113, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h000002e5, 4'd6, 27'h00000253, 4'd0, 27'h00000211, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h000000fc, 4'd8, 27'h0000031e, 4'd12, 27'h000001da, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd8, 27'h0000004d, 4'd12, 27'h0000018d, 4'd2, 27'h00000125, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd5, 27'h00000228, 4'd13, 27'h00000201, 4'd5, 27'h00000043, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd9, 27'h00000358, 4'd14, 27'h00000192, 4'd11, 27'h00000388, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000168, 4'd1, 27'h000001d4, 4'd0, 27'h000002c5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000003a8, 4'd2, 27'h000001bb, 4'd5, 27'h0000003a, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000023c, 4'd2, 27'h00000175, 4'd14, 27'h000001e5, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h00000173, 4'd8, 27'h000000d0, 4'd4, 27'h000000b6, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h000002d0, 4'd9, 27'h0000018a, 4'd5, 27'h0000021c, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd12, 27'h00000004, 4'd7, 27'h0000011f, 4'd14, 27'h0000016e, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd14, 27'h0000000a, 4'd12, 27'h000002f3, 4'd0, 27'h00000225, 32'h00000400,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd13, 27'h0000008e, 4'd14, 27'h00000057, 4'd5, 27'h0000010b, 32'hfffffc00,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd0,  4'd0, 27'h00000000, 4'd0, 27'h00000000, 4'd0, 27'h00000000, 32'h00000000,
  1'd1,  4'd11, 27'h00000097, 4'd11, 27'h00000177, 4'd10, 27'h000000b9, 32'h00000400};
