-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
IW/DcW6CbkGF+f2xGdKiMTNz851TXsWVVJXXzI2a2F6wDJ5OWaBrjZdiUwYOf3wc
L9UGKkEk5TK4og3nnXG2UyamclXJ94nyPf2mRUmlI7GYJxoskpEaU1815sI/lPM6
R420BAqbufgzAF54ZP35QuKmMKimqgudTp1YghWoZcc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1012)

`protect DATA_BLOCK
QQb5rt+z5Ir6N+kvCAa/Jz3ABgqz42NnJRSPPHFOV8soefkhM1mosM4MjAkGwpfO
5PA6U9TatmFedqLl0BgJlyNISZtgUEFsItsWq81ms3hqh3Zg3kJ0cQ5RIf7aOBtS
FEC5qs0YUWrTTl6GJZzoCkOCLbiWT3yN+WpL6aZLXzMtu76911uymd2wPbuCURKC
qZNfYA6nNnJXqFKTFVlZa+eCKvmmAQLNxv4rCx8xTHrnEDXzZIBErdfZFZJaTMwu
dbwrayd/ss/E4xEgNDju469TK6A/G72zFSsm/sqYO5VI3AA/qN9Lyp8W/CCR1jYN
p1o9Drdetr6hQjhB246rKMFF/rV04Vojq99MudkTJEHlVoOrqWjf9WUGnsiCoimg
BeC3no3A4WUAk2Nac3OjEO2yBkjQ/+mqIw+DOFHfYu47KAWOJk5mjkuLQqctMEs6
x8v6UoQZvp0oT1tmYOZ17cLTsSNjqcjd145FOYveUIDfe7a78zWDmvO2W6wl/Kxk
P3oXbtXkKtaqAnVBXxXXvg6qm5ptlYgJ6r4i9+bI2BBDWUnfCpCUKYfCghDynraW
yFt64D6ID15ueILlmKXgr79H3K4wfx2gmsVC+VkWgFq04n5BLg3rCTpcf0Pm513M
TOKWhyVHplSXbnOLOUZRflIgBCk3lKPyELTqNzh7w/dY2bE6vSx4vi78ASknwfT7
hKufQ06UacgfB4ZCK1JmjT7XfJ+iYZwPImIPrR1xqaTFgdVU2/sdR/Q+qPxglsEI
D+Ud+NJg5MGBboKWe0zesbHjecXj/r3BnN9tPB120dhb908+yLb0TG0AZCxunL2U
OiUyD7ObEpRnHcQn7IzOt9vSFhTeuEs5xuG2W9lV/a+fdIb1bH1bxe1zGrQ0zLkj
H+Mthvm+6Pd1yjbdt1GixUAk+WTC/lxROst526B15uDemF4qbem8MJX+13lrGIm7
/fKtGt6S09KNLiwzm2HgdasykPX65LTwsIjCqVoHfLqMyEWwwyV0z5XokpKGdQB1
iuiy+HPPL9hT7PArCLT5QW6P2k733nn9lMNgNKt+QfDiJaVM1zN/Zh/D0TJP6s1t
a6kNkJ5+0+Xzg3oTlBw52/av5guD0b+v8kQFw0GvOOYyFhJyRjGm1Dccg4FJ167n
LUwkIUJup6m/JrgUClCugVK1YIkQF9+KY5R160fgBQsa+Xuv2HUzsQrbQE/3Cyls
iqPo2ceRsX39azZUpADezs7MS4Fofws1y3vsZ8F4LGU/9xpNZxmaS7WdXfWMAe2C
BxtZ4Js/Dmbwm/37ktS7LJizN9LoCVihnTC2YqIyeSD1CTC3OApNnq0JIIJDL8uz
fNkA1ozPEk2pU3s7EwPJopgIVFdz4ecc9Qj3RJWy9Ow=
`protect END_PROTECTED