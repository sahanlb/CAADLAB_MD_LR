-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
L6J7DB34Z/+IPFD3K24gST7gqVj764MYOZ7shqCiMkF8in8n9ISLEu5p3h0O3vuG
Zers/N2aMHfu2EF7tOkToCC9kyuNH+ZOKIQO3IPIjH/naDf3Vcd4dNtibTuA7cFr
cmQyQQ0neW3P0jeQLYUuAXg2kaWx3xPsOHaIl9RRGEi7TRGa/nhnWg==
--pragma protect end_key_block
--pragma protect digest_block
XjB1P1G34tr1T00fF51h6Mhhp+Y=
--pragma protect end_digest_block
--pragma protect data_block
4K0Gz7MYbHCr++8mRFqG3m2xxR4O2BdiGMqjcgnzFt/MMNs8dMsIyIgb9Al+i0Uj
4rMbUtenDIJ2M0KW/+Q+nlyxQZbTte+rulbuSAX8F1qEHs9y82FvvtyhDsYvE2wo
x42G0T4gM4OK9Ob3QUYcmpijuEyGdSW/HBrA2h8XS14jSdSDEUqyxgaFrMxoAg7x
1Z9PWe+wXbpcpmtikbIRFmB8on7zmmRbXy+SA/OJx0255VG6PkWbBXsBzuIm0NjZ
4KG1xUeF3EXYaJq3L5RjhFsi8PehJKxd/anYhWB28tLIXmdTmhAROmddthE3HeMF
E0x3S2gmzLmU46aofnJew3+A0NdQxrLehdBjr89UyYQhQ1DQLDOE62RZzMw8Beit
HYWwRyQKmu2jIWLkaq1pY+Jw98R24P3mOi7SKvPT+sA34QzvrXDc3aPGoWIvn050
jmV+YyA/5ZR1tRhLGs2Xz22YdsDSkZ3dDJU72PeiVA016X7vb/i0HB1xJfVe7jb1
fHjGXR/V2zYDOK1EEFhUyubm+M/wWS5sNINyMp2BfEfhQ5wSNFsJwQpOaL5FmwAW
LQWHXlDjq6CHzWygkKORNandqF2FQAetzUZFb6KsF+UMYATUSRjOV42qvJHEmFg6
5g5ufhsE5WfGX9661HrRUAspfjHEDG2R2LFzpYYjA/6qUG5wvUJnb98cYQb8TTdR
kpKnlgxY4BAl0TVJQswS2De0vpEho4ERC0dneCnxvMFdwQzU7mppwbdHVaQRZAzP
4AKD5RXFdrUavEv5fBpGzz1Fq1mMSWhfxXIBO1SYCRnkKMh1Lh0OBiQ+ebDG53lB
PFgzFJE0SHL5VcLqIbQllYvZo8KvsP3c9hWPnyOJTZBmwD5Ks0CiseGAzvLqoeLK
X1qGy+PLBYMAFQoc4Mz3Idw2ZCiQyAOcPY+FKr4T06l3pbaC9rjA+OdS9q2mRNk8
/vigKB4uKQcLhyePdeEyoKEDhimzq8sX4sWfmb6E14BT1XBS62rPkIOcDojroWxK
pMOo4Mc8enDN+zoBbDQIRiMI99kQtPlsSsYiHxvLkXsYHIay0rkUCAWGo7RQRyUB
uJNWBqI3EMxuKDI8wkpd8bZakkelxt0xl/BBA1Bn6ylysJGcLGG7o/KpdR8n661E
F6TxycocKTh4QgQa6pJV3gUpaL8aphB+3H3fZ1h5mRBweDnqcQB2amN38t47vMFU
DtQmbTxOAD7xygf4+9qz3yAjMkV2iGe3avoLg5nf+8PeS20xfz+igQ0xchXVVup2
Y7fzub56vwiqBxdr3j1hT4R7dZiGlGnBHY6K4woP1EdUTLDW7yAuHTatYqFnxTEB
EynZ/e9DFGcEqh1q92ICxUfIljQd8yFd4u4S0eCnQ07LIqy5GR+YwuJZKi3kJf5k
zTWSeTZsf0NkwbyLCChgzeBuJLG3ToXBN9zwMN9rS73ravge7hLZ4IjlK4XojNX4
eQZgKJZpB8z6K+7jU8dUwbE7KnQnIifgPhQSLwUDn9JI8L1YF6COxkXLmiBxZZr1
Yn2GHzVxH+RZODavFfRYb99D2ZMcWyiZ4qYbM+DysPXe/RKDQqG4e20C4u1VDi46
3q2iHHgcZF+dZZVVNOt4KDSjHVMCBzNlFIIf4NOgruVrjZGTRGz1bWgjYaECE9Kp
HW5VVyEEdv3r4O1OaOsN5W0Qs3DN7z2qyGbkkfPXtJD9QQXOYDz69zi185F41K8v
Id0LmaXUun8mih50rpn0GfRe+6OApDgN7IIz7nSYBBz6FidUKL3aBfiUN2NLI511
8JiSTTObSjRuRgzmIl8P8UecYNztxnIQ77ItXWp7B421idw5McYdZ5qDlVwGyeGK
qD5eUyjhfmayjVVXUZRjZPhE63+3EV1M2WLja2VH0hPVcWEgCaeYKYDAHGGJc+hB
1zqBpdzi+R0nzmrvNvbMe1MjGKremSm8hR27NSg519gl3Gqu3vtbl/vqf9BB4vJy
t+aXLfvP/x8qCVBXufsi2BBssOYzNyDFNUyj2UIJM57ME/SHcF70yMENsUDjHjyI
gWi9oOVNxJB2Oitjao6hKCCrLf9sDGwQN2knYM00kYIJ7txZ41IlxBgasTQpR5Az
NeQ9/riLLkd8eYHwWyo0T6Y/f6WX1q7JlNrKxdh37Fyh4tmUqgcGda3AfC54FfuX
F8IpilFH6xSSiwWDaRhBouyQZqXQ0UMT4srWk3F5gOsenx+jcLkstGRCzM5rhj7X
3jI4umEJ2Hq9zEjQydIEMrpbuUwWggPWB7iqk1lXW6XlmJYUTt9m1UwqStQINyUX
8rZe14+/zUYK5cZVaN/oZ263ecXlQvWV3ZzvrOATHXE7gee6sHsViC718r6ZiRa/
Y/b+QpQa5wW+M6Jv6aYishUGdCotq3DmEkUBhakHuoDJnP2MVyzC9tuH99VWc/iV
FD/jXMQx6d3VpZfC1UqFGczS57ro4VbpFaoFVKi8E9tav/6VpI+b7EmDFtUnHzKz
4o76g+h9QJdm1TcSbzTA8NlDqokfMHnmkK0SmSwudyVVIDWHjkgFHdR6A3saSyKA
DnKsSrma2fNjNvC3UZ3avvOqgY+vwsJ9oceZMpJjni+C9wmUmHeW4WXWLQdGLtTU
ZZbwzZmzyGPtSWMJgZlCBYpjv6vZblNIrHX+VPHMe77Kqfg1aFSyNToAmIbnNxEK
evJlvt70+dzo7KD+GarI1eVrHYJikPIUV4isPT421pVRz51ommOKnwvOSlqymQHj
ibfRWx8TOMB5poDvxbQ2OU2GnecM+ub/Ta5aMoq71x84LqSNQAt54EJtk6i8V6zS
JzCzDVEBCWdOnSnEh8AzGssMCKsrK3+lO01XO6d2YvdsEpvM6EHke6u1VZktgLeu
Kx8T4sYFbM1yODWaiNXgk6O5EoiK7IxRhSdpDLozLbF2hvlAIV9hfiznjzvMsdL0
1D4v9q2YQhQH4soUamHInAJDmzY79qWXHHq9D+1tD8qvQBvQSVDqdVYNYdTv80jk
GMkjUpGwX+/7W0bCePLtF1Wh6XPoKR3rdOs9fwoQjLlc9Hioxi46g72ZwgEbdMrn
nGTaImPpy9EqDBo99iA5Mrg2NAWMluLK9+kolBsWEJGpJS5XO20cdhb1UkOymjGh
/YfgYIakSESGRShgJEXc6NYGtteGNLIuBHzcMZUD/lRQtqufGzEqKdjwVPDHyui2
CCo1PEaiReYRrP+X5yKZnIrDvbgzrmtNHwdE8DQ+h5VItLaXxCiRHuZSEdb/Tl1W
5322HBnoL80qOutitGwjLICpWzOPcXHPU1MLzjStBjqtiigxv/FN5w7JNqjq4un3
G/kvkWUZoJCnFpAI9VzRfV6KObegFa4iU07/w9fhJPdSZ0zoxXr2e0+CpwkOjY6I
hwPaAQY+GxvAkUvI0KIaizZ37ZTtsu4E26WxgrhPBJdo0WPyCTFm+gSFh4KOo9+z
J08curNxuOTvr4FvVhmj5dmkgS+yMupI11U98iXp2uI68OQWn9yBnXOQXTsonSGY
LTN1RNOtLrXJfVXbgb4eO30hD2rWSctbvrBAItAWyPs9QahML+uJngahRILt8QHr
LfQ8huHk9C4lpq2OigH3iE4RBLX3yeTa2BqNIyKy/tZ39NTtK+wszBOfYV4O7dR0
mKHy4LSmDrcO2oEOczFUskXK4LO8kvkZZ8psPcz2tku4xCFp5uxlHRvqwE/5gsM9
OxFUkSuRd9HzYlsc0W9iiYpSNL8l3rHQCV4HPTpH9DSyMV570tYGGpLcPItt8uGE
+nwaP9YjNvON3QWuhSFNPIUGkWBC0nQWmuKy+qpQpxGNwT1i9sYOspyk+vSudkNd
TnFoB1JJYrDaHSveuwtcc3mBQljdNQmAGjx5n6obytmdP7jhi8pFQulKY5UpBb4J
Ra6INMnkBxxO3VJ+PdmtzXo6D59xdcGlZJlH6fpmspLmSfMMyXq4JGHEPqj/y+l4
2YNvXByvWOYuwdWLa3kzs2+8ONO4HdX0qYAE3jngG9N1TIbc0bSeS+GRSo1AG3fv
+3C8MqR7cnAPLjtMwo1X4F4r4g+dDngDTN0/b0T6aX2OkQDKRsvX8xfvvFMsGZ1d
um1Ib6GKT7v5JpDun8c8q/m+GZtci+DshuSLCSGlju0m6ErKRU7J6JwKvL4MMG9x
RI5xSQn/b6+myyUOoZT3SgHJQ0UVar4g7WUvwEzNP8ktHPPkr52a0YBWL31yNdb5
vlVXqrSwm2cxVYCIXQJa9UmxlyE3CGJCoZJMb9t3WDpK7OoKj2t2KyyofVqKusI+
SZjjCGRbohgzJxx4y5vI92JEJH4D9+eU5WZ4Hu0qqC39/CXmK0GR2KZ3eLkRwTSy
8M0VolOmpwwrcEqIViel4ew6A7a0R4ICDT2sB2SPVyoth86L9q/YJj8Ogc/lHKre
r3Jc6YGh1dpCyMP0jxxei2LWZ16hfzfU0h+haDuTzpOw1KFjzXadrynPM8VhTYsE
CH3oZ0WSNWyoNNOjBR8juS9l3pRRZLm7j2Khp1VTgN5ZNjT8CP9gIiYA6wIuzO5X
6xnosRnfwfawRvipLxCRHnktOxcc+5SoJpG1iuRHh6L+4h/ZkJiPGqKGCmIx2/xr
B5MBD68yPJF7hBWiF4aK0dKADro8M7sLNet3VnUQqKY2lZANxtiWxQw71D5bCQ//
A5rCFTCLhcZJHlOVA1AfpiKBe51Zotdp8k6XdAgCYQopltI3HdrxFLi0vbeY/R0u
yHBBhbyF10TuA3Icz4WHEJpw6y4QEK/sqhcuwRaZzthotn8F7Sy2Qjw7MIp6Dxfy
OL3hoy4CXoGGdVMgQjBKC8r6JaenNo2AezBOE5/Idx5E//7CB+hRVIzW+25W7sD2
k2pTGwGLCDxsCSGLrLlIUutICNXDLwb+wKm9hiNPkBB5HLpl08MJn4Sz/yrlm4+g
Qu0QD+eXG5teDYoIgNDRwo07OTyjAk5pleB4hrpJ83WTq5IKIFPTZ0jvIg+et7F7
y0JhnWJ7hk/q2whVnQnJ1+557A78UI1nTSy3rKQ48Qj+z8D4b3OyJQFbuTNGXHRA
DoGkVDwWMO5YKloBSPaGjq2hZHHBbahdTO5DvHTgUgU770kpjSkgJ0Bk3m0Xeo/E
7EBabg7MxmdDsNCDyYnSVdZJROSt18x0RlAWXBEc7YMigTfJZzpeaZ/bZm1NIeej
Fi9r9IXtGXvo+hmK7oF4NqZcBs5lzgiSWZbAyiHh8UhnQTG2+vA80aOPiwwdoUHg
SB5yZ/g2knP4xj5B1xc16wjjOgDBleBEaNaXwSxXvUS1l4sAI0WTonUesO1/NFKA
VdeWbe2YjEDWtft9MxgPsrE9CZp8a0qVVPcRUYZkzK7cvlhe4jxVXxAtK1qOIWkn
NgVnu/tWC/KrM5yjjIyFW5w2soeNko2vhJE4RNaDJoEZrOYSckJVMR+GpLfCYDdz
/BpDWimFXTxz0duoS6Ddr0QOQBs3LcwDFxhqdjHC03i0q8pGfK5IVp9uKnQMlBTW
LANyu17F1IzHLDvapcReqZrG/hG23AZKEgKvntRL3nv0GM6zjYY+4v5Kz/GCZXJ5
CF62DIUQzYVqXGqbByW4XYBzO0PVt102w4iywQewhvRDRxzQeOwotetX+6WZawgm
3i5X4NHgjMWbBVR9i+olgd1p13BDfXxZPeaB1hFPtMfOCGV5xvjjpRrAT1YodgLc
DbH2WLw/+1w6xOF3ONlAeL12qJ9aFEJ6JLMc3czKEwgcQInJtDUSmpW+YIfkqrf4
3ZgweSiQqviqfH5KWuOaZ2XoLLzqSX/G6L3n6/X3UMzLf/ksRVlfEjoNR/U4etJn
ZU0Y3or1Ff6k05khu9ltfIjSas3TV1hIjlrHNcv0PtaGMGar0iJr74VDRd0pdvpI
gXA8oCyPLrsyr8GlUfEzbbZq/54tUGXmp3xDWlPJrgsqRRIWUMvsKIdWk+gPW2Cx
MnJ12FK1+SQvtGNTsvrzoNc8kmCVUlgRTl/fRGmKDHZAsS51uzMhu8JNoCAtQCMD
dw5E4dqCzNHoxMhTW6dAgsaVtgfamqm0hEkY8FL8uDDzXN7vByzejbA1wglsyb4X
tC5xe3djwiWV5RjpqafmCuTAp1yTZyt2mXL50nOGCHlFJTDqdlc/WXs8if1+zgBY
YL3dHbI7fDwRIsEQKRcyg19zbRtf/12LPTR8KVA9AX2lBioDZRzm5z7iIE6G++JL
rBQTL1gb21I9u9FTnjM1WjSKNfyV2xFZMEuZL3mjAmSphNuSRAdELPaTQ/htPziT
Dvu+5OTqei/2pVG72rXuq/zpW7xAxeTjgE1M2EPhEdmBvgFrkXbcjaZg24F5du36
EKhACKw2CYQ/2c40QEPxgHdJgCGt89xSuNI2VB9ky2XZw5e8Yqv3t/t3NeDie2Ew
tPktmUvTNoERW1ddkX/rE/o9B6Rhl2B6rx9kzF55llTAIdHcSNjSqfm5Y1cq8Jof
hF80QAX65ZtBr07VVEnFFeKjsRvS1Ju7fy9YtluPcx34+CYwQUJvdICpBU1mB2Py
BKL2peUryE1oD4WnYADdU6iV3uZ86hDmPSzZudkkoSrgSywXw2HLfOa2UoVe5HWc
GGizjEfExxpsG6VAQvQSM+NbU1/vL7J6vL/5mEUiZhsWhwzxgY43O1OMIy/CJASB
QvcPuBbhShGl+xZGOe2qJwatvqz50yPF8hxIhpQerzOncnNZDq4olS3J15sMs4bi
3eBxQRlHDRm4L6Nm4kAiexJDwzZbnP+rPUYd7SoMS73+6AafoFU7i84I21uepynD
W3fHiSV9le+Up1f1E7MHKmIODzRHuLZKREk8d3S6UIvnfZxb8DRAWaVbpSasPjgM
IEWvIJhPPG6cFrEiXHAPaRr52D4TwnUca7UUnIpxmPWR+TRDBN4LdS4FJLc60+op
hgPafrvlgMrS3QBQXZ4f3OPpPyeDdvQYcXOdrOXTbfyglmOO15btLYmbvjtTgH6l
kEZfCaZdla4+ZwkcspmWNtQd9gXuwRFLAe9wTsDjNETKBCjsRJmIU43+gvOau73j
mtwgRsIvEo10rcLgf0n2aQtO8Ju3VB3ng2PwIj6ijgu4VW0JwbmFZCL6yLnlHa9D
8IFnFDHNQE1tsLhSFQtbgWulEgu2SB2fqePKAQEqAdys8WuTWCaYYXsIZHWDPXwf
WsFAV2qk+31RInpGse0GqSclpBpK7x3tJ2dSweui3vm+GCLbFi0zEShBP3tPfIik
1ToSOn2lx3WsyLOjVOOUlyY93nMUR3IEqudBy/TxBn2m/3bSAFFGzLAZsDvyu+Rl
3GM5omKUXUG+8aSNpTK/yJ8qOBlLSV+CSzRg4P8eBN3iV6oDJ4K1pkX4Z/uh5UVL
b5RtCRD7tfjrJpQwhPh8Ey3LNVV9hOptk/iqZwJAN4QnrhmtlNWaZNe+j+1/HmB/
kDz2Fsh0lepo9dVIjzFEM0/tJCLK/DXRwxs8Na3/Du2QwBqGJ59JcKfHGcRbZ8tw
Y+kCQwuaKDZw6rlAQzmCTQ==
--pragma protect end_data_block
--pragma protect digest_block
4p2Q+X2lmm36hqtxcvYKF8sZa30=
--pragma protect end_digest_block
--pragma protect end_protected
