localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTX_CHK = {
  {32'h439dee52, 32'hc2938702} /* (31, 31, 31) {real, imag} */,
  {32'hc30daf0d, 32'h4332027c} /* (31, 31, 30) {real, imag} */,
  {32'h41362f1c, 32'hc213848f} /* (31, 31, 29) {real, imag} */,
  {32'h42119b1d, 32'h41a57278} /* (31, 31, 28) {real, imag} */,
  {32'hc1c19ccd, 32'h419e7756} /* (31, 31, 27) {real, imag} */,
  {32'hc0fabd28, 32'h40531204} /* (31, 31, 26) {real, imag} */,
  {32'h4034c462, 32'hc1a033b4} /* (31, 31, 25) {real, imag} */,
  {32'h40aeb782, 32'h41dd0b00} /* (31, 31, 24) {real, imag} */,
  {32'h40befc4c, 32'h416eb4a8} /* (31, 31, 23) {real, imag} */,
  {32'hc0a1aa6b, 32'h3fe88044} /* (31, 31, 22) {real, imag} */,
  {32'hc13e7cb9, 32'hbffc6964} /* (31, 31, 21) {real, imag} */,
  {32'h40b9e30e, 32'hc0d4cb9f} /* (31, 31, 20) {real, imag} */,
  {32'h40754597, 32'hc1920d4f} /* (31, 31, 19) {real, imag} */,
  {32'hc113965f, 32'h411959cb} /* (31, 31, 18) {real, imag} */,
  {32'h3fce1af4, 32'hc1359f0a} /* (31, 31, 17) {real, imag} */,
  {32'hc0956dda, 32'hc068c794} /* (31, 31, 16) {real, imag} */,
  {32'hc03376be, 32'hc0ebb03b} /* (31, 31, 15) {real, imag} */,
  {32'h3f9663be, 32'hc0bf7cac} /* (31, 31, 14) {real, imag} */,
  {32'hc18ff067, 32'hc11a0dd8} /* (31, 31, 13) {real, imag} */,
  {32'h4162982f, 32'hc184c0fc} /* (31, 31, 12) {real, imag} */,
  {32'hc0b47e5f, 32'hc0d40cf9} /* (31, 31, 11) {real, imag} */,
  {32'h4030aed2, 32'h3fdba0ce} /* (31, 31, 10) {real, imag} */,
  {32'hc18af551, 32'h3f9eae88} /* (31, 31, 9) {real, imag} */,
  {32'hc1806408, 32'h40ce4434} /* (31, 31, 8) {real, imag} */,
  {32'h409b413c, 32'h416214f5} /* (31, 31, 7) {real, imag} */,
  {32'hbfb810a0, 32'hbfffde38} /* (31, 31, 6) {real, imag} */,
  {32'hc1d80064, 32'hc05a9e8c} /* (31, 31, 5) {real, imag} */,
  {32'h421a1c02, 32'h410caad7} /* (31, 31, 4) {real, imag} */,
  {32'hc11bf57e, 32'hc125fb3a} /* (31, 31, 3) {real, imag} */,
  {32'hc2ef09e9, 32'hc1182aed} /* (31, 31, 2) {real, imag} */,
  {32'h438493cc, 32'h42b80d32} /* (31, 31, 1) {real, imag} */,
  {32'h4326c852, 32'hc2bb7234} /* (31, 31, 0) {real, imag} */,
  {32'hc3499a5c, 32'hc2bd7840} /* (31, 30, 31) {real, imag} */,
  {32'h42dd3696, 32'hc0d124e8} /* (31, 30, 30) {real, imag} */,
  {32'hc1a0ac18, 32'h4200c31b} /* (31, 30, 29) {real, imag} */,
  {32'hc1b6511c, 32'hc12337df} /* (31, 30, 28) {real, imag} */,
  {32'h41530186, 32'hc0737260} /* (31, 30, 27) {real, imag} */,
  {32'h40897e56, 32'hc12ed806} /* (31, 30, 26) {real, imag} */,
  {32'hc12bb2f7, 32'h414b5111} /* (31, 30, 25) {real, imag} */,
  {32'h41ef2bee, 32'hc0d2222c} /* (31, 30, 24) {real, imag} */,
  {32'hc118dfc2, 32'hc13158fd} /* (31, 30, 23) {real, imag} */,
  {32'hbfd9caf4, 32'hbd9b3b10} /* (31, 30, 22) {real, imag} */,
  {32'hbfb4c15e, 32'hc0e9df0e} /* (31, 30, 21) {real, imag} */,
  {32'h40dc355c, 32'hc0cdd14b} /* (31, 30, 20) {real, imag} */,
  {32'h40409b1c, 32'h3fcf5d8a} /* (31, 30, 19) {real, imag} */,
  {32'h41095751, 32'hc148427a} /* (31, 30, 18) {real, imag} */,
  {32'hc106fac4, 32'h401b8682} /* (31, 30, 17) {real, imag} */,
  {32'hbee31124, 32'h3f4d4240} /* (31, 30, 16) {real, imag} */,
  {32'h4109e9f6, 32'h3fc4be64} /* (31, 30, 15) {real, imag} */,
  {32'hc06ba101, 32'h3fe6c780} /* (31, 30, 14) {real, imag} */,
  {32'h4162f04c, 32'hc0819754} /* (31, 30, 13) {real, imag} */,
  {32'hbfa3ec68, 32'hbfae130e} /* (31, 30, 12) {real, imag} */,
  {32'h4162f668, 32'h40e1515c} /* (31, 30, 11) {real, imag} */,
  {32'hc172f0ec, 32'h3f0e8310} /* (31, 30, 10) {real, imag} */,
  {32'h412b479c, 32'hc00c3dfa} /* (31, 30, 9) {real, imag} */,
  {32'h419b96c1, 32'h40fb7fe6} /* (31, 30, 8) {real, imag} */,
  {32'hc08a9e1e, 32'h409fd663} /* (31, 30, 7) {real, imag} */,
  {32'h40ea6cf8, 32'hc1038de6} /* (31, 30, 6) {real, imag} */,
  {32'h41ed2bd4, 32'hbf8c53b0} /* (31, 30, 5) {real, imag} */,
  {32'hc23fda9e, 32'hc24d1a50} /* (31, 30, 4) {real, imag} */,
  {32'h3facdf70, 32'hc0aeaf80} /* (31, 30, 3) {real, imag} */,
  {32'h43019d18, 32'h42949812} /* (31, 30, 2) {real, imag} */,
  {32'hc36f6960, 32'h424168f2} /* (31, 30, 1) {real, imag} */,
  {32'hc3276984, 32'h41ad4ce4} /* (31, 30, 0) {real, imag} */,
  {32'h421bedbb, 32'h3f2e9a40} /* (31, 29, 31) {real, imag} */,
  {32'hc1bbf5ae, 32'h41b43a34} /* (31, 29, 30) {real, imag} */,
  {32'h41bd52ca, 32'h413569dc} /* (31, 29, 29) {real, imag} */,
  {32'hc0cf0708, 32'hc0cfc6d6} /* (31, 29, 28) {real, imag} */,
  {32'hc1cfc8b4, 32'hc17dcb73} /* (31, 29, 27) {real, imag} */,
  {32'hc08a434c, 32'hc0b4a165} /* (31, 29, 26) {real, imag} */,
  {32'hc11072bd, 32'hc083d25f} /* (31, 29, 25) {real, imag} */,
  {32'h4113b4ba, 32'h41430222} /* (31, 29, 24) {real, imag} */,
  {32'hc05561a2, 32'hc0c77273} /* (31, 29, 23) {real, imag} */,
  {32'hc13e0bff, 32'h40f308ea} /* (31, 29, 22) {real, imag} */,
  {32'h4077c029, 32'h411e2e57} /* (31, 29, 21) {real, imag} */,
  {32'hc11260de, 32'h4076e638} /* (31, 29, 20) {real, imag} */,
  {32'hc0e67c76, 32'h40c9adce} /* (31, 29, 19) {real, imag} */,
  {32'h410b7d17, 32'hc1381d17} /* (31, 29, 18) {real, imag} */,
  {32'hbffbca76, 32'h402ced04} /* (31, 29, 17) {real, imag} */,
  {32'hc03d577a, 32'hc0831819} /* (31, 29, 16) {real, imag} */,
  {32'h40a39150, 32'h4061ab12} /* (31, 29, 15) {real, imag} */,
  {32'h417cc18b, 32'h415345b8} /* (31, 29, 14) {real, imag} */,
  {32'h3ffeee6c, 32'h3f9dff84} /* (31, 29, 13) {real, imag} */,
  {32'hc029770b, 32'hbfeb5224} /* (31, 29, 12) {real, imag} */,
  {32'h3e90a1b8, 32'h418a7893} /* (31, 29, 11) {real, imag} */,
  {32'h405ce6d2, 32'hc0cb54ff} /* (31, 29, 10) {real, imag} */,
  {32'hc101ca50, 32'hbff97fac} /* (31, 29, 9) {real, imag} */,
  {32'h405299b0, 32'hc0d6086c} /* (31, 29, 8) {real, imag} */,
  {32'h40730f8c, 32'h3facd130} /* (31, 29, 7) {real, imag} */,
  {32'hc0028ff6, 32'h4081c2d8} /* (31, 29, 6) {real, imag} */,
  {32'hc0adcfd6, 32'h411d4a9e} /* (31, 29, 5) {real, imag} */,
  {32'h40ce45fe, 32'hc187ec76} /* (31, 29, 4) {real, imag} */,
  {32'h41e8cefa, 32'hbf8fbcf8} /* (31, 29, 3) {real, imag} */,
  {32'h41b3963e, 32'h420d7a5d} /* (31, 29, 2) {real, imag} */,
  {32'hc23608b6, 32'hc1f72bdf} /* (31, 29, 1) {real, imag} */,
  {32'h408c0d34, 32'hc1a5b2a1} /* (31, 29, 0) {real, imag} */,
  {32'h428b97f5, 32'hc25b3f8b} /* (31, 28, 31) {real, imag} */,
  {32'hc21d270a, 32'h420f271f} /* (31, 28, 30) {real, imag} */,
  {32'h40c4b08c, 32'hc180d07c} /* (31, 28, 29) {real, imag} */,
  {32'hbeeed220, 32'hc1ce1884} /* (31, 28, 28) {real, imag} */,
  {32'h4149c876, 32'h41bf98cf} /* (31, 28, 27) {real, imag} */,
  {32'hbfdb1d20, 32'hc105cabc} /* (31, 28, 26) {real, imag} */,
  {32'h413c07ec, 32'hc1346270} /* (31, 28, 25) {real, imag} */,
  {32'hc10fa1f5, 32'hc05ddcf8} /* (31, 28, 24) {real, imag} */,
  {32'hc07d92de, 32'hc0f2a6ac} /* (31, 28, 23) {real, imag} */,
  {32'hc1483aa2, 32'hc0882314} /* (31, 28, 22) {real, imag} */,
  {32'h41255d38, 32'h407b0a90} /* (31, 28, 21) {real, imag} */,
  {32'h40e4a678, 32'h41449646} /* (31, 28, 20) {real, imag} */,
  {32'h416dec7a, 32'h4019efa9} /* (31, 28, 19) {real, imag} */,
  {32'h40b4afc2, 32'hc043539c} /* (31, 28, 18) {real, imag} */,
  {32'hc02c984a, 32'h40a09fa2} /* (31, 28, 17) {real, imag} */,
  {32'h3e8a9b1c, 32'h405ee748} /* (31, 28, 16) {real, imag} */,
  {32'h40645e95, 32'hc150588b} /* (31, 28, 15) {real, imag} */,
  {32'h408576ca, 32'h4095ebf1} /* (31, 28, 14) {real, imag} */,
  {32'h40cb28c2, 32'h3f0655f8} /* (31, 28, 13) {real, imag} */,
  {32'h419eb55e, 32'h41329cf9} /* (31, 28, 12) {real, imag} */,
  {32'hc12e4620, 32'hc0c0408f} /* (31, 28, 11) {real, imag} */,
  {32'h40f950e0, 32'hc1609340} /* (31, 28, 10) {real, imag} */,
  {32'hc10443ac, 32'hbfd3453e} /* (31, 28, 9) {real, imag} */,
  {32'hc00fe500, 32'h40c56b6c} /* (31, 28, 8) {real, imag} */,
  {32'hc107ea4e, 32'hbfe26a54} /* (31, 28, 7) {real, imag} */,
  {32'hc121d585, 32'h40fb82a8} /* (31, 28, 6) {real, imag} */,
  {32'hc18bfcda, 32'h41851f03} /* (31, 28, 5) {real, imag} */,
  {32'h41e042af, 32'hc0f156a7} /* (31, 28, 4) {real, imag} */,
  {32'hc10fbb80, 32'hbdb66200} /* (31, 28, 3) {real, imag} */,
  {32'hc28cd4ce, 32'h40824a68} /* (31, 28, 2) {real, imag} */,
  {32'h419c4ad8, 32'hc2311866} /* (31, 28, 1) {real, imag} */,
  {32'h427929bb, 32'hc1778e14} /* (31, 28, 0) {real, imag} */,
  {32'hc21ae460, 32'h420d72c8} /* (31, 27, 31) {real, imag} */,
  {32'h421e150c, 32'hc1a2426c} /* (31, 27, 30) {real, imag} */,
  {32'hc1b6e6c7, 32'h40d9bee6} /* (31, 27, 29) {real, imag} */,
  {32'hc1cdd508, 32'h40b3407b} /* (31, 27, 28) {real, imag} */,
  {32'h3fc7fd20, 32'hc123aa34} /* (31, 27, 27) {real, imag} */,
  {32'h4185fe23, 32'hc0e9b1fe} /* (31, 27, 26) {real, imag} */,
  {32'h41464126, 32'h41a5b9b8} /* (31, 27, 25) {real, imag} */,
  {32'hbfb1666c, 32'hc13e995e} /* (31, 27, 24) {real, imag} */,
  {32'h3fda6cb6, 32'hc12e0e2d} /* (31, 27, 23) {real, imag} */,
  {32'h40506fff, 32'hc103cb71} /* (31, 27, 22) {real, imag} */,
  {32'hc15aee64, 32'h40aa447c} /* (31, 27, 21) {real, imag} */,
  {32'h409ad9ac, 32'hc0a615b6} /* (31, 27, 20) {real, imag} */,
  {32'hc0778f8c, 32'hc0907087} /* (31, 27, 19) {real, imag} */,
  {32'hc0f14d14, 32'hc094ddf8} /* (31, 27, 18) {real, imag} */,
  {32'hc070d2ba, 32'h40cfe692} /* (31, 27, 17) {real, imag} */,
  {32'hc13eb538, 32'h3d5e6d00} /* (31, 27, 16) {real, imag} */,
  {32'hc04538e9, 32'h403481fc} /* (31, 27, 15) {real, imag} */,
  {32'h3f48afe8, 32'hc08b4f34} /* (31, 27, 14) {real, imag} */,
  {32'h40f76658, 32'h4009a787} /* (31, 27, 13) {real, imag} */,
  {32'h415b75a4, 32'h41322510} /* (31, 27, 12) {real, imag} */,
  {32'hc0744fbb, 32'hc14768a9} /* (31, 27, 11) {real, imag} */,
  {32'h40c89cda, 32'h411036b4} /* (31, 27, 10) {real, imag} */,
  {32'h401d31ad, 32'hbfe35210} /* (31, 27, 9) {real, imag} */,
  {32'hc0850512, 32'h3eab8fb0} /* (31, 27, 8) {real, imag} */,
  {32'hc11f7293, 32'hc146d03c} /* (31, 27, 7) {real, imag} */,
  {32'h405a5d36, 32'hc05d2658} /* (31, 27, 6) {real, imag} */,
  {32'h41b5ed08, 32'h40219d04} /* (31, 27, 5) {real, imag} */,
  {32'hbff8d7b2, 32'h4193d560} /* (31, 27, 4) {real, imag} */,
  {32'hc00cb030, 32'h40dec44c} /* (31, 27, 3) {real, imag} */,
  {32'h410b8b90, 32'h41894173} /* (31, 27, 2) {real, imag} */,
  {32'hc24af712, 32'h4050c9e2} /* (31, 27, 1) {real, imag} */,
  {32'hc23893cf, 32'hc0d2dc80} /* (31, 27, 0) {real, imag} */,
  {32'hc18981a3, 32'h4088c332} /* (31, 26, 31) {real, imag} */,
  {32'hbff42db6, 32'h41ba80eb} /* (31, 26, 30) {real, imag} */,
  {32'h40a03cb0, 32'hc031741e} /* (31, 26, 29) {real, imag} */,
  {32'hc01133dc, 32'hc0c43be0} /* (31, 26, 28) {real, imag} */,
  {32'h413e0844, 32'hc139b7c6} /* (31, 26, 27) {real, imag} */,
  {32'hc0e9ead0, 32'h3f2e1798} /* (31, 26, 26) {real, imag} */,
  {32'hc16b66f3, 32'hc13550c5} /* (31, 26, 25) {real, imag} */,
  {32'h415cb0f2, 32'hc109e8af} /* (31, 26, 24) {real, imag} */,
  {32'h40894cfb, 32'h3e1c0a00} /* (31, 26, 23) {real, imag} */,
  {32'hc0d41c83, 32'h4101bad7} /* (31, 26, 22) {real, imag} */,
  {32'hbf7641e8, 32'hbe1e9700} /* (31, 26, 21) {real, imag} */,
  {32'hc1192283, 32'hbf03d8ac} /* (31, 26, 20) {real, imag} */,
  {32'hc108d089, 32'h41282d26} /* (31, 26, 19) {real, imag} */,
  {32'h40281c76, 32'h41447cdf} /* (31, 26, 18) {real, imag} */,
  {32'h40acefb7, 32'hc0db3ad6} /* (31, 26, 17) {real, imag} */,
  {32'h4063b9c0, 32'hbfd28bf4} /* (31, 26, 16) {real, imag} */,
  {32'hc0b10418, 32'h412579d2} /* (31, 26, 15) {real, imag} */,
  {32'h3f2bda52, 32'hc0f84644} /* (31, 26, 14) {real, imag} */,
  {32'hc1300fbd, 32'h3f5b33f8} /* (31, 26, 13) {real, imag} */,
  {32'hc131d34a, 32'h3f00427a} /* (31, 26, 12) {real, imag} */,
  {32'h4122b3a2, 32'h41495768} /* (31, 26, 11) {real, imag} */,
  {32'h3fa39282, 32'h41210a6a} /* (31, 26, 10) {real, imag} */,
  {32'hc09a798c, 32'h4165a3df} /* (31, 26, 9) {real, imag} */,
  {32'h40ae60dc, 32'hc0d95abe} /* (31, 26, 8) {real, imag} */,
  {32'hbfe73422, 32'h4073e94a} /* (31, 26, 7) {real, imag} */,
  {32'h40f3b8d0, 32'hc185d8c4} /* (31, 26, 6) {real, imag} */,
  {32'hc0a40e4c, 32'hc0c78610} /* (31, 26, 5) {real, imag} */,
  {32'hc0379818, 32'hc0532e6a} /* (31, 26, 4) {real, imag} */,
  {32'h415501e8, 32'hbf1024a0} /* (31, 26, 3) {real, imag} */,
  {32'hc1793ef2, 32'h4192f0bd} /* (31, 26, 2) {real, imag} */,
  {32'hc11e14ac, 32'hc1990a00} /* (31, 26, 1) {real, imag} */,
  {32'h418b9ecc, 32'h41094da7} /* (31, 26, 0) {real, imag} */,
  {32'hc0fba278, 32'hbfdf8b58} /* (31, 25, 31) {real, imag} */,
  {32'h41293268, 32'h41165ef5} /* (31, 25, 30) {real, imag} */,
  {32'h411f2e3e, 32'hbebc42c0} /* (31, 25, 29) {real, imag} */,
  {32'h409e1d5e, 32'h3f280c30} /* (31, 25, 28) {real, imag} */,
  {32'h4109c6b4, 32'h3eac5f60} /* (31, 25, 27) {real, imag} */,
  {32'h40c1bab5, 32'h40331082} /* (31, 25, 26) {real, imag} */,
  {32'h3f9a2034, 32'h3fb470e4} /* (31, 25, 25) {real, imag} */,
  {32'hc0b78ca5, 32'hc0ac7309} /* (31, 25, 24) {real, imag} */,
  {32'hc0d4eccd, 32'h4110d042} /* (31, 25, 23) {real, imag} */,
  {32'h40f8dbc1, 32'hbd141200} /* (31, 25, 22) {real, imag} */,
  {32'h4136823c, 32'hbff50374} /* (31, 25, 21) {real, imag} */,
  {32'hbff19626, 32'h40b1cac9} /* (31, 25, 20) {real, imag} */,
  {32'hc0cdd438, 32'h4032e3e0} /* (31, 25, 19) {real, imag} */,
  {32'hc0f39be6, 32'hc1110df6} /* (31, 25, 18) {real, imag} */,
  {32'h4019860d, 32'hc0b0dd6d} /* (31, 25, 17) {real, imag} */,
  {32'h4005a819, 32'h4034fd79} /* (31, 25, 16) {real, imag} */,
  {32'h4166fd63, 32'hc0b8346a} /* (31, 25, 15) {real, imag} */,
  {32'hc0a0c473, 32'hc0c0fea0} /* (31, 25, 14) {real, imag} */,
  {32'hbfe83328, 32'hc0e44fbc} /* (31, 25, 13) {real, imag} */,
  {32'hc10a01ef, 32'h409af006} /* (31, 25, 12) {real, imag} */,
  {32'hbf88a6e0, 32'hc123dc38} /* (31, 25, 11) {real, imag} */,
  {32'hc08df467, 32'hbf1b1934} /* (31, 25, 10) {real, imag} */,
  {32'h411f2d74, 32'hc04b695e} /* (31, 25, 9) {real, imag} */,
  {32'hc0c2e356, 32'hc13c8bcd} /* (31, 25, 8) {real, imag} */,
  {32'h40c79370, 32'h3feb8a66} /* (31, 25, 7) {real, imag} */,
  {32'h410a5bc2, 32'hc0d82780} /* (31, 25, 6) {real, imag} */,
  {32'hc0f785e5, 32'h40ce5842} /* (31, 25, 5) {real, imag} */,
  {32'hc15baf1b, 32'hbfc9e580} /* (31, 25, 4) {real, imag} */,
  {32'h3fe7df34, 32'h3f780128} /* (31, 25, 3) {real, imag} */,
  {32'hc0b13a1e, 32'h40a653c2} /* (31, 25, 2) {real, imag} */,
  {32'h40e7ff8e, 32'hbe5a9460} /* (31, 25, 1) {real, imag} */,
  {32'h41bc68b9, 32'hc15dbf4f} /* (31, 25, 0) {real, imag} */,
  {32'hc19a969c, 32'h416db412} /* (31, 24, 31) {real, imag} */,
  {32'h41594f0e, 32'hc214167c} /* (31, 24, 30) {real, imag} */,
  {32'hc1c4b78b, 32'h3fee5298} /* (31, 24, 29) {real, imag} */,
  {32'h40c2184c, 32'hc0c9c841} /* (31, 24, 28) {real, imag} */,
  {32'h3fe6175a, 32'hc0ee92c0} /* (31, 24, 27) {real, imag} */,
  {32'h412f152f, 32'hc0974dd7} /* (31, 24, 26) {real, imag} */,
  {32'hc0145f40, 32'h413bd7cf} /* (31, 24, 25) {real, imag} */,
  {32'h3fd70de0, 32'h40f56abe} /* (31, 24, 24) {real, imag} */,
  {32'h4028504e, 32'h40878ba2} /* (31, 24, 23) {real, imag} */,
  {32'hbfab4bc4, 32'hc1115521} /* (31, 24, 22) {real, imag} */,
  {32'hc0d49f56, 32'hc0ccf1b2} /* (31, 24, 21) {real, imag} */,
  {32'hbe836b80, 32'hc1115e94} /* (31, 24, 20) {real, imag} */,
  {32'h4088d7d6, 32'h3fe0e870} /* (31, 24, 19) {real, imag} */,
  {32'h3fe91e8c, 32'hc00c5802} /* (31, 24, 18) {real, imag} */,
  {32'hbf8ba3a0, 32'h3faa554a} /* (31, 24, 17) {real, imag} */,
  {32'hbfc52614, 32'h40526313} /* (31, 24, 16) {real, imag} */,
  {32'h410095c5, 32'hc15d26c9} /* (31, 24, 15) {real, imag} */,
  {32'hc0b90fcc, 32'hc09af45e} /* (31, 24, 14) {real, imag} */,
  {32'hc039c6be, 32'hc031a2e4} /* (31, 24, 13) {real, imag} */,
  {32'hbffdd8d0, 32'hc075aaaa} /* (31, 24, 12) {real, imag} */,
  {32'hc0e4b441, 32'hbf97b2cf} /* (31, 24, 11) {real, imag} */,
  {32'h409babf0, 32'h40d466b6} /* (31, 24, 10) {real, imag} */,
  {32'h4037007c, 32'hc10f0ba4} /* (31, 24, 9) {real, imag} */,
  {32'hc0c92ac2, 32'h40377b80} /* (31, 24, 8) {real, imag} */,
  {32'h40f2cd22, 32'h3e4eb150} /* (31, 24, 7) {real, imag} */,
  {32'hc15ea0ef, 32'h3f97d3d0} /* (31, 24, 6) {real, imag} */,
  {32'h409bef4b, 32'hc060721f} /* (31, 24, 5) {real, imag} */,
  {32'hc15f86e0, 32'hc11cb912} /* (31, 24, 4) {real, imag} */,
  {32'hc0e482e0, 32'hbf6ce152} /* (31, 24, 3) {real, imag} */,
  {32'h42084781, 32'h4075c13c} /* (31, 24, 2) {real, imag} */,
  {32'hc1d0e843, 32'h41a4fb94} /* (31, 24, 1) {real, imag} */,
  {32'hc1914c26, 32'hbcc21600} /* (31, 24, 0) {real, imag} */,
  {32'h40cc622c, 32'h3f985c98} /* (31, 23, 31) {real, imag} */,
  {32'hc07f7808, 32'h4184fa9e} /* (31, 23, 30) {real, imag} */,
  {32'hc1d21346, 32'hc0896349} /* (31, 23, 29) {real, imag} */,
  {32'h4198b11b, 32'h3f4e8150} /* (31, 23, 28) {real, imag} */,
  {32'hc073cc42, 32'h3e0c8420} /* (31, 23, 27) {real, imag} */,
  {32'hc12282da, 32'h407e8882} /* (31, 23, 26) {real, imag} */,
  {32'h41712da5, 32'h40c8d34e} /* (31, 23, 25) {real, imag} */,
  {32'hc0f0dc44, 32'h413d8d9c} /* (31, 23, 24) {real, imag} */,
  {32'h4068b5d8, 32'h4135b0c7} /* (31, 23, 23) {real, imag} */,
  {32'h404ac83a, 32'hc01e7aaa} /* (31, 23, 22) {real, imag} */,
  {32'h408f7852, 32'h3f232ec4} /* (31, 23, 21) {real, imag} */,
  {32'hbffbc24e, 32'h41422173} /* (31, 23, 20) {real, imag} */,
  {32'h4185fe52, 32'h3e3170a0} /* (31, 23, 19) {real, imag} */,
  {32'h40e63a16, 32'h3fc2c578} /* (31, 23, 18) {real, imag} */,
  {32'h3fefa734, 32'h4037f21d} /* (31, 23, 17) {real, imag} */,
  {32'h3feb3254, 32'h3fe06e7c} /* (31, 23, 16) {real, imag} */,
  {32'h41194d99, 32'h403ecb92} /* (31, 23, 15) {real, imag} */,
  {32'hc0c72524, 32'h3fb68b96} /* (31, 23, 14) {real, imag} */,
  {32'hc148ab2c, 32'h40948950} /* (31, 23, 13) {real, imag} */,
  {32'h3fad2ad0, 32'h408c6ea8} /* (31, 23, 12) {real, imag} */,
  {32'h40e4eb5c, 32'h40ede0ce} /* (31, 23, 11) {real, imag} */,
  {32'h3da1e380, 32'hc0928605} /* (31, 23, 10) {real, imag} */,
  {32'hc0174a9c, 32'hbfbcfafe} /* (31, 23, 9) {real, imag} */,
  {32'h400aae08, 32'h3fede7f4} /* (31, 23, 8) {real, imag} */,
  {32'h402eeba3, 32'hbd242480} /* (31, 23, 7) {real, imag} */,
  {32'h4088c8e4, 32'hc0e7a1cc} /* (31, 23, 6) {real, imag} */,
  {32'h40f5c4d8, 32'h40fe20d1} /* (31, 23, 5) {real, imag} */,
  {32'h418b52f8, 32'hc10fa040} /* (31, 23, 4) {real, imag} */,
  {32'h4153cc2b, 32'hc0251eb4} /* (31, 23, 3) {real, imag} */,
  {32'h403bd282, 32'hc0f5aaae} /* (31, 23, 2) {real, imag} */,
  {32'hbf951e64, 32'hc1b06eab} /* (31, 23, 1) {real, imag} */,
  {32'h3ee423a0, 32'hc1298906} /* (31, 23, 0) {real, imag} */,
  {32'h417b2137, 32'h4062948a} /* (31, 22, 31) {real, imag} */,
  {32'h3f292820, 32'h41099ad6} /* (31, 22, 30) {real, imag} */,
  {32'h416fcaff, 32'h409234fb} /* (31, 22, 29) {real, imag} */,
  {32'hbf821650, 32'hc0d04090} /* (31, 22, 28) {real, imag} */,
  {32'h3ec17f20, 32'h40a459bc} /* (31, 22, 27) {real, imag} */,
  {32'hc0b2ae8a, 32'h41280efc} /* (31, 22, 26) {real, imag} */,
  {32'h410499a7, 32'hc11ac8ae} /* (31, 22, 25) {real, imag} */,
  {32'hc04b8329, 32'h409ed2ac} /* (31, 22, 24) {real, imag} */,
  {32'h40c99dcc, 32'hc1266e8c} /* (31, 22, 23) {real, imag} */,
  {32'hc11be0ba, 32'h3f267df0} /* (31, 22, 22) {real, imag} */,
  {32'hc0a0c3c1, 32'h4084d479} /* (31, 22, 21) {real, imag} */,
  {32'hc0d003ac, 32'hc142e57a} /* (31, 22, 20) {real, imag} */,
  {32'h3f1332f0, 32'hc1526b2c} /* (31, 22, 19) {real, imag} */,
  {32'hbfbeac1c, 32'h3f158a18} /* (31, 22, 18) {real, imag} */,
  {32'hbf0d18d3, 32'h3f15a1f8} /* (31, 22, 17) {real, imag} */,
  {32'hc0478fae, 32'hc03b0c29} /* (31, 22, 16) {real, imag} */,
  {32'hc0b83a84, 32'h402bd4e2} /* (31, 22, 15) {real, imag} */,
  {32'h40c9545a, 32'h40ffc24c} /* (31, 22, 14) {real, imag} */,
  {32'h3ff29148, 32'h4135247e} /* (31, 22, 13) {real, imag} */,
  {32'hc0cdc24c, 32'hc161f6d6} /* (31, 22, 12) {real, imag} */,
  {32'hc1591886, 32'h40b57960} /* (31, 22, 11) {real, imag} */,
  {32'h413605f8, 32'h4028a82e} /* (31, 22, 10) {real, imag} */,
  {32'hc18732e3, 32'hc112e901} /* (31, 22, 9) {real, imag} */,
  {32'hc0565b06, 32'h3fb05448} /* (31, 22, 8) {real, imag} */,
  {32'hc03f5fa4, 32'h40ebcc2c} /* (31, 22, 7) {real, imag} */,
  {32'hbfed302c, 32'hc1073d2c} /* (31, 22, 6) {real, imag} */,
  {32'hc04ce049, 32'h41529c58} /* (31, 22, 5) {real, imag} */,
  {32'h417aab8a, 32'h405d56f4} /* (31, 22, 4) {real, imag} */,
  {32'hbf15a9f0, 32'hc076f8b6} /* (31, 22, 3) {real, imag} */,
  {32'h3fc85468, 32'hc0409008} /* (31, 22, 2) {real, imag} */,
  {32'hc037182e, 32'hc155751c} /* (31, 22, 1) {real, imag} */,
  {32'hc11b69de, 32'hbff16ea6} /* (31, 22, 0) {real, imag} */,
  {32'hc021a8e4, 32'hc04a40bc} /* (31, 21, 31) {real, imag} */,
  {32'hc0c33bf4, 32'hc06b53c8} /* (31, 21, 30) {real, imag} */,
  {32'h4088b553, 32'h3fc2f370} /* (31, 21, 29) {real, imag} */,
  {32'h40a5fa2a, 32'hc15776c7} /* (31, 21, 28) {real, imag} */,
  {32'h4107d1fd, 32'h40fb2ea3} /* (31, 21, 27) {real, imag} */,
  {32'h3febae20, 32'hc09bf936} /* (31, 21, 26) {real, imag} */,
  {32'hc0e31f3a, 32'h4113480f} /* (31, 21, 25) {real, imag} */,
  {32'h40c1b487, 32'h3f2dbd94} /* (31, 21, 24) {real, imag} */,
  {32'hc02c9ad2, 32'h3ff942dc} /* (31, 21, 23) {real, imag} */,
  {32'h419546ee, 32'hc0fefc90} /* (31, 21, 22) {real, imag} */,
  {32'h40b1c0c8, 32'hc17db588} /* (31, 21, 21) {real, imag} */,
  {32'hc0e8ec32, 32'h41cddde0} /* (31, 21, 20) {real, imag} */,
  {32'hc124ae6e, 32'h40c3f882} /* (31, 21, 19) {real, imag} */,
  {32'hc146cd51, 32'h3f82daf4} /* (31, 21, 18) {real, imag} */,
  {32'h3f1997e4, 32'h400a0578} /* (31, 21, 17) {real, imag} */,
  {32'h3f7b1668, 32'hbf85a969} /* (31, 21, 16) {real, imag} */,
  {32'h3fe6146c, 32'hc055fabb} /* (31, 21, 15) {real, imag} */,
  {32'hbec0bd30, 32'h4106079f} /* (31, 21, 14) {real, imag} */,
  {32'hc07dc950, 32'h4176c5f8} /* (31, 21, 13) {real, imag} */,
  {32'hc0be6374, 32'hc0dbb608} /* (31, 21, 12) {real, imag} */,
  {32'h4112f17d, 32'hc1639db0} /* (31, 21, 11) {real, imag} */,
  {32'hbed09060, 32'h3f7aff60} /* (31, 21, 10) {real, imag} */,
  {32'h3fcf8258, 32'hc182107c} /* (31, 21, 9) {real, imag} */,
  {32'h408376c0, 32'h4100dec2} /* (31, 21, 8) {real, imag} */,
  {32'hc1814fd7, 32'hc0888f4e} /* (31, 21, 7) {real, imag} */,
  {32'hc04356a4, 32'h40823a46} /* (31, 21, 6) {real, imag} */,
  {32'hbf60ec54, 32'hbe7ca8c0} /* (31, 21, 5) {real, imag} */,
  {32'hc105a598, 32'hc1154e42} /* (31, 21, 4) {real, imag} */,
  {32'h4020c944, 32'hc0ad8e7a} /* (31, 21, 3) {real, imag} */,
  {32'hc0653658, 32'hc1437cfc} /* (31, 21, 2) {real, imag} */,
  {32'h4028efb0, 32'h40cc6be4} /* (31, 21, 1) {real, imag} */,
  {32'h400acf98, 32'h40b02c98} /* (31, 21, 0) {real, imag} */,
  {32'hc0543cf8, 32'hc13f0ac8} /* (31, 20, 31) {real, imag} */,
  {32'hc1589a43, 32'h3fa4cdc4} /* (31, 20, 30) {real, imag} */,
  {32'hc0d64c01, 32'hbe86f570} /* (31, 20, 29) {real, imag} */,
  {32'h3fd80b50, 32'h4084a77d} /* (31, 20, 28) {real, imag} */,
  {32'h3ee9c1c0, 32'h40009b30} /* (31, 20, 27) {real, imag} */,
  {32'h3eb58d80, 32'h40ba8861} /* (31, 20, 26) {real, imag} */,
  {32'hc108fbc3, 32'h4124c18d} /* (31, 20, 25) {real, imag} */,
  {32'h407f55dc, 32'hc11a0719} /* (31, 20, 24) {real, imag} */,
  {32'hbd8d6120, 32'h416156ec} /* (31, 20, 23) {real, imag} */,
  {32'h40b589ae, 32'hc1156562} /* (31, 20, 22) {real, imag} */,
  {32'h40cceeb6, 32'h409d76f5} /* (31, 20, 21) {real, imag} */,
  {32'hc0a4d572, 32'hc09b5ac0} /* (31, 20, 20) {real, imag} */,
  {32'hc178413e, 32'hc09d2f8d} /* (31, 20, 19) {real, imag} */,
  {32'h4027b070, 32'hc10028b7} /* (31, 20, 18) {real, imag} */,
  {32'hc0f92e4c, 32'hc095de98} /* (31, 20, 17) {real, imag} */,
  {32'h408742f1, 32'h40311834} /* (31, 20, 16) {real, imag} */,
  {32'h40bde3ee, 32'h40968084} /* (31, 20, 15) {real, imag} */,
  {32'hc16de012, 32'h3f174a9c} /* (31, 20, 14) {real, imag} */,
  {32'hc1850658, 32'h40763ff8} /* (31, 20, 13) {real, imag} */,
  {32'hc0e45933, 32'hc121384f} /* (31, 20, 12) {real, imag} */,
  {32'h4118e874, 32'hc109367a} /* (31, 20, 11) {real, imag} */,
  {32'hbf83b0a0, 32'hc1078050} /* (31, 20, 10) {real, imag} */,
  {32'h3fccdd22, 32'h3f9f3a48} /* (31, 20, 9) {real, imag} */,
  {32'hc0d0279e, 32'h413709e2} /* (31, 20, 8) {real, imag} */,
  {32'h3f15e1c8, 32'hc1682ee6} /* (31, 20, 7) {real, imag} */,
  {32'hbe894928, 32'h4096d987} /* (31, 20, 6) {real, imag} */,
  {32'h409d1826, 32'h40db0090} /* (31, 20, 5) {real, imag} */,
  {32'hc10a7620, 32'h4173d52d} /* (31, 20, 4) {real, imag} */,
  {32'h40aad024, 32'h3fe399a8} /* (31, 20, 3) {real, imag} */,
  {32'h411c4160, 32'hc10a4e9d} /* (31, 20, 2) {real, imag} */,
  {32'h4000ec8a, 32'h40a1efa1} /* (31, 20, 1) {real, imag} */,
  {32'h406c86e8, 32'hbfdee5a0} /* (31, 20, 0) {real, imag} */,
  {32'h40d81b6a, 32'h3fb1fd74} /* (31, 19, 31) {real, imag} */,
  {32'h3fab63d0, 32'h3f62140e} /* (31, 19, 30) {real, imag} */,
  {32'hc0464b7b, 32'hc0ab7c00} /* (31, 19, 29) {real, imag} */,
  {32'hc0ef1cd4, 32'hbec9b078} /* (31, 19, 28) {real, imag} */,
  {32'hc11c26dd, 32'h3fa4c24c} /* (31, 19, 27) {real, imag} */,
  {32'hc0347838, 32'hbfabb318} /* (31, 19, 26) {real, imag} */,
  {32'h4117f0f1, 32'h3f192d38} /* (31, 19, 25) {real, imag} */,
  {32'hc13c521a, 32'h3fffaf34} /* (31, 19, 24) {real, imag} */,
  {32'h41251077, 32'h40a3cb33} /* (31, 19, 23) {real, imag} */,
  {32'h3f9e061c, 32'hc017175f} /* (31, 19, 22) {real, imag} */,
  {32'hc11ccd3e, 32'hc09bca84} /* (31, 19, 21) {real, imag} */,
  {32'hc083d163, 32'hbe81be44} /* (31, 19, 20) {real, imag} */,
  {32'hc14929d3, 32'h4042d611} /* (31, 19, 19) {real, imag} */,
  {32'h40a60478, 32'hbe84a4ac} /* (31, 19, 18) {real, imag} */,
  {32'hc0ad712a, 32'h3f0bea74} /* (31, 19, 17) {real, imag} */,
  {32'hbfae0778, 32'hc1266b70} /* (31, 19, 16) {real, imag} */,
  {32'h40966334, 32'h41027db3} /* (31, 19, 15) {real, imag} */,
  {32'h41971075, 32'h40c809a3} /* (31, 19, 14) {real, imag} */,
  {32'h4169b856, 32'hc0d57d13} /* (31, 19, 13) {real, imag} */,
  {32'h4092d966, 32'h3f33c830} /* (31, 19, 12) {real, imag} */,
  {32'hc00bea62, 32'h411ebb67} /* (31, 19, 11) {real, imag} */,
  {32'hbde82a60, 32'h4070add0} /* (31, 19, 10) {real, imag} */,
  {32'h402e39ce, 32'h401df376} /* (31, 19, 9) {real, imag} */,
  {32'hc064bd6c, 32'h40ed93fc} /* (31, 19, 8) {real, imag} */,
  {32'hbefd8678, 32'h3fe37ce8} /* (31, 19, 7) {real, imag} */,
  {32'h409b2502, 32'h4127c662} /* (31, 19, 6) {real, imag} */,
  {32'h3f68bb7a, 32'h411442a4} /* (31, 19, 5) {real, imag} */,
  {32'h3da664c0, 32'hc020a082} /* (31, 19, 4) {real, imag} */,
  {32'h411e1c76, 32'h3e0577a8} /* (31, 19, 3) {real, imag} */,
  {32'hc166f562, 32'hc04fa33c} /* (31, 19, 2) {real, imag} */,
  {32'hc0d80b49, 32'h40a4a311} /* (31, 19, 1) {real, imag} */,
  {32'hc0fe0ebe, 32'h3f9b3684} /* (31, 19, 0) {real, imag} */,
  {32'h4101bf84, 32'h408b7d9b} /* (31, 18, 31) {real, imag} */,
  {32'h40a93009, 32'hbffe9298} /* (31, 18, 30) {real, imag} */,
  {32'h4103903f, 32'hc0acb238} /* (31, 18, 29) {real, imag} */,
  {32'h3fca79ae, 32'h40ef80ca} /* (31, 18, 28) {real, imag} */,
  {32'h412b6264, 32'hc117f7ec} /* (31, 18, 27) {real, imag} */,
  {32'hc13b58ff, 32'hbfccc574} /* (31, 18, 26) {real, imag} */,
  {32'hc133f133, 32'hc1b296e0} /* (31, 18, 25) {real, imag} */,
  {32'h40bb7a3a, 32'h3f017220} /* (31, 18, 24) {real, imag} */,
  {32'h412f36b2, 32'hc0682970} /* (31, 18, 23) {real, imag} */,
  {32'h411751a8, 32'hc031307c} /* (31, 18, 22) {real, imag} */,
  {32'hc09bceac, 32'h3fe3da30} /* (31, 18, 21) {real, imag} */,
  {32'h3db1bcc0, 32'hc027ea2e} /* (31, 18, 20) {real, imag} */,
  {32'h40501aa2, 32'hc163deb6} /* (31, 18, 19) {real, imag} */,
  {32'h3ef086c0, 32'h414eb670} /* (31, 18, 18) {real, imag} */,
  {32'hc097802f, 32'h3fc7bf90} /* (31, 18, 17) {real, imag} */,
  {32'hc020b9a0, 32'hc104032c} /* (31, 18, 16) {real, imag} */,
  {32'hc0b7c90e, 32'h400fe72c} /* (31, 18, 15) {real, imag} */,
  {32'hc0925510, 32'hbdba12a0} /* (31, 18, 14) {real, imag} */,
  {32'hc04ca990, 32'hc1735c1c} /* (31, 18, 13) {real, imag} */,
  {32'hc111509c, 32'hc008059a} /* (31, 18, 12) {real, imag} */,
  {32'h3f9be65a, 32'h40a3716b} /* (31, 18, 11) {real, imag} */,
  {32'h413a0946, 32'hc178b440} /* (31, 18, 10) {real, imag} */,
  {32'hc1074454, 32'hc04751d2} /* (31, 18, 9) {real, imag} */,
  {32'h401acde2, 32'h40f27ffb} /* (31, 18, 8) {real, imag} */,
  {32'h405e656c, 32'hc0860b01} /* (31, 18, 7) {real, imag} */,
  {32'h416e40ac, 32'hc0b2cdec} /* (31, 18, 6) {real, imag} */,
  {32'hc161b329, 32'hc0c17294} /* (31, 18, 5) {real, imag} */,
  {32'hc1365b50, 32'h4019b62d} /* (31, 18, 4) {real, imag} */,
  {32'hc0ac0c12, 32'h40276470} /* (31, 18, 3) {real, imag} */,
  {32'h40bc42c3, 32'hc0bb78df} /* (31, 18, 2) {real, imag} */,
  {32'hc0f35f1a, 32'h402968e9} /* (31, 18, 1) {real, imag} */,
  {32'hc04ce2f7, 32'h40742a7a} /* (31, 18, 0) {real, imag} */,
  {32'h4074a53b, 32'hc084cc7a} /* (31, 17, 31) {real, imag} */,
  {32'hbe5bfb60, 32'h407ef370} /* (31, 17, 30) {real, imag} */,
  {32'h3f814068, 32'hc025de1e} /* (31, 17, 29) {real, imag} */,
  {32'h3f53b3e0, 32'hc06e7580} /* (31, 17, 28) {real, imag} */,
  {32'h401487ef, 32'hbfc3c96c} /* (31, 17, 27) {real, imag} */,
  {32'h40ae9c56, 32'hc02f9e12} /* (31, 17, 26) {real, imag} */,
  {32'h40a9fbe4, 32'h41122d20} /* (31, 17, 25) {real, imag} */,
  {32'hc0ef167a, 32'hbefa0940} /* (31, 17, 24) {real, imag} */,
  {32'h40a20942, 32'hc05f8dbe} /* (31, 17, 23) {real, imag} */,
  {32'hc08b75ea, 32'h3f9200e4} /* (31, 17, 22) {real, imag} */,
  {32'h4105b139, 32'h40274b7c} /* (31, 17, 21) {real, imag} */,
  {32'h406ae666, 32'hc115cad1} /* (31, 17, 20) {real, imag} */,
  {32'hc08f8b84, 32'h40981a4e} /* (31, 17, 19) {real, imag} */,
  {32'h4000daef, 32'hc1426d7a} /* (31, 17, 18) {real, imag} */,
  {32'hbf318148, 32'h40788808} /* (31, 17, 17) {real, imag} */,
  {32'h3f0a84ac, 32'hbfecb748} /* (31, 17, 16) {real, imag} */,
  {32'h4045f59a, 32'h40f8547c} /* (31, 17, 15) {real, imag} */,
  {32'hc09f0069, 32'hc103ae12} /* (31, 17, 14) {real, imag} */,
  {32'h3dce6b00, 32'h408753f7} /* (31, 17, 13) {real, imag} */,
  {32'h3fd23c7f, 32'hc10f67df} /* (31, 17, 12) {real, imag} */,
  {32'h40cbbabb, 32'h40bb11bf} /* (31, 17, 11) {real, imag} */,
  {32'h3fdd7938, 32'hc0d890eb} /* (31, 17, 10) {real, imag} */,
  {32'h405ad27c, 32'h40ef4fdd} /* (31, 17, 9) {real, imag} */,
  {32'hbfdbea20, 32'hbfb0d2f8} /* (31, 17, 8) {real, imag} */,
  {32'hc0a5a7ee, 32'h408fa31e} /* (31, 17, 7) {real, imag} */,
  {32'h40ec48b5, 32'hc0833c0f} /* (31, 17, 6) {real, imag} */,
  {32'h40191868, 32'hc0442bb2} /* (31, 17, 5) {real, imag} */,
  {32'h402f87ac, 32'h4085e8a5} /* (31, 17, 4) {real, imag} */,
  {32'hbfbe9c4c, 32'h411a840d} /* (31, 17, 3) {real, imag} */,
  {32'h3f619fd8, 32'h401e5058} /* (31, 17, 2) {real, imag} */,
  {32'hc112b414, 32'hc00fe061} /* (31, 17, 1) {real, imag} */,
  {32'hc08948b2, 32'h409a678d} /* (31, 17, 0) {real, imag} */,
  {32'h40335242, 32'h40335c43} /* (31, 16, 31) {real, imag} */,
  {32'hc0b771b3, 32'h40042732} /* (31, 16, 30) {real, imag} */,
  {32'h41001190, 32'h4028a1b2} /* (31, 16, 29) {real, imag} */,
  {32'h402a207f, 32'h40bb70a8} /* (31, 16, 28) {real, imag} */,
  {32'h3f687118, 32'h3f25d780} /* (31, 16, 27) {real, imag} */,
  {32'h409c574a, 32'hbfb9b54e} /* (31, 16, 26) {real, imag} */,
  {32'h4010fa58, 32'hc0892f70} /* (31, 16, 25) {real, imag} */,
  {32'h40a255bf, 32'h412c6e22} /* (31, 16, 24) {real, imag} */,
  {32'hc02eae0c, 32'hc0c97008} /* (31, 16, 23) {real, imag} */,
  {32'hc0d2f68a, 32'h407cd688} /* (31, 16, 22) {real, imag} */,
  {32'h3fc7a490, 32'hc092958d} /* (31, 16, 21) {real, imag} */,
  {32'h404599f2, 32'h3ffa860c} /* (31, 16, 20) {real, imag} */,
  {32'h4071a6bb, 32'hc01ccfed} /* (31, 16, 19) {real, imag} */,
  {32'h40fc737d, 32'h3f5cece8} /* (31, 16, 18) {real, imag} */,
  {32'hc0ab9d15, 32'hc0149a13} /* (31, 16, 17) {real, imag} */,
  {32'hc0a670fc, 32'h00000000} /* (31, 16, 16) {real, imag} */,
  {32'hc0ab9d15, 32'h40149a13} /* (31, 16, 15) {real, imag} */,
  {32'h40fc737d, 32'hbf5cece8} /* (31, 16, 14) {real, imag} */,
  {32'h4071a6bb, 32'h401ccfed} /* (31, 16, 13) {real, imag} */,
  {32'h404599f2, 32'hbffa860c} /* (31, 16, 12) {real, imag} */,
  {32'h3fc7a490, 32'h4092958d} /* (31, 16, 11) {real, imag} */,
  {32'hc0d2f68a, 32'hc07cd688} /* (31, 16, 10) {real, imag} */,
  {32'hc02eae0c, 32'h40c97008} /* (31, 16, 9) {real, imag} */,
  {32'h40a255bf, 32'hc12c6e22} /* (31, 16, 8) {real, imag} */,
  {32'h4010fa58, 32'h40892f70} /* (31, 16, 7) {real, imag} */,
  {32'h409c574a, 32'h3fb9b54e} /* (31, 16, 6) {real, imag} */,
  {32'h3f687118, 32'hbf25d780} /* (31, 16, 5) {real, imag} */,
  {32'h402a207f, 32'hc0bb70a8} /* (31, 16, 4) {real, imag} */,
  {32'h41001190, 32'hc028a1b2} /* (31, 16, 3) {real, imag} */,
  {32'hc0b771b3, 32'hc0042732} /* (31, 16, 2) {real, imag} */,
  {32'h40335242, 32'hc0335c43} /* (31, 16, 1) {real, imag} */,
  {32'hc16215fa, 32'h00000000} /* (31, 16, 0) {real, imag} */,
  {32'hc112b414, 32'h400fe061} /* (31, 15, 31) {real, imag} */,
  {32'h3f619fd8, 32'hc01e5058} /* (31, 15, 30) {real, imag} */,
  {32'hbfbe9c4c, 32'hc11a840d} /* (31, 15, 29) {real, imag} */,
  {32'h402f87ac, 32'hc085e8a5} /* (31, 15, 28) {real, imag} */,
  {32'h40191868, 32'h40442bb2} /* (31, 15, 27) {real, imag} */,
  {32'h40ec48b5, 32'h40833c0f} /* (31, 15, 26) {real, imag} */,
  {32'hc0a5a7ee, 32'hc08fa31e} /* (31, 15, 25) {real, imag} */,
  {32'hbfdbea20, 32'h3fb0d2f8} /* (31, 15, 24) {real, imag} */,
  {32'h405ad27c, 32'hc0ef4fdd} /* (31, 15, 23) {real, imag} */,
  {32'h3fdd7938, 32'h40d890eb} /* (31, 15, 22) {real, imag} */,
  {32'h40cbbabb, 32'hc0bb11bf} /* (31, 15, 21) {real, imag} */,
  {32'h3fd23c7f, 32'h410f67df} /* (31, 15, 20) {real, imag} */,
  {32'h3dce6b00, 32'hc08753f7} /* (31, 15, 19) {real, imag} */,
  {32'hc09f0069, 32'h4103ae12} /* (31, 15, 18) {real, imag} */,
  {32'h4045f59a, 32'hc0f8547c} /* (31, 15, 17) {real, imag} */,
  {32'h3f0a84ac, 32'h3fecb748} /* (31, 15, 16) {real, imag} */,
  {32'hbf318148, 32'hc0788808} /* (31, 15, 15) {real, imag} */,
  {32'h4000daef, 32'h41426d7a} /* (31, 15, 14) {real, imag} */,
  {32'hc08f8b84, 32'hc0981a4e} /* (31, 15, 13) {real, imag} */,
  {32'h406ae666, 32'h4115cad1} /* (31, 15, 12) {real, imag} */,
  {32'h4105b139, 32'hc0274b7c} /* (31, 15, 11) {real, imag} */,
  {32'hc08b75ea, 32'hbf9200e4} /* (31, 15, 10) {real, imag} */,
  {32'h40a20942, 32'h405f8dbe} /* (31, 15, 9) {real, imag} */,
  {32'hc0ef167a, 32'h3efa0940} /* (31, 15, 8) {real, imag} */,
  {32'h40a9fbe4, 32'hc1122d20} /* (31, 15, 7) {real, imag} */,
  {32'h40ae9c56, 32'h402f9e12} /* (31, 15, 6) {real, imag} */,
  {32'h401487ef, 32'h3fc3c96c} /* (31, 15, 5) {real, imag} */,
  {32'h3f53b3e0, 32'h406e7580} /* (31, 15, 4) {real, imag} */,
  {32'h3f814068, 32'h4025de1e} /* (31, 15, 3) {real, imag} */,
  {32'hbe5bfb60, 32'hc07ef370} /* (31, 15, 2) {real, imag} */,
  {32'h4074a53b, 32'h4084cc7a} /* (31, 15, 1) {real, imag} */,
  {32'hc08948b2, 32'hc09a678d} /* (31, 15, 0) {real, imag} */,
  {32'hc0f35f1a, 32'hc02968e9} /* (31, 14, 31) {real, imag} */,
  {32'h40bc42c3, 32'h40bb78df} /* (31, 14, 30) {real, imag} */,
  {32'hc0ac0c12, 32'hc0276470} /* (31, 14, 29) {real, imag} */,
  {32'hc1365b50, 32'hc019b62d} /* (31, 14, 28) {real, imag} */,
  {32'hc161b329, 32'h40c17294} /* (31, 14, 27) {real, imag} */,
  {32'h416e40ac, 32'h40b2cdec} /* (31, 14, 26) {real, imag} */,
  {32'h405e656c, 32'h40860b01} /* (31, 14, 25) {real, imag} */,
  {32'h401acde2, 32'hc0f27ffb} /* (31, 14, 24) {real, imag} */,
  {32'hc1074454, 32'h404751d2} /* (31, 14, 23) {real, imag} */,
  {32'h413a0946, 32'h4178b440} /* (31, 14, 22) {real, imag} */,
  {32'h3f9be65a, 32'hc0a3716b} /* (31, 14, 21) {real, imag} */,
  {32'hc111509c, 32'h4008059a} /* (31, 14, 20) {real, imag} */,
  {32'hc04ca990, 32'h41735c1c} /* (31, 14, 19) {real, imag} */,
  {32'hc0925510, 32'h3dba12a0} /* (31, 14, 18) {real, imag} */,
  {32'hc0b7c90e, 32'hc00fe72c} /* (31, 14, 17) {real, imag} */,
  {32'hc020b9a0, 32'h4104032c} /* (31, 14, 16) {real, imag} */,
  {32'hc097802f, 32'hbfc7bf90} /* (31, 14, 15) {real, imag} */,
  {32'h3ef086c0, 32'hc14eb670} /* (31, 14, 14) {real, imag} */,
  {32'h40501aa2, 32'h4163deb6} /* (31, 14, 13) {real, imag} */,
  {32'h3db1bcc0, 32'h4027ea2e} /* (31, 14, 12) {real, imag} */,
  {32'hc09bceac, 32'hbfe3da30} /* (31, 14, 11) {real, imag} */,
  {32'h411751a8, 32'h4031307c} /* (31, 14, 10) {real, imag} */,
  {32'h412f36b2, 32'h40682970} /* (31, 14, 9) {real, imag} */,
  {32'h40bb7a3a, 32'hbf017220} /* (31, 14, 8) {real, imag} */,
  {32'hc133f133, 32'h41b296e0} /* (31, 14, 7) {real, imag} */,
  {32'hc13b58ff, 32'h3fccc574} /* (31, 14, 6) {real, imag} */,
  {32'h412b6264, 32'h4117f7ec} /* (31, 14, 5) {real, imag} */,
  {32'h3fca79ae, 32'hc0ef80ca} /* (31, 14, 4) {real, imag} */,
  {32'h4103903f, 32'h40acb238} /* (31, 14, 3) {real, imag} */,
  {32'h40a93009, 32'h3ffe9298} /* (31, 14, 2) {real, imag} */,
  {32'h4101bf84, 32'hc08b7d9b} /* (31, 14, 1) {real, imag} */,
  {32'hc04ce2f7, 32'hc0742a7a} /* (31, 14, 0) {real, imag} */,
  {32'hc0d80b49, 32'hc0a4a311} /* (31, 13, 31) {real, imag} */,
  {32'hc166f562, 32'h404fa33c} /* (31, 13, 30) {real, imag} */,
  {32'h411e1c76, 32'hbe0577a8} /* (31, 13, 29) {real, imag} */,
  {32'h3da664c0, 32'h4020a082} /* (31, 13, 28) {real, imag} */,
  {32'h3f68bb7a, 32'hc11442a4} /* (31, 13, 27) {real, imag} */,
  {32'h409b2502, 32'hc127c662} /* (31, 13, 26) {real, imag} */,
  {32'hbefd8678, 32'hbfe37ce8} /* (31, 13, 25) {real, imag} */,
  {32'hc064bd6c, 32'hc0ed93fc} /* (31, 13, 24) {real, imag} */,
  {32'h402e39ce, 32'hc01df376} /* (31, 13, 23) {real, imag} */,
  {32'hbde82a60, 32'hc070add0} /* (31, 13, 22) {real, imag} */,
  {32'hc00bea62, 32'hc11ebb67} /* (31, 13, 21) {real, imag} */,
  {32'h4092d966, 32'hbf33c830} /* (31, 13, 20) {real, imag} */,
  {32'h4169b856, 32'h40d57d13} /* (31, 13, 19) {real, imag} */,
  {32'h41971075, 32'hc0c809a3} /* (31, 13, 18) {real, imag} */,
  {32'h40966334, 32'hc1027db3} /* (31, 13, 17) {real, imag} */,
  {32'hbfae0778, 32'h41266b70} /* (31, 13, 16) {real, imag} */,
  {32'hc0ad712a, 32'hbf0bea74} /* (31, 13, 15) {real, imag} */,
  {32'h40a60478, 32'h3e84a4ac} /* (31, 13, 14) {real, imag} */,
  {32'hc14929d3, 32'hc042d611} /* (31, 13, 13) {real, imag} */,
  {32'hc083d163, 32'h3e81be44} /* (31, 13, 12) {real, imag} */,
  {32'hc11ccd3e, 32'h409bca84} /* (31, 13, 11) {real, imag} */,
  {32'h3f9e061c, 32'h4017175f} /* (31, 13, 10) {real, imag} */,
  {32'h41251077, 32'hc0a3cb33} /* (31, 13, 9) {real, imag} */,
  {32'hc13c521a, 32'hbfffaf34} /* (31, 13, 8) {real, imag} */,
  {32'h4117f0f1, 32'hbf192d38} /* (31, 13, 7) {real, imag} */,
  {32'hc0347838, 32'h3fabb318} /* (31, 13, 6) {real, imag} */,
  {32'hc11c26dd, 32'hbfa4c24c} /* (31, 13, 5) {real, imag} */,
  {32'hc0ef1cd4, 32'h3ec9b078} /* (31, 13, 4) {real, imag} */,
  {32'hc0464b7b, 32'h40ab7c00} /* (31, 13, 3) {real, imag} */,
  {32'h3fab63d0, 32'hbf62140e} /* (31, 13, 2) {real, imag} */,
  {32'h40d81b6a, 32'hbfb1fd74} /* (31, 13, 1) {real, imag} */,
  {32'hc0fe0ebe, 32'hbf9b3684} /* (31, 13, 0) {real, imag} */,
  {32'h4000ec8a, 32'hc0a1efa1} /* (31, 12, 31) {real, imag} */,
  {32'h411c4160, 32'h410a4e9d} /* (31, 12, 30) {real, imag} */,
  {32'h40aad024, 32'hbfe399a8} /* (31, 12, 29) {real, imag} */,
  {32'hc10a7620, 32'hc173d52d} /* (31, 12, 28) {real, imag} */,
  {32'h409d1826, 32'hc0db0090} /* (31, 12, 27) {real, imag} */,
  {32'hbe894928, 32'hc096d987} /* (31, 12, 26) {real, imag} */,
  {32'h3f15e1c8, 32'h41682ee6} /* (31, 12, 25) {real, imag} */,
  {32'hc0d0279e, 32'hc13709e2} /* (31, 12, 24) {real, imag} */,
  {32'h3fccdd22, 32'hbf9f3a48} /* (31, 12, 23) {real, imag} */,
  {32'hbf83b0a0, 32'h41078050} /* (31, 12, 22) {real, imag} */,
  {32'h4118e874, 32'h4109367a} /* (31, 12, 21) {real, imag} */,
  {32'hc0e45933, 32'h4121384f} /* (31, 12, 20) {real, imag} */,
  {32'hc1850658, 32'hc0763ff8} /* (31, 12, 19) {real, imag} */,
  {32'hc16de012, 32'hbf174a9c} /* (31, 12, 18) {real, imag} */,
  {32'h40bde3ee, 32'hc0968084} /* (31, 12, 17) {real, imag} */,
  {32'h408742f1, 32'hc0311834} /* (31, 12, 16) {real, imag} */,
  {32'hc0f92e4c, 32'h4095de98} /* (31, 12, 15) {real, imag} */,
  {32'h4027b070, 32'h410028b7} /* (31, 12, 14) {real, imag} */,
  {32'hc178413e, 32'h409d2f8d} /* (31, 12, 13) {real, imag} */,
  {32'hc0a4d572, 32'h409b5ac0} /* (31, 12, 12) {real, imag} */,
  {32'h40cceeb6, 32'hc09d76f5} /* (31, 12, 11) {real, imag} */,
  {32'h40b589ae, 32'h41156562} /* (31, 12, 10) {real, imag} */,
  {32'hbd8d6120, 32'hc16156ec} /* (31, 12, 9) {real, imag} */,
  {32'h407f55dc, 32'h411a0719} /* (31, 12, 8) {real, imag} */,
  {32'hc108fbc3, 32'hc124c18d} /* (31, 12, 7) {real, imag} */,
  {32'h3eb58d80, 32'hc0ba8861} /* (31, 12, 6) {real, imag} */,
  {32'h3ee9c1c0, 32'hc0009b30} /* (31, 12, 5) {real, imag} */,
  {32'h3fd80b50, 32'hc084a77d} /* (31, 12, 4) {real, imag} */,
  {32'hc0d64c01, 32'h3e86f570} /* (31, 12, 3) {real, imag} */,
  {32'hc1589a43, 32'hbfa4cdc4} /* (31, 12, 2) {real, imag} */,
  {32'hc0543cf8, 32'h413f0ac8} /* (31, 12, 1) {real, imag} */,
  {32'h406c86e8, 32'h3fdee5a0} /* (31, 12, 0) {real, imag} */,
  {32'h4028efb0, 32'hc0cc6be4} /* (31, 11, 31) {real, imag} */,
  {32'hc0653658, 32'h41437cfc} /* (31, 11, 30) {real, imag} */,
  {32'h4020c944, 32'h40ad8e7a} /* (31, 11, 29) {real, imag} */,
  {32'hc105a598, 32'h41154e42} /* (31, 11, 28) {real, imag} */,
  {32'hbf60ec54, 32'h3e7ca8c0} /* (31, 11, 27) {real, imag} */,
  {32'hc04356a4, 32'hc0823a46} /* (31, 11, 26) {real, imag} */,
  {32'hc1814fd7, 32'h40888f4e} /* (31, 11, 25) {real, imag} */,
  {32'h408376c0, 32'hc100dec2} /* (31, 11, 24) {real, imag} */,
  {32'h3fcf8258, 32'h4182107c} /* (31, 11, 23) {real, imag} */,
  {32'hbed09060, 32'hbf7aff60} /* (31, 11, 22) {real, imag} */,
  {32'h4112f17d, 32'h41639db0} /* (31, 11, 21) {real, imag} */,
  {32'hc0be6374, 32'h40dbb608} /* (31, 11, 20) {real, imag} */,
  {32'hc07dc950, 32'hc176c5f8} /* (31, 11, 19) {real, imag} */,
  {32'hbec0bd30, 32'hc106079f} /* (31, 11, 18) {real, imag} */,
  {32'h3fe6146c, 32'h4055fabb} /* (31, 11, 17) {real, imag} */,
  {32'h3f7b1668, 32'h3f85a969} /* (31, 11, 16) {real, imag} */,
  {32'h3f1997e4, 32'hc00a0578} /* (31, 11, 15) {real, imag} */,
  {32'hc146cd51, 32'hbf82daf4} /* (31, 11, 14) {real, imag} */,
  {32'hc124ae6e, 32'hc0c3f882} /* (31, 11, 13) {real, imag} */,
  {32'hc0e8ec32, 32'hc1cddde0} /* (31, 11, 12) {real, imag} */,
  {32'h40b1c0c8, 32'h417db588} /* (31, 11, 11) {real, imag} */,
  {32'h419546ee, 32'h40fefc90} /* (31, 11, 10) {real, imag} */,
  {32'hc02c9ad2, 32'hbff942dc} /* (31, 11, 9) {real, imag} */,
  {32'h40c1b487, 32'hbf2dbd94} /* (31, 11, 8) {real, imag} */,
  {32'hc0e31f3a, 32'hc113480f} /* (31, 11, 7) {real, imag} */,
  {32'h3febae20, 32'h409bf936} /* (31, 11, 6) {real, imag} */,
  {32'h4107d1fd, 32'hc0fb2ea3} /* (31, 11, 5) {real, imag} */,
  {32'h40a5fa2a, 32'h415776c7} /* (31, 11, 4) {real, imag} */,
  {32'h4088b553, 32'hbfc2f370} /* (31, 11, 3) {real, imag} */,
  {32'hc0c33bf4, 32'h406b53c8} /* (31, 11, 2) {real, imag} */,
  {32'hc021a8e4, 32'h404a40bc} /* (31, 11, 1) {real, imag} */,
  {32'h400acf98, 32'hc0b02c98} /* (31, 11, 0) {real, imag} */,
  {32'hc037182e, 32'h4155751c} /* (31, 10, 31) {real, imag} */,
  {32'h3fc85468, 32'h40409008} /* (31, 10, 30) {real, imag} */,
  {32'hbf15a9f0, 32'h4076f8b6} /* (31, 10, 29) {real, imag} */,
  {32'h417aab8a, 32'hc05d56f4} /* (31, 10, 28) {real, imag} */,
  {32'hc04ce049, 32'hc1529c58} /* (31, 10, 27) {real, imag} */,
  {32'hbfed302c, 32'h41073d2c} /* (31, 10, 26) {real, imag} */,
  {32'hc03f5fa4, 32'hc0ebcc2c} /* (31, 10, 25) {real, imag} */,
  {32'hc0565b06, 32'hbfb05448} /* (31, 10, 24) {real, imag} */,
  {32'hc18732e3, 32'h4112e901} /* (31, 10, 23) {real, imag} */,
  {32'h413605f8, 32'hc028a82e} /* (31, 10, 22) {real, imag} */,
  {32'hc1591886, 32'hc0b57960} /* (31, 10, 21) {real, imag} */,
  {32'hc0cdc24c, 32'h4161f6d6} /* (31, 10, 20) {real, imag} */,
  {32'h3ff29148, 32'hc135247e} /* (31, 10, 19) {real, imag} */,
  {32'h40c9545a, 32'hc0ffc24c} /* (31, 10, 18) {real, imag} */,
  {32'hc0b83a84, 32'hc02bd4e2} /* (31, 10, 17) {real, imag} */,
  {32'hc0478fae, 32'h403b0c29} /* (31, 10, 16) {real, imag} */,
  {32'hbf0d18d3, 32'hbf15a1f8} /* (31, 10, 15) {real, imag} */,
  {32'hbfbeac1c, 32'hbf158a18} /* (31, 10, 14) {real, imag} */,
  {32'h3f1332f0, 32'h41526b2c} /* (31, 10, 13) {real, imag} */,
  {32'hc0d003ac, 32'h4142e57a} /* (31, 10, 12) {real, imag} */,
  {32'hc0a0c3c1, 32'hc084d479} /* (31, 10, 11) {real, imag} */,
  {32'hc11be0ba, 32'hbf267df0} /* (31, 10, 10) {real, imag} */,
  {32'h40c99dcc, 32'h41266e8c} /* (31, 10, 9) {real, imag} */,
  {32'hc04b8329, 32'hc09ed2ac} /* (31, 10, 8) {real, imag} */,
  {32'h410499a7, 32'h411ac8ae} /* (31, 10, 7) {real, imag} */,
  {32'hc0b2ae8a, 32'hc1280efc} /* (31, 10, 6) {real, imag} */,
  {32'h3ec17f20, 32'hc0a459bc} /* (31, 10, 5) {real, imag} */,
  {32'hbf821650, 32'h40d04090} /* (31, 10, 4) {real, imag} */,
  {32'h416fcaff, 32'hc09234fb} /* (31, 10, 3) {real, imag} */,
  {32'h3f292820, 32'hc1099ad6} /* (31, 10, 2) {real, imag} */,
  {32'h417b2137, 32'hc062948a} /* (31, 10, 1) {real, imag} */,
  {32'hc11b69de, 32'h3ff16ea6} /* (31, 10, 0) {real, imag} */,
  {32'hbf951e64, 32'h41b06eab} /* (31, 9, 31) {real, imag} */,
  {32'h403bd282, 32'h40f5aaae} /* (31, 9, 30) {real, imag} */,
  {32'h4153cc2b, 32'h40251eb4} /* (31, 9, 29) {real, imag} */,
  {32'h418b52f8, 32'h410fa040} /* (31, 9, 28) {real, imag} */,
  {32'h40f5c4d8, 32'hc0fe20d1} /* (31, 9, 27) {real, imag} */,
  {32'h4088c8e4, 32'h40e7a1cc} /* (31, 9, 26) {real, imag} */,
  {32'h402eeba3, 32'h3d242480} /* (31, 9, 25) {real, imag} */,
  {32'h400aae08, 32'hbfede7f4} /* (31, 9, 24) {real, imag} */,
  {32'hc0174a9c, 32'h3fbcfafe} /* (31, 9, 23) {real, imag} */,
  {32'h3da1e380, 32'h40928605} /* (31, 9, 22) {real, imag} */,
  {32'h40e4eb5c, 32'hc0ede0ce} /* (31, 9, 21) {real, imag} */,
  {32'h3fad2ad0, 32'hc08c6ea8} /* (31, 9, 20) {real, imag} */,
  {32'hc148ab2c, 32'hc0948950} /* (31, 9, 19) {real, imag} */,
  {32'hc0c72524, 32'hbfb68b96} /* (31, 9, 18) {real, imag} */,
  {32'h41194d99, 32'hc03ecb92} /* (31, 9, 17) {real, imag} */,
  {32'h3feb3254, 32'hbfe06e7c} /* (31, 9, 16) {real, imag} */,
  {32'h3fefa734, 32'hc037f21d} /* (31, 9, 15) {real, imag} */,
  {32'h40e63a16, 32'hbfc2c578} /* (31, 9, 14) {real, imag} */,
  {32'h4185fe52, 32'hbe3170a0} /* (31, 9, 13) {real, imag} */,
  {32'hbffbc24e, 32'hc1422173} /* (31, 9, 12) {real, imag} */,
  {32'h408f7852, 32'hbf232ec4} /* (31, 9, 11) {real, imag} */,
  {32'h404ac83a, 32'h401e7aaa} /* (31, 9, 10) {real, imag} */,
  {32'h4068b5d8, 32'hc135b0c7} /* (31, 9, 9) {real, imag} */,
  {32'hc0f0dc44, 32'hc13d8d9c} /* (31, 9, 8) {real, imag} */,
  {32'h41712da5, 32'hc0c8d34e} /* (31, 9, 7) {real, imag} */,
  {32'hc12282da, 32'hc07e8882} /* (31, 9, 6) {real, imag} */,
  {32'hc073cc42, 32'hbe0c8420} /* (31, 9, 5) {real, imag} */,
  {32'h4198b11b, 32'hbf4e8150} /* (31, 9, 4) {real, imag} */,
  {32'hc1d21346, 32'h40896349} /* (31, 9, 3) {real, imag} */,
  {32'hc07f7808, 32'hc184fa9e} /* (31, 9, 2) {real, imag} */,
  {32'h40cc622c, 32'hbf985c98} /* (31, 9, 1) {real, imag} */,
  {32'h3ee423a0, 32'h41298906} /* (31, 9, 0) {real, imag} */,
  {32'hc1d0e843, 32'hc1a4fb94} /* (31, 8, 31) {real, imag} */,
  {32'h42084781, 32'hc075c13c} /* (31, 8, 30) {real, imag} */,
  {32'hc0e482e0, 32'h3f6ce152} /* (31, 8, 29) {real, imag} */,
  {32'hc15f86e0, 32'h411cb912} /* (31, 8, 28) {real, imag} */,
  {32'h409bef4b, 32'h4060721f} /* (31, 8, 27) {real, imag} */,
  {32'hc15ea0ef, 32'hbf97d3d0} /* (31, 8, 26) {real, imag} */,
  {32'h40f2cd22, 32'hbe4eb150} /* (31, 8, 25) {real, imag} */,
  {32'hc0c92ac2, 32'hc0377b80} /* (31, 8, 24) {real, imag} */,
  {32'h4037007c, 32'h410f0ba4} /* (31, 8, 23) {real, imag} */,
  {32'h409babf0, 32'hc0d466b6} /* (31, 8, 22) {real, imag} */,
  {32'hc0e4b441, 32'h3f97b2cf} /* (31, 8, 21) {real, imag} */,
  {32'hbffdd8d0, 32'h4075aaaa} /* (31, 8, 20) {real, imag} */,
  {32'hc039c6be, 32'h4031a2e4} /* (31, 8, 19) {real, imag} */,
  {32'hc0b90fcc, 32'h409af45e} /* (31, 8, 18) {real, imag} */,
  {32'h410095c5, 32'h415d26c9} /* (31, 8, 17) {real, imag} */,
  {32'hbfc52614, 32'hc0526313} /* (31, 8, 16) {real, imag} */,
  {32'hbf8ba3a0, 32'hbfaa554a} /* (31, 8, 15) {real, imag} */,
  {32'h3fe91e8c, 32'h400c5802} /* (31, 8, 14) {real, imag} */,
  {32'h4088d7d6, 32'hbfe0e870} /* (31, 8, 13) {real, imag} */,
  {32'hbe836b80, 32'h41115e94} /* (31, 8, 12) {real, imag} */,
  {32'hc0d49f56, 32'h40ccf1b2} /* (31, 8, 11) {real, imag} */,
  {32'hbfab4bc4, 32'h41115521} /* (31, 8, 10) {real, imag} */,
  {32'h4028504e, 32'hc0878ba2} /* (31, 8, 9) {real, imag} */,
  {32'h3fd70de0, 32'hc0f56abe} /* (31, 8, 8) {real, imag} */,
  {32'hc0145f40, 32'hc13bd7cf} /* (31, 8, 7) {real, imag} */,
  {32'h412f152f, 32'h40974dd7} /* (31, 8, 6) {real, imag} */,
  {32'h3fe6175a, 32'h40ee92c0} /* (31, 8, 5) {real, imag} */,
  {32'h40c2184c, 32'h40c9c841} /* (31, 8, 4) {real, imag} */,
  {32'hc1c4b78b, 32'hbfee5298} /* (31, 8, 3) {real, imag} */,
  {32'h41594f0e, 32'h4214167c} /* (31, 8, 2) {real, imag} */,
  {32'hc19a969c, 32'hc16db412} /* (31, 8, 1) {real, imag} */,
  {32'hc1914c26, 32'h3cc21600} /* (31, 8, 0) {real, imag} */,
  {32'h40e7ff8e, 32'h3e5a9460} /* (31, 7, 31) {real, imag} */,
  {32'hc0b13a1e, 32'hc0a653c2} /* (31, 7, 30) {real, imag} */,
  {32'h3fe7df34, 32'hbf780128} /* (31, 7, 29) {real, imag} */,
  {32'hc15baf1b, 32'h3fc9e580} /* (31, 7, 28) {real, imag} */,
  {32'hc0f785e5, 32'hc0ce5842} /* (31, 7, 27) {real, imag} */,
  {32'h410a5bc2, 32'h40d82780} /* (31, 7, 26) {real, imag} */,
  {32'h40c79370, 32'hbfeb8a66} /* (31, 7, 25) {real, imag} */,
  {32'hc0c2e356, 32'h413c8bcd} /* (31, 7, 24) {real, imag} */,
  {32'h411f2d74, 32'h404b695e} /* (31, 7, 23) {real, imag} */,
  {32'hc08df467, 32'h3f1b1934} /* (31, 7, 22) {real, imag} */,
  {32'hbf88a6e0, 32'h4123dc38} /* (31, 7, 21) {real, imag} */,
  {32'hc10a01ef, 32'hc09af006} /* (31, 7, 20) {real, imag} */,
  {32'hbfe83328, 32'h40e44fbc} /* (31, 7, 19) {real, imag} */,
  {32'hc0a0c473, 32'h40c0fea0} /* (31, 7, 18) {real, imag} */,
  {32'h4166fd63, 32'h40b8346a} /* (31, 7, 17) {real, imag} */,
  {32'h4005a819, 32'hc034fd79} /* (31, 7, 16) {real, imag} */,
  {32'h4019860d, 32'h40b0dd6d} /* (31, 7, 15) {real, imag} */,
  {32'hc0f39be6, 32'h41110df6} /* (31, 7, 14) {real, imag} */,
  {32'hc0cdd438, 32'hc032e3e0} /* (31, 7, 13) {real, imag} */,
  {32'hbff19626, 32'hc0b1cac9} /* (31, 7, 12) {real, imag} */,
  {32'h4136823c, 32'h3ff50374} /* (31, 7, 11) {real, imag} */,
  {32'h40f8dbc1, 32'h3d141200} /* (31, 7, 10) {real, imag} */,
  {32'hc0d4eccd, 32'hc110d042} /* (31, 7, 9) {real, imag} */,
  {32'hc0b78ca5, 32'h40ac7309} /* (31, 7, 8) {real, imag} */,
  {32'h3f9a2034, 32'hbfb470e4} /* (31, 7, 7) {real, imag} */,
  {32'h40c1bab5, 32'hc0331082} /* (31, 7, 6) {real, imag} */,
  {32'h4109c6b4, 32'hbeac5f60} /* (31, 7, 5) {real, imag} */,
  {32'h409e1d5e, 32'hbf280c30} /* (31, 7, 4) {real, imag} */,
  {32'h411f2e3e, 32'h3ebc42c0} /* (31, 7, 3) {real, imag} */,
  {32'h41293268, 32'hc1165ef5} /* (31, 7, 2) {real, imag} */,
  {32'hc0fba278, 32'h3fdf8b58} /* (31, 7, 1) {real, imag} */,
  {32'h41bc68b9, 32'h415dbf4f} /* (31, 7, 0) {real, imag} */,
  {32'hc11e14ac, 32'h41990a00} /* (31, 6, 31) {real, imag} */,
  {32'hc1793ef2, 32'hc192f0bd} /* (31, 6, 30) {real, imag} */,
  {32'h415501e8, 32'h3f1024a0} /* (31, 6, 29) {real, imag} */,
  {32'hc0379818, 32'h40532e6a} /* (31, 6, 28) {real, imag} */,
  {32'hc0a40e4c, 32'h40c78610} /* (31, 6, 27) {real, imag} */,
  {32'h40f3b8d0, 32'h4185d8c4} /* (31, 6, 26) {real, imag} */,
  {32'hbfe73422, 32'hc073e94a} /* (31, 6, 25) {real, imag} */,
  {32'h40ae60dc, 32'h40d95abe} /* (31, 6, 24) {real, imag} */,
  {32'hc09a798c, 32'hc165a3df} /* (31, 6, 23) {real, imag} */,
  {32'h3fa39282, 32'hc1210a6a} /* (31, 6, 22) {real, imag} */,
  {32'h4122b3a2, 32'hc1495768} /* (31, 6, 21) {real, imag} */,
  {32'hc131d34a, 32'hbf00427a} /* (31, 6, 20) {real, imag} */,
  {32'hc1300fbd, 32'hbf5b33f8} /* (31, 6, 19) {real, imag} */,
  {32'h3f2bda52, 32'h40f84644} /* (31, 6, 18) {real, imag} */,
  {32'hc0b10418, 32'hc12579d2} /* (31, 6, 17) {real, imag} */,
  {32'h4063b9c0, 32'h3fd28bf4} /* (31, 6, 16) {real, imag} */,
  {32'h40acefb7, 32'h40db3ad6} /* (31, 6, 15) {real, imag} */,
  {32'h40281c76, 32'hc1447cdf} /* (31, 6, 14) {real, imag} */,
  {32'hc108d089, 32'hc1282d26} /* (31, 6, 13) {real, imag} */,
  {32'hc1192283, 32'h3f03d8ac} /* (31, 6, 12) {real, imag} */,
  {32'hbf7641e8, 32'h3e1e9700} /* (31, 6, 11) {real, imag} */,
  {32'hc0d41c83, 32'hc101bad7} /* (31, 6, 10) {real, imag} */,
  {32'h40894cfb, 32'hbe1c0a00} /* (31, 6, 9) {real, imag} */,
  {32'h415cb0f2, 32'h4109e8af} /* (31, 6, 8) {real, imag} */,
  {32'hc16b66f3, 32'h413550c5} /* (31, 6, 7) {real, imag} */,
  {32'hc0e9ead0, 32'hbf2e1798} /* (31, 6, 6) {real, imag} */,
  {32'h413e0844, 32'h4139b7c6} /* (31, 6, 5) {real, imag} */,
  {32'hc01133dc, 32'h40c43be0} /* (31, 6, 4) {real, imag} */,
  {32'h40a03cb0, 32'h4031741e} /* (31, 6, 3) {real, imag} */,
  {32'hbff42db6, 32'hc1ba80eb} /* (31, 6, 2) {real, imag} */,
  {32'hc18981a3, 32'hc088c332} /* (31, 6, 1) {real, imag} */,
  {32'h418b9ecc, 32'hc1094da7} /* (31, 6, 0) {real, imag} */,
  {32'hc24af712, 32'hc050c9e2} /* (31, 5, 31) {real, imag} */,
  {32'h410b8b90, 32'hc1894173} /* (31, 5, 30) {real, imag} */,
  {32'hc00cb030, 32'hc0dec44c} /* (31, 5, 29) {real, imag} */,
  {32'hbff8d7b2, 32'hc193d560} /* (31, 5, 28) {real, imag} */,
  {32'h41b5ed08, 32'hc0219d04} /* (31, 5, 27) {real, imag} */,
  {32'h405a5d36, 32'h405d2658} /* (31, 5, 26) {real, imag} */,
  {32'hc11f7293, 32'h4146d03c} /* (31, 5, 25) {real, imag} */,
  {32'hc0850512, 32'hbeab8fb0} /* (31, 5, 24) {real, imag} */,
  {32'h401d31ad, 32'h3fe35210} /* (31, 5, 23) {real, imag} */,
  {32'h40c89cda, 32'hc11036b4} /* (31, 5, 22) {real, imag} */,
  {32'hc0744fbb, 32'h414768a9} /* (31, 5, 21) {real, imag} */,
  {32'h415b75a4, 32'hc1322510} /* (31, 5, 20) {real, imag} */,
  {32'h40f76658, 32'hc009a787} /* (31, 5, 19) {real, imag} */,
  {32'h3f48afe8, 32'h408b4f34} /* (31, 5, 18) {real, imag} */,
  {32'hc04538e9, 32'hc03481fc} /* (31, 5, 17) {real, imag} */,
  {32'hc13eb538, 32'hbd5e6d00} /* (31, 5, 16) {real, imag} */,
  {32'hc070d2ba, 32'hc0cfe692} /* (31, 5, 15) {real, imag} */,
  {32'hc0f14d14, 32'h4094ddf8} /* (31, 5, 14) {real, imag} */,
  {32'hc0778f8c, 32'h40907087} /* (31, 5, 13) {real, imag} */,
  {32'h409ad9ac, 32'h40a615b6} /* (31, 5, 12) {real, imag} */,
  {32'hc15aee64, 32'hc0aa447c} /* (31, 5, 11) {real, imag} */,
  {32'h40506fff, 32'h4103cb71} /* (31, 5, 10) {real, imag} */,
  {32'h3fda6cb6, 32'h412e0e2d} /* (31, 5, 9) {real, imag} */,
  {32'hbfb1666c, 32'h413e995e} /* (31, 5, 8) {real, imag} */,
  {32'h41464126, 32'hc1a5b9b8} /* (31, 5, 7) {real, imag} */,
  {32'h4185fe23, 32'h40e9b1fe} /* (31, 5, 6) {real, imag} */,
  {32'h3fc7fd20, 32'h4123aa34} /* (31, 5, 5) {real, imag} */,
  {32'hc1cdd508, 32'hc0b3407b} /* (31, 5, 4) {real, imag} */,
  {32'hc1b6e6c7, 32'hc0d9bee6} /* (31, 5, 3) {real, imag} */,
  {32'h421e150c, 32'h41a2426c} /* (31, 5, 2) {real, imag} */,
  {32'hc21ae460, 32'hc20d72c8} /* (31, 5, 1) {real, imag} */,
  {32'hc23893cf, 32'h40d2dc80} /* (31, 5, 0) {real, imag} */,
  {32'h419c4ad8, 32'h42311866} /* (31, 4, 31) {real, imag} */,
  {32'hc28cd4ce, 32'hc0824a68} /* (31, 4, 30) {real, imag} */,
  {32'hc10fbb80, 32'h3db66200} /* (31, 4, 29) {real, imag} */,
  {32'h41e042af, 32'h40f156a7} /* (31, 4, 28) {real, imag} */,
  {32'hc18bfcda, 32'hc1851f03} /* (31, 4, 27) {real, imag} */,
  {32'hc121d585, 32'hc0fb82a8} /* (31, 4, 26) {real, imag} */,
  {32'hc107ea4e, 32'h3fe26a54} /* (31, 4, 25) {real, imag} */,
  {32'hc00fe500, 32'hc0c56b6c} /* (31, 4, 24) {real, imag} */,
  {32'hc10443ac, 32'h3fd3453e} /* (31, 4, 23) {real, imag} */,
  {32'h40f950e0, 32'h41609340} /* (31, 4, 22) {real, imag} */,
  {32'hc12e4620, 32'h40c0408f} /* (31, 4, 21) {real, imag} */,
  {32'h419eb55e, 32'hc1329cf9} /* (31, 4, 20) {real, imag} */,
  {32'h40cb28c2, 32'hbf0655f8} /* (31, 4, 19) {real, imag} */,
  {32'h408576ca, 32'hc095ebf1} /* (31, 4, 18) {real, imag} */,
  {32'h40645e95, 32'h4150588b} /* (31, 4, 17) {real, imag} */,
  {32'h3e8a9b1c, 32'hc05ee748} /* (31, 4, 16) {real, imag} */,
  {32'hc02c984a, 32'hc0a09fa2} /* (31, 4, 15) {real, imag} */,
  {32'h40b4afc2, 32'h4043539c} /* (31, 4, 14) {real, imag} */,
  {32'h416dec7a, 32'hc019efa9} /* (31, 4, 13) {real, imag} */,
  {32'h40e4a678, 32'hc1449646} /* (31, 4, 12) {real, imag} */,
  {32'h41255d38, 32'hc07b0a90} /* (31, 4, 11) {real, imag} */,
  {32'hc1483aa2, 32'h40882314} /* (31, 4, 10) {real, imag} */,
  {32'hc07d92de, 32'h40f2a6ac} /* (31, 4, 9) {real, imag} */,
  {32'hc10fa1f5, 32'h405ddcf8} /* (31, 4, 8) {real, imag} */,
  {32'h413c07ec, 32'h41346270} /* (31, 4, 7) {real, imag} */,
  {32'hbfdb1d20, 32'h4105cabc} /* (31, 4, 6) {real, imag} */,
  {32'h4149c876, 32'hc1bf98cf} /* (31, 4, 5) {real, imag} */,
  {32'hbeeed220, 32'h41ce1884} /* (31, 4, 4) {real, imag} */,
  {32'h40c4b08c, 32'h4180d07c} /* (31, 4, 3) {real, imag} */,
  {32'hc21d270a, 32'hc20f271f} /* (31, 4, 2) {real, imag} */,
  {32'h428b97f5, 32'h425b3f8b} /* (31, 4, 1) {real, imag} */,
  {32'h427929bb, 32'h41778e14} /* (31, 4, 0) {real, imag} */,
  {32'hc23608b6, 32'h41f72bdf} /* (31, 3, 31) {real, imag} */,
  {32'h41b3963e, 32'hc20d7a5d} /* (31, 3, 30) {real, imag} */,
  {32'h41e8cefa, 32'h3f8fbcf8} /* (31, 3, 29) {real, imag} */,
  {32'h40ce45fe, 32'h4187ec76} /* (31, 3, 28) {real, imag} */,
  {32'hc0adcfd6, 32'hc11d4a9e} /* (31, 3, 27) {real, imag} */,
  {32'hc0028ff6, 32'hc081c2d8} /* (31, 3, 26) {real, imag} */,
  {32'h40730f8c, 32'hbfacd130} /* (31, 3, 25) {real, imag} */,
  {32'h405299b0, 32'h40d6086c} /* (31, 3, 24) {real, imag} */,
  {32'hc101ca50, 32'h3ff97fac} /* (31, 3, 23) {real, imag} */,
  {32'h405ce6d2, 32'h40cb54ff} /* (31, 3, 22) {real, imag} */,
  {32'h3e90a1b8, 32'hc18a7893} /* (31, 3, 21) {real, imag} */,
  {32'hc029770b, 32'h3feb5224} /* (31, 3, 20) {real, imag} */,
  {32'h3ffeee6c, 32'hbf9dff84} /* (31, 3, 19) {real, imag} */,
  {32'h417cc18b, 32'hc15345b8} /* (31, 3, 18) {real, imag} */,
  {32'h40a39150, 32'hc061ab12} /* (31, 3, 17) {real, imag} */,
  {32'hc03d577a, 32'h40831819} /* (31, 3, 16) {real, imag} */,
  {32'hbffbca76, 32'hc02ced04} /* (31, 3, 15) {real, imag} */,
  {32'h410b7d17, 32'h41381d17} /* (31, 3, 14) {real, imag} */,
  {32'hc0e67c76, 32'hc0c9adce} /* (31, 3, 13) {real, imag} */,
  {32'hc11260de, 32'hc076e638} /* (31, 3, 12) {real, imag} */,
  {32'h4077c029, 32'hc11e2e57} /* (31, 3, 11) {real, imag} */,
  {32'hc13e0bff, 32'hc0f308ea} /* (31, 3, 10) {real, imag} */,
  {32'hc05561a2, 32'h40c77273} /* (31, 3, 9) {real, imag} */,
  {32'h4113b4ba, 32'hc1430222} /* (31, 3, 8) {real, imag} */,
  {32'hc11072bd, 32'h4083d25f} /* (31, 3, 7) {real, imag} */,
  {32'hc08a434c, 32'h40b4a165} /* (31, 3, 6) {real, imag} */,
  {32'hc1cfc8b4, 32'h417dcb73} /* (31, 3, 5) {real, imag} */,
  {32'hc0cf0708, 32'h40cfc6d6} /* (31, 3, 4) {real, imag} */,
  {32'h41bd52ca, 32'hc13569dc} /* (31, 3, 3) {real, imag} */,
  {32'hc1bbf5ae, 32'hc1b43a34} /* (31, 3, 2) {real, imag} */,
  {32'h421bedbb, 32'hbf2e9a40} /* (31, 3, 1) {real, imag} */,
  {32'h408c0d34, 32'h41a5b2a1} /* (31, 3, 0) {real, imag} */,
  {32'hc36f6960, 32'hc24168f2} /* (31, 2, 31) {real, imag} */,
  {32'h43019d18, 32'hc2949812} /* (31, 2, 30) {real, imag} */,
  {32'h3facdf70, 32'h40aeaf80} /* (31, 2, 29) {real, imag} */,
  {32'hc23fda9e, 32'h424d1a50} /* (31, 2, 28) {real, imag} */,
  {32'h41ed2bd4, 32'h3f8c53b0} /* (31, 2, 27) {real, imag} */,
  {32'h40ea6cf8, 32'h41038de6} /* (31, 2, 26) {real, imag} */,
  {32'hc08a9e1e, 32'hc09fd663} /* (31, 2, 25) {real, imag} */,
  {32'h419b96c1, 32'hc0fb7fe6} /* (31, 2, 24) {real, imag} */,
  {32'h412b479c, 32'h400c3dfa} /* (31, 2, 23) {real, imag} */,
  {32'hc172f0ec, 32'hbf0e8310} /* (31, 2, 22) {real, imag} */,
  {32'h4162f668, 32'hc0e1515c} /* (31, 2, 21) {real, imag} */,
  {32'hbfa3ec68, 32'h3fae130e} /* (31, 2, 20) {real, imag} */,
  {32'h4162f04c, 32'h40819754} /* (31, 2, 19) {real, imag} */,
  {32'hc06ba101, 32'hbfe6c780} /* (31, 2, 18) {real, imag} */,
  {32'h4109e9f6, 32'hbfc4be64} /* (31, 2, 17) {real, imag} */,
  {32'hbee31124, 32'hbf4d4240} /* (31, 2, 16) {real, imag} */,
  {32'hc106fac4, 32'hc01b8682} /* (31, 2, 15) {real, imag} */,
  {32'h41095751, 32'h4148427a} /* (31, 2, 14) {real, imag} */,
  {32'h40409b1c, 32'hbfcf5d8a} /* (31, 2, 13) {real, imag} */,
  {32'h40dc355c, 32'h40cdd14b} /* (31, 2, 12) {real, imag} */,
  {32'hbfb4c15e, 32'h40e9df0e} /* (31, 2, 11) {real, imag} */,
  {32'hbfd9caf4, 32'h3d9b3b10} /* (31, 2, 10) {real, imag} */,
  {32'hc118dfc2, 32'h413158fd} /* (31, 2, 9) {real, imag} */,
  {32'h41ef2bee, 32'h40d2222c} /* (31, 2, 8) {real, imag} */,
  {32'hc12bb2f7, 32'hc14b5111} /* (31, 2, 7) {real, imag} */,
  {32'h40897e56, 32'h412ed806} /* (31, 2, 6) {real, imag} */,
  {32'h41530186, 32'h40737260} /* (31, 2, 5) {real, imag} */,
  {32'hc1b6511c, 32'h412337df} /* (31, 2, 4) {real, imag} */,
  {32'hc1a0ac18, 32'hc200c31b} /* (31, 2, 3) {real, imag} */,
  {32'h42dd3696, 32'h40d124e8} /* (31, 2, 2) {real, imag} */,
  {32'hc3499a5c, 32'h42bd7840} /* (31, 2, 1) {real, imag} */,
  {32'hc3276984, 32'hc1ad4ce4} /* (31, 2, 0) {real, imag} */,
  {32'h438493cc, 32'hc2b80d32} /* (31, 1, 31) {real, imag} */,
  {32'hc2ef09e9, 32'h41182aed} /* (31, 1, 30) {real, imag} */,
  {32'hc11bf57e, 32'h4125fb3a} /* (31, 1, 29) {real, imag} */,
  {32'h421a1c02, 32'hc10caad7} /* (31, 1, 28) {real, imag} */,
  {32'hc1d80064, 32'h405a9e8c} /* (31, 1, 27) {real, imag} */,
  {32'hbfb810a0, 32'h3fffde38} /* (31, 1, 26) {real, imag} */,
  {32'h409b413c, 32'hc16214f5} /* (31, 1, 25) {real, imag} */,
  {32'hc1806408, 32'hc0ce4434} /* (31, 1, 24) {real, imag} */,
  {32'hc18af551, 32'hbf9eae88} /* (31, 1, 23) {real, imag} */,
  {32'h4030aed2, 32'hbfdba0ce} /* (31, 1, 22) {real, imag} */,
  {32'hc0b47e5f, 32'h40d40cf9} /* (31, 1, 21) {real, imag} */,
  {32'h4162982f, 32'h4184c0fc} /* (31, 1, 20) {real, imag} */,
  {32'hc18ff067, 32'h411a0dd8} /* (31, 1, 19) {real, imag} */,
  {32'h3f9663be, 32'h40bf7cac} /* (31, 1, 18) {real, imag} */,
  {32'hc03376be, 32'h40ebb03b} /* (31, 1, 17) {real, imag} */,
  {32'hc0956dda, 32'h4068c794} /* (31, 1, 16) {real, imag} */,
  {32'h3fce1af4, 32'h41359f0a} /* (31, 1, 15) {real, imag} */,
  {32'hc113965f, 32'hc11959cb} /* (31, 1, 14) {real, imag} */,
  {32'h40754597, 32'h41920d4f} /* (31, 1, 13) {real, imag} */,
  {32'h40b9e30e, 32'h40d4cb9f} /* (31, 1, 12) {real, imag} */,
  {32'hc13e7cb9, 32'h3ffc6964} /* (31, 1, 11) {real, imag} */,
  {32'hc0a1aa6b, 32'hbfe88044} /* (31, 1, 10) {real, imag} */,
  {32'h40befc4c, 32'hc16eb4a8} /* (31, 1, 9) {real, imag} */,
  {32'h40aeb782, 32'hc1dd0b00} /* (31, 1, 8) {real, imag} */,
  {32'h4034c462, 32'h41a033b4} /* (31, 1, 7) {real, imag} */,
  {32'hc0fabd28, 32'hc0531204} /* (31, 1, 6) {real, imag} */,
  {32'hc1c19ccd, 32'hc19e7756} /* (31, 1, 5) {real, imag} */,
  {32'h42119b1d, 32'hc1a57278} /* (31, 1, 4) {real, imag} */,
  {32'h41362f1c, 32'h4213848f} /* (31, 1, 3) {real, imag} */,
  {32'hc30daf0d, 32'hc332027c} /* (31, 1, 2) {real, imag} */,
  {32'h439dee52, 32'h42938702} /* (31, 1, 1) {real, imag} */,
  {32'h4326c852, 32'h42bb7234} /* (31, 1, 0) {real, imag} */,
  {32'h42e591e2, 32'hc302af47} /* (31, 0, 31) {real, imag} */,
  {32'hc2939901, 32'h42f35c40} /* (31, 0, 30) {real, imag} */,
  {32'hc0728870, 32'h419941c4} /* (31, 0, 29) {real, imag} */,
  {32'hc180970b, 32'h408278d0} /* (31, 0, 28) {real, imag} */,
  {32'h4026e590, 32'hbf8108d8} /* (31, 0, 27) {real, imag} */,
  {32'hc17c997b, 32'h40382b37} /* (31, 0, 26) {real, imag} */,
  {32'hc1105c1e, 32'hc1c942cd} /* (31, 0, 25) {real, imag} */,
  {32'h407e83b0, 32'h400c4b38} /* (31, 0, 24) {real, imag} */,
  {32'hc1460724, 32'h40e9cb32} /* (31, 0, 23) {real, imag} */,
  {32'h4097e8f4, 32'hc12d2e0a} /* (31, 0, 22) {real, imag} */,
  {32'hc1881b3d, 32'h4014ba00} /* (31, 0, 21) {real, imag} */,
  {32'hc12edbb8, 32'hbf78b388} /* (31, 0, 20) {real, imag} */,
  {32'hc05cd052, 32'hc13145fc} /* (31, 0, 19) {real, imag} */,
  {32'h40f135b3, 32'h4024c5c0} /* (31, 0, 18) {real, imag} */,
  {32'h3f4ba7d8, 32'h40e49236} /* (31, 0, 17) {real, imag} */,
  {32'h40cc8415, 32'h00000000} /* (31, 0, 16) {real, imag} */,
  {32'h3f4ba7d8, 32'hc0e49236} /* (31, 0, 15) {real, imag} */,
  {32'h40f135b3, 32'hc024c5c0} /* (31, 0, 14) {real, imag} */,
  {32'hc05cd052, 32'h413145fc} /* (31, 0, 13) {real, imag} */,
  {32'hc12edbb8, 32'h3f78b388} /* (31, 0, 12) {real, imag} */,
  {32'hc1881b3d, 32'hc014ba00} /* (31, 0, 11) {real, imag} */,
  {32'h4097e8f4, 32'h412d2e0a} /* (31, 0, 10) {real, imag} */,
  {32'hc1460724, 32'hc0e9cb32} /* (31, 0, 9) {real, imag} */,
  {32'h407e83b0, 32'hc00c4b38} /* (31, 0, 8) {real, imag} */,
  {32'hc1105c1e, 32'h41c942cd} /* (31, 0, 7) {real, imag} */,
  {32'hc17c997b, 32'hc0382b37} /* (31, 0, 6) {real, imag} */,
  {32'h4026e590, 32'h3f8108d8} /* (31, 0, 5) {real, imag} */,
  {32'hc180970b, 32'hc08278d0} /* (31, 0, 4) {real, imag} */,
  {32'hc0728870, 32'hc19941c4} /* (31, 0, 3) {real, imag} */,
  {32'hc2939901, 32'hc2f35c40} /* (31, 0, 2) {real, imag} */,
  {32'h42e591e2, 32'h4302af47} /* (31, 0, 1) {real, imag} */,
  {32'h3fa82280, 32'h00000000} /* (31, 0, 0) {real, imag} */,
  {32'h44421f17, 32'hc3a27cc4} /* (30, 31, 31) {real, imag} */,
  {32'hc39e4521, 32'h43b0ccd0} /* (30, 31, 30) {real, imag} */,
  {32'hc1d471d1, 32'hc2625256} /* (30, 31, 29) {real, imag} */,
  {32'h4219e16e, 32'hc0417f90} /* (30, 31, 28) {real, imag} */,
  {32'hc2b8d91a, 32'h4213a988} /* (30, 31, 27) {real, imag} */,
  {32'hc1b2c782, 32'hc1b59bb4} /* (30, 31, 26) {real, imag} */,
  {32'hc17184f2, 32'hc193b1cb} /* (30, 31, 25) {real, imag} */,
  {32'h3f863858, 32'h42527a4a} /* (30, 31, 24) {real, imag} */,
  {32'h4198db4c, 32'hc139a8f2} /* (30, 31, 23) {real, imag} */,
  {32'hc13f4064, 32'hc07e9342} /* (30, 31, 22) {real, imag} */,
  {32'hbf325a50, 32'h4129db26} /* (30, 31, 21) {real, imag} */,
  {32'h4179c11e, 32'h409b6199} /* (30, 31, 20) {real, imag} */,
  {32'h408fc74a, 32'hc195c9ad} /* (30, 31, 19) {real, imag} */,
  {32'hc079a088, 32'h40e6a9ed} /* (30, 31, 18) {real, imag} */,
  {32'hc1589c5c, 32'h3f88bd24} /* (30, 31, 17) {real, imag} */,
  {32'h3fea57ea, 32'hbe916758} /* (30, 31, 16) {real, imag} */,
  {32'h4063144b, 32'h40a5d5b4} /* (30, 31, 15) {real, imag} */,
  {32'hc1454006, 32'hc18c791b} /* (30, 31, 14) {real, imag} */,
  {32'h40a4a62a, 32'hc0207b78} /* (30, 31, 13) {real, imag} */,
  {32'h412f6794, 32'hbf1b6f90} /* (30, 31, 12) {real, imag} */,
  {32'hc0f7277c, 32'hc215520f} /* (30, 31, 11) {real, imag} */,
  {32'h41265ee8, 32'h41541d05} /* (30, 31, 10) {real, imag} */,
  {32'hc16073d7, 32'h3fe6efc4} /* (30, 31, 9) {real, imag} */,
  {32'hc1244c3c, 32'hc20901d8} /* (30, 31, 8) {real, imag} */,
  {32'h41816a50, 32'h42075831} /* (30, 31, 7) {real, imag} */,
  {32'hc1896380, 32'h41993bbc} /* (30, 31, 6) {real, imag} */,
  {32'hc29085d0, 32'h405918e3} /* (30, 31, 5) {real, imag} */,
  {32'h4258ebff, 32'hc15a0434} /* (30, 31, 4) {real, imag} */,
  {32'hc1b856be, 32'hc00f5720} /* (30, 31, 3) {real, imag} */,
  {32'hc368e09c, 32'hc1c6c33f} /* (30, 31, 2) {real, imag} */,
  {32'h440cc7f4, 32'h431c48f1} /* (30, 31, 1) {real, imag} */,
  {32'h43ea7508, 32'hc2dc2030} /* (30, 31, 0) {real, imag} */,
  {32'hc3cc7bde, 32'hc314ae16} /* (30, 30, 31) {real, imag} */,
  {32'h43604551, 32'h41a7d804} /* (30, 30, 30) {real, imag} */,
  {32'hc213b24c, 32'h421ef420} /* (30, 30, 29) {real, imag} */,
  {32'hc24a1882, 32'hc101c8f0} /* (30, 30, 28) {real, imag} */,
  {32'h424c8b2c, 32'hc144d83c} /* (30, 30, 27) {real, imag} */,
  {32'h4033ab24, 32'hc14a03fe} /* (30, 30, 26) {real, imag} */,
  {32'h40e13ed8, 32'h41aea44b} /* (30, 30, 25) {real, imag} */,
  {32'h4114623a, 32'hc04c80cc} /* (30, 30, 24) {real, imag} */,
  {32'h4190a162, 32'hc000af9b} /* (30, 30, 23) {real, imag} */,
  {32'h3d01ad00, 32'h41288ab8} /* (30, 30, 22) {real, imag} */,
  {32'h41d159aa, 32'hc20343f8} /* (30, 30, 21) {real, imag} */,
  {32'h3f15ef50, 32'h41491cc6} /* (30, 30, 20) {real, imag} */,
  {32'hc1296c5a, 32'h3f36d1be} /* (30, 30, 19) {real, imag} */,
  {32'hbeff0570, 32'h3f91b640} /* (30, 30, 18) {real, imag} */,
  {32'hc10ddf8d, 32'hc0248edc} /* (30, 30, 17) {real, imag} */,
  {32'h402f37a3, 32'hc078583c} /* (30, 30, 16) {real, imag} */,
  {32'h411e51fd, 32'h40ece93b} /* (30, 30, 15) {real, imag} */,
  {32'hc091d9f6, 32'h417a90a0} /* (30, 30, 14) {real, imag} */,
  {32'hc01dc810, 32'h40afe492} /* (30, 30, 13) {real, imag} */,
  {32'hc04d99d1, 32'hc1707dc8} /* (30, 30, 12) {real, imag} */,
  {32'hc0a974d3, 32'h4173507e} /* (30, 30, 11) {real, imag} */,
  {32'hc125b02e, 32'hc08b10c2} /* (30, 30, 10) {real, imag} */,
  {32'h3f4a5ee0, 32'hc0cd3253} /* (30, 30, 9) {real, imag} */,
  {32'h422e19b9, 32'h41264456} /* (30, 30, 8) {real, imag} */,
  {32'hc135bba6, 32'h40e836ca} /* (30, 30, 7) {real, imag} */,
  {32'h418ee529, 32'hc10e4f4a} /* (30, 30, 6) {real, imag} */,
  {32'h4236c4f6, 32'h411f778e} /* (30, 30, 5) {real, imag} */,
  {32'hc24c6cd7, 32'hc2b5afd4} /* (30, 30, 4) {real, imag} */,
  {32'h42171962, 32'hc03e4ad4} /* (30, 30, 3) {real, imag} */,
  {32'h439c9632, 32'h42f2ba10} /* (30, 30, 2) {real, imag} */,
  {32'hc41425c8, 32'h428b522d} /* (30, 30, 1) {real, imag} */,
  {32'hc3a6596a, 32'h42016126} /* (30, 30, 0) {real, imag} */,
  {32'h42621b78, 32'hc25d548c} /* (30, 29, 31) {real, imag} */,
  {32'hc0d39334, 32'h428bb6a3} /* (30, 29, 30) {real, imag} */,
  {32'h41d4574d, 32'hc0410af0} /* (30, 29, 29) {real, imag} */,
  {32'hc0e8d1cc, 32'hc195f5e1} /* (30, 29, 28) {real, imag} */,
  {32'hc1ddf5c5, 32'hc18f1870} /* (30, 29, 27) {real, imag} */,
  {32'hbf7a5d40, 32'hc098577e} /* (30, 29, 26) {real, imag} */,
  {32'h41bd5a26, 32'hc105a390} /* (30, 29, 25) {real, imag} */,
  {32'hc0625cf7, 32'h40abeb4c} /* (30, 29, 24) {real, imag} */,
  {32'h4095c2aa, 32'hc0c7d443} /* (30, 29, 23) {real, imag} */,
  {32'hc191b68a, 32'h417e70c3} /* (30, 29, 22) {real, imag} */,
  {32'hc1164c3f, 32'hc14198a1} /* (30, 29, 21) {real, imag} */,
  {32'hc0a2c39c, 32'h40e08925} /* (30, 29, 20) {real, imag} */,
  {32'h414d5ac8, 32'hc11b256e} /* (30, 29, 19) {real, imag} */,
  {32'hbf84a0f0, 32'h3fb25bc0} /* (30, 29, 18) {real, imag} */,
  {32'h4025959d, 32'hc06b5d44} /* (30, 29, 17) {real, imag} */,
  {32'hbd51b640, 32'h417fa722} /* (30, 29, 16) {real, imag} */,
  {32'h40b20d94, 32'h409062ce} /* (30, 29, 15) {real, imag} */,
  {32'h3ffa41db, 32'hbfb0baf8} /* (30, 29, 14) {real, imag} */,
  {32'hc0adddc2, 32'hc0e6501a} /* (30, 29, 13) {real, imag} */,
  {32'hc17ad778, 32'hc01371e4} /* (30, 29, 12) {real, imag} */,
  {32'hc14dbfc9, 32'hc08d0915} /* (30, 29, 11) {real, imag} */,
  {32'hbc7cf580, 32'hc12c0f0b} /* (30, 29, 10) {real, imag} */,
  {32'h3f5d1d40, 32'hc040569c} /* (30, 29, 9) {real, imag} */,
  {32'hc11da3a4, 32'h3eede760} /* (30, 29, 8) {real, imag} */,
  {32'hc11fd18d, 32'hc1177b6e} /* (30, 29, 7) {real, imag} */,
  {32'h402cf338, 32'h409d30f0} /* (30, 29, 6) {real, imag} */,
  {32'h40b148a3, 32'h419bf8b4} /* (30, 29, 5) {real, imag} */,
  {32'h402db324, 32'hc1acd2ee} /* (30, 29, 4) {real, imag} */,
  {32'h4138d2b4, 32'hc138d840} /* (30, 29, 3) {real, imag} */,
  {32'h426322f8, 32'h429a2415} /* (30, 29, 2) {real, imag} */,
  {32'hc2b6eec5, 32'hc29606d2} /* (30, 29, 1) {real, imag} */,
  {32'hc13fa95e, 32'hc197dbf8} /* (30, 29, 0) {real, imag} */,
  {32'h4300b95a, 32'hc28a6147} /* (30, 28, 31) {real, imag} */,
  {32'hc2212f4a, 32'h42918674} /* (30, 28, 30) {real, imag} */,
  {32'h40c3c42e, 32'hc186919d} /* (30, 28, 29) {real, imag} */,
  {32'hc00600f4, 32'hc1ecb9e9} /* (30, 28, 28) {real, imag} */,
  {32'h417df056, 32'h41d8f569} /* (30, 28, 27) {real, imag} */,
  {32'hbeca2cf0, 32'h410da080} /* (30, 28, 26) {real, imag} */,
  {32'h41a79a69, 32'hc1e04ac4} /* (30, 28, 25) {real, imag} */,
  {32'hbf91c210, 32'hc0f111a4} /* (30, 28, 24) {real, imag} */,
  {32'h419798d1, 32'h3f754592} /* (30, 28, 23) {real, imag} */,
  {32'hc19261bf, 32'hc1c50aba} /* (30, 28, 22) {real, imag} */,
  {32'h41351043, 32'h40f0734c} /* (30, 28, 21) {real, imag} */,
  {32'hbe7523d0, 32'h4132ec21} /* (30, 28, 20) {real, imag} */,
  {32'h41043fae, 32'h4081e9d0} /* (30, 28, 19) {real, imag} */,
  {32'hc06cddf0, 32'h402f1f6c} /* (30, 28, 18) {real, imag} */,
  {32'h407835ca, 32'h3f77d3c0} /* (30, 28, 17) {real, imag} */,
  {32'hc12f5a5c, 32'h3f50cb5e} /* (30, 28, 16) {real, imag} */,
  {32'h40a4b966, 32'h4023b0fc} /* (30, 28, 15) {real, imag} */,
  {32'h403b39a8, 32'hc127093e} /* (30, 28, 14) {real, imag} */,
  {32'h4073f710, 32'hc05b3409} /* (30, 28, 13) {real, imag} */,
  {32'h4052ee7b, 32'h412a1db6} /* (30, 28, 12) {real, imag} */,
  {32'hc18f906e, 32'hc111c2d4} /* (30, 28, 11) {real, imag} */,
  {32'h417cc0b4, 32'h400e9a2c} /* (30, 28, 10) {real, imag} */,
  {32'h41388d6a, 32'hc0aed6cc} /* (30, 28, 9) {real, imag} */,
  {32'hc0147ad1, 32'h4040b6f4} /* (30, 28, 8) {real, imag} */,
  {32'hc1670735, 32'h40855dcf} /* (30, 28, 7) {real, imag} */,
  {32'hbdd56980, 32'hbeebd640} /* (30, 28, 6) {real, imag} */,
  {32'hc1f31231, 32'h414c2f3e} /* (30, 28, 5) {real, imag} */,
  {32'h420456f6, 32'hc1bfa27a} /* (30, 28, 4) {real, imag} */,
  {32'hc0f43d2a, 32'hc1eaa4fc} /* (30, 28, 3) {real, imag} */,
  {32'hc2be70cc, 32'h4068fcf0} /* (30, 28, 2) {real, imag} */,
  {32'h42608b95, 32'hc2820672} /* (30, 28, 1) {real, imag} */,
  {32'h4288bf4e, 32'hc1a9079d} /* (30, 28, 0) {real, imag} */,
  {32'hc2685825, 32'h4284576e} /* (30, 27, 31) {real, imag} */,
  {32'h424840ea, 32'hc2197758} /* (30, 27, 30) {real, imag} */,
  {32'hc087ca4c, 32'h3df14fc0} /* (30, 27, 29) {real, imag} */,
  {32'hc19401c5, 32'h419075ac} /* (30, 27, 28) {real, imag} */,
  {32'hc16ecd65, 32'hc18397dc} /* (30, 27, 27) {real, imag} */,
  {32'h4188efa0, 32'h3fd322ec} /* (30, 27, 26) {real, imag} */,
  {32'h415540df, 32'h41760a79} /* (30, 27, 25) {real, imag} */,
  {32'hc11cf8d5, 32'hc15de052} /* (30, 27, 24) {real, imag} */,
  {32'h4084106e, 32'hc1856184} /* (30, 27, 23) {real, imag} */,
  {32'hbfd81dea, 32'hc0722fb6} /* (30, 27, 22) {real, imag} */,
  {32'hc1a9fc6d, 32'hc02c69c4} /* (30, 27, 21) {real, imag} */,
  {32'hc03c5990, 32'hc17987d1} /* (30, 27, 20) {real, imag} */,
  {32'h40fa1402, 32'hbec4d0c0} /* (30, 27, 19) {real, imag} */,
  {32'h3fc183de, 32'hc0e235ca} /* (30, 27, 18) {real, imag} */,
  {32'hc09e57c3, 32'hbfc5a6f4} /* (30, 27, 17) {real, imag} */,
  {32'hc044c6d9, 32'hc0597a15} /* (30, 27, 16) {real, imag} */,
  {32'hc0820c95, 32'h3fdb1ac2} /* (30, 27, 15) {real, imag} */,
  {32'hc107ba82, 32'h3f37e630} /* (30, 27, 14) {real, imag} */,
  {32'h40924e91, 32'h405b4768} /* (30, 27, 13) {real, imag} */,
  {32'hc09a1fad, 32'h407e8696} /* (30, 27, 12) {real, imag} */,
  {32'h40b9d914, 32'h3f669868} /* (30, 27, 11) {real, imag} */,
  {32'h3fce1470, 32'h41e86c70} /* (30, 27, 10) {real, imag} */,
  {32'hc1513b06, 32'h4108c0c7} /* (30, 27, 9) {real, imag} */,
  {32'hc0201f6e, 32'hc18ab02e} /* (30, 27, 8) {real, imag} */,
  {32'hc1b76f45, 32'hc130e778} /* (30, 27, 7) {real, imag} */,
  {32'hc0f84284, 32'hc01ea044} /* (30, 27, 6) {real, imag} */,
  {32'h41d5bf3b, 32'h400f45c6} /* (30, 27, 5) {real, imag} */,
  {32'h4124fc64, 32'hc1545c23} /* (30, 27, 4) {real, imag} */,
  {32'h4092d792, 32'h40928776} /* (30, 27, 3) {real, imag} */,
  {32'h41b82820, 32'h420b0019} /* (30, 27, 2) {real, imag} */,
  {32'hc29f0a5e, 32'h4150e478} /* (30, 27, 1) {real, imag} */,
  {32'hc291a4a3, 32'hc0eb5d26} /* (30, 27, 0) {real, imag} */,
  {32'hc21b5ed5, 32'h4112e702} /* (30, 26, 31) {real, imag} */,
  {32'h403392c0, 32'h414b219a} /* (30, 26, 30) {real, imag} */,
  {32'hc11d94b9, 32'hc104dd62} /* (30, 26, 29) {real, imag} */,
  {32'h4158ef52, 32'hbf82cc2c} /* (30, 26, 28) {real, imag} */,
  {32'h41b200d6, 32'hc12e0121} /* (30, 26, 27) {real, imag} */,
  {32'hc180f4e0, 32'hc166e546} /* (30, 26, 26) {real, imag} */,
  {32'h4013c534, 32'hc123cba9} /* (30, 26, 25) {real, imag} */,
  {32'h4090d4ec, 32'hc064432c} /* (30, 26, 24) {real, imag} */,
  {32'hc16c06c4, 32'hc108b9da} /* (30, 26, 23) {real, imag} */,
  {32'h40723bd8, 32'h4188211b} /* (30, 26, 22) {real, imag} */,
  {32'h40362000, 32'h40de3954} /* (30, 26, 21) {real, imag} */,
  {32'hc15475ce, 32'h40b759a2} /* (30, 26, 20) {real, imag} */,
  {32'h4089b9b2, 32'hc0d2a89b} /* (30, 26, 19) {real, imag} */,
  {32'h403d65c1, 32'hc09ffa9c} /* (30, 26, 18) {real, imag} */,
  {32'hc0cf65f8, 32'hc0865fbc} /* (30, 26, 17) {real, imag} */,
  {32'h41006c63, 32'h40cb91b6} /* (30, 26, 16) {real, imag} */,
  {32'hc00535b6, 32'h4128c4b4} /* (30, 26, 15) {real, imag} */,
  {32'h41813200, 32'hc12d4bfe} /* (30, 26, 14) {real, imag} */,
  {32'hc1a4ee8c, 32'h416aadce} /* (30, 26, 13) {real, imag} */,
  {32'hc182fe59, 32'hc0c346d2} /* (30, 26, 12) {real, imag} */,
  {32'hc1160f55, 32'hbff131b8} /* (30, 26, 11) {real, imag} */,
  {32'h40641684, 32'h3fe6d9a0} /* (30, 26, 10) {real, imag} */,
  {32'hbf8a9284, 32'h408fc940} /* (30, 26, 9) {real, imag} */,
  {32'h418ad94a, 32'h4169030b} /* (30, 26, 8) {real, imag} */,
  {32'h3f8cef84, 32'h3fa59848} /* (30, 26, 7) {real, imag} */,
  {32'h4131d327, 32'hc1ae08e8} /* (30, 26, 6) {real, imag} */,
  {32'h3fb770f2, 32'hc10c30b1} /* (30, 26, 5) {real, imag} */,
  {32'hbfd80430, 32'h3fe085c0} /* (30, 26, 4) {real, imag} */,
  {32'h405b73e8, 32'h41a8213e} /* (30, 26, 3) {real, imag} */,
  {32'hc19e0e33, 32'hc0b3dfed} /* (30, 26, 2) {real, imag} */,
  {32'hc1a87fe7, 32'hc217ef32} /* (30, 26, 1) {real, imag} */,
  {32'h41bb76e3, 32'hc045bf5b} /* (30, 26, 0) {real, imag} */,
  {32'hc0bd6db2, 32'hc16ef9e3} /* (30, 25, 31) {real, imag} */,
  {32'h419e2ee1, 32'h4179c2d0} /* (30, 25, 30) {real, imag} */,
  {32'h40850b90, 32'h4112043d} /* (30, 25, 29) {real, imag} */,
  {32'h40501f4c, 32'hc03cfb98} /* (30, 25, 28) {real, imag} */,
  {32'h415786f6, 32'hc11063f8} /* (30, 25, 27) {real, imag} */,
  {32'h40843dea, 32'h40c64d82} /* (30, 25, 26) {real, imag} */,
  {32'h4031f4d7, 32'h4095bfd4} /* (30, 25, 25) {real, imag} */,
  {32'h4131bb08, 32'hc012e5c4} /* (30, 25, 24) {real, imag} */,
  {32'h400fd6ac, 32'h3fe7c2e8} /* (30, 25, 23) {real, imag} */,
  {32'h412d0b25, 32'hc115a868} /* (30, 25, 22) {real, imag} */,
  {32'h404641d6, 32'hc011d657} /* (30, 25, 21) {real, imag} */,
  {32'h404c8518, 32'h40575962} /* (30, 25, 20) {real, imag} */,
  {32'h411ceef9, 32'h3ff26084} /* (30, 25, 19) {real, imag} */,
  {32'hc11ff05d, 32'hbfc78734} /* (30, 25, 18) {real, imag} */,
  {32'hc07a5d28, 32'h40566ab7} /* (30, 25, 17) {real, imag} */,
  {32'h4131ac6d, 32'h3fd6d25a} /* (30, 25, 16) {real, imag} */,
  {32'hc11caaf4, 32'hbf228cfc} /* (30, 25, 15) {real, imag} */,
  {32'h4075cd34, 32'hbffa7830} /* (30, 25, 14) {real, imag} */,
  {32'h40bcceba, 32'h4103d585} /* (30, 25, 13) {real, imag} */,
  {32'hc171bda8, 32'hbfc918b8} /* (30, 25, 12) {real, imag} */,
  {32'h41623703, 32'hc03635cb} /* (30, 25, 11) {real, imag} */,
  {32'hc089818a, 32'h408bd4d5} /* (30, 25, 10) {real, imag} */,
  {32'h411dc2e9, 32'hc12bfa4d} /* (30, 25, 9) {real, imag} */,
  {32'hc05c959c, 32'hbf56a23c} /* (30, 25, 8) {real, imag} */,
  {32'hc18697da, 32'h3ff39020} /* (30, 25, 7) {real, imag} */,
  {32'h414798e6, 32'hc1a581d0} /* (30, 25, 6) {real, imag} */,
  {32'hc144aa52, 32'h41234d83} /* (30, 25, 5) {real, imag} */,
  {32'hc1c44bba, 32'h3e9fae30} /* (30, 25, 4) {real, imag} */,
  {32'h40ee91b0, 32'hc1255a68} /* (30, 25, 3) {real, imag} */,
  {32'hc18689a4, 32'h416a6674} /* (30, 25, 2) {real, imag} */,
  {32'h40d1cba9, 32'hc135a8d2} /* (30, 25, 1) {real, imag} */,
  {32'h41c6a4ad, 32'hc0b5171e} /* (30, 25, 0) {real, imag} */,
  {32'hc1b32438, 32'h41edf06f} /* (30, 24, 31) {real, imag} */,
  {32'h419b5584, 32'hc22504e6} /* (30, 24, 30) {real, imag} */,
  {32'hc13001c4, 32'hc1702912} /* (30, 24, 29) {real, imag} */,
  {32'hc19471d2, 32'hc1078619} /* (30, 24, 28) {real, imag} */,
  {32'h412c15fa, 32'hc0807bad} /* (30, 24, 27) {real, imag} */,
  {32'h40252170, 32'hc126649a} /* (30, 24, 26) {real, imag} */,
  {32'hc0f95c26, 32'hc15e36ea} /* (30, 24, 25) {real, imag} */,
  {32'hc104fe0f, 32'h3ffb56b6} /* (30, 24, 24) {real, imag} */,
  {32'hc1165bf5, 32'h414aefe6} /* (30, 24, 23) {real, imag} */,
  {32'h40426b7e, 32'hc18358a9} /* (30, 24, 22) {real, imag} */,
  {32'hbf20c910, 32'hc04e748c} /* (30, 24, 21) {real, imag} */,
  {32'hc163c9f2, 32'hc08388ee} /* (30, 24, 20) {real, imag} */,
  {32'hc0137ce0, 32'h410a1193} /* (30, 24, 19) {real, imag} */,
  {32'hc00e7770, 32'h4181f9c7} /* (30, 24, 18) {real, imag} */,
  {32'hc0fce68a, 32'h3ffbb210} /* (30, 24, 17) {real, imag} */,
  {32'hc1382322, 32'hc0970fcc} /* (30, 24, 16) {real, imag} */,
  {32'h418c39fe, 32'hc05d06e5} /* (30, 24, 15) {real, imag} */,
  {32'hbfee6366, 32'hc0edcf2f} /* (30, 24, 14) {real, imag} */,
  {32'h412380d8, 32'hbfaf3668} /* (30, 24, 13) {real, imag} */,
  {32'h406492b8, 32'h40abb85a} /* (30, 24, 12) {real, imag} */,
  {32'h403a114e, 32'h414b43ca} /* (30, 24, 11) {real, imag} */,
  {32'h407c39da, 32'h413a9878} /* (30, 24, 10) {real, imag} */,
  {32'hc0884798, 32'hc0348eb0} /* (30, 24, 9) {real, imag} */,
  {32'h408cefeb, 32'h402c7548} /* (30, 24, 8) {real, imag} */,
  {32'h400a2bb4, 32'h414e5c8b} /* (30, 24, 7) {real, imag} */,
  {32'h401f7754, 32'hc11d7536} /* (30, 24, 6) {real, imag} */,
  {32'hc09ae594, 32'hc0ff5602} /* (30, 24, 5) {real, imag} */,
  {32'hc0158e38, 32'hc15515d3} /* (30, 24, 4) {real, imag} */,
  {32'hc13f5af0, 32'h41987ff3} /* (30, 24, 3) {real, imag} */,
  {32'h4210b064, 32'hbeac1720} /* (30, 24, 2) {real, imag} */,
  {32'hc20c8f3f, 32'h41b22d7c} /* (30, 24, 1) {real, imag} */,
  {32'hc21f2882, 32'hbfed2c20} /* (30, 24, 0) {real, imag} */,
  {32'h41d45051, 32'hc09e398e} /* (30, 23, 31) {real, imag} */,
  {32'hc1f117be, 32'h41c2bc3e} /* (30, 23, 30) {real, imag} */,
  {32'hc1c37583, 32'h414abf67} /* (30, 23, 29) {real, imag} */,
  {32'h4074c8e1, 32'hc13d72f0} /* (30, 23, 28) {real, imag} */,
  {32'h40c5e35f, 32'hc181f461} /* (30, 23, 27) {real, imag} */,
  {32'hbfce00d2, 32'h40630438} /* (30, 23, 26) {real, imag} */,
  {32'h40de55f9, 32'h418ce627} /* (30, 23, 25) {real, imag} */,
  {32'hc00fb214, 32'hc083d40c} /* (30, 23, 24) {real, imag} */,
  {32'h412f055c, 32'hc0158a74} /* (30, 23, 23) {real, imag} */,
  {32'hc0aa0f40, 32'h411abc9b} /* (30, 23, 22) {real, imag} */,
  {32'hc0e77c3a, 32'hbf7765c0} /* (30, 23, 21) {real, imag} */,
  {32'h40f27e2a, 32'h4187b336} /* (30, 23, 20) {real, imag} */,
  {32'hc103398a, 32'h3f65778c} /* (30, 23, 19) {real, imag} */,
  {32'hc178098c, 32'hc1264943} /* (30, 23, 18) {real, imag} */,
  {32'hc083cfec, 32'hbfd10ef0} /* (30, 23, 17) {real, imag} */,
  {32'h40bc6a7a, 32'h3e84cc40} /* (30, 23, 16) {real, imag} */,
  {32'h4041f254, 32'hbf3a6898} /* (30, 23, 15) {real, imag} */,
  {32'h40b73258, 32'h418cbd82} /* (30, 23, 14) {real, imag} */,
  {32'hc1197830, 32'h4060e2ab} /* (30, 23, 13) {real, imag} */,
  {32'h4187d16d, 32'h411eea4b} /* (30, 23, 12) {real, imag} */,
  {32'h4104c942, 32'hc13ee5ad} /* (30, 23, 11) {real, imag} */,
  {32'h40a59cd6, 32'hc12737c6} /* (30, 23, 10) {real, imag} */,
  {32'hc0575508, 32'h40fba745} /* (30, 23, 9) {real, imag} */,
  {32'hc17965c9, 32'h41b694d7} /* (30, 23, 8) {real, imag} */,
  {32'h4078e610, 32'h41184bdd} /* (30, 23, 7) {real, imag} */,
  {32'h4131e7da, 32'hc114b30d} /* (30, 23, 6) {real, imag} */,
  {32'hc15e196a, 32'h415292ae} /* (30, 23, 5) {real, imag} */,
  {32'hbff5d16e, 32'hc0d2beca} /* (30, 23, 4) {real, imag} */,
  {32'hc18f4920, 32'hc1b1f972} /* (30, 23, 3) {real, imag} */,
  {32'h40c232de, 32'h40439528} /* (30, 23, 2) {real, imag} */,
  {32'hc18ed06e, 32'hc138c11c} /* (30, 23, 1) {real, imag} */,
  {32'h405a2068, 32'hc0fc53fe} /* (30, 23, 0) {real, imag} */,
  {32'hc115bedf, 32'hbfda6bac} /* (30, 22, 31) {real, imag} */,
  {32'hc16ef0b4, 32'h41927529} /* (30, 22, 30) {real, imag} */,
  {32'h409b1c70, 32'hc106a8e6} /* (30, 22, 29) {real, imag} */,
  {32'hc0c79b4a, 32'hbaa9a000} /* (30, 22, 28) {real, imag} */,
  {32'hc108b1d6, 32'h4100da76} /* (30, 22, 27) {real, imag} */,
  {32'hc07ea1aa, 32'h41a8ad98} /* (30, 22, 26) {real, imag} */,
  {32'h4139ce38, 32'hc15d0a30} /* (30, 22, 25) {real, imag} */,
  {32'h40cf3be3, 32'h41220cc7} /* (30, 22, 24) {real, imag} */,
  {32'h41074a44, 32'hbfd47fa0} /* (30, 22, 23) {real, imag} */,
  {32'hc0e6cd6b, 32'hc1484332} /* (30, 22, 22) {real, imag} */,
  {32'h408059c2, 32'hc0842ad2} /* (30, 22, 21) {real, imag} */,
  {32'hc19ec2e5, 32'hc0baa276} /* (30, 22, 20) {real, imag} */,
  {32'h41f1c158, 32'h41157f1e} /* (30, 22, 19) {real, imag} */,
  {32'hc002409c, 32'hc084bffa} /* (30, 22, 18) {real, imag} */,
  {32'hc087a3f2, 32'hc10cb621} /* (30, 22, 17) {real, imag} */,
  {32'hc0e0bd61, 32'hbf547bb8} /* (30, 22, 16) {real, imag} */,
  {32'h3fb31994, 32'hc07661a1} /* (30, 22, 15) {real, imag} */,
  {32'h40e1b281, 32'h414b7c42} /* (30, 22, 14) {real, imag} */,
  {32'h41b60d69, 32'hc09ea928} /* (30, 22, 13) {real, imag} */,
  {32'h40c0898e, 32'hc1a1188e} /* (30, 22, 12) {real, imag} */,
  {32'hc1bb61aa, 32'h3fb3b9c8} /* (30, 22, 11) {real, imag} */,
  {32'h407562e6, 32'h41bdb0e8} /* (30, 22, 10) {real, imag} */,
  {32'hc10af730, 32'h40647bf4} /* (30, 22, 9) {real, imag} */,
  {32'hc16f821e, 32'h408b15bb} /* (30, 22, 8) {real, imag} */,
  {32'hc01d5bce, 32'h41072227} /* (30, 22, 7) {real, imag} */,
  {32'h405e485a, 32'h4096c279} /* (30, 22, 6) {real, imag} */,
  {32'h40b7f15a, 32'hc0520ca5} /* (30, 22, 5) {real, imag} */,
  {32'h40cbc290, 32'h413c59b2} /* (30, 22, 4) {real, imag} */,
  {32'h40dfc0dd, 32'h3f71c478} /* (30, 22, 3) {real, imag} */,
  {32'h417e9c1b, 32'h410fdf20} /* (30, 22, 2) {real, imag} */,
  {32'hbf037ded, 32'hc1a44a5a} /* (30, 22, 1) {real, imag} */,
  {32'hc01c8662, 32'h414188d2} /* (30, 22, 0) {real, imag} */,
  {32'hc0a86b2d, 32'h412e839f} /* (30, 21, 31) {real, imag} */,
  {32'hc1306b0b, 32'hc17655dd} /* (30, 21, 30) {real, imag} */,
  {32'h4166c75a, 32'h4115b272} /* (30, 21, 29) {real, imag} */,
  {32'h408902ec, 32'h40ed00c0} /* (30, 21, 28) {real, imag} */,
  {32'h4095f5da, 32'hbf3e0370} /* (30, 21, 27) {real, imag} */,
  {32'hc0fb842a, 32'h40830f5e} /* (30, 21, 26) {real, imag} */,
  {32'h4114cd2e, 32'h40a2297d} /* (30, 21, 25) {real, imag} */,
  {32'hc02822ee, 32'h40ef4c10} /* (30, 21, 24) {real, imag} */,
  {32'hc1865044, 32'hc0d73561} /* (30, 21, 23) {real, imag} */,
  {32'h412996e6, 32'hc094882b} /* (30, 21, 22) {real, imag} */,
  {32'h40ee4c9c, 32'h412a0132} /* (30, 21, 21) {real, imag} */,
  {32'hbe7da970, 32'hc122ba80} /* (30, 21, 20) {real, imag} */,
  {32'h40974a51, 32'hc08229ca} /* (30, 21, 19) {real, imag} */,
  {32'hc10a1767, 32'hbeeda5a0} /* (30, 21, 18) {real, imag} */,
  {32'h412225ef, 32'h40f7a1cf} /* (30, 21, 17) {real, imag} */,
  {32'hc121d6bd, 32'hc05e3d58} /* (30, 21, 16) {real, imag} */,
  {32'h3fb2293a, 32'hc120ddea} /* (30, 21, 15) {real, imag} */,
  {32'h4132d10a, 32'h40b726ca} /* (30, 21, 14) {real, imag} */,
  {32'hc185f5ac, 32'hc0696e77} /* (30, 21, 13) {real, imag} */,
  {32'h415c7672, 32'hc112ad82} /* (30, 21, 12) {real, imag} */,
  {32'h412abc1b, 32'hc109efe8} /* (30, 21, 11) {real, imag} */,
  {32'hc19c0043, 32'h40bf8a0a} /* (30, 21, 10) {real, imag} */,
  {32'hbf8bba78, 32'h4158f721} /* (30, 21, 9) {real, imag} */,
  {32'hc0517870, 32'hc14f13ea} /* (30, 21, 8) {real, imag} */,
  {32'hbfd8f9c0, 32'h3f000590} /* (30, 21, 7) {real, imag} */,
  {32'hc14121f4, 32'hc1507525} /* (30, 21, 6) {real, imag} */,
  {32'hc076c9ca, 32'h405341f0} /* (30, 21, 5) {real, imag} */,
  {32'h4147f48e, 32'h406e1e7c} /* (30, 21, 4) {real, imag} */,
  {32'h4111fee8, 32'hc1007700} /* (30, 21, 3) {real, imag} */,
  {32'h416f55f6, 32'hc178a8f4} /* (30, 21, 2) {real, imag} */,
  {32'hc080c062, 32'h415a124a} /* (30, 21, 1) {real, imag} */,
  {32'hc065903f, 32'h41c4ca47} /* (30, 21, 0) {real, imag} */,
  {32'h40974fb8, 32'hc0fff5ea} /* (30, 20, 31) {real, imag} */,
  {32'hbf8edd60, 32'h3fab7942} /* (30, 20, 30) {real, imag} */,
  {32'h4126259e, 32'hc075d25e} /* (30, 20, 29) {real, imag} */,
  {32'h3e8a7468, 32'h40a2f9da} /* (30, 20, 28) {real, imag} */,
  {32'hc13419bb, 32'h40f45c2b} /* (30, 20, 27) {real, imag} */,
  {32'h4180dc04, 32'hbf281340} /* (30, 20, 26) {real, imag} */,
  {32'h3b609000, 32'hc0e1ea44} /* (30, 20, 25) {real, imag} */,
  {32'hc10e824e, 32'hc0e3533d} /* (30, 20, 24) {real, imag} */,
  {32'hc0a3d86e, 32'hbf35e280} /* (30, 20, 23) {real, imag} */,
  {32'hc1083ca8, 32'h3f17b748} /* (30, 20, 22) {real, imag} */,
  {32'hc111c2c6, 32'hc11d05c4} /* (30, 20, 21) {real, imag} */,
  {32'h4159882a, 32'hc0922226} /* (30, 20, 20) {real, imag} */,
  {32'hc10e083b, 32'hbf1470a0} /* (30, 20, 19) {real, imag} */,
  {32'hbfe756a8, 32'hc00a09d8} /* (30, 20, 18) {real, imag} */,
  {32'h4062f340, 32'hc065f8f4} /* (30, 20, 17) {real, imag} */,
  {32'h3f72f122, 32'hc10aa61c} /* (30, 20, 16) {real, imag} */,
  {32'h411949e6, 32'hc139ea26} /* (30, 20, 15) {real, imag} */,
  {32'hc116e3ec, 32'h414224ac} /* (30, 20, 14) {real, imag} */,
  {32'hc18527cb, 32'h4173b049} /* (30, 20, 13) {real, imag} */,
  {32'hc153098a, 32'h3f788d78} /* (30, 20, 12) {real, imag} */,
  {32'h416e7ce5, 32'hc039e252} /* (30, 20, 11) {real, imag} */,
  {32'h4172e13f, 32'hc09bed08} /* (30, 20, 10) {real, imag} */,
  {32'hbef258e8, 32'hc0da4104} /* (30, 20, 9) {real, imag} */,
  {32'h3fd39486, 32'h40ad0cbe} /* (30, 20, 8) {real, imag} */,
  {32'hc09df638, 32'hbea424e0} /* (30, 20, 7) {real, imag} */,
  {32'h3fe87a52, 32'h41a7dd56} /* (30, 20, 6) {real, imag} */,
  {32'hc0b879f2, 32'hc0f347be} /* (30, 20, 5) {real, imag} */,
  {32'hc09e51a3, 32'hc0f8a863} /* (30, 20, 4) {real, imag} */,
  {32'h4103396c, 32'h4155d77a} /* (30, 20, 3) {real, imag} */,
  {32'hc004b48c, 32'hc18d2cd6} /* (30, 20, 2) {real, imag} */,
  {32'hbe98e780, 32'h3fca38d0} /* (30, 20, 1) {real, imag} */,
  {32'hbff31310, 32'h41008ecd} /* (30, 20, 0) {real, imag} */,
  {32'h419f5b05, 32'hc041d768} /* (30, 19, 31) {real, imag} */,
  {32'hc13997fa, 32'h400ecb58} /* (30, 19, 30) {real, imag} */,
  {32'h41202240, 32'h3fcee400} /* (30, 19, 29) {real, imag} */,
  {32'hc035ec2c, 32'h418124ab} /* (30, 19, 28) {real, imag} */,
  {32'hc155d369, 32'hc14d0fc2} /* (30, 19, 27) {real, imag} */,
  {32'h416a3900, 32'hbfaf1604} /* (30, 19, 26) {real, imag} */,
  {32'h408516c0, 32'hc17c4d68} /* (30, 19, 25) {real, imag} */,
  {32'hc1330781, 32'hbefd7ff0} /* (30, 19, 24) {real, imag} */,
  {32'hc0a75752, 32'h3f924640} /* (30, 19, 23) {real, imag} */,
  {32'hc022d9c8, 32'h40ed85c4} /* (30, 19, 22) {real, imag} */,
  {32'hc11393e8, 32'hc1175cd8} /* (30, 19, 21) {real, imag} */,
  {32'hc18d1bd9, 32'hc0220d74} /* (30, 19, 20) {real, imag} */,
  {32'hbec1b110, 32'hc0aa2195} /* (30, 19, 19) {real, imag} */,
  {32'h41055c05, 32'h401b5b10} /* (30, 19, 18) {real, imag} */,
  {32'h4155e640, 32'h4190fc78} /* (30, 19, 17) {real, imag} */,
  {32'h40f074f6, 32'h3f1f3a9e} /* (30, 19, 16) {real, imag} */,
  {32'hc15af2d2, 32'h410300fe} /* (30, 19, 15) {real, imag} */,
  {32'hc19cba2f, 32'h3ec57a50} /* (30, 19, 14) {real, imag} */,
  {32'hc118983d, 32'h401c37c0} /* (30, 19, 13) {real, imag} */,
  {32'hc07d7d3d, 32'h40ba843c} /* (30, 19, 12) {real, imag} */,
  {32'h409cdb3c, 32'h40853084} /* (30, 19, 11) {real, imag} */,
  {32'h41180f00, 32'h3f45b310} /* (30, 19, 10) {real, imag} */,
  {32'hbf91fa60, 32'hc087d1c2} /* (30, 19, 9) {real, imag} */,
  {32'hbf245f10, 32'hc08f7e29} /* (30, 19, 8) {real, imag} */,
  {32'h3ebed5e0, 32'hc11aa37d} /* (30, 19, 7) {real, imag} */,
  {32'h400fd739, 32'h41bd360d} /* (30, 19, 6) {real, imag} */,
  {32'hc1256ae2, 32'h40af55e4} /* (30, 19, 5) {real, imag} */,
  {32'h40f81470, 32'h40946000} /* (30, 19, 4) {real, imag} */,
  {32'h40a09dc6, 32'h406f6e92} /* (30, 19, 3) {real, imag} */,
  {32'hc149915e, 32'hbf13b010} /* (30, 19, 2) {real, imag} */,
  {32'hc112dc48, 32'h4122d0d4} /* (30, 19, 1) {real, imag} */,
  {32'h406d2d6f, 32'hc0b4e4e6} /* (30, 19, 0) {real, imag} */,
  {32'hbea90890, 32'h4145f24a} /* (30, 18, 31) {real, imag} */,
  {32'hbff30368, 32'hc035d37e} /* (30, 18, 30) {real, imag} */,
  {32'hbf92ac84, 32'hc0c5b661} /* (30, 18, 29) {real, imag} */,
  {32'hc17d7086, 32'h4183fc4b} /* (30, 18, 28) {real, imag} */,
  {32'h4107fc74, 32'hc015fe68} /* (30, 18, 27) {real, imag} */,
  {32'h4188589a, 32'hc0d9d81e} /* (30, 18, 26) {real, imag} */,
  {32'h40955823, 32'h400630e8} /* (30, 18, 25) {real, imag} */,
  {32'h41743b75, 32'hc0de26dc} /* (30, 18, 24) {real, imag} */,
  {32'hc0b5e323, 32'h412e52a5} /* (30, 18, 23) {real, imag} */,
  {32'hc17ee23c, 32'h3fc0d8c5} /* (30, 18, 22) {real, imag} */,
  {32'hbf7dbfe0, 32'h4028926c} /* (30, 18, 21) {real, imag} */,
  {32'hc0c1b471, 32'h3fc64d88} /* (30, 18, 20) {real, imag} */,
  {32'hc1219672, 32'h408ee620} /* (30, 18, 19) {real, imag} */,
  {32'h4162530a, 32'h408bf508} /* (30, 18, 18) {real, imag} */,
  {32'h4038d8b5, 32'hc0b04b3c} /* (30, 18, 17) {real, imag} */,
  {32'h40ff8645, 32'h40fe86b8} /* (30, 18, 16) {real, imag} */,
  {32'h403cad34, 32'h40408fb1} /* (30, 18, 15) {real, imag} */,
  {32'hc16271c9, 32'hc186eee4} /* (30, 18, 14) {real, imag} */,
  {32'hbec54308, 32'hc1983775} /* (30, 18, 13) {real, imag} */,
  {32'hc0feadc7, 32'h40947ffa} /* (30, 18, 12) {real, imag} */,
  {32'hbfd960a5, 32'h405c0ab0} /* (30, 18, 11) {real, imag} */,
  {32'hc0ef2772, 32'hc02e0dee} /* (30, 18, 10) {real, imag} */,
  {32'hc0d6e280, 32'hc0138d8c} /* (30, 18, 9) {real, imag} */,
  {32'h418c7b1b, 32'hbe5addb0} /* (30, 18, 8) {real, imag} */,
  {32'h4114ddde, 32'hbf87ef20} /* (30, 18, 7) {real, imag} */,
  {32'h41891ebe, 32'h408c3e6d} /* (30, 18, 6) {real, imag} */,
  {32'h3dab6fc0, 32'hc0dddc99} /* (30, 18, 5) {real, imag} */,
  {32'hc0075a94, 32'h40229434} /* (30, 18, 4) {real, imag} */,
  {32'h3f4c1550, 32'hc01afcd6} /* (30, 18, 3) {real, imag} */,
  {32'h403dbca2, 32'hbfe26840} /* (30, 18, 2) {real, imag} */,
  {32'h3eb4dc6e, 32'h4195ee2a} /* (30, 18, 1) {real, imag} */,
  {32'h4143c66e, 32'h418cb16e} /* (30, 18, 0) {real, imag} */,
  {32'h3ef5d9e8, 32'hc0be077b} /* (30, 17, 31) {real, imag} */,
  {32'hbc2d1c00, 32'h415bc9cc} /* (30, 17, 30) {real, imag} */,
  {32'hc132531d, 32'h3fdc54fd} /* (30, 17, 29) {real, imag} */,
  {32'h41122e44, 32'hbfda470e} /* (30, 17, 28) {real, imag} */,
  {32'hc0bf6420, 32'hc0db4af5} /* (30, 17, 27) {real, imag} */,
  {32'h40405ef0, 32'hc099a0b0} /* (30, 17, 26) {real, imag} */,
  {32'hc10ccc96, 32'h40927e63} /* (30, 17, 25) {real, imag} */,
  {32'hc146ef75, 32'hc16db41a} /* (30, 17, 24) {real, imag} */,
  {32'h40108484, 32'hbfcf85f6} /* (30, 17, 23) {real, imag} */,
  {32'hc01d41be, 32'h410236cf} /* (30, 17, 22) {real, imag} */,
  {32'h41a40fa8, 32'hc0cc3151} /* (30, 17, 21) {real, imag} */,
  {32'h40e3ff33, 32'hc0466fc9} /* (30, 17, 20) {real, imag} */,
  {32'hbfc3c7b0, 32'h408ce660} /* (30, 17, 19) {real, imag} */,
  {32'hc108d9e7, 32'h4010f5da} /* (30, 17, 18) {real, imag} */,
  {32'h402a6ccf, 32'h4036414a} /* (30, 17, 17) {real, imag} */,
  {32'h40f30b59, 32'h40ca2682} /* (30, 17, 16) {real, imag} */,
  {32'hbfbc9c93, 32'hc0c8a377} /* (30, 17, 15) {real, imag} */,
  {32'h3f935bfa, 32'hc0779ed0} /* (30, 17, 14) {real, imag} */,
  {32'hc16b7a1c, 32'h40aca59c} /* (30, 17, 13) {real, imag} */,
  {32'h40e9525c, 32'h40c0ca8b} /* (30, 17, 12) {real, imag} */,
  {32'hc0671c92, 32'hc08017d3} /* (30, 17, 11) {real, imag} */,
  {32'h40792392, 32'hc119945e} /* (30, 17, 10) {real, imag} */,
  {32'hbf5cac5c, 32'h3eba2900} /* (30, 17, 9) {real, imag} */,
  {32'h41102d09, 32'h4071bdab} /* (30, 17, 8) {real, imag} */,
  {32'hc059c5ae, 32'hc122ab8c} /* (30, 17, 7) {real, imag} */,
  {32'h410b9547, 32'hbf8c4bfa} /* (30, 17, 6) {real, imag} */,
  {32'h4078cdac, 32'h3fa9b848} /* (30, 17, 5) {real, imag} */,
  {32'h3fa8eb47, 32'hc0bd9e08} /* (30, 17, 4) {real, imag} */,
  {32'h403b9036, 32'hc053a2a5} /* (30, 17, 3) {real, imag} */,
  {32'h401b0bc8, 32'h41b07e06} /* (30, 17, 2) {real, imag} */,
  {32'hbfd137f0, 32'hc09cd7f2} /* (30, 17, 1) {real, imag} */,
  {32'h3f09f38c, 32'h40d5801a} /* (30, 17, 0) {real, imag} */,
  {32'h40855a50, 32'hc05820f9} /* (30, 16, 31) {real, imag} */,
  {32'hc06d626a, 32'h40178731} /* (30, 16, 30) {real, imag} */,
  {32'hc018b504, 32'hc0f21dd4} /* (30, 16, 29) {real, imag} */,
  {32'hbf94f03c, 32'hc0f2a4c2} /* (30, 16, 28) {real, imag} */,
  {32'hc067764c, 32'hbee2a50c} /* (30, 16, 27) {real, imag} */,
  {32'h3fd310e4, 32'h412c6029} /* (30, 16, 26) {real, imag} */,
  {32'hc102bbac, 32'h3ea6c600} /* (30, 16, 25) {real, imag} */,
  {32'h40903a62, 32'h3f9cd470} /* (30, 16, 24) {real, imag} */,
  {32'hbf3ec850, 32'h40820317} /* (30, 16, 23) {real, imag} */,
  {32'h4154fde2, 32'hc108832a} /* (30, 16, 22) {real, imag} */,
  {32'h40f2aa30, 32'h409a1ede} /* (30, 16, 21) {real, imag} */,
  {32'h40a56bb6, 32'h410877d8} /* (30, 16, 20) {real, imag} */,
  {32'hc1136893, 32'h4188f6b7} /* (30, 16, 19) {real, imag} */,
  {32'hc02e362e, 32'h409d9e36} /* (30, 16, 18) {real, imag} */,
  {32'hc0c14c16, 32'hc0b02e4e} /* (30, 16, 17) {real, imag} */,
  {32'hbffce92c, 32'h00000000} /* (30, 16, 16) {real, imag} */,
  {32'hc0c14c16, 32'h40b02e4e} /* (30, 16, 15) {real, imag} */,
  {32'hc02e362e, 32'hc09d9e36} /* (30, 16, 14) {real, imag} */,
  {32'hc1136893, 32'hc188f6b7} /* (30, 16, 13) {real, imag} */,
  {32'h40a56bb6, 32'hc10877d8} /* (30, 16, 12) {real, imag} */,
  {32'h40f2aa30, 32'hc09a1ede} /* (30, 16, 11) {real, imag} */,
  {32'h4154fde2, 32'h4108832a} /* (30, 16, 10) {real, imag} */,
  {32'hbf3ec850, 32'hc0820317} /* (30, 16, 9) {real, imag} */,
  {32'h40903a62, 32'hbf9cd470} /* (30, 16, 8) {real, imag} */,
  {32'hc102bbac, 32'hbea6c600} /* (30, 16, 7) {real, imag} */,
  {32'h3fd310e4, 32'hc12c6029} /* (30, 16, 6) {real, imag} */,
  {32'hc067764c, 32'h3ee2a50c} /* (30, 16, 5) {real, imag} */,
  {32'hbf94f03c, 32'h40f2a4c2} /* (30, 16, 4) {real, imag} */,
  {32'hc018b504, 32'h40f21dd4} /* (30, 16, 3) {real, imag} */,
  {32'hc06d626a, 32'hc0178731} /* (30, 16, 2) {real, imag} */,
  {32'h40855a50, 32'h405820f9} /* (30, 16, 1) {real, imag} */,
  {32'hbe8f9638, 32'h00000000} /* (30, 16, 0) {real, imag} */,
  {32'hbfd137f0, 32'h409cd7f2} /* (30, 15, 31) {real, imag} */,
  {32'h401b0bc8, 32'hc1b07e06} /* (30, 15, 30) {real, imag} */,
  {32'h403b9036, 32'h4053a2a5} /* (30, 15, 29) {real, imag} */,
  {32'h3fa8eb47, 32'h40bd9e08} /* (30, 15, 28) {real, imag} */,
  {32'h4078cdac, 32'hbfa9b848} /* (30, 15, 27) {real, imag} */,
  {32'h410b9547, 32'h3f8c4bfa} /* (30, 15, 26) {real, imag} */,
  {32'hc059c5ae, 32'h4122ab8c} /* (30, 15, 25) {real, imag} */,
  {32'h41102d09, 32'hc071bdab} /* (30, 15, 24) {real, imag} */,
  {32'hbf5cac5c, 32'hbeba2900} /* (30, 15, 23) {real, imag} */,
  {32'h40792392, 32'h4119945e} /* (30, 15, 22) {real, imag} */,
  {32'hc0671c92, 32'h408017d3} /* (30, 15, 21) {real, imag} */,
  {32'h40e9525c, 32'hc0c0ca8b} /* (30, 15, 20) {real, imag} */,
  {32'hc16b7a1c, 32'hc0aca59c} /* (30, 15, 19) {real, imag} */,
  {32'h3f935bfa, 32'h40779ed0} /* (30, 15, 18) {real, imag} */,
  {32'hbfbc9c93, 32'h40c8a377} /* (30, 15, 17) {real, imag} */,
  {32'h40f30b59, 32'hc0ca2682} /* (30, 15, 16) {real, imag} */,
  {32'h402a6ccf, 32'hc036414a} /* (30, 15, 15) {real, imag} */,
  {32'hc108d9e7, 32'hc010f5da} /* (30, 15, 14) {real, imag} */,
  {32'hbfc3c7b0, 32'hc08ce660} /* (30, 15, 13) {real, imag} */,
  {32'h40e3ff33, 32'h40466fc9} /* (30, 15, 12) {real, imag} */,
  {32'h41a40fa8, 32'h40cc3151} /* (30, 15, 11) {real, imag} */,
  {32'hc01d41be, 32'hc10236cf} /* (30, 15, 10) {real, imag} */,
  {32'h40108484, 32'h3fcf85f6} /* (30, 15, 9) {real, imag} */,
  {32'hc146ef75, 32'h416db41a} /* (30, 15, 8) {real, imag} */,
  {32'hc10ccc96, 32'hc0927e63} /* (30, 15, 7) {real, imag} */,
  {32'h40405ef0, 32'h4099a0b0} /* (30, 15, 6) {real, imag} */,
  {32'hc0bf6420, 32'h40db4af5} /* (30, 15, 5) {real, imag} */,
  {32'h41122e44, 32'h3fda470e} /* (30, 15, 4) {real, imag} */,
  {32'hc132531d, 32'hbfdc54fd} /* (30, 15, 3) {real, imag} */,
  {32'hbc2d1c00, 32'hc15bc9cc} /* (30, 15, 2) {real, imag} */,
  {32'h3ef5d9e8, 32'h40be077b} /* (30, 15, 1) {real, imag} */,
  {32'h3f09f38c, 32'hc0d5801a} /* (30, 15, 0) {real, imag} */,
  {32'h3eb4dc6e, 32'hc195ee2a} /* (30, 14, 31) {real, imag} */,
  {32'h403dbca2, 32'h3fe26840} /* (30, 14, 30) {real, imag} */,
  {32'h3f4c1550, 32'h401afcd6} /* (30, 14, 29) {real, imag} */,
  {32'hc0075a94, 32'hc0229434} /* (30, 14, 28) {real, imag} */,
  {32'h3dab6fc0, 32'h40dddc99} /* (30, 14, 27) {real, imag} */,
  {32'h41891ebe, 32'hc08c3e6d} /* (30, 14, 26) {real, imag} */,
  {32'h4114ddde, 32'h3f87ef20} /* (30, 14, 25) {real, imag} */,
  {32'h418c7b1b, 32'h3e5addb0} /* (30, 14, 24) {real, imag} */,
  {32'hc0d6e280, 32'h40138d8c} /* (30, 14, 23) {real, imag} */,
  {32'hc0ef2772, 32'h402e0dee} /* (30, 14, 22) {real, imag} */,
  {32'hbfd960a5, 32'hc05c0ab0} /* (30, 14, 21) {real, imag} */,
  {32'hc0feadc7, 32'hc0947ffa} /* (30, 14, 20) {real, imag} */,
  {32'hbec54308, 32'h41983775} /* (30, 14, 19) {real, imag} */,
  {32'hc16271c9, 32'h4186eee4} /* (30, 14, 18) {real, imag} */,
  {32'h403cad34, 32'hc0408fb1} /* (30, 14, 17) {real, imag} */,
  {32'h40ff8645, 32'hc0fe86b8} /* (30, 14, 16) {real, imag} */,
  {32'h4038d8b5, 32'h40b04b3c} /* (30, 14, 15) {real, imag} */,
  {32'h4162530a, 32'hc08bf508} /* (30, 14, 14) {real, imag} */,
  {32'hc1219672, 32'hc08ee620} /* (30, 14, 13) {real, imag} */,
  {32'hc0c1b471, 32'hbfc64d88} /* (30, 14, 12) {real, imag} */,
  {32'hbf7dbfe0, 32'hc028926c} /* (30, 14, 11) {real, imag} */,
  {32'hc17ee23c, 32'hbfc0d8c5} /* (30, 14, 10) {real, imag} */,
  {32'hc0b5e323, 32'hc12e52a5} /* (30, 14, 9) {real, imag} */,
  {32'h41743b75, 32'h40de26dc} /* (30, 14, 8) {real, imag} */,
  {32'h40955823, 32'hc00630e8} /* (30, 14, 7) {real, imag} */,
  {32'h4188589a, 32'h40d9d81e} /* (30, 14, 6) {real, imag} */,
  {32'h4107fc74, 32'h4015fe68} /* (30, 14, 5) {real, imag} */,
  {32'hc17d7086, 32'hc183fc4b} /* (30, 14, 4) {real, imag} */,
  {32'hbf92ac84, 32'h40c5b661} /* (30, 14, 3) {real, imag} */,
  {32'hbff30368, 32'h4035d37e} /* (30, 14, 2) {real, imag} */,
  {32'hbea90890, 32'hc145f24a} /* (30, 14, 1) {real, imag} */,
  {32'h4143c66e, 32'hc18cb16e} /* (30, 14, 0) {real, imag} */,
  {32'hc112dc48, 32'hc122d0d4} /* (30, 13, 31) {real, imag} */,
  {32'hc149915e, 32'h3f13b010} /* (30, 13, 30) {real, imag} */,
  {32'h40a09dc6, 32'hc06f6e92} /* (30, 13, 29) {real, imag} */,
  {32'h40f81470, 32'hc0946000} /* (30, 13, 28) {real, imag} */,
  {32'hc1256ae2, 32'hc0af55e4} /* (30, 13, 27) {real, imag} */,
  {32'h400fd739, 32'hc1bd360d} /* (30, 13, 26) {real, imag} */,
  {32'h3ebed5e0, 32'h411aa37d} /* (30, 13, 25) {real, imag} */,
  {32'hbf245f10, 32'h408f7e29} /* (30, 13, 24) {real, imag} */,
  {32'hbf91fa60, 32'h4087d1c2} /* (30, 13, 23) {real, imag} */,
  {32'h41180f00, 32'hbf45b310} /* (30, 13, 22) {real, imag} */,
  {32'h409cdb3c, 32'hc0853084} /* (30, 13, 21) {real, imag} */,
  {32'hc07d7d3d, 32'hc0ba843c} /* (30, 13, 20) {real, imag} */,
  {32'hc118983d, 32'hc01c37c0} /* (30, 13, 19) {real, imag} */,
  {32'hc19cba2f, 32'hbec57a50} /* (30, 13, 18) {real, imag} */,
  {32'hc15af2d2, 32'hc10300fe} /* (30, 13, 17) {real, imag} */,
  {32'h40f074f6, 32'hbf1f3a9e} /* (30, 13, 16) {real, imag} */,
  {32'h4155e640, 32'hc190fc78} /* (30, 13, 15) {real, imag} */,
  {32'h41055c05, 32'hc01b5b10} /* (30, 13, 14) {real, imag} */,
  {32'hbec1b110, 32'h40aa2195} /* (30, 13, 13) {real, imag} */,
  {32'hc18d1bd9, 32'h40220d74} /* (30, 13, 12) {real, imag} */,
  {32'hc11393e8, 32'h41175cd8} /* (30, 13, 11) {real, imag} */,
  {32'hc022d9c8, 32'hc0ed85c4} /* (30, 13, 10) {real, imag} */,
  {32'hc0a75752, 32'hbf924640} /* (30, 13, 9) {real, imag} */,
  {32'hc1330781, 32'h3efd7ff0} /* (30, 13, 8) {real, imag} */,
  {32'h408516c0, 32'h417c4d68} /* (30, 13, 7) {real, imag} */,
  {32'h416a3900, 32'h3faf1604} /* (30, 13, 6) {real, imag} */,
  {32'hc155d369, 32'h414d0fc2} /* (30, 13, 5) {real, imag} */,
  {32'hc035ec2c, 32'hc18124ab} /* (30, 13, 4) {real, imag} */,
  {32'h41202240, 32'hbfcee400} /* (30, 13, 3) {real, imag} */,
  {32'hc13997fa, 32'hc00ecb58} /* (30, 13, 2) {real, imag} */,
  {32'h419f5b05, 32'h4041d768} /* (30, 13, 1) {real, imag} */,
  {32'h406d2d6f, 32'h40b4e4e6} /* (30, 13, 0) {real, imag} */,
  {32'hbe98e780, 32'hbfca38d0} /* (30, 12, 31) {real, imag} */,
  {32'hc004b48c, 32'h418d2cd6} /* (30, 12, 30) {real, imag} */,
  {32'h4103396c, 32'hc155d77a} /* (30, 12, 29) {real, imag} */,
  {32'hc09e51a3, 32'h40f8a863} /* (30, 12, 28) {real, imag} */,
  {32'hc0b879f2, 32'h40f347be} /* (30, 12, 27) {real, imag} */,
  {32'h3fe87a52, 32'hc1a7dd56} /* (30, 12, 26) {real, imag} */,
  {32'hc09df638, 32'h3ea424e0} /* (30, 12, 25) {real, imag} */,
  {32'h3fd39486, 32'hc0ad0cbe} /* (30, 12, 24) {real, imag} */,
  {32'hbef258e8, 32'h40da4104} /* (30, 12, 23) {real, imag} */,
  {32'h4172e13f, 32'h409bed08} /* (30, 12, 22) {real, imag} */,
  {32'h416e7ce5, 32'h4039e252} /* (30, 12, 21) {real, imag} */,
  {32'hc153098a, 32'hbf788d78} /* (30, 12, 20) {real, imag} */,
  {32'hc18527cb, 32'hc173b049} /* (30, 12, 19) {real, imag} */,
  {32'hc116e3ec, 32'hc14224ac} /* (30, 12, 18) {real, imag} */,
  {32'h411949e6, 32'h4139ea26} /* (30, 12, 17) {real, imag} */,
  {32'h3f72f122, 32'h410aa61c} /* (30, 12, 16) {real, imag} */,
  {32'h4062f340, 32'h4065f8f4} /* (30, 12, 15) {real, imag} */,
  {32'hbfe756a8, 32'h400a09d8} /* (30, 12, 14) {real, imag} */,
  {32'hc10e083b, 32'h3f1470a0} /* (30, 12, 13) {real, imag} */,
  {32'h4159882a, 32'h40922226} /* (30, 12, 12) {real, imag} */,
  {32'hc111c2c6, 32'h411d05c4} /* (30, 12, 11) {real, imag} */,
  {32'hc1083ca8, 32'hbf17b748} /* (30, 12, 10) {real, imag} */,
  {32'hc0a3d86e, 32'h3f35e280} /* (30, 12, 9) {real, imag} */,
  {32'hc10e824e, 32'h40e3533d} /* (30, 12, 8) {real, imag} */,
  {32'h3b609000, 32'h40e1ea44} /* (30, 12, 7) {real, imag} */,
  {32'h4180dc04, 32'h3f281340} /* (30, 12, 6) {real, imag} */,
  {32'hc13419bb, 32'hc0f45c2b} /* (30, 12, 5) {real, imag} */,
  {32'h3e8a7468, 32'hc0a2f9da} /* (30, 12, 4) {real, imag} */,
  {32'h4126259e, 32'h4075d25e} /* (30, 12, 3) {real, imag} */,
  {32'hbf8edd60, 32'hbfab7942} /* (30, 12, 2) {real, imag} */,
  {32'h40974fb8, 32'h40fff5ea} /* (30, 12, 1) {real, imag} */,
  {32'hbff31310, 32'hc1008ecd} /* (30, 12, 0) {real, imag} */,
  {32'hc080c062, 32'hc15a124a} /* (30, 11, 31) {real, imag} */,
  {32'h416f55f6, 32'h4178a8f4} /* (30, 11, 30) {real, imag} */,
  {32'h4111fee8, 32'h41007700} /* (30, 11, 29) {real, imag} */,
  {32'h4147f48e, 32'hc06e1e7c} /* (30, 11, 28) {real, imag} */,
  {32'hc076c9ca, 32'hc05341f0} /* (30, 11, 27) {real, imag} */,
  {32'hc14121f4, 32'h41507525} /* (30, 11, 26) {real, imag} */,
  {32'hbfd8f9c0, 32'hbf000590} /* (30, 11, 25) {real, imag} */,
  {32'hc0517870, 32'h414f13ea} /* (30, 11, 24) {real, imag} */,
  {32'hbf8bba78, 32'hc158f721} /* (30, 11, 23) {real, imag} */,
  {32'hc19c0043, 32'hc0bf8a0a} /* (30, 11, 22) {real, imag} */,
  {32'h412abc1b, 32'h4109efe8} /* (30, 11, 21) {real, imag} */,
  {32'h415c7672, 32'h4112ad82} /* (30, 11, 20) {real, imag} */,
  {32'hc185f5ac, 32'h40696e77} /* (30, 11, 19) {real, imag} */,
  {32'h4132d10a, 32'hc0b726ca} /* (30, 11, 18) {real, imag} */,
  {32'h3fb2293a, 32'h4120ddea} /* (30, 11, 17) {real, imag} */,
  {32'hc121d6bd, 32'h405e3d58} /* (30, 11, 16) {real, imag} */,
  {32'h412225ef, 32'hc0f7a1cf} /* (30, 11, 15) {real, imag} */,
  {32'hc10a1767, 32'h3eeda5a0} /* (30, 11, 14) {real, imag} */,
  {32'h40974a51, 32'h408229ca} /* (30, 11, 13) {real, imag} */,
  {32'hbe7da970, 32'h4122ba80} /* (30, 11, 12) {real, imag} */,
  {32'h40ee4c9c, 32'hc12a0132} /* (30, 11, 11) {real, imag} */,
  {32'h412996e6, 32'h4094882b} /* (30, 11, 10) {real, imag} */,
  {32'hc1865044, 32'h40d73561} /* (30, 11, 9) {real, imag} */,
  {32'hc02822ee, 32'hc0ef4c10} /* (30, 11, 8) {real, imag} */,
  {32'h4114cd2e, 32'hc0a2297d} /* (30, 11, 7) {real, imag} */,
  {32'hc0fb842a, 32'hc0830f5e} /* (30, 11, 6) {real, imag} */,
  {32'h4095f5da, 32'h3f3e0370} /* (30, 11, 5) {real, imag} */,
  {32'h408902ec, 32'hc0ed00c0} /* (30, 11, 4) {real, imag} */,
  {32'h4166c75a, 32'hc115b272} /* (30, 11, 3) {real, imag} */,
  {32'hc1306b0b, 32'h417655dd} /* (30, 11, 2) {real, imag} */,
  {32'hc0a86b2d, 32'hc12e839f} /* (30, 11, 1) {real, imag} */,
  {32'hc065903f, 32'hc1c4ca47} /* (30, 11, 0) {real, imag} */,
  {32'hbf037ded, 32'h41a44a5a} /* (30, 10, 31) {real, imag} */,
  {32'h417e9c1b, 32'hc10fdf20} /* (30, 10, 30) {real, imag} */,
  {32'h40dfc0dd, 32'hbf71c478} /* (30, 10, 29) {real, imag} */,
  {32'h40cbc290, 32'hc13c59b2} /* (30, 10, 28) {real, imag} */,
  {32'h40b7f15a, 32'h40520ca5} /* (30, 10, 27) {real, imag} */,
  {32'h405e485a, 32'hc096c279} /* (30, 10, 26) {real, imag} */,
  {32'hc01d5bce, 32'hc1072227} /* (30, 10, 25) {real, imag} */,
  {32'hc16f821e, 32'hc08b15bb} /* (30, 10, 24) {real, imag} */,
  {32'hc10af730, 32'hc0647bf4} /* (30, 10, 23) {real, imag} */,
  {32'h407562e6, 32'hc1bdb0e8} /* (30, 10, 22) {real, imag} */,
  {32'hc1bb61aa, 32'hbfb3b9c8} /* (30, 10, 21) {real, imag} */,
  {32'h40c0898e, 32'h41a1188e} /* (30, 10, 20) {real, imag} */,
  {32'h41b60d69, 32'h409ea928} /* (30, 10, 19) {real, imag} */,
  {32'h40e1b281, 32'hc14b7c42} /* (30, 10, 18) {real, imag} */,
  {32'h3fb31994, 32'h407661a1} /* (30, 10, 17) {real, imag} */,
  {32'hc0e0bd61, 32'h3f547bb8} /* (30, 10, 16) {real, imag} */,
  {32'hc087a3f2, 32'h410cb621} /* (30, 10, 15) {real, imag} */,
  {32'hc002409c, 32'h4084bffa} /* (30, 10, 14) {real, imag} */,
  {32'h41f1c158, 32'hc1157f1e} /* (30, 10, 13) {real, imag} */,
  {32'hc19ec2e5, 32'h40baa276} /* (30, 10, 12) {real, imag} */,
  {32'h408059c2, 32'h40842ad2} /* (30, 10, 11) {real, imag} */,
  {32'hc0e6cd6b, 32'h41484332} /* (30, 10, 10) {real, imag} */,
  {32'h41074a44, 32'h3fd47fa0} /* (30, 10, 9) {real, imag} */,
  {32'h40cf3be3, 32'hc1220cc7} /* (30, 10, 8) {real, imag} */,
  {32'h4139ce38, 32'h415d0a30} /* (30, 10, 7) {real, imag} */,
  {32'hc07ea1aa, 32'hc1a8ad98} /* (30, 10, 6) {real, imag} */,
  {32'hc108b1d6, 32'hc100da76} /* (30, 10, 5) {real, imag} */,
  {32'hc0c79b4a, 32'h3aa9a000} /* (30, 10, 4) {real, imag} */,
  {32'h409b1c70, 32'h4106a8e6} /* (30, 10, 3) {real, imag} */,
  {32'hc16ef0b4, 32'hc1927529} /* (30, 10, 2) {real, imag} */,
  {32'hc115bedf, 32'h3fda6bac} /* (30, 10, 1) {real, imag} */,
  {32'hc01c8662, 32'hc14188d2} /* (30, 10, 0) {real, imag} */,
  {32'hc18ed06e, 32'h4138c11c} /* (30, 9, 31) {real, imag} */,
  {32'h40c232de, 32'hc0439528} /* (30, 9, 30) {real, imag} */,
  {32'hc18f4920, 32'h41b1f972} /* (30, 9, 29) {real, imag} */,
  {32'hbff5d16e, 32'h40d2beca} /* (30, 9, 28) {real, imag} */,
  {32'hc15e196a, 32'hc15292ae} /* (30, 9, 27) {real, imag} */,
  {32'h4131e7da, 32'h4114b30d} /* (30, 9, 26) {real, imag} */,
  {32'h4078e610, 32'hc1184bdd} /* (30, 9, 25) {real, imag} */,
  {32'hc17965c9, 32'hc1b694d7} /* (30, 9, 24) {real, imag} */,
  {32'hc0575508, 32'hc0fba745} /* (30, 9, 23) {real, imag} */,
  {32'h40a59cd6, 32'h412737c6} /* (30, 9, 22) {real, imag} */,
  {32'h4104c942, 32'h413ee5ad} /* (30, 9, 21) {real, imag} */,
  {32'h4187d16d, 32'hc11eea4b} /* (30, 9, 20) {real, imag} */,
  {32'hc1197830, 32'hc060e2ab} /* (30, 9, 19) {real, imag} */,
  {32'h40b73258, 32'hc18cbd82} /* (30, 9, 18) {real, imag} */,
  {32'h4041f254, 32'h3f3a6898} /* (30, 9, 17) {real, imag} */,
  {32'h40bc6a7a, 32'hbe84cc40} /* (30, 9, 16) {real, imag} */,
  {32'hc083cfec, 32'h3fd10ef0} /* (30, 9, 15) {real, imag} */,
  {32'hc178098c, 32'h41264943} /* (30, 9, 14) {real, imag} */,
  {32'hc103398a, 32'hbf65778c} /* (30, 9, 13) {real, imag} */,
  {32'h40f27e2a, 32'hc187b336} /* (30, 9, 12) {real, imag} */,
  {32'hc0e77c3a, 32'h3f7765c0} /* (30, 9, 11) {real, imag} */,
  {32'hc0aa0f40, 32'hc11abc9b} /* (30, 9, 10) {real, imag} */,
  {32'h412f055c, 32'h40158a74} /* (30, 9, 9) {real, imag} */,
  {32'hc00fb214, 32'h4083d40c} /* (30, 9, 8) {real, imag} */,
  {32'h40de55f9, 32'hc18ce627} /* (30, 9, 7) {real, imag} */,
  {32'hbfce00d2, 32'hc0630438} /* (30, 9, 6) {real, imag} */,
  {32'h40c5e35f, 32'h4181f461} /* (30, 9, 5) {real, imag} */,
  {32'h4074c8e1, 32'h413d72f0} /* (30, 9, 4) {real, imag} */,
  {32'hc1c37583, 32'hc14abf67} /* (30, 9, 3) {real, imag} */,
  {32'hc1f117be, 32'hc1c2bc3e} /* (30, 9, 2) {real, imag} */,
  {32'h41d45051, 32'h409e398e} /* (30, 9, 1) {real, imag} */,
  {32'h405a2068, 32'h40fc53fe} /* (30, 9, 0) {real, imag} */,
  {32'hc20c8f3f, 32'hc1b22d7c} /* (30, 8, 31) {real, imag} */,
  {32'h4210b064, 32'h3eac1720} /* (30, 8, 30) {real, imag} */,
  {32'hc13f5af0, 32'hc1987ff3} /* (30, 8, 29) {real, imag} */,
  {32'hc0158e38, 32'h415515d3} /* (30, 8, 28) {real, imag} */,
  {32'hc09ae594, 32'h40ff5602} /* (30, 8, 27) {real, imag} */,
  {32'h401f7754, 32'h411d7536} /* (30, 8, 26) {real, imag} */,
  {32'h400a2bb4, 32'hc14e5c8b} /* (30, 8, 25) {real, imag} */,
  {32'h408cefeb, 32'hc02c7548} /* (30, 8, 24) {real, imag} */,
  {32'hc0884798, 32'h40348eb0} /* (30, 8, 23) {real, imag} */,
  {32'h407c39da, 32'hc13a9878} /* (30, 8, 22) {real, imag} */,
  {32'h403a114e, 32'hc14b43ca} /* (30, 8, 21) {real, imag} */,
  {32'h406492b8, 32'hc0abb85a} /* (30, 8, 20) {real, imag} */,
  {32'h412380d8, 32'h3faf3668} /* (30, 8, 19) {real, imag} */,
  {32'hbfee6366, 32'h40edcf2f} /* (30, 8, 18) {real, imag} */,
  {32'h418c39fe, 32'h405d06e5} /* (30, 8, 17) {real, imag} */,
  {32'hc1382322, 32'h40970fcc} /* (30, 8, 16) {real, imag} */,
  {32'hc0fce68a, 32'hbffbb210} /* (30, 8, 15) {real, imag} */,
  {32'hc00e7770, 32'hc181f9c7} /* (30, 8, 14) {real, imag} */,
  {32'hc0137ce0, 32'hc10a1193} /* (30, 8, 13) {real, imag} */,
  {32'hc163c9f2, 32'h408388ee} /* (30, 8, 12) {real, imag} */,
  {32'hbf20c910, 32'h404e748c} /* (30, 8, 11) {real, imag} */,
  {32'h40426b7e, 32'h418358a9} /* (30, 8, 10) {real, imag} */,
  {32'hc1165bf5, 32'hc14aefe6} /* (30, 8, 9) {real, imag} */,
  {32'hc104fe0f, 32'hbffb56b6} /* (30, 8, 8) {real, imag} */,
  {32'hc0f95c26, 32'h415e36ea} /* (30, 8, 7) {real, imag} */,
  {32'h40252170, 32'h4126649a} /* (30, 8, 6) {real, imag} */,
  {32'h412c15fa, 32'h40807bad} /* (30, 8, 5) {real, imag} */,
  {32'hc19471d2, 32'h41078619} /* (30, 8, 4) {real, imag} */,
  {32'hc13001c4, 32'h41702912} /* (30, 8, 3) {real, imag} */,
  {32'h419b5584, 32'h422504e6} /* (30, 8, 2) {real, imag} */,
  {32'hc1b32438, 32'hc1edf06f} /* (30, 8, 1) {real, imag} */,
  {32'hc21f2882, 32'h3fed2c20} /* (30, 8, 0) {real, imag} */,
  {32'h40d1cba9, 32'h4135a8d2} /* (30, 7, 31) {real, imag} */,
  {32'hc18689a4, 32'hc16a6674} /* (30, 7, 30) {real, imag} */,
  {32'h40ee91b0, 32'h41255a68} /* (30, 7, 29) {real, imag} */,
  {32'hc1c44bba, 32'hbe9fae30} /* (30, 7, 28) {real, imag} */,
  {32'hc144aa52, 32'hc1234d83} /* (30, 7, 27) {real, imag} */,
  {32'h414798e6, 32'h41a581d0} /* (30, 7, 26) {real, imag} */,
  {32'hc18697da, 32'hbff39020} /* (30, 7, 25) {real, imag} */,
  {32'hc05c959c, 32'h3f56a23c} /* (30, 7, 24) {real, imag} */,
  {32'h411dc2e9, 32'h412bfa4d} /* (30, 7, 23) {real, imag} */,
  {32'hc089818a, 32'hc08bd4d5} /* (30, 7, 22) {real, imag} */,
  {32'h41623703, 32'h403635cb} /* (30, 7, 21) {real, imag} */,
  {32'hc171bda8, 32'h3fc918b8} /* (30, 7, 20) {real, imag} */,
  {32'h40bcceba, 32'hc103d585} /* (30, 7, 19) {real, imag} */,
  {32'h4075cd34, 32'h3ffa7830} /* (30, 7, 18) {real, imag} */,
  {32'hc11caaf4, 32'h3f228cfc} /* (30, 7, 17) {real, imag} */,
  {32'h4131ac6d, 32'hbfd6d25a} /* (30, 7, 16) {real, imag} */,
  {32'hc07a5d28, 32'hc0566ab7} /* (30, 7, 15) {real, imag} */,
  {32'hc11ff05d, 32'h3fc78734} /* (30, 7, 14) {real, imag} */,
  {32'h411ceef9, 32'hbff26084} /* (30, 7, 13) {real, imag} */,
  {32'h404c8518, 32'hc0575962} /* (30, 7, 12) {real, imag} */,
  {32'h404641d6, 32'h4011d657} /* (30, 7, 11) {real, imag} */,
  {32'h412d0b25, 32'h4115a868} /* (30, 7, 10) {real, imag} */,
  {32'h400fd6ac, 32'hbfe7c2e8} /* (30, 7, 9) {real, imag} */,
  {32'h4131bb08, 32'h4012e5c4} /* (30, 7, 8) {real, imag} */,
  {32'h4031f4d7, 32'hc095bfd4} /* (30, 7, 7) {real, imag} */,
  {32'h40843dea, 32'hc0c64d82} /* (30, 7, 6) {real, imag} */,
  {32'h415786f6, 32'h411063f8} /* (30, 7, 5) {real, imag} */,
  {32'h40501f4c, 32'h403cfb98} /* (30, 7, 4) {real, imag} */,
  {32'h40850b90, 32'hc112043d} /* (30, 7, 3) {real, imag} */,
  {32'h419e2ee1, 32'hc179c2d0} /* (30, 7, 2) {real, imag} */,
  {32'hc0bd6db2, 32'h416ef9e3} /* (30, 7, 1) {real, imag} */,
  {32'h41c6a4ad, 32'h40b5171e} /* (30, 7, 0) {real, imag} */,
  {32'hc1a87fe7, 32'h4217ef32} /* (30, 6, 31) {real, imag} */,
  {32'hc19e0e33, 32'h40b3dfed} /* (30, 6, 30) {real, imag} */,
  {32'h405b73e8, 32'hc1a8213e} /* (30, 6, 29) {real, imag} */,
  {32'hbfd80430, 32'hbfe085c0} /* (30, 6, 28) {real, imag} */,
  {32'h3fb770f2, 32'h410c30b1} /* (30, 6, 27) {real, imag} */,
  {32'h4131d327, 32'h41ae08e8} /* (30, 6, 26) {real, imag} */,
  {32'h3f8cef84, 32'hbfa59848} /* (30, 6, 25) {real, imag} */,
  {32'h418ad94a, 32'hc169030b} /* (30, 6, 24) {real, imag} */,
  {32'hbf8a9284, 32'hc08fc940} /* (30, 6, 23) {real, imag} */,
  {32'h40641684, 32'hbfe6d9a0} /* (30, 6, 22) {real, imag} */,
  {32'hc1160f55, 32'h3ff131b8} /* (30, 6, 21) {real, imag} */,
  {32'hc182fe59, 32'h40c346d2} /* (30, 6, 20) {real, imag} */,
  {32'hc1a4ee8c, 32'hc16aadce} /* (30, 6, 19) {real, imag} */,
  {32'h41813200, 32'h412d4bfe} /* (30, 6, 18) {real, imag} */,
  {32'hc00535b6, 32'hc128c4b4} /* (30, 6, 17) {real, imag} */,
  {32'h41006c63, 32'hc0cb91b6} /* (30, 6, 16) {real, imag} */,
  {32'hc0cf65f8, 32'h40865fbc} /* (30, 6, 15) {real, imag} */,
  {32'h403d65c1, 32'h409ffa9c} /* (30, 6, 14) {real, imag} */,
  {32'h4089b9b2, 32'h40d2a89b} /* (30, 6, 13) {real, imag} */,
  {32'hc15475ce, 32'hc0b759a2} /* (30, 6, 12) {real, imag} */,
  {32'h40362000, 32'hc0de3954} /* (30, 6, 11) {real, imag} */,
  {32'h40723bd8, 32'hc188211b} /* (30, 6, 10) {real, imag} */,
  {32'hc16c06c4, 32'h4108b9da} /* (30, 6, 9) {real, imag} */,
  {32'h4090d4ec, 32'h4064432c} /* (30, 6, 8) {real, imag} */,
  {32'h4013c534, 32'h4123cba9} /* (30, 6, 7) {real, imag} */,
  {32'hc180f4e0, 32'h4166e546} /* (30, 6, 6) {real, imag} */,
  {32'h41b200d6, 32'h412e0121} /* (30, 6, 5) {real, imag} */,
  {32'h4158ef52, 32'h3f82cc2c} /* (30, 6, 4) {real, imag} */,
  {32'hc11d94b9, 32'h4104dd62} /* (30, 6, 3) {real, imag} */,
  {32'h403392c0, 32'hc14b219a} /* (30, 6, 2) {real, imag} */,
  {32'hc21b5ed5, 32'hc112e702} /* (30, 6, 1) {real, imag} */,
  {32'h41bb76e3, 32'h4045bf5b} /* (30, 6, 0) {real, imag} */,
  {32'hc29f0a5e, 32'hc150e478} /* (30, 5, 31) {real, imag} */,
  {32'h41b82820, 32'hc20b0019} /* (30, 5, 30) {real, imag} */,
  {32'h4092d792, 32'hc0928776} /* (30, 5, 29) {real, imag} */,
  {32'h4124fc64, 32'h41545c23} /* (30, 5, 28) {real, imag} */,
  {32'h41d5bf3b, 32'hc00f45c6} /* (30, 5, 27) {real, imag} */,
  {32'hc0f84284, 32'h401ea044} /* (30, 5, 26) {real, imag} */,
  {32'hc1b76f45, 32'h4130e778} /* (30, 5, 25) {real, imag} */,
  {32'hc0201f6e, 32'h418ab02e} /* (30, 5, 24) {real, imag} */,
  {32'hc1513b06, 32'hc108c0c7} /* (30, 5, 23) {real, imag} */,
  {32'h3fce1470, 32'hc1e86c70} /* (30, 5, 22) {real, imag} */,
  {32'h40b9d914, 32'hbf669868} /* (30, 5, 21) {real, imag} */,
  {32'hc09a1fad, 32'hc07e8696} /* (30, 5, 20) {real, imag} */,
  {32'h40924e91, 32'hc05b4768} /* (30, 5, 19) {real, imag} */,
  {32'hc107ba82, 32'hbf37e630} /* (30, 5, 18) {real, imag} */,
  {32'hc0820c95, 32'hbfdb1ac2} /* (30, 5, 17) {real, imag} */,
  {32'hc044c6d9, 32'h40597a15} /* (30, 5, 16) {real, imag} */,
  {32'hc09e57c3, 32'h3fc5a6f4} /* (30, 5, 15) {real, imag} */,
  {32'h3fc183de, 32'h40e235ca} /* (30, 5, 14) {real, imag} */,
  {32'h40fa1402, 32'h3ec4d0c0} /* (30, 5, 13) {real, imag} */,
  {32'hc03c5990, 32'h417987d1} /* (30, 5, 12) {real, imag} */,
  {32'hc1a9fc6d, 32'h402c69c4} /* (30, 5, 11) {real, imag} */,
  {32'hbfd81dea, 32'h40722fb6} /* (30, 5, 10) {real, imag} */,
  {32'h4084106e, 32'h41856184} /* (30, 5, 9) {real, imag} */,
  {32'hc11cf8d5, 32'h415de052} /* (30, 5, 8) {real, imag} */,
  {32'h415540df, 32'hc1760a79} /* (30, 5, 7) {real, imag} */,
  {32'h4188efa0, 32'hbfd322ec} /* (30, 5, 6) {real, imag} */,
  {32'hc16ecd65, 32'h418397dc} /* (30, 5, 5) {real, imag} */,
  {32'hc19401c5, 32'hc19075ac} /* (30, 5, 4) {real, imag} */,
  {32'hc087ca4c, 32'hbdf14fc0} /* (30, 5, 3) {real, imag} */,
  {32'h424840ea, 32'h42197758} /* (30, 5, 2) {real, imag} */,
  {32'hc2685825, 32'hc284576e} /* (30, 5, 1) {real, imag} */,
  {32'hc291a4a3, 32'h40eb5d26} /* (30, 5, 0) {real, imag} */,
  {32'h42608b95, 32'h42820672} /* (30, 4, 31) {real, imag} */,
  {32'hc2be70cc, 32'hc068fcf0} /* (30, 4, 30) {real, imag} */,
  {32'hc0f43d2a, 32'h41eaa4fc} /* (30, 4, 29) {real, imag} */,
  {32'h420456f6, 32'h41bfa27a} /* (30, 4, 28) {real, imag} */,
  {32'hc1f31231, 32'hc14c2f3e} /* (30, 4, 27) {real, imag} */,
  {32'hbdd56980, 32'h3eebd640} /* (30, 4, 26) {real, imag} */,
  {32'hc1670735, 32'hc0855dcf} /* (30, 4, 25) {real, imag} */,
  {32'hc0147ad1, 32'hc040b6f4} /* (30, 4, 24) {real, imag} */,
  {32'h41388d6a, 32'h40aed6cc} /* (30, 4, 23) {real, imag} */,
  {32'h417cc0b4, 32'hc00e9a2c} /* (30, 4, 22) {real, imag} */,
  {32'hc18f906e, 32'h4111c2d4} /* (30, 4, 21) {real, imag} */,
  {32'h4052ee7b, 32'hc12a1db6} /* (30, 4, 20) {real, imag} */,
  {32'h4073f710, 32'h405b3409} /* (30, 4, 19) {real, imag} */,
  {32'h403b39a8, 32'h4127093e} /* (30, 4, 18) {real, imag} */,
  {32'h40a4b966, 32'hc023b0fc} /* (30, 4, 17) {real, imag} */,
  {32'hc12f5a5c, 32'hbf50cb5e} /* (30, 4, 16) {real, imag} */,
  {32'h407835ca, 32'hbf77d3c0} /* (30, 4, 15) {real, imag} */,
  {32'hc06cddf0, 32'hc02f1f6c} /* (30, 4, 14) {real, imag} */,
  {32'h41043fae, 32'hc081e9d0} /* (30, 4, 13) {real, imag} */,
  {32'hbe7523d0, 32'hc132ec21} /* (30, 4, 12) {real, imag} */,
  {32'h41351043, 32'hc0f0734c} /* (30, 4, 11) {real, imag} */,
  {32'hc19261bf, 32'h41c50aba} /* (30, 4, 10) {real, imag} */,
  {32'h419798d1, 32'hbf754592} /* (30, 4, 9) {real, imag} */,
  {32'hbf91c210, 32'h40f111a4} /* (30, 4, 8) {real, imag} */,
  {32'h41a79a69, 32'h41e04ac4} /* (30, 4, 7) {real, imag} */,
  {32'hbeca2cf0, 32'hc10da080} /* (30, 4, 6) {real, imag} */,
  {32'h417df056, 32'hc1d8f569} /* (30, 4, 5) {real, imag} */,
  {32'hc00600f4, 32'h41ecb9e9} /* (30, 4, 4) {real, imag} */,
  {32'h40c3c42e, 32'h4186919d} /* (30, 4, 3) {real, imag} */,
  {32'hc2212f4a, 32'hc2918674} /* (30, 4, 2) {real, imag} */,
  {32'h4300b95a, 32'h428a6147} /* (30, 4, 1) {real, imag} */,
  {32'h4288bf4e, 32'h41a9079d} /* (30, 4, 0) {real, imag} */,
  {32'hc2b6eec5, 32'h429606d2} /* (30, 3, 31) {real, imag} */,
  {32'h426322f8, 32'hc29a2415} /* (30, 3, 30) {real, imag} */,
  {32'h4138d2b4, 32'h4138d840} /* (30, 3, 29) {real, imag} */,
  {32'h402db324, 32'h41acd2ee} /* (30, 3, 28) {real, imag} */,
  {32'h40b148a3, 32'hc19bf8b4} /* (30, 3, 27) {real, imag} */,
  {32'h402cf338, 32'hc09d30f0} /* (30, 3, 26) {real, imag} */,
  {32'hc11fd18d, 32'h41177b6e} /* (30, 3, 25) {real, imag} */,
  {32'hc11da3a4, 32'hbeede760} /* (30, 3, 24) {real, imag} */,
  {32'h3f5d1d40, 32'h4040569c} /* (30, 3, 23) {real, imag} */,
  {32'hbc7cf580, 32'h412c0f0b} /* (30, 3, 22) {real, imag} */,
  {32'hc14dbfc9, 32'h408d0915} /* (30, 3, 21) {real, imag} */,
  {32'hc17ad778, 32'h401371e4} /* (30, 3, 20) {real, imag} */,
  {32'hc0adddc2, 32'h40e6501a} /* (30, 3, 19) {real, imag} */,
  {32'h3ffa41db, 32'h3fb0baf8} /* (30, 3, 18) {real, imag} */,
  {32'h40b20d94, 32'hc09062ce} /* (30, 3, 17) {real, imag} */,
  {32'hbd51b640, 32'hc17fa722} /* (30, 3, 16) {real, imag} */,
  {32'h4025959d, 32'h406b5d44} /* (30, 3, 15) {real, imag} */,
  {32'hbf84a0f0, 32'hbfb25bc0} /* (30, 3, 14) {real, imag} */,
  {32'h414d5ac8, 32'h411b256e} /* (30, 3, 13) {real, imag} */,
  {32'hc0a2c39c, 32'hc0e08925} /* (30, 3, 12) {real, imag} */,
  {32'hc1164c3f, 32'h414198a1} /* (30, 3, 11) {real, imag} */,
  {32'hc191b68a, 32'hc17e70c3} /* (30, 3, 10) {real, imag} */,
  {32'h4095c2aa, 32'h40c7d443} /* (30, 3, 9) {real, imag} */,
  {32'hc0625cf7, 32'hc0abeb4c} /* (30, 3, 8) {real, imag} */,
  {32'h41bd5a26, 32'h4105a390} /* (30, 3, 7) {real, imag} */,
  {32'hbf7a5d40, 32'h4098577e} /* (30, 3, 6) {real, imag} */,
  {32'hc1ddf5c5, 32'h418f1870} /* (30, 3, 5) {real, imag} */,
  {32'hc0e8d1cc, 32'h4195f5e1} /* (30, 3, 4) {real, imag} */,
  {32'h41d4574d, 32'h40410af0} /* (30, 3, 3) {real, imag} */,
  {32'hc0d39334, 32'hc28bb6a3} /* (30, 3, 2) {real, imag} */,
  {32'h42621b78, 32'h425d548c} /* (30, 3, 1) {real, imag} */,
  {32'hc13fa95e, 32'h4197dbf8} /* (30, 3, 0) {real, imag} */,
  {32'hc41425c8, 32'hc28b522d} /* (30, 2, 31) {real, imag} */,
  {32'h439c9632, 32'hc2f2ba10} /* (30, 2, 30) {real, imag} */,
  {32'h42171962, 32'h403e4ad4} /* (30, 2, 29) {real, imag} */,
  {32'hc24c6cd7, 32'h42b5afd4} /* (30, 2, 28) {real, imag} */,
  {32'h4236c4f6, 32'hc11f778e} /* (30, 2, 27) {real, imag} */,
  {32'h418ee529, 32'h410e4f4a} /* (30, 2, 26) {real, imag} */,
  {32'hc135bba6, 32'hc0e836ca} /* (30, 2, 25) {real, imag} */,
  {32'h422e19b9, 32'hc1264456} /* (30, 2, 24) {real, imag} */,
  {32'h3f4a5ee0, 32'h40cd3253} /* (30, 2, 23) {real, imag} */,
  {32'hc125b02e, 32'h408b10c2} /* (30, 2, 22) {real, imag} */,
  {32'hc0a974d3, 32'hc173507e} /* (30, 2, 21) {real, imag} */,
  {32'hc04d99d1, 32'h41707dc8} /* (30, 2, 20) {real, imag} */,
  {32'hc01dc810, 32'hc0afe492} /* (30, 2, 19) {real, imag} */,
  {32'hc091d9f6, 32'hc17a90a0} /* (30, 2, 18) {real, imag} */,
  {32'h411e51fd, 32'hc0ece93b} /* (30, 2, 17) {real, imag} */,
  {32'h402f37a3, 32'h4078583c} /* (30, 2, 16) {real, imag} */,
  {32'hc10ddf8d, 32'h40248edc} /* (30, 2, 15) {real, imag} */,
  {32'hbeff0570, 32'hbf91b640} /* (30, 2, 14) {real, imag} */,
  {32'hc1296c5a, 32'hbf36d1be} /* (30, 2, 13) {real, imag} */,
  {32'h3f15ef50, 32'hc1491cc6} /* (30, 2, 12) {real, imag} */,
  {32'h41d159aa, 32'h420343f8} /* (30, 2, 11) {real, imag} */,
  {32'h3d01ad00, 32'hc1288ab8} /* (30, 2, 10) {real, imag} */,
  {32'h4190a162, 32'h4000af9b} /* (30, 2, 9) {real, imag} */,
  {32'h4114623a, 32'h404c80cc} /* (30, 2, 8) {real, imag} */,
  {32'h40e13ed8, 32'hc1aea44b} /* (30, 2, 7) {real, imag} */,
  {32'h4033ab24, 32'h414a03fe} /* (30, 2, 6) {real, imag} */,
  {32'h424c8b2c, 32'h4144d83c} /* (30, 2, 5) {real, imag} */,
  {32'hc24a1882, 32'h4101c8f0} /* (30, 2, 4) {real, imag} */,
  {32'hc213b24c, 32'hc21ef420} /* (30, 2, 3) {real, imag} */,
  {32'h43604551, 32'hc1a7d804} /* (30, 2, 2) {real, imag} */,
  {32'hc3cc7bde, 32'h4314ae16} /* (30, 2, 1) {real, imag} */,
  {32'hc3a6596a, 32'hc2016126} /* (30, 2, 0) {real, imag} */,
  {32'h440cc7f4, 32'hc31c48f1} /* (30, 1, 31) {real, imag} */,
  {32'hc368e09c, 32'h41c6c33f} /* (30, 1, 30) {real, imag} */,
  {32'hc1b856be, 32'h400f5720} /* (30, 1, 29) {real, imag} */,
  {32'h4258ebff, 32'h415a0434} /* (30, 1, 28) {real, imag} */,
  {32'hc29085d0, 32'hc05918e3} /* (30, 1, 27) {real, imag} */,
  {32'hc1896380, 32'hc1993bbc} /* (30, 1, 26) {real, imag} */,
  {32'h41816a50, 32'hc2075831} /* (30, 1, 25) {real, imag} */,
  {32'hc1244c3c, 32'h420901d8} /* (30, 1, 24) {real, imag} */,
  {32'hc16073d7, 32'hbfe6efc4} /* (30, 1, 23) {real, imag} */,
  {32'h41265ee8, 32'hc1541d05} /* (30, 1, 22) {real, imag} */,
  {32'hc0f7277c, 32'h4215520f} /* (30, 1, 21) {real, imag} */,
  {32'h412f6794, 32'h3f1b6f90} /* (30, 1, 20) {real, imag} */,
  {32'h40a4a62a, 32'h40207b78} /* (30, 1, 19) {real, imag} */,
  {32'hc1454006, 32'h418c791b} /* (30, 1, 18) {real, imag} */,
  {32'h4063144b, 32'hc0a5d5b4} /* (30, 1, 17) {real, imag} */,
  {32'h3fea57ea, 32'h3e916758} /* (30, 1, 16) {real, imag} */,
  {32'hc1589c5c, 32'hbf88bd24} /* (30, 1, 15) {real, imag} */,
  {32'hc079a088, 32'hc0e6a9ed} /* (30, 1, 14) {real, imag} */,
  {32'h408fc74a, 32'h4195c9ad} /* (30, 1, 13) {real, imag} */,
  {32'h4179c11e, 32'hc09b6199} /* (30, 1, 12) {real, imag} */,
  {32'hbf325a50, 32'hc129db26} /* (30, 1, 11) {real, imag} */,
  {32'hc13f4064, 32'h407e9342} /* (30, 1, 10) {real, imag} */,
  {32'h4198db4c, 32'h4139a8f2} /* (30, 1, 9) {real, imag} */,
  {32'h3f863858, 32'hc2527a4a} /* (30, 1, 8) {real, imag} */,
  {32'hc17184f2, 32'h4193b1cb} /* (30, 1, 7) {real, imag} */,
  {32'hc1b2c782, 32'h41b59bb4} /* (30, 1, 6) {real, imag} */,
  {32'hc2b8d91a, 32'hc213a988} /* (30, 1, 5) {real, imag} */,
  {32'h4219e16e, 32'h40417f90} /* (30, 1, 4) {real, imag} */,
  {32'hc1d471d1, 32'h42625256} /* (30, 1, 3) {real, imag} */,
  {32'hc39e4521, 32'hc3b0ccd0} /* (30, 1, 2) {real, imag} */,
  {32'h44421f17, 32'h43a27cc4} /* (30, 1, 1) {real, imag} */,
  {32'h43ea7508, 32'h42dc2030} /* (30, 1, 0) {real, imag} */,
  {32'h4396b5b5, 32'hc387eb1d} /* (30, 0, 31) {real, imag} */,
  {32'hc2a3310d, 32'h4359e4c2} /* (30, 0, 30) {real, imag} */,
  {32'hc18f67ac, 32'h40b3bea8} /* (30, 0, 29) {real, imag} */,
  {32'hc0a79b62, 32'h42183828} /* (30, 0, 28) {real, imag} */,
  {32'hc204d0e0, 32'hc108d736} /* (30, 0, 27) {real, imag} */,
  {32'hc155bc83, 32'hc0f3985c} /* (30, 0, 26) {real, imag} */,
  {32'hc1bf91c0, 32'hc1a5d6ba} /* (30, 0, 25) {real, imag} */,
  {32'hc1a00882, 32'h41d7d573} /* (30, 0, 24) {real, imag} */,
  {32'hc0393eb2, 32'h41a244c4} /* (30, 0, 23) {real, imag} */,
  {32'h40971eed, 32'hc08b66a1} /* (30, 0, 22) {real, imag} */,
  {32'hbfbb1660, 32'hc01b0dd0} /* (30, 0, 21) {real, imag} */,
  {32'hbfb55350, 32'hc12081c7} /* (30, 0, 20) {real, imag} */,
  {32'h3fb7e9bc, 32'hc037545b} /* (30, 0, 19) {real, imag} */,
  {32'h40cf8ec4, 32'h4097dd0a} /* (30, 0, 18) {real, imag} */,
  {32'h416a8982, 32'h3fb28282} /* (30, 0, 17) {real, imag} */,
  {32'hc1272180, 32'h00000000} /* (30, 0, 16) {real, imag} */,
  {32'h416a8982, 32'hbfb28282} /* (30, 0, 15) {real, imag} */,
  {32'h40cf8ec4, 32'hc097dd0a} /* (30, 0, 14) {real, imag} */,
  {32'h3fb7e9bc, 32'h4037545b} /* (30, 0, 13) {real, imag} */,
  {32'hbfb55350, 32'h412081c7} /* (30, 0, 12) {real, imag} */,
  {32'hbfbb1660, 32'h401b0dd0} /* (30, 0, 11) {real, imag} */,
  {32'h40971eed, 32'h408b66a1} /* (30, 0, 10) {real, imag} */,
  {32'hc0393eb2, 32'hc1a244c4} /* (30, 0, 9) {real, imag} */,
  {32'hc1a00882, 32'hc1d7d573} /* (30, 0, 8) {real, imag} */,
  {32'hc1bf91c0, 32'h41a5d6ba} /* (30, 0, 7) {real, imag} */,
  {32'hc155bc83, 32'h40f3985c} /* (30, 0, 6) {real, imag} */,
  {32'hc204d0e0, 32'h4108d736} /* (30, 0, 5) {real, imag} */,
  {32'hc0a79b62, 32'hc2183828} /* (30, 0, 4) {real, imag} */,
  {32'hc18f67ac, 32'hc0b3bea8} /* (30, 0, 3) {real, imag} */,
  {32'hc2a3310d, 32'hc359e4c2} /* (30, 0, 2) {real, imag} */,
  {32'h4396b5b5, 32'h4387eb1d} /* (30, 0, 1) {real, imag} */,
  {32'h42a338ba, 32'h00000000} /* (30, 0, 0) {real, imag} */,
  {32'h446981a4, 32'hc3c56bdc} /* (29, 31, 31) {real, imag} */,
  {32'hc3c0cccc, 32'h43e3363a} /* (29, 31, 30) {real, imag} */,
  {32'hc1c6232c, 32'hc2449552} /* (29, 31, 29) {real, imag} */,
  {32'h423cf852, 32'hc20e7a8a} /* (29, 31, 28) {real, imag} */,
  {32'hc28d7d19, 32'h42062d79} /* (29, 31, 27) {real, imag} */,
  {32'hc123bcfc, 32'hc155cc87} /* (29, 31, 26) {real, imag} */,
  {32'hc1303fd2, 32'hc100b5bc} /* (29, 31, 25) {real, imag} */,
  {32'hc0d3e927, 32'h41e2fc62} /* (29, 31, 24) {real, imag} */,
  {32'hc12c2cae, 32'hc0d8be7f} /* (29, 31, 23) {real, imag} */,
  {32'hc1d014ec, 32'hbf6fafe0} /* (29, 31, 22) {real, imag} */,
  {32'h40a2a97c, 32'h4177e64d} /* (29, 31, 21) {real, imag} */,
  {32'h40a18aee, 32'hc09d66f0} /* (29, 31, 20) {real, imag} */,
  {32'h40637cec, 32'h40f46b4a} /* (29, 31, 19) {real, imag} */,
  {32'h410d20a3, 32'h413c3204} /* (29, 31, 18) {real, imag} */,
  {32'h4068306e, 32'hc0309a0e} /* (29, 31, 17) {real, imag} */,
  {32'hc0ea626f, 32'h4110d995} /* (29, 31, 16) {real, imag} */,
  {32'h3fa3cfd8, 32'hbf8d225c} /* (29, 31, 15) {real, imag} */,
  {32'hc18de0e5, 32'hc0b41b40} /* (29, 31, 14) {real, imag} */,
  {32'h413f87fc, 32'hc039c239} /* (29, 31, 13) {real, imag} */,
  {32'hc0b5c04e, 32'hc0b27d7b} /* (29, 31, 12) {real, imag} */,
  {32'hc09a43f6, 32'hc1b2db66} /* (29, 31, 11) {real, imag} */,
  {32'h4135fd69, 32'h40eb686f} /* (29, 31, 10) {real, imag} */,
  {32'h409f221c, 32'h403c9a68} /* (29, 31, 9) {real, imag} */,
  {32'h4060bee0, 32'hc1c062bd} /* (29, 31, 8) {real, imag} */,
  {32'h3f6d8b00, 32'h423a28f8} /* (29, 31, 7) {real, imag} */,
  {32'hc1966796, 32'hc07de660} /* (29, 31, 6) {real, imag} */,
  {32'hc2e9e5bc, 32'hc234c304} /* (29, 31, 5) {real, imag} */,
  {32'h4245a46a, 32'hc2800d1f} /* (29, 31, 4) {real, imag} */,
  {32'hc0b4d694, 32'h4186f9a0} /* (29, 31, 3) {real, imag} */,
  {32'hc38976e2, 32'hc0729c18} /* (29, 31, 2) {real, imag} */,
  {32'h4420b567, 32'h434716e8} /* (29, 31, 1) {real, imag} */,
  {32'h440e6846, 32'hc2b994f4} /* (29, 31, 0) {real, imag} */,
  {32'hc3e4ca54, 32'hc303ee06} /* (29, 30, 31) {real, imag} */,
  {32'h4388fdd2, 32'h429f5e9c} /* (29, 30, 30) {real, imag} */,
  {32'hc1bd1c38, 32'h41a3899d} /* (29, 30, 29) {real, imag} */,
  {32'hc263036c, 32'h4175a0d6} /* (29, 30, 28) {real, imag} */,
  {32'h421b7092, 32'hc13f1c97} /* (29, 30, 27) {real, imag} */,
  {32'h3f8e2640, 32'hc1725786} /* (29, 30, 26) {real, imag} */,
  {32'h4154c7f0, 32'h411d8360} /* (29, 30, 25) {real, imag} */,
  {32'hc0ad2634, 32'hc10bf4a1} /* (29, 30, 24) {real, imag} */,
  {32'h41698acd, 32'hc0a2cc1f} /* (29, 30, 23) {real, imag} */,
  {32'hc1801f2f, 32'hc18c7bd0} /* (29, 30, 22) {real, imag} */,
  {32'h41528e85, 32'hc126298e} /* (29, 30, 21) {real, imag} */,
  {32'h3fe7d760, 32'hc12baf6c} /* (29, 30, 20) {real, imag} */,
  {32'h4097fee6, 32'h417c5bf3} /* (29, 30, 19) {real, imag} */,
  {32'h4071c924, 32'hc0d8a92f} /* (29, 30, 18) {real, imag} */,
  {32'hc09ed663, 32'h40e248c8} /* (29, 30, 17) {real, imag} */,
  {32'h40d61933, 32'h40d684e9} /* (29, 30, 16) {real, imag} */,
  {32'hbf9e136e, 32'hc0d03fb5} /* (29, 30, 15) {real, imag} */,
  {32'h4107b257, 32'h3e742080} /* (29, 30, 14) {real, imag} */,
  {32'hc03966c4, 32'h41368f86} /* (29, 30, 13) {real, imag} */,
  {32'hc18e3ab9, 32'hc161cc11} /* (29, 30, 12) {real, imag} */,
  {32'h413accce, 32'h4132d43e} /* (29, 30, 11) {real, imag} */,
  {32'h4122f6ad, 32'hc19941f3} /* (29, 30, 10) {real, imag} */,
  {32'hc0edcd34, 32'h403a5248} /* (29, 30, 9) {real, imag} */,
  {32'h4219f172, 32'h41ab32ee} /* (29, 30, 8) {real, imag} */,
  {32'hc027b968, 32'hc1f3f13f} /* (29, 30, 7) {real, imag} */,
  {32'h410ebeba, 32'hc11c4232} /* (29, 30, 6) {real, imag} */,
  {32'h424bd6e6, 32'h41cd27c1} /* (29, 30, 5) {real, imag} */,
  {32'hc20df8e2, 32'hc29fef6e} /* (29, 30, 4) {real, imag} */,
  {32'h40fbede4, 32'h41550b5a} /* (29, 30, 3) {real, imag} */,
  {32'h43ccf7ac, 32'h43103bce} /* (29, 30, 2) {real, imag} */,
  {32'hc435e489, 32'h41c80b8a} /* (29, 30, 1) {real, imag} */,
  {32'hc3be597d, 32'h426894af} /* (29, 30, 0) {real, imag} */,
  {32'h428333fa, 32'hc2f13afc} /* (29, 29, 31) {real, imag} */,
  {32'hc045ee4c, 32'h429b7f9e} /* (29, 29, 30) {real, imag} */,
  {32'h41803b05, 32'hc16188aa} /* (29, 29, 29) {real, imag} */,
  {32'hc142324c, 32'hc1fb9454} /* (29, 29, 28) {real, imag} */,
  {32'hbed47b00, 32'hc082952c} /* (29, 29, 27) {real, imag} */,
  {32'hc1c935f0, 32'h41a53013} /* (29, 29, 26) {real, imag} */,
  {32'h41da5811, 32'hc09c433c} /* (29, 29, 25) {real, imag} */,
  {32'hc08a70d2, 32'h3f0cb730} /* (29, 29, 24) {real, imag} */,
  {32'h40dc5bac, 32'h3f83dc8a} /* (29, 29, 23) {real, imag} */,
  {32'h406a5ab8, 32'h40c01e90} /* (29, 29, 22) {real, imag} */,
  {32'hbfd2d808, 32'h3f689cf0} /* (29, 29, 21) {real, imag} */,
  {32'h4136dc91, 32'hc1813486} /* (29, 29, 20) {real, imag} */,
  {32'h40d5aaa8, 32'h40287e92} /* (29, 29, 19) {real, imag} */,
  {32'h3fea1162, 32'hc0b16024} /* (29, 29, 18) {real, imag} */,
  {32'h40bcc4aa, 32'h410420a1} /* (29, 29, 17) {real, imag} */,
  {32'hc039534a, 32'h4058d5d9} /* (29, 29, 16) {real, imag} */,
  {32'h40007b5c, 32'hc0477155} /* (29, 29, 15) {real, imag} */,
  {32'hc094c728, 32'h3d994f20} /* (29, 29, 14) {real, imag} */,
  {32'hc1335c07, 32'hc1061542} /* (29, 29, 13) {real, imag} */,
  {32'h40acb71a, 32'hc1336d6a} /* (29, 29, 12) {real, imag} */,
  {32'hc1ef964a, 32'hbfb34a00} /* (29, 29, 11) {real, imag} */,
  {32'h40b7213a, 32'h3f4ccad8} /* (29, 29, 10) {real, imag} */,
  {32'h4112f84d, 32'hbfd7fa70} /* (29, 29, 9) {real, imag} */,
  {32'hc14bbb9a, 32'h41b5f5b2} /* (29, 29, 8) {real, imag} */,
  {32'hc1043f86, 32'hc11607ae} /* (29, 29, 7) {real, imag} */,
  {32'hc0b11c4a, 32'hc1043564} /* (29, 29, 6) {real, imag} */,
  {32'hc0bb6a7c, 32'h421dc348} /* (29, 29, 5) {real, imag} */,
  {32'h417d76fd, 32'hc1e46c6a} /* (29, 29, 4) {real, imag} */,
  {32'h401a5a4c, 32'hc17a681b} /* (29, 29, 3) {real, imag} */,
  {32'h4285dcc3, 32'h429d31b6} /* (29, 29, 2) {real, imag} */,
  {32'hc2f54d4c, 32'hc29403bf} /* (29, 29, 1) {real, imag} */,
  {32'h41039992, 32'h3f912a38} /* (29, 29, 0) {real, imag} */,
  {32'h43204205, 32'hc28c80a3} /* (29, 28, 31) {real, imag} */,
  {32'hc212ba78, 32'h427ea0c2} /* (29, 28, 30) {real, imag} */,
  {32'h40f6001b, 32'h40b49028} /* (29, 28, 29) {real, imag} */,
  {32'h41cd952e, 32'hc14ac78e} /* (29, 28, 28) {real, imag} */,
  {32'h3fa7d09a, 32'h41d82390} /* (29, 28, 27) {real, imag} */,
  {32'hc04db624, 32'hc147aaed} /* (29, 28, 26) {real, imag} */,
  {32'h410d7a3c, 32'h41388083} /* (29, 28, 25) {real, imag} */,
  {32'hc11b468f, 32'h413e9f39} /* (29, 28, 24) {real, imag} */,
  {32'h40c0acc6, 32'h417ff297} /* (29, 28, 23) {real, imag} */,
  {32'hbfe8f344, 32'hc11e8616} /* (29, 28, 22) {real, imag} */,
  {32'h4020e28b, 32'hc16666ec} /* (29, 28, 21) {real, imag} */,
  {32'hc12d7468, 32'h4123988c} /* (29, 28, 20) {real, imag} */,
  {32'h40b01119, 32'h4178d3d8} /* (29, 28, 19) {real, imag} */,
  {32'hc09c403e, 32'hc07cb684} /* (29, 28, 18) {real, imag} */,
  {32'hc1214475, 32'h3f01c6e8} /* (29, 28, 17) {real, imag} */,
  {32'hc0a28a79, 32'h3f975a39} /* (29, 28, 16) {real, imag} */,
  {32'h412dada3, 32'h3f72dfa8} /* (29, 28, 15) {real, imag} */,
  {32'hc1bb638d, 32'h40535941} /* (29, 28, 14) {real, imag} */,
  {32'h4100ccfc, 32'h41386b56} /* (29, 28, 13) {real, imag} */,
  {32'hc0896b6e, 32'h41055abe} /* (29, 28, 12) {real, imag} */,
  {32'h3ff7d138, 32'h40ded278} /* (29, 28, 11) {real, imag} */,
  {32'h402a60fc, 32'h40b751f0} /* (29, 28, 10) {real, imag} */,
  {32'hc1821620, 32'h419be7ae} /* (29, 28, 9) {real, imag} */,
  {32'hc1431488, 32'hbf5d0a88} /* (29, 28, 8) {real, imag} */,
  {32'hc0eea136, 32'hbefc1050} /* (29, 28, 7) {real, imag} */,
  {32'h40b52336, 32'hc145bc19} /* (29, 28, 6) {real, imag} */,
  {32'hc26983fa, 32'hc1a5379e} /* (29, 28, 5) {real, imag} */,
  {32'h420c07fc, 32'h4036ad34} /* (29, 28, 4) {real, imag} */,
  {32'hc209de3a, 32'hc26e653c} /* (29, 28, 3) {real, imag} */,
  {32'hc299d5af, 32'h41fd2350} /* (29, 28, 2) {real, imag} */,
  {32'h42a757d7, 32'hc29cd0ce} /* (29, 28, 1) {real, imag} */,
  {32'h4253fc1a, 32'hc2071e66} /* (29, 28, 0) {real, imag} */,
  {32'hc291ac68, 32'h425e705c} /* (29, 27, 31) {real, imag} */,
  {32'h42246168, 32'h3f14cae0} /* (29, 27, 30) {real, imag} */,
  {32'h40c611ae, 32'h414938be} /* (29, 27, 29) {real, imag} */,
  {32'hc17e69bd, 32'h41038b41} /* (29, 27, 28) {real, imag} */,
  {32'hbf6208c0, 32'hc217000c} /* (29, 27, 27) {real, imag} */,
  {32'hc0b21746, 32'h413ccb46} /* (29, 27, 26) {real, imag} */,
  {32'h40aea345, 32'hc0449fa8} /* (29, 27, 25) {real, imag} */,
  {32'h40d950e5, 32'hbf751580} /* (29, 27, 24) {real, imag} */,
  {32'hc0112d60, 32'hbf93a558} /* (29, 27, 23) {real, imag} */,
  {32'hc186ab3e, 32'h40d4db47} /* (29, 27, 22) {real, imag} */,
  {32'h400a1da1, 32'h40dddeef} /* (29, 27, 21) {real, imag} */,
  {32'h4012dcda, 32'h3eab1660} /* (29, 27, 20) {real, imag} */,
  {32'hc0b3532a, 32'h406486fe} /* (29, 27, 19) {real, imag} */,
  {32'h4006e269, 32'h40a38b44} /* (29, 27, 18) {real, imag} */,
  {32'hbfe742d0, 32'hc09da836} /* (29, 27, 17) {real, imag} */,
  {32'h403405a2, 32'h40a23b46} /* (29, 27, 16) {real, imag} */,
  {32'h40b5f004, 32'hc09008ce} /* (29, 27, 15) {real, imag} */,
  {32'h405646e2, 32'hc00d6d65} /* (29, 27, 14) {real, imag} */,
  {32'h40dbbbea, 32'hbef22748} /* (29, 27, 13) {real, imag} */,
  {32'hc05a8138, 32'hc0b65176} /* (29, 27, 12) {real, imag} */,
  {32'h419ed5c1, 32'h40407660} /* (29, 27, 11) {real, imag} */,
  {32'h40693fec, 32'hc1ce8117} /* (29, 27, 10) {real, imag} */,
  {32'hc0eb3758, 32'h410f080e} /* (29, 27, 9) {real, imag} */,
  {32'hc0d9e0a2, 32'hbe59dd10} /* (29, 27, 8) {real, imag} */,
  {32'hc19da539, 32'hc121be85} /* (29, 27, 7) {real, imag} */,
  {32'h40b46253, 32'h417f8d9c} /* (29, 27, 6) {real, imag} */,
  {32'h4214df07, 32'hc1315bc9} /* (29, 27, 5) {real, imag} */,
  {32'hc1ab6320, 32'hc16612d7} /* (29, 27, 4) {real, imag} */,
  {32'h41574e96, 32'h41bddeb1} /* (29, 27, 3) {real, imag} */,
  {32'h40e5522e, 32'h41d81c36} /* (29, 27, 2) {real, imag} */,
  {32'hc2da22bc, 32'h419b92e9} /* (29, 27, 1) {real, imag} */,
  {32'hc279715a, 32'h4206368c} /* (29, 27, 0) {real, imag} */,
  {32'hc1d80c40, 32'hc15e2120} /* (29, 26, 31) {real, imag} */,
  {32'hbba0a800, 32'h4025bc9c} /* (29, 26, 30) {real, imag} */,
  {32'h408fcf25, 32'h3dc405c0} /* (29, 26, 29) {real, imag} */,
  {32'h41824f82, 32'h40cbf979} /* (29, 26, 28) {real, imag} */,
  {32'h40f182c8, 32'hbff41818} /* (29, 26, 27) {real, imag} */,
  {32'hbe8aae40, 32'hc070b19c} /* (29, 26, 26) {real, imag} */,
  {32'h41c3cc15, 32'hc12f472b} /* (29, 26, 25) {real, imag} */,
  {32'h3fea60de, 32'hc06e0e0c} /* (29, 26, 24) {real, imag} */,
  {32'h408476ac, 32'hc080ba64} /* (29, 26, 23) {real, imag} */,
  {32'h40c7ee34, 32'h4079e334} /* (29, 26, 22) {real, imag} */,
  {32'h3fe8176c, 32'hc1826d5e} /* (29, 26, 21) {real, imag} */,
  {32'h41600a5e, 32'hc16b9e9c} /* (29, 26, 20) {real, imag} */,
  {32'h41592c34, 32'hc0fc256f} /* (29, 26, 19) {real, imag} */,
  {32'hc1880b34, 32'hc0e35262} /* (29, 26, 18) {real, imag} */,
  {32'hc13061fd, 32'h410a2db6} /* (29, 26, 17) {real, imag} */,
  {32'h3fa3ecf0, 32'hc1007e58} /* (29, 26, 16) {real, imag} */,
  {32'hc103dbce, 32'hc0e069c6} /* (29, 26, 15) {real, imag} */,
  {32'h41433878, 32'hc0999570} /* (29, 26, 14) {real, imag} */,
  {32'h413a5d3a, 32'h41c160c0} /* (29, 26, 13) {real, imag} */,
  {32'hbfeaee8c, 32'h40a95d83} /* (29, 26, 12) {real, imag} */,
  {32'hc197e075, 32'h411f4a16} /* (29, 26, 11) {real, imag} */,
  {32'hc10d7024, 32'hc0aee5ef} /* (29, 26, 10) {real, imag} */,
  {32'h418e5da6, 32'h40f2fce8} /* (29, 26, 9) {real, imag} */,
  {32'hc1146fa1, 32'hc1dfc1da} /* (29, 26, 8) {real, imag} */,
  {32'h415d6bcc, 32'hc1ef1faa} /* (29, 26, 7) {real, imag} */,
  {32'hc13ce9f8, 32'h4065b973} /* (29, 26, 6) {real, imag} */,
  {32'hc207fe74, 32'hc06fb05f} /* (29, 26, 5) {real, imag} */,
  {32'hc0420a48, 32'h41b2fc21} /* (29, 26, 4) {real, imag} */,
  {32'h3dbbb3a0, 32'hbf86d348} /* (29, 26, 3) {real, imag} */,
  {32'h4180d86e, 32'hc1a2ee15} /* (29, 26, 2) {real, imag} */,
  {32'h415e14bc, 32'hc1ca7d0e} /* (29, 26, 1) {real, imag} */,
  {32'h411ef882, 32'hc138a253} /* (29, 26, 0) {real, imag} */,
  {32'h4237f53c, 32'hbfa91360} /* (29, 25, 31) {real, imag} */,
  {32'h41408744, 32'h40f15334} /* (29, 25, 30) {real, imag} */,
  {32'hc1bfa8c2, 32'h4136ea50} /* (29, 25, 29) {real, imag} */,
  {32'h3f4acd60, 32'h408a06cd} /* (29, 25, 28) {real, imag} */,
  {32'h408c9a26, 32'h41d92f99} /* (29, 25, 27) {real, imag} */,
  {32'h41cd13f4, 32'h4167a1ca} /* (29, 25, 26) {real, imag} */,
  {32'hc0695e04, 32'h412a0862} /* (29, 25, 25) {real, imag} */,
  {32'hc0ad8f49, 32'h4054b929} /* (29, 25, 24) {real, imag} */,
  {32'h4146f770, 32'hc14e263c} /* (29, 25, 23) {real, imag} */,
  {32'hc100e071, 32'h4064a56b} /* (29, 25, 22) {real, imag} */,
  {32'hc10b6491, 32'hc1822dce} /* (29, 25, 21) {real, imag} */,
  {32'h408b8dea, 32'h3fde3984} /* (29, 25, 20) {real, imag} */,
  {32'hc1684bb8, 32'hc06cff98} /* (29, 25, 19) {real, imag} */,
  {32'hbfaad8a4, 32'h40c4e83c} /* (29, 25, 18) {real, imag} */,
  {32'hbeb7fe10, 32'h4017c0e0} /* (29, 25, 17) {real, imag} */,
  {32'h403b379a, 32'h4106b1d8} /* (29, 25, 16) {real, imag} */,
  {32'hc1813f4c, 32'h41264641} /* (29, 25, 15) {real, imag} */,
  {32'h4127c3a6, 32'hc08110bc} /* (29, 25, 14) {real, imag} */,
  {32'h41260a35, 32'hc0befc9a} /* (29, 25, 13) {real, imag} */,
  {32'h40fe2e4d, 32'hbf091f00} /* (29, 25, 12) {real, imag} */,
  {32'hc072c9fc, 32'hc12a4c4f} /* (29, 25, 11) {real, imag} */,
  {32'hc0ceef20, 32'hc1a8d10e} /* (29, 25, 10) {real, imag} */,
  {32'h3d7d6300, 32'h412a06d7} /* (29, 25, 9) {real, imag} */,
  {32'hbf08042a, 32'h40b8d04b} /* (29, 25, 8) {real, imag} */,
  {32'hc17df12b, 32'hc0daeb8b} /* (29, 25, 7) {real, imag} */,
  {32'hc0b9af4a, 32'hbd3e1700} /* (29, 25, 6) {real, imag} */,
  {32'h41285846, 32'hc1b0d7c9} /* (29, 25, 5) {real, imag} */,
  {32'hc1a1fc78, 32'h40b4d244} /* (29, 25, 4) {real, imag} */,
  {32'hc122feaf, 32'hbfa7a23c} /* (29, 25, 3) {real, imag} */,
  {32'hc1938f1c, 32'hc1dc0515} /* (29, 25, 2) {real, imag} */,
  {32'hc067bc7e, 32'h410ce8fa} /* (29, 25, 1) {real, imag} */,
  {32'h421315c2, 32'h4055a24c} /* (29, 25, 0) {real, imag} */,
  {32'hc18c2148, 32'h422ca212} /* (29, 24, 31) {real, imag} */,
  {32'hc0aafe14, 32'h4163f56f} /* (29, 24, 30) {real, imag} */,
  {32'h41d554d8, 32'hc1a2e601} /* (29, 24, 29) {real, imag} */,
  {32'hc0be2ea7, 32'h4107af7c} /* (29, 24, 28) {real, imag} */,
  {32'h410896a8, 32'hc175af81} /* (29, 24, 27) {real, imag} */,
  {32'hc13d9f33, 32'hc16cfabc} /* (29, 24, 26) {real, imag} */,
  {32'hc16f64fa, 32'hc0140df7} /* (29, 24, 25) {real, imag} */,
  {32'h4073bfb0, 32'hc0baa950} /* (29, 24, 24) {real, imag} */,
  {32'hc119ed08, 32'h40f5475e} /* (29, 24, 23) {real, imag} */,
  {32'h411fbc46, 32'h412f67fa} /* (29, 24, 22) {real, imag} */,
  {32'hbf0bec78, 32'hc1d2b48e} /* (29, 24, 21) {real, imag} */,
  {32'hc0607c02, 32'hc0eb9c1a} /* (29, 24, 20) {real, imag} */,
  {32'h41bcf1e7, 32'hc08f413a} /* (29, 24, 19) {real, imag} */,
  {32'hbf552eb0, 32'h4102907d} /* (29, 24, 18) {real, imag} */,
  {32'h41063393, 32'hbe4d4fc0} /* (29, 24, 17) {real, imag} */,
  {32'h411d3ae3, 32'hc0edb3e6} /* (29, 24, 16) {real, imag} */,
  {32'hbe16f480, 32'hc0686fa6} /* (29, 24, 15) {real, imag} */,
  {32'h415324bd, 32'h415adac9} /* (29, 24, 14) {real, imag} */,
  {32'hc13528bb, 32'hc0810c29} /* (29, 24, 13) {real, imag} */,
  {32'hc0fd21e6, 32'h40e07c79} /* (29, 24, 12) {real, imag} */,
  {32'h4178ce4c, 32'hc1647cee} /* (29, 24, 11) {real, imag} */,
  {32'h41af30de, 32'h41220684} /* (29, 24, 10) {real, imag} */,
  {32'hc0e78150, 32'h400e0fab} /* (29, 24, 9) {real, imag} */,
  {32'h3f940f90, 32'hbf9534b0} /* (29, 24, 8) {real, imag} */,
  {32'hc12d3a13, 32'h41b215bc} /* (29, 24, 7) {real, imag} */,
  {32'h41451a58, 32'h4101e3a0} /* (29, 24, 6) {real, imag} */,
  {32'hc16bd34d, 32'h40854d50} /* (29, 24, 5) {real, imag} */,
  {32'h411dc24c, 32'h40e2ce16} /* (29, 24, 4) {real, imag} */,
  {32'hbfd55d70, 32'h41bddbb4} /* (29, 24, 3) {real, imag} */,
  {32'h41d44fbc, 32'hc19a93fd} /* (29, 24, 2) {real, imag} */,
  {32'hc273bd9a, 32'h4226fe51} /* (29, 24, 1) {real, imag} */,
  {32'hc1866be3, 32'h40ecc587} /* (29, 24, 0) {real, imag} */,
  {32'h41ce3aae, 32'h402618c0} /* (29, 23, 31) {real, imag} */,
  {32'hc1c02127, 32'h41834bcc} /* (29, 23, 30) {real, imag} */,
  {32'hc148c264, 32'hc03ee9ba} /* (29, 23, 29) {real, imag} */,
  {32'h3fb6dd06, 32'h3fc9c147} /* (29, 23, 28) {real, imag} */,
  {32'h409fd260, 32'hc1cd0b14} /* (29, 23, 27) {real, imag} */,
  {32'h40ed125e, 32'h3fb22ba9} /* (29, 23, 26) {real, imag} */,
  {32'hc0605c1a, 32'h40fa94a6} /* (29, 23, 25) {real, imag} */,
  {32'h41632176, 32'h40e07702} /* (29, 23, 24) {real, imag} */,
  {32'hc10b4b9e, 32'h3dad58c0} /* (29, 23, 23) {real, imag} */,
  {32'hc1baa175, 32'hc056bba8} /* (29, 23, 22) {real, imag} */,
  {32'h3e3a46b0, 32'h40da6d4f} /* (29, 23, 21) {real, imag} */,
  {32'h411cbcc0, 32'hc12104bd} /* (29, 23, 20) {real, imag} */,
  {32'hc15e9694, 32'hc1854fae} /* (29, 23, 19) {real, imag} */,
  {32'hc0ed99bb, 32'hc1885a56} /* (29, 23, 18) {real, imag} */,
  {32'hc06e75a7, 32'hc0d9ecc3} /* (29, 23, 17) {real, imag} */,
  {32'h415f7688, 32'h40fac36d} /* (29, 23, 16) {real, imag} */,
  {32'hc10b350c, 32'h4107cac0} /* (29, 23, 15) {real, imag} */,
  {32'h4149cf49, 32'hc0ae3d66} /* (29, 23, 14) {real, imag} */,
  {32'h4153fefe, 32'hc1ab96ae} /* (29, 23, 13) {real, imag} */,
  {32'hc0d79ffe, 32'h418e8cc6} /* (29, 23, 12) {real, imag} */,
  {32'hc14f2d0e, 32'h4109a696} /* (29, 23, 11) {real, imag} */,
  {32'hc1f04259, 32'h413d588e} /* (29, 23, 10) {real, imag} */,
  {32'hc0d53f06, 32'hc155ebef} /* (29, 23, 9) {real, imag} */,
  {32'h4083e961, 32'h410b2d18} /* (29, 23, 8) {real, imag} */,
  {32'hc1392f02, 32'hc05ce680} /* (29, 23, 7) {real, imag} */,
  {32'hc02a9e82, 32'hc15dbb75} /* (29, 23, 6) {real, imag} */,
  {32'hc151f940, 32'hc094e59e} /* (29, 23, 5) {real, imag} */,
  {32'hbf6141d8, 32'hc1efc942} /* (29, 23, 4) {real, imag} */,
  {32'h4100e1f9, 32'h3e1a2040} /* (29, 23, 3) {real, imag} */,
  {32'h41f00e87, 32'h407b6408} /* (29, 23, 2) {real, imag} */,
  {32'hc21d4b78, 32'hc12fedfd} /* (29, 23, 1) {real, imag} */,
  {32'hc15b22aa, 32'h41933602} /* (29, 23, 0) {real, imag} */,
  {32'h3f74b9b0, 32'h3ffec1f8} /* (29, 22, 31) {real, imag} */,
  {32'h3ff663b8, 32'hc06dcbda} /* (29, 22, 30) {real, imag} */,
  {32'hc1a8222c, 32'h3f882e0e} /* (29, 22, 29) {real, imag} */,
  {32'hc1a5fbab, 32'h418ca5de} /* (29, 22, 28) {real, imag} */,
  {32'hc1242e18, 32'hc00cda36} /* (29, 22, 27) {real, imag} */,
  {32'h41165c5e, 32'h414ad827} /* (29, 22, 26) {real, imag} */,
  {32'h414935dc, 32'h41538068} /* (29, 22, 25) {real, imag} */,
  {32'hc0d98cdb, 32'hc10b345d} /* (29, 22, 24) {real, imag} */,
  {32'hc10ad5a8, 32'hc07ea94f} /* (29, 22, 23) {real, imag} */,
  {32'h40896bcc, 32'hc138ed01} /* (29, 22, 22) {real, imag} */,
  {32'h417b1dd4, 32'hc086643c} /* (29, 22, 21) {real, imag} */,
  {32'h40ac7e6a, 32'hc17c905a} /* (29, 22, 20) {real, imag} */,
  {32'hc19a7738, 32'hc0357cd4} /* (29, 22, 19) {real, imag} */,
  {32'h41ac238a, 32'h3f06ee38} /* (29, 22, 18) {real, imag} */,
  {32'h4170d46d, 32'h40dc259e} /* (29, 22, 17) {real, imag} */,
  {32'hc14fa086, 32'hc0d3c999} /* (29, 22, 16) {real, imag} */,
  {32'h3eedba88, 32'hc07e5fa2} /* (29, 22, 15) {real, imag} */,
  {32'h400a3a04, 32'hc0de0e08} /* (29, 22, 14) {real, imag} */,
  {32'h4100663a, 32'h414d31a0} /* (29, 22, 13) {real, imag} */,
  {32'h4125c536, 32'h41151ed2} /* (29, 22, 12) {real, imag} */,
  {32'h408d77a2, 32'h40f7c95c} /* (29, 22, 11) {real, imag} */,
  {32'h4006baee, 32'hc1abb94a} /* (29, 22, 10) {real, imag} */,
  {32'hc1749658, 32'hc0b99fe2} /* (29, 22, 9) {real, imag} */,
  {32'hc04c0f8a, 32'h41b1cc43} /* (29, 22, 8) {real, imag} */,
  {32'h410fb50b, 32'hc1147ef8} /* (29, 22, 7) {real, imag} */,
  {32'h408dd4ca, 32'h4161c73e} /* (29, 22, 6) {real, imag} */,
  {32'h4182ceb2, 32'h41545c67} /* (29, 22, 5) {real, imag} */,
  {32'h403d040a, 32'hbf4f1120} /* (29, 22, 4) {real, imag} */,
  {32'h411fd5c0, 32'hc1431c44} /* (29, 22, 3) {real, imag} */,
  {32'h4088d53f, 32'h410a0253} /* (29, 22, 2) {real, imag} */,
  {32'h41893280, 32'hc0e251be} /* (29, 22, 1) {real, imag} */,
  {32'hc1840ff1, 32'hc0c2fdb9} /* (29, 22, 0) {real, imag} */,
  {32'hc02d1db6, 32'h41e8f050} /* (29, 21, 31) {real, imag} */,
  {32'hc08ca481, 32'hc201279d} /* (29, 21, 30) {real, imag} */,
  {32'hc031742e, 32'hc0a5b40a} /* (29, 21, 29) {real, imag} */,
  {32'hc17e4fe0, 32'hc18673a6} /* (29, 21, 28) {real, imag} */,
  {32'hc110ef5f, 32'hc18a923c} /* (29, 21, 27) {real, imag} */,
  {32'hc16a89be, 32'hc15f8912} /* (29, 21, 26) {real, imag} */,
  {32'hbfb14d3e, 32'hc0b2f829} /* (29, 21, 25) {real, imag} */,
  {32'h40ae3a98, 32'hc12fe429} /* (29, 21, 24) {real, imag} */,
  {32'h41cd18fc, 32'hc022d232} /* (29, 21, 23) {real, imag} */,
  {32'h418d3517, 32'h4035bba6} /* (29, 21, 22) {real, imag} */,
  {32'hc0f9ada9, 32'h400e350a} /* (29, 21, 21) {real, imag} */,
  {32'h40f09d21, 32'h40e4a33d} /* (29, 21, 20) {real, imag} */,
  {32'hc114815e, 32'h40309f50} /* (29, 21, 19) {real, imag} */,
  {32'hc0538ea9, 32'h41810ee0} /* (29, 21, 18) {real, imag} */,
  {32'hc18a0f4c, 32'hc09d8042} /* (29, 21, 17) {real, imag} */,
  {32'hc0a74d4e, 32'h4047046c} /* (29, 21, 16) {real, imag} */,
  {32'h3f34fd70, 32'hc0a68cac} /* (29, 21, 15) {real, imag} */,
  {32'hc135e27a, 32'h411b7e1e} /* (29, 21, 14) {real, imag} */,
  {32'h4161e42e, 32'h3f168420} /* (29, 21, 13) {real, imag} */,
  {32'h41015a29, 32'h40fcdc92} /* (29, 21, 12) {real, imag} */,
  {32'h41071699, 32'h4188a7f0} /* (29, 21, 11) {real, imag} */,
  {32'hc1b02278, 32'hc0d1fb2a} /* (29, 21, 10) {real, imag} */,
  {32'hc0bb9e5e, 32'hc11154d4} /* (29, 21, 9) {real, imag} */,
  {32'hc1198ce8, 32'h4058c814} /* (29, 21, 8) {real, imag} */,
  {32'h41408d4c, 32'hc0c57db5} /* (29, 21, 7) {real, imag} */,
  {32'hc140c734, 32'hc11f8e09} /* (29, 21, 6) {real, imag} */,
  {32'h400de658, 32'h4180de65} /* (29, 21, 5) {real, imag} */,
  {32'h415fd46e, 32'hc0378fbf} /* (29, 21, 4) {real, imag} */,
  {32'h41357124, 32'h402d3ed4} /* (29, 21, 3) {real, imag} */,
  {32'h4081b80b, 32'hc155cd53} /* (29, 21, 2) {real, imag} */,
  {32'hc0f1669e, 32'h4137be2a} /* (29, 21, 1) {real, imag} */,
  {32'hc1c8c8d5, 32'h41e190a6} /* (29, 21, 0) {real, imag} */,
  {32'h40847005, 32'h4009a964} /* (29, 20, 31) {real, imag} */,
  {32'hc1967eae, 32'h3f168e10} /* (29, 20, 30) {real, imag} */,
  {32'h4001bb26, 32'hc099f5d0} /* (29, 20, 29) {real, imag} */,
  {32'hc046f93c, 32'h413bc80d} /* (29, 20, 28) {real, imag} */,
  {32'h3eb310d8, 32'hc1010fb9} /* (29, 20, 27) {real, imag} */,
  {32'h409ad192, 32'h3ffc850e} /* (29, 20, 26) {real, imag} */,
  {32'hc12c6ea6, 32'h4136ffd2} /* (29, 20, 25) {real, imag} */,
  {32'hc19d60be, 32'hbfaf4ba0} /* (29, 20, 24) {real, imag} */,
  {32'h40999126, 32'h400b8296} /* (29, 20, 23) {real, imag} */,
  {32'hc1548e53, 32'hc0059a5c} /* (29, 20, 22) {real, imag} */,
  {32'h4121d2d3, 32'h4185c4bf} /* (29, 20, 21) {real, imag} */,
  {32'hc0913716, 32'hc16658ad} /* (29, 20, 20) {real, imag} */,
  {32'h40b32ed5, 32'h40f687fc} /* (29, 20, 19) {real, imag} */,
  {32'hc107228e, 32'h409da82e} /* (29, 20, 18) {real, imag} */,
  {32'h409fb6de, 32'hc0434418} /* (29, 20, 17) {real, imag} */,
  {32'hc0a0e8e4, 32'hbebc7b30} /* (29, 20, 16) {real, imag} */,
  {32'hbff1b190, 32'h3fe90a0c} /* (29, 20, 15) {real, imag} */,
  {32'h40ff429a, 32'hc0eea53f} /* (29, 20, 14) {real, imag} */,
  {32'h3f22587f, 32'hc0e58bcc} /* (29, 20, 13) {real, imag} */,
  {32'h405aa03d, 32'hc0ec6b61} /* (29, 20, 12) {real, imag} */,
  {32'hc1451336, 32'hc131647c} /* (29, 20, 11) {real, imag} */,
  {32'hc08abd26, 32'h419835cc} /* (29, 20, 10) {real, imag} */,
  {32'hc18be8cd, 32'h3fd7e876} /* (29, 20, 9) {real, imag} */,
  {32'h402a7c00, 32'hc068fc05} /* (29, 20, 8) {real, imag} */,
  {32'hc0f58c0c, 32'h4141bfd4} /* (29, 20, 7) {real, imag} */,
  {32'h404dbab0, 32'hc1096148} /* (29, 20, 6) {real, imag} */,
  {32'h3fb7ef96, 32'h412d2b92} /* (29, 20, 5) {real, imag} */,
  {32'h41b97dd8, 32'h3f3fae98} /* (29, 20, 4) {real, imag} */,
  {32'hc09eff65, 32'hc1841617} /* (29, 20, 3) {real, imag} */,
  {32'h40cf02d0, 32'hc084ae80} /* (29, 20, 2) {real, imag} */,
  {32'h40ecb2d6, 32'hc1211ae9} /* (29, 20, 1) {real, imag} */,
  {32'hc0856e92, 32'h40affb60} /* (29, 20, 0) {real, imag} */,
  {32'h40d4a2ee, 32'hc117d557} /* (29, 19, 31) {real, imag} */,
  {32'h3ed770fc, 32'h418ba3cd} /* (29, 19, 30) {real, imag} */,
  {32'h412cb908, 32'h40de57a6} /* (29, 19, 29) {real, imag} */,
  {32'h412547c9, 32'hbed9a290} /* (29, 19, 28) {real, imag} */,
  {32'hc18caf56, 32'h4126147f} /* (29, 19, 27) {real, imag} */,
  {32'h40867b7c, 32'hbfd1cc44} /* (29, 19, 26) {real, imag} */,
  {32'h401b16a4, 32'h40299531} /* (29, 19, 25) {real, imag} */,
  {32'hc0eba2e8, 32'hbf924400} /* (29, 19, 24) {real, imag} */,
  {32'hc17e61ae, 32'h3ffce973} /* (29, 19, 23) {real, imag} */,
  {32'hc100cf90, 32'hc0a9573e} /* (29, 19, 22) {real, imag} */,
  {32'hc07d5ab4, 32'h408848ca} /* (29, 19, 21) {real, imag} */,
  {32'h41169ef8, 32'h41340c84} /* (29, 19, 20) {real, imag} */,
  {32'h40c973af, 32'h40c4c7bb} /* (29, 19, 19) {real, imag} */,
  {32'h41849638, 32'h4071d478} /* (29, 19, 18) {real, imag} */,
  {32'hbfb505dc, 32'hc1a54efe} /* (29, 19, 17) {real, imag} */,
  {32'hbfd0d4c0, 32'h4066795e} /* (29, 19, 16) {real, imag} */,
  {32'hc080ecc7, 32'h411a0e5c} /* (29, 19, 15) {real, imag} */,
  {32'hc0f1bd1f, 32'h40728fd4} /* (29, 19, 14) {real, imag} */,
  {32'h405e8208, 32'h3ec06b20} /* (29, 19, 13) {real, imag} */,
  {32'hbfbdbbd4, 32'hc106436c} /* (29, 19, 12) {real, imag} */,
  {32'h41698bfc, 32'hc11ae316} /* (29, 19, 11) {real, imag} */,
  {32'hc08feb33, 32'h4133276c} /* (29, 19, 10) {real, imag} */,
  {32'h4148dc6a, 32'hc19cab74} /* (29, 19, 9) {real, imag} */,
  {32'h40b87803, 32'h407f2c93} /* (29, 19, 8) {real, imag} */,
  {32'hc065fabc, 32'h410e6d62} /* (29, 19, 7) {real, imag} */,
  {32'h4187376e, 32'h408685e3} /* (29, 19, 6) {real, imag} */,
  {32'h4051b777, 32'hc03b4199} /* (29, 19, 5) {real, imag} */,
  {32'h405b3e8a, 32'h400be55c} /* (29, 19, 4) {real, imag} */,
  {32'hc16aabeb, 32'hc1635331} /* (29, 19, 3) {real, imag} */,
  {32'h416358bc, 32'h40eed2cc} /* (29, 19, 2) {real, imag} */,
  {32'hbf22fcb0, 32'hbfd95910} /* (29, 19, 1) {real, imag} */,
  {32'h41a12d44, 32'hc1445c50} /* (29, 19, 0) {real, imag} */,
  {32'hc0fa2e6d, 32'h410707ee} /* (29, 18, 31) {real, imag} */,
  {32'hbfa467bc, 32'hc0ff90b0} /* (29, 18, 30) {real, imag} */,
  {32'hc1232008, 32'hc136105d} /* (29, 18, 29) {real, imag} */,
  {32'hc152f3f5, 32'hc148d664} /* (29, 18, 28) {real, imag} */,
  {32'hc1724c12, 32'hc0c658ea} /* (29, 18, 27) {real, imag} */,
  {32'h40ad07bc, 32'hc0f2cf76} /* (29, 18, 26) {real, imag} */,
  {32'hc19ef27f, 32'hc1363de2} /* (29, 18, 25) {real, imag} */,
  {32'h40ad8112, 32'h40aaf467} /* (29, 18, 24) {real, imag} */,
  {32'h41c8eb5d, 32'h4181a58b} /* (29, 18, 23) {real, imag} */,
  {32'hc0d60cb1, 32'h419a111f} /* (29, 18, 22) {real, imag} */,
  {32'hc0d3f290, 32'hc1215912} /* (29, 18, 21) {real, imag} */,
  {32'hc1806a97, 32'h41005194} /* (29, 18, 20) {real, imag} */,
  {32'h411b7695, 32'h411f1686} /* (29, 18, 19) {real, imag} */,
  {32'hc0daf0ef, 32'h40804178} /* (29, 18, 18) {real, imag} */,
  {32'hbfb157b4, 32'h40f9927c} /* (29, 18, 17) {real, imag} */,
  {32'h410a6f9c, 32'h409b0381} /* (29, 18, 16) {real, imag} */,
  {32'hbfa1cfba, 32'hc07bf516} /* (29, 18, 15) {real, imag} */,
  {32'h41047f12, 32'h3fbfbe30} /* (29, 18, 14) {real, imag} */,
  {32'hbfb2b52e, 32'h3fee57c8} /* (29, 18, 13) {real, imag} */,
  {32'h40123474, 32'h40ecdd78} /* (29, 18, 12) {real, imag} */,
  {32'hbf9302e3, 32'h41af83af} /* (29, 18, 11) {real, imag} */,
  {32'h41200cc8, 32'h3fc34d1a} /* (29, 18, 10) {real, imag} */,
  {32'hbf82a664, 32'h3db603d0} /* (29, 18, 9) {real, imag} */,
  {32'h4082645b, 32'h3f84a8a0} /* (29, 18, 8) {real, imag} */,
  {32'hc0b68c7a, 32'hc096c349} /* (29, 18, 7) {real, imag} */,
  {32'hc1074b84, 32'h412ba979} /* (29, 18, 6) {real, imag} */,
  {32'h410dbc0c, 32'hc11b8340} /* (29, 18, 5) {real, imag} */,
  {32'h3f1bf610, 32'h3f922038} /* (29, 18, 4) {real, imag} */,
  {32'h40a8f0e9, 32'h4186260c} /* (29, 18, 3) {real, imag} */,
  {32'hc0316950, 32'h40746d44} /* (29, 18, 2) {real, imag} */,
  {32'hc0bacb3a, 32'h40c76a52} /* (29, 18, 1) {real, imag} */,
  {32'hc0aa0964, 32'h416009d4} /* (29, 18, 0) {real, imag} */,
  {32'h40ab920e, 32'hc0b73a0e} /* (29, 17, 31) {real, imag} */,
  {32'h3fc38797, 32'h402d04a4} /* (29, 17, 30) {real, imag} */,
  {32'h40c82168, 32'h3f7ba950} /* (29, 17, 29) {real, imag} */,
  {32'hbfe184d4, 32'h40f05478} /* (29, 17, 28) {real, imag} */,
  {32'hc1135174, 32'hbc8d9140} /* (29, 17, 27) {real, imag} */,
  {32'hc10c1689, 32'hc04a48bc} /* (29, 17, 26) {real, imag} */,
  {32'h4051e19f, 32'h402d99e6} /* (29, 17, 25) {real, imag} */,
  {32'h3f741c9a, 32'h41152ed5} /* (29, 17, 24) {real, imag} */,
  {32'hc0db7497, 32'h40dfe5a6} /* (29, 17, 23) {real, imag} */,
  {32'hc0ec8c82, 32'hbf1f1510} /* (29, 17, 22) {real, imag} */,
  {32'h4182d0aa, 32'hc04da594} /* (29, 17, 21) {real, imag} */,
  {32'h413c3036, 32'h418f8754} /* (29, 17, 20) {real, imag} */,
  {32'hbf8cd7e4, 32'h40be1c3a} /* (29, 17, 19) {real, imag} */,
  {32'h3f8800bc, 32'h402f6958} /* (29, 17, 18) {real, imag} */,
  {32'hc095f09a, 32'h3f905943} /* (29, 17, 17) {real, imag} */,
  {32'hc0423242, 32'h40d7c8c1} /* (29, 17, 16) {real, imag} */,
  {32'hbe155bc0, 32'h3fdc3074} /* (29, 17, 15) {real, imag} */,
  {32'h4111214b, 32'h4070ae3d} /* (29, 17, 14) {real, imag} */,
  {32'h41170064, 32'h40b6ba7e} /* (29, 17, 13) {real, imag} */,
  {32'hc11e7f3b, 32'hc0ac8158} /* (29, 17, 12) {real, imag} */,
  {32'h413fc9da, 32'hbe3c8950} /* (29, 17, 11) {real, imag} */,
  {32'hc0bc3cca, 32'hc09ab975} /* (29, 17, 10) {real, imag} */,
  {32'hbff08154, 32'h41279397} /* (29, 17, 9) {real, imag} */,
  {32'h4125993c, 32'hc196bb08} /* (29, 17, 8) {real, imag} */,
  {32'h4151aa62, 32'h40445adf} /* (29, 17, 7) {real, imag} */,
  {32'h40b6eef4, 32'hc19484af} /* (29, 17, 6) {real, imag} */,
  {32'h403ea870, 32'h3ebab560} /* (29, 17, 5) {real, imag} */,
  {32'hc1081ff2, 32'h410713df} /* (29, 17, 4) {real, imag} */,
  {32'h40a8ab0c, 32'hc141c69a} /* (29, 17, 3) {real, imag} */,
  {32'h414daac1, 32'h404bfdf2} /* (29, 17, 2) {real, imag} */,
  {32'hc078e9f0, 32'hc108e117} /* (29, 17, 1) {real, imag} */,
  {32'h408800ae, 32'hc0031845} /* (29, 17, 0) {real, imag} */,
  {32'hbf155428, 32'hc039a658} /* (29, 16, 31) {real, imag} */,
  {32'h411e2693, 32'h4095f4bc} /* (29, 16, 30) {real, imag} */,
  {32'hbf7f918e, 32'hc0df2856} /* (29, 16, 29) {real, imag} */,
  {32'hbf650b2c, 32'hc0559718} /* (29, 16, 28) {real, imag} */,
  {32'h4120a2a8, 32'h40e37287} /* (29, 16, 27) {real, imag} */,
  {32'hc08276d9, 32'hbf9b1aa8} /* (29, 16, 26) {real, imag} */,
  {32'hbfbd5c3f, 32'h411015cc} /* (29, 16, 25) {real, imag} */,
  {32'hc115e63a, 32'hc03b1ea2} /* (29, 16, 24) {real, imag} */,
  {32'h416812e0, 32'h415865a5} /* (29, 16, 23) {real, imag} */,
  {32'hc0fa732f, 32'h3fa336c4} /* (29, 16, 22) {real, imag} */,
  {32'hc1305132, 32'hc1033e4f} /* (29, 16, 21) {real, imag} */,
  {32'hbfae88b0, 32'hc0ea9dac} /* (29, 16, 20) {real, imag} */,
  {32'hc09d1c89, 32'h403a2b30} /* (29, 16, 19) {real, imag} */,
  {32'h418ec182, 32'hc0739af2} /* (29, 16, 18) {real, imag} */,
  {32'h4019de53, 32'hc06537fe} /* (29, 16, 17) {real, imag} */,
  {32'hbfc1b8d5, 32'h00000000} /* (29, 16, 16) {real, imag} */,
  {32'h4019de53, 32'h406537fe} /* (29, 16, 15) {real, imag} */,
  {32'h418ec182, 32'h40739af2} /* (29, 16, 14) {real, imag} */,
  {32'hc09d1c89, 32'hc03a2b30} /* (29, 16, 13) {real, imag} */,
  {32'hbfae88b0, 32'h40ea9dac} /* (29, 16, 12) {real, imag} */,
  {32'hc1305132, 32'h41033e4f} /* (29, 16, 11) {real, imag} */,
  {32'hc0fa732f, 32'hbfa336c4} /* (29, 16, 10) {real, imag} */,
  {32'h416812e0, 32'hc15865a5} /* (29, 16, 9) {real, imag} */,
  {32'hc115e63a, 32'h403b1ea2} /* (29, 16, 8) {real, imag} */,
  {32'hbfbd5c3f, 32'hc11015cc} /* (29, 16, 7) {real, imag} */,
  {32'hc08276d9, 32'h3f9b1aa8} /* (29, 16, 6) {real, imag} */,
  {32'h4120a2a8, 32'hc0e37287} /* (29, 16, 5) {real, imag} */,
  {32'hbf650b2c, 32'h40559718} /* (29, 16, 4) {real, imag} */,
  {32'hbf7f918e, 32'h40df2856} /* (29, 16, 3) {real, imag} */,
  {32'h411e2693, 32'hc095f4bc} /* (29, 16, 2) {real, imag} */,
  {32'hbf155428, 32'h4039a658} /* (29, 16, 1) {real, imag} */,
  {32'h411952a2, 32'h00000000} /* (29, 16, 0) {real, imag} */,
  {32'hc078e9f0, 32'h4108e117} /* (29, 15, 31) {real, imag} */,
  {32'h414daac1, 32'hc04bfdf2} /* (29, 15, 30) {real, imag} */,
  {32'h40a8ab0c, 32'h4141c69a} /* (29, 15, 29) {real, imag} */,
  {32'hc1081ff2, 32'hc10713df} /* (29, 15, 28) {real, imag} */,
  {32'h403ea870, 32'hbebab560} /* (29, 15, 27) {real, imag} */,
  {32'h40b6eef4, 32'h419484af} /* (29, 15, 26) {real, imag} */,
  {32'h4151aa62, 32'hc0445adf} /* (29, 15, 25) {real, imag} */,
  {32'h4125993c, 32'h4196bb08} /* (29, 15, 24) {real, imag} */,
  {32'hbff08154, 32'hc1279397} /* (29, 15, 23) {real, imag} */,
  {32'hc0bc3cca, 32'h409ab975} /* (29, 15, 22) {real, imag} */,
  {32'h413fc9da, 32'h3e3c8950} /* (29, 15, 21) {real, imag} */,
  {32'hc11e7f3b, 32'h40ac8158} /* (29, 15, 20) {real, imag} */,
  {32'h41170064, 32'hc0b6ba7e} /* (29, 15, 19) {real, imag} */,
  {32'h4111214b, 32'hc070ae3d} /* (29, 15, 18) {real, imag} */,
  {32'hbe155bc0, 32'hbfdc3074} /* (29, 15, 17) {real, imag} */,
  {32'hc0423242, 32'hc0d7c8c1} /* (29, 15, 16) {real, imag} */,
  {32'hc095f09a, 32'hbf905943} /* (29, 15, 15) {real, imag} */,
  {32'h3f8800bc, 32'hc02f6958} /* (29, 15, 14) {real, imag} */,
  {32'hbf8cd7e4, 32'hc0be1c3a} /* (29, 15, 13) {real, imag} */,
  {32'h413c3036, 32'hc18f8754} /* (29, 15, 12) {real, imag} */,
  {32'h4182d0aa, 32'h404da594} /* (29, 15, 11) {real, imag} */,
  {32'hc0ec8c82, 32'h3f1f1510} /* (29, 15, 10) {real, imag} */,
  {32'hc0db7497, 32'hc0dfe5a6} /* (29, 15, 9) {real, imag} */,
  {32'h3f741c9a, 32'hc1152ed5} /* (29, 15, 8) {real, imag} */,
  {32'h4051e19f, 32'hc02d99e6} /* (29, 15, 7) {real, imag} */,
  {32'hc10c1689, 32'h404a48bc} /* (29, 15, 6) {real, imag} */,
  {32'hc1135174, 32'h3c8d9140} /* (29, 15, 5) {real, imag} */,
  {32'hbfe184d4, 32'hc0f05478} /* (29, 15, 4) {real, imag} */,
  {32'h40c82168, 32'hbf7ba950} /* (29, 15, 3) {real, imag} */,
  {32'h3fc38797, 32'hc02d04a4} /* (29, 15, 2) {real, imag} */,
  {32'h40ab920e, 32'h40b73a0e} /* (29, 15, 1) {real, imag} */,
  {32'h408800ae, 32'h40031845} /* (29, 15, 0) {real, imag} */,
  {32'hc0bacb3a, 32'hc0c76a52} /* (29, 14, 31) {real, imag} */,
  {32'hc0316950, 32'hc0746d44} /* (29, 14, 30) {real, imag} */,
  {32'h40a8f0e9, 32'hc186260c} /* (29, 14, 29) {real, imag} */,
  {32'h3f1bf610, 32'hbf922038} /* (29, 14, 28) {real, imag} */,
  {32'h410dbc0c, 32'h411b8340} /* (29, 14, 27) {real, imag} */,
  {32'hc1074b84, 32'hc12ba979} /* (29, 14, 26) {real, imag} */,
  {32'hc0b68c7a, 32'h4096c349} /* (29, 14, 25) {real, imag} */,
  {32'h4082645b, 32'hbf84a8a0} /* (29, 14, 24) {real, imag} */,
  {32'hbf82a664, 32'hbdb603d0} /* (29, 14, 23) {real, imag} */,
  {32'h41200cc8, 32'hbfc34d1a} /* (29, 14, 22) {real, imag} */,
  {32'hbf9302e3, 32'hc1af83af} /* (29, 14, 21) {real, imag} */,
  {32'h40123474, 32'hc0ecdd78} /* (29, 14, 20) {real, imag} */,
  {32'hbfb2b52e, 32'hbfee57c8} /* (29, 14, 19) {real, imag} */,
  {32'h41047f12, 32'hbfbfbe30} /* (29, 14, 18) {real, imag} */,
  {32'hbfa1cfba, 32'h407bf516} /* (29, 14, 17) {real, imag} */,
  {32'h410a6f9c, 32'hc09b0381} /* (29, 14, 16) {real, imag} */,
  {32'hbfb157b4, 32'hc0f9927c} /* (29, 14, 15) {real, imag} */,
  {32'hc0daf0ef, 32'hc0804178} /* (29, 14, 14) {real, imag} */,
  {32'h411b7695, 32'hc11f1686} /* (29, 14, 13) {real, imag} */,
  {32'hc1806a97, 32'hc1005194} /* (29, 14, 12) {real, imag} */,
  {32'hc0d3f290, 32'h41215912} /* (29, 14, 11) {real, imag} */,
  {32'hc0d60cb1, 32'hc19a111f} /* (29, 14, 10) {real, imag} */,
  {32'h41c8eb5d, 32'hc181a58b} /* (29, 14, 9) {real, imag} */,
  {32'h40ad8112, 32'hc0aaf467} /* (29, 14, 8) {real, imag} */,
  {32'hc19ef27f, 32'h41363de2} /* (29, 14, 7) {real, imag} */,
  {32'h40ad07bc, 32'h40f2cf76} /* (29, 14, 6) {real, imag} */,
  {32'hc1724c12, 32'h40c658ea} /* (29, 14, 5) {real, imag} */,
  {32'hc152f3f5, 32'h4148d664} /* (29, 14, 4) {real, imag} */,
  {32'hc1232008, 32'h4136105d} /* (29, 14, 3) {real, imag} */,
  {32'hbfa467bc, 32'h40ff90b0} /* (29, 14, 2) {real, imag} */,
  {32'hc0fa2e6d, 32'hc10707ee} /* (29, 14, 1) {real, imag} */,
  {32'hc0aa0964, 32'hc16009d4} /* (29, 14, 0) {real, imag} */,
  {32'hbf22fcb0, 32'h3fd95910} /* (29, 13, 31) {real, imag} */,
  {32'h416358bc, 32'hc0eed2cc} /* (29, 13, 30) {real, imag} */,
  {32'hc16aabeb, 32'h41635331} /* (29, 13, 29) {real, imag} */,
  {32'h405b3e8a, 32'hc00be55c} /* (29, 13, 28) {real, imag} */,
  {32'h4051b777, 32'h403b4199} /* (29, 13, 27) {real, imag} */,
  {32'h4187376e, 32'hc08685e3} /* (29, 13, 26) {real, imag} */,
  {32'hc065fabc, 32'hc10e6d62} /* (29, 13, 25) {real, imag} */,
  {32'h40b87803, 32'hc07f2c93} /* (29, 13, 24) {real, imag} */,
  {32'h4148dc6a, 32'h419cab74} /* (29, 13, 23) {real, imag} */,
  {32'hc08feb33, 32'hc133276c} /* (29, 13, 22) {real, imag} */,
  {32'h41698bfc, 32'h411ae316} /* (29, 13, 21) {real, imag} */,
  {32'hbfbdbbd4, 32'h4106436c} /* (29, 13, 20) {real, imag} */,
  {32'h405e8208, 32'hbec06b20} /* (29, 13, 19) {real, imag} */,
  {32'hc0f1bd1f, 32'hc0728fd4} /* (29, 13, 18) {real, imag} */,
  {32'hc080ecc7, 32'hc11a0e5c} /* (29, 13, 17) {real, imag} */,
  {32'hbfd0d4c0, 32'hc066795e} /* (29, 13, 16) {real, imag} */,
  {32'hbfb505dc, 32'h41a54efe} /* (29, 13, 15) {real, imag} */,
  {32'h41849638, 32'hc071d478} /* (29, 13, 14) {real, imag} */,
  {32'h40c973af, 32'hc0c4c7bb} /* (29, 13, 13) {real, imag} */,
  {32'h41169ef8, 32'hc1340c84} /* (29, 13, 12) {real, imag} */,
  {32'hc07d5ab4, 32'hc08848ca} /* (29, 13, 11) {real, imag} */,
  {32'hc100cf90, 32'h40a9573e} /* (29, 13, 10) {real, imag} */,
  {32'hc17e61ae, 32'hbffce973} /* (29, 13, 9) {real, imag} */,
  {32'hc0eba2e8, 32'h3f924400} /* (29, 13, 8) {real, imag} */,
  {32'h401b16a4, 32'hc0299531} /* (29, 13, 7) {real, imag} */,
  {32'h40867b7c, 32'h3fd1cc44} /* (29, 13, 6) {real, imag} */,
  {32'hc18caf56, 32'hc126147f} /* (29, 13, 5) {real, imag} */,
  {32'h412547c9, 32'h3ed9a290} /* (29, 13, 4) {real, imag} */,
  {32'h412cb908, 32'hc0de57a6} /* (29, 13, 3) {real, imag} */,
  {32'h3ed770fc, 32'hc18ba3cd} /* (29, 13, 2) {real, imag} */,
  {32'h40d4a2ee, 32'h4117d557} /* (29, 13, 1) {real, imag} */,
  {32'h41a12d44, 32'h41445c50} /* (29, 13, 0) {real, imag} */,
  {32'h40ecb2d6, 32'h41211ae9} /* (29, 12, 31) {real, imag} */,
  {32'h40cf02d0, 32'h4084ae80} /* (29, 12, 30) {real, imag} */,
  {32'hc09eff65, 32'h41841617} /* (29, 12, 29) {real, imag} */,
  {32'h41b97dd8, 32'hbf3fae98} /* (29, 12, 28) {real, imag} */,
  {32'h3fb7ef96, 32'hc12d2b92} /* (29, 12, 27) {real, imag} */,
  {32'h404dbab0, 32'h41096148} /* (29, 12, 26) {real, imag} */,
  {32'hc0f58c0c, 32'hc141bfd4} /* (29, 12, 25) {real, imag} */,
  {32'h402a7c00, 32'h4068fc05} /* (29, 12, 24) {real, imag} */,
  {32'hc18be8cd, 32'hbfd7e876} /* (29, 12, 23) {real, imag} */,
  {32'hc08abd26, 32'hc19835cc} /* (29, 12, 22) {real, imag} */,
  {32'hc1451336, 32'h4131647c} /* (29, 12, 21) {real, imag} */,
  {32'h405aa03d, 32'h40ec6b61} /* (29, 12, 20) {real, imag} */,
  {32'h3f22587f, 32'h40e58bcc} /* (29, 12, 19) {real, imag} */,
  {32'h40ff429a, 32'h40eea53f} /* (29, 12, 18) {real, imag} */,
  {32'hbff1b190, 32'hbfe90a0c} /* (29, 12, 17) {real, imag} */,
  {32'hc0a0e8e4, 32'h3ebc7b30} /* (29, 12, 16) {real, imag} */,
  {32'h409fb6de, 32'h40434418} /* (29, 12, 15) {real, imag} */,
  {32'hc107228e, 32'hc09da82e} /* (29, 12, 14) {real, imag} */,
  {32'h40b32ed5, 32'hc0f687fc} /* (29, 12, 13) {real, imag} */,
  {32'hc0913716, 32'h416658ad} /* (29, 12, 12) {real, imag} */,
  {32'h4121d2d3, 32'hc185c4bf} /* (29, 12, 11) {real, imag} */,
  {32'hc1548e53, 32'h40059a5c} /* (29, 12, 10) {real, imag} */,
  {32'h40999126, 32'hc00b8296} /* (29, 12, 9) {real, imag} */,
  {32'hc19d60be, 32'h3faf4ba0} /* (29, 12, 8) {real, imag} */,
  {32'hc12c6ea6, 32'hc136ffd2} /* (29, 12, 7) {real, imag} */,
  {32'h409ad192, 32'hbffc850e} /* (29, 12, 6) {real, imag} */,
  {32'h3eb310d8, 32'h41010fb9} /* (29, 12, 5) {real, imag} */,
  {32'hc046f93c, 32'hc13bc80d} /* (29, 12, 4) {real, imag} */,
  {32'h4001bb26, 32'h4099f5d0} /* (29, 12, 3) {real, imag} */,
  {32'hc1967eae, 32'hbf168e10} /* (29, 12, 2) {real, imag} */,
  {32'h40847005, 32'hc009a964} /* (29, 12, 1) {real, imag} */,
  {32'hc0856e92, 32'hc0affb60} /* (29, 12, 0) {real, imag} */,
  {32'hc0f1669e, 32'hc137be2a} /* (29, 11, 31) {real, imag} */,
  {32'h4081b80b, 32'h4155cd53} /* (29, 11, 30) {real, imag} */,
  {32'h41357124, 32'hc02d3ed4} /* (29, 11, 29) {real, imag} */,
  {32'h415fd46e, 32'h40378fbf} /* (29, 11, 28) {real, imag} */,
  {32'h400de658, 32'hc180de65} /* (29, 11, 27) {real, imag} */,
  {32'hc140c734, 32'h411f8e09} /* (29, 11, 26) {real, imag} */,
  {32'h41408d4c, 32'h40c57db5} /* (29, 11, 25) {real, imag} */,
  {32'hc1198ce8, 32'hc058c814} /* (29, 11, 24) {real, imag} */,
  {32'hc0bb9e5e, 32'h411154d4} /* (29, 11, 23) {real, imag} */,
  {32'hc1b02278, 32'h40d1fb2a} /* (29, 11, 22) {real, imag} */,
  {32'h41071699, 32'hc188a7f0} /* (29, 11, 21) {real, imag} */,
  {32'h41015a29, 32'hc0fcdc92} /* (29, 11, 20) {real, imag} */,
  {32'h4161e42e, 32'hbf168420} /* (29, 11, 19) {real, imag} */,
  {32'hc135e27a, 32'hc11b7e1e} /* (29, 11, 18) {real, imag} */,
  {32'h3f34fd70, 32'h40a68cac} /* (29, 11, 17) {real, imag} */,
  {32'hc0a74d4e, 32'hc047046c} /* (29, 11, 16) {real, imag} */,
  {32'hc18a0f4c, 32'h409d8042} /* (29, 11, 15) {real, imag} */,
  {32'hc0538ea9, 32'hc1810ee0} /* (29, 11, 14) {real, imag} */,
  {32'hc114815e, 32'hc0309f50} /* (29, 11, 13) {real, imag} */,
  {32'h40f09d21, 32'hc0e4a33d} /* (29, 11, 12) {real, imag} */,
  {32'hc0f9ada9, 32'hc00e350a} /* (29, 11, 11) {real, imag} */,
  {32'h418d3517, 32'hc035bba6} /* (29, 11, 10) {real, imag} */,
  {32'h41cd18fc, 32'h4022d232} /* (29, 11, 9) {real, imag} */,
  {32'h40ae3a98, 32'h412fe429} /* (29, 11, 8) {real, imag} */,
  {32'hbfb14d3e, 32'h40b2f829} /* (29, 11, 7) {real, imag} */,
  {32'hc16a89be, 32'h415f8912} /* (29, 11, 6) {real, imag} */,
  {32'hc110ef5f, 32'h418a923c} /* (29, 11, 5) {real, imag} */,
  {32'hc17e4fe0, 32'h418673a6} /* (29, 11, 4) {real, imag} */,
  {32'hc031742e, 32'h40a5b40a} /* (29, 11, 3) {real, imag} */,
  {32'hc08ca481, 32'h4201279d} /* (29, 11, 2) {real, imag} */,
  {32'hc02d1db6, 32'hc1e8f050} /* (29, 11, 1) {real, imag} */,
  {32'hc1c8c8d5, 32'hc1e190a6} /* (29, 11, 0) {real, imag} */,
  {32'h41893280, 32'h40e251be} /* (29, 10, 31) {real, imag} */,
  {32'h4088d53f, 32'hc10a0253} /* (29, 10, 30) {real, imag} */,
  {32'h411fd5c0, 32'h41431c44} /* (29, 10, 29) {real, imag} */,
  {32'h403d040a, 32'h3f4f1120} /* (29, 10, 28) {real, imag} */,
  {32'h4182ceb2, 32'hc1545c67} /* (29, 10, 27) {real, imag} */,
  {32'h408dd4ca, 32'hc161c73e} /* (29, 10, 26) {real, imag} */,
  {32'h410fb50b, 32'h41147ef8} /* (29, 10, 25) {real, imag} */,
  {32'hc04c0f8a, 32'hc1b1cc43} /* (29, 10, 24) {real, imag} */,
  {32'hc1749658, 32'h40b99fe2} /* (29, 10, 23) {real, imag} */,
  {32'h4006baee, 32'h41abb94a} /* (29, 10, 22) {real, imag} */,
  {32'h408d77a2, 32'hc0f7c95c} /* (29, 10, 21) {real, imag} */,
  {32'h4125c536, 32'hc1151ed2} /* (29, 10, 20) {real, imag} */,
  {32'h4100663a, 32'hc14d31a0} /* (29, 10, 19) {real, imag} */,
  {32'h400a3a04, 32'h40de0e08} /* (29, 10, 18) {real, imag} */,
  {32'h3eedba88, 32'h407e5fa2} /* (29, 10, 17) {real, imag} */,
  {32'hc14fa086, 32'h40d3c999} /* (29, 10, 16) {real, imag} */,
  {32'h4170d46d, 32'hc0dc259e} /* (29, 10, 15) {real, imag} */,
  {32'h41ac238a, 32'hbf06ee38} /* (29, 10, 14) {real, imag} */,
  {32'hc19a7738, 32'h40357cd4} /* (29, 10, 13) {real, imag} */,
  {32'h40ac7e6a, 32'h417c905a} /* (29, 10, 12) {real, imag} */,
  {32'h417b1dd4, 32'h4086643c} /* (29, 10, 11) {real, imag} */,
  {32'h40896bcc, 32'h4138ed01} /* (29, 10, 10) {real, imag} */,
  {32'hc10ad5a8, 32'h407ea94f} /* (29, 10, 9) {real, imag} */,
  {32'hc0d98cdb, 32'h410b345d} /* (29, 10, 8) {real, imag} */,
  {32'h414935dc, 32'hc1538068} /* (29, 10, 7) {real, imag} */,
  {32'h41165c5e, 32'hc14ad827} /* (29, 10, 6) {real, imag} */,
  {32'hc1242e18, 32'h400cda36} /* (29, 10, 5) {real, imag} */,
  {32'hc1a5fbab, 32'hc18ca5de} /* (29, 10, 4) {real, imag} */,
  {32'hc1a8222c, 32'hbf882e0e} /* (29, 10, 3) {real, imag} */,
  {32'h3ff663b8, 32'h406dcbda} /* (29, 10, 2) {real, imag} */,
  {32'h3f74b9b0, 32'hbffec1f8} /* (29, 10, 1) {real, imag} */,
  {32'hc1840ff1, 32'h40c2fdb9} /* (29, 10, 0) {real, imag} */,
  {32'hc21d4b78, 32'h412fedfd} /* (29, 9, 31) {real, imag} */,
  {32'h41f00e87, 32'hc07b6408} /* (29, 9, 30) {real, imag} */,
  {32'h4100e1f9, 32'hbe1a2040} /* (29, 9, 29) {real, imag} */,
  {32'hbf6141d8, 32'h41efc942} /* (29, 9, 28) {real, imag} */,
  {32'hc151f940, 32'h4094e59e} /* (29, 9, 27) {real, imag} */,
  {32'hc02a9e82, 32'h415dbb75} /* (29, 9, 26) {real, imag} */,
  {32'hc1392f02, 32'h405ce680} /* (29, 9, 25) {real, imag} */,
  {32'h4083e961, 32'hc10b2d18} /* (29, 9, 24) {real, imag} */,
  {32'hc0d53f06, 32'h4155ebef} /* (29, 9, 23) {real, imag} */,
  {32'hc1f04259, 32'hc13d588e} /* (29, 9, 22) {real, imag} */,
  {32'hc14f2d0e, 32'hc109a696} /* (29, 9, 21) {real, imag} */,
  {32'hc0d79ffe, 32'hc18e8cc6} /* (29, 9, 20) {real, imag} */,
  {32'h4153fefe, 32'h41ab96ae} /* (29, 9, 19) {real, imag} */,
  {32'h4149cf49, 32'h40ae3d66} /* (29, 9, 18) {real, imag} */,
  {32'hc10b350c, 32'hc107cac0} /* (29, 9, 17) {real, imag} */,
  {32'h415f7688, 32'hc0fac36d} /* (29, 9, 16) {real, imag} */,
  {32'hc06e75a7, 32'h40d9ecc3} /* (29, 9, 15) {real, imag} */,
  {32'hc0ed99bb, 32'h41885a56} /* (29, 9, 14) {real, imag} */,
  {32'hc15e9694, 32'h41854fae} /* (29, 9, 13) {real, imag} */,
  {32'h411cbcc0, 32'h412104bd} /* (29, 9, 12) {real, imag} */,
  {32'h3e3a46b0, 32'hc0da6d4f} /* (29, 9, 11) {real, imag} */,
  {32'hc1baa175, 32'h4056bba8} /* (29, 9, 10) {real, imag} */,
  {32'hc10b4b9e, 32'hbdad58c0} /* (29, 9, 9) {real, imag} */,
  {32'h41632176, 32'hc0e07702} /* (29, 9, 8) {real, imag} */,
  {32'hc0605c1a, 32'hc0fa94a6} /* (29, 9, 7) {real, imag} */,
  {32'h40ed125e, 32'hbfb22ba9} /* (29, 9, 6) {real, imag} */,
  {32'h409fd260, 32'h41cd0b14} /* (29, 9, 5) {real, imag} */,
  {32'h3fb6dd06, 32'hbfc9c147} /* (29, 9, 4) {real, imag} */,
  {32'hc148c264, 32'h403ee9ba} /* (29, 9, 3) {real, imag} */,
  {32'hc1c02127, 32'hc1834bcc} /* (29, 9, 2) {real, imag} */,
  {32'h41ce3aae, 32'hc02618c0} /* (29, 9, 1) {real, imag} */,
  {32'hc15b22aa, 32'hc1933602} /* (29, 9, 0) {real, imag} */,
  {32'hc273bd9a, 32'hc226fe51} /* (29, 8, 31) {real, imag} */,
  {32'h41d44fbc, 32'h419a93fd} /* (29, 8, 30) {real, imag} */,
  {32'hbfd55d70, 32'hc1bddbb4} /* (29, 8, 29) {real, imag} */,
  {32'h411dc24c, 32'hc0e2ce16} /* (29, 8, 28) {real, imag} */,
  {32'hc16bd34d, 32'hc0854d50} /* (29, 8, 27) {real, imag} */,
  {32'h41451a58, 32'hc101e3a0} /* (29, 8, 26) {real, imag} */,
  {32'hc12d3a13, 32'hc1b215bc} /* (29, 8, 25) {real, imag} */,
  {32'h3f940f90, 32'h3f9534b0} /* (29, 8, 24) {real, imag} */,
  {32'hc0e78150, 32'hc00e0fab} /* (29, 8, 23) {real, imag} */,
  {32'h41af30de, 32'hc1220684} /* (29, 8, 22) {real, imag} */,
  {32'h4178ce4c, 32'h41647cee} /* (29, 8, 21) {real, imag} */,
  {32'hc0fd21e6, 32'hc0e07c79} /* (29, 8, 20) {real, imag} */,
  {32'hc13528bb, 32'h40810c29} /* (29, 8, 19) {real, imag} */,
  {32'h415324bd, 32'hc15adac9} /* (29, 8, 18) {real, imag} */,
  {32'hbe16f480, 32'h40686fa6} /* (29, 8, 17) {real, imag} */,
  {32'h411d3ae3, 32'h40edb3e6} /* (29, 8, 16) {real, imag} */,
  {32'h41063393, 32'h3e4d4fc0} /* (29, 8, 15) {real, imag} */,
  {32'hbf552eb0, 32'hc102907d} /* (29, 8, 14) {real, imag} */,
  {32'h41bcf1e7, 32'h408f413a} /* (29, 8, 13) {real, imag} */,
  {32'hc0607c02, 32'h40eb9c1a} /* (29, 8, 12) {real, imag} */,
  {32'hbf0bec78, 32'h41d2b48e} /* (29, 8, 11) {real, imag} */,
  {32'h411fbc46, 32'hc12f67fa} /* (29, 8, 10) {real, imag} */,
  {32'hc119ed08, 32'hc0f5475e} /* (29, 8, 9) {real, imag} */,
  {32'h4073bfb0, 32'h40baa950} /* (29, 8, 8) {real, imag} */,
  {32'hc16f64fa, 32'h40140df7} /* (29, 8, 7) {real, imag} */,
  {32'hc13d9f33, 32'h416cfabc} /* (29, 8, 6) {real, imag} */,
  {32'h410896a8, 32'h4175af81} /* (29, 8, 5) {real, imag} */,
  {32'hc0be2ea7, 32'hc107af7c} /* (29, 8, 4) {real, imag} */,
  {32'h41d554d8, 32'h41a2e601} /* (29, 8, 3) {real, imag} */,
  {32'hc0aafe14, 32'hc163f56f} /* (29, 8, 2) {real, imag} */,
  {32'hc18c2148, 32'hc22ca212} /* (29, 8, 1) {real, imag} */,
  {32'hc1866be3, 32'hc0ecc587} /* (29, 8, 0) {real, imag} */,
  {32'hc067bc7e, 32'hc10ce8fa} /* (29, 7, 31) {real, imag} */,
  {32'hc1938f1c, 32'h41dc0515} /* (29, 7, 30) {real, imag} */,
  {32'hc122feaf, 32'h3fa7a23c} /* (29, 7, 29) {real, imag} */,
  {32'hc1a1fc78, 32'hc0b4d244} /* (29, 7, 28) {real, imag} */,
  {32'h41285846, 32'h41b0d7c9} /* (29, 7, 27) {real, imag} */,
  {32'hc0b9af4a, 32'h3d3e1700} /* (29, 7, 26) {real, imag} */,
  {32'hc17df12b, 32'h40daeb8b} /* (29, 7, 25) {real, imag} */,
  {32'hbf08042a, 32'hc0b8d04b} /* (29, 7, 24) {real, imag} */,
  {32'h3d7d6300, 32'hc12a06d7} /* (29, 7, 23) {real, imag} */,
  {32'hc0ceef20, 32'h41a8d10e} /* (29, 7, 22) {real, imag} */,
  {32'hc072c9fc, 32'h412a4c4f} /* (29, 7, 21) {real, imag} */,
  {32'h40fe2e4d, 32'h3f091f00} /* (29, 7, 20) {real, imag} */,
  {32'h41260a35, 32'h40befc9a} /* (29, 7, 19) {real, imag} */,
  {32'h4127c3a6, 32'h408110bc} /* (29, 7, 18) {real, imag} */,
  {32'hc1813f4c, 32'hc1264641} /* (29, 7, 17) {real, imag} */,
  {32'h403b379a, 32'hc106b1d8} /* (29, 7, 16) {real, imag} */,
  {32'hbeb7fe10, 32'hc017c0e0} /* (29, 7, 15) {real, imag} */,
  {32'hbfaad8a4, 32'hc0c4e83c} /* (29, 7, 14) {real, imag} */,
  {32'hc1684bb8, 32'h406cff98} /* (29, 7, 13) {real, imag} */,
  {32'h408b8dea, 32'hbfde3984} /* (29, 7, 12) {real, imag} */,
  {32'hc10b6491, 32'h41822dce} /* (29, 7, 11) {real, imag} */,
  {32'hc100e071, 32'hc064a56b} /* (29, 7, 10) {real, imag} */,
  {32'h4146f770, 32'h414e263c} /* (29, 7, 9) {real, imag} */,
  {32'hc0ad8f49, 32'hc054b929} /* (29, 7, 8) {real, imag} */,
  {32'hc0695e04, 32'hc12a0862} /* (29, 7, 7) {real, imag} */,
  {32'h41cd13f4, 32'hc167a1ca} /* (29, 7, 6) {real, imag} */,
  {32'h408c9a26, 32'hc1d92f99} /* (29, 7, 5) {real, imag} */,
  {32'h3f4acd60, 32'hc08a06cd} /* (29, 7, 4) {real, imag} */,
  {32'hc1bfa8c2, 32'hc136ea50} /* (29, 7, 3) {real, imag} */,
  {32'h41408744, 32'hc0f15334} /* (29, 7, 2) {real, imag} */,
  {32'h4237f53c, 32'h3fa91360} /* (29, 7, 1) {real, imag} */,
  {32'h421315c2, 32'hc055a24c} /* (29, 7, 0) {real, imag} */,
  {32'h415e14bc, 32'h41ca7d0e} /* (29, 6, 31) {real, imag} */,
  {32'h4180d86e, 32'h41a2ee15} /* (29, 6, 30) {real, imag} */,
  {32'h3dbbb3a0, 32'h3f86d348} /* (29, 6, 29) {real, imag} */,
  {32'hc0420a48, 32'hc1b2fc21} /* (29, 6, 28) {real, imag} */,
  {32'hc207fe74, 32'h406fb05f} /* (29, 6, 27) {real, imag} */,
  {32'hc13ce9f8, 32'hc065b973} /* (29, 6, 26) {real, imag} */,
  {32'h415d6bcc, 32'h41ef1faa} /* (29, 6, 25) {real, imag} */,
  {32'hc1146fa1, 32'h41dfc1da} /* (29, 6, 24) {real, imag} */,
  {32'h418e5da6, 32'hc0f2fce8} /* (29, 6, 23) {real, imag} */,
  {32'hc10d7024, 32'h40aee5ef} /* (29, 6, 22) {real, imag} */,
  {32'hc197e075, 32'hc11f4a16} /* (29, 6, 21) {real, imag} */,
  {32'hbfeaee8c, 32'hc0a95d83} /* (29, 6, 20) {real, imag} */,
  {32'h413a5d3a, 32'hc1c160c0} /* (29, 6, 19) {real, imag} */,
  {32'h41433878, 32'h40999570} /* (29, 6, 18) {real, imag} */,
  {32'hc103dbce, 32'h40e069c6} /* (29, 6, 17) {real, imag} */,
  {32'h3fa3ecf0, 32'h41007e58} /* (29, 6, 16) {real, imag} */,
  {32'hc13061fd, 32'hc10a2db6} /* (29, 6, 15) {real, imag} */,
  {32'hc1880b34, 32'h40e35262} /* (29, 6, 14) {real, imag} */,
  {32'h41592c34, 32'h40fc256f} /* (29, 6, 13) {real, imag} */,
  {32'h41600a5e, 32'h416b9e9c} /* (29, 6, 12) {real, imag} */,
  {32'h3fe8176c, 32'h41826d5e} /* (29, 6, 11) {real, imag} */,
  {32'h40c7ee34, 32'hc079e334} /* (29, 6, 10) {real, imag} */,
  {32'h408476ac, 32'h4080ba64} /* (29, 6, 9) {real, imag} */,
  {32'h3fea60de, 32'h406e0e0c} /* (29, 6, 8) {real, imag} */,
  {32'h41c3cc15, 32'h412f472b} /* (29, 6, 7) {real, imag} */,
  {32'hbe8aae40, 32'h4070b19c} /* (29, 6, 6) {real, imag} */,
  {32'h40f182c8, 32'h3ff41818} /* (29, 6, 5) {real, imag} */,
  {32'h41824f82, 32'hc0cbf979} /* (29, 6, 4) {real, imag} */,
  {32'h408fcf25, 32'hbdc405c0} /* (29, 6, 3) {real, imag} */,
  {32'hbba0a800, 32'hc025bc9c} /* (29, 6, 2) {real, imag} */,
  {32'hc1d80c40, 32'h415e2120} /* (29, 6, 1) {real, imag} */,
  {32'h411ef882, 32'h4138a253} /* (29, 6, 0) {real, imag} */,
  {32'hc2da22bc, 32'hc19b92e9} /* (29, 5, 31) {real, imag} */,
  {32'h40e5522e, 32'hc1d81c36} /* (29, 5, 30) {real, imag} */,
  {32'h41574e96, 32'hc1bddeb1} /* (29, 5, 29) {real, imag} */,
  {32'hc1ab6320, 32'h416612d7} /* (29, 5, 28) {real, imag} */,
  {32'h4214df07, 32'h41315bc9} /* (29, 5, 27) {real, imag} */,
  {32'h40b46253, 32'hc17f8d9c} /* (29, 5, 26) {real, imag} */,
  {32'hc19da539, 32'h4121be85} /* (29, 5, 25) {real, imag} */,
  {32'hc0d9e0a2, 32'h3e59dd10} /* (29, 5, 24) {real, imag} */,
  {32'hc0eb3758, 32'hc10f080e} /* (29, 5, 23) {real, imag} */,
  {32'h40693fec, 32'h41ce8117} /* (29, 5, 22) {real, imag} */,
  {32'h419ed5c1, 32'hc0407660} /* (29, 5, 21) {real, imag} */,
  {32'hc05a8138, 32'h40b65176} /* (29, 5, 20) {real, imag} */,
  {32'h40dbbbea, 32'h3ef22748} /* (29, 5, 19) {real, imag} */,
  {32'h405646e2, 32'h400d6d65} /* (29, 5, 18) {real, imag} */,
  {32'h40b5f004, 32'h409008ce} /* (29, 5, 17) {real, imag} */,
  {32'h403405a2, 32'hc0a23b46} /* (29, 5, 16) {real, imag} */,
  {32'hbfe742d0, 32'h409da836} /* (29, 5, 15) {real, imag} */,
  {32'h4006e269, 32'hc0a38b44} /* (29, 5, 14) {real, imag} */,
  {32'hc0b3532a, 32'hc06486fe} /* (29, 5, 13) {real, imag} */,
  {32'h4012dcda, 32'hbeab1660} /* (29, 5, 12) {real, imag} */,
  {32'h400a1da1, 32'hc0dddeef} /* (29, 5, 11) {real, imag} */,
  {32'hc186ab3e, 32'hc0d4db47} /* (29, 5, 10) {real, imag} */,
  {32'hc0112d60, 32'h3f93a558} /* (29, 5, 9) {real, imag} */,
  {32'h40d950e5, 32'h3f751580} /* (29, 5, 8) {real, imag} */,
  {32'h40aea345, 32'h40449fa8} /* (29, 5, 7) {real, imag} */,
  {32'hc0b21746, 32'hc13ccb46} /* (29, 5, 6) {real, imag} */,
  {32'hbf6208c0, 32'h4217000c} /* (29, 5, 5) {real, imag} */,
  {32'hc17e69bd, 32'hc1038b41} /* (29, 5, 4) {real, imag} */,
  {32'h40c611ae, 32'hc14938be} /* (29, 5, 3) {real, imag} */,
  {32'h42246168, 32'hbf14cae0} /* (29, 5, 2) {real, imag} */,
  {32'hc291ac68, 32'hc25e705c} /* (29, 5, 1) {real, imag} */,
  {32'hc279715a, 32'hc206368c} /* (29, 5, 0) {real, imag} */,
  {32'h42a757d7, 32'h429cd0ce} /* (29, 4, 31) {real, imag} */,
  {32'hc299d5af, 32'hc1fd2350} /* (29, 4, 30) {real, imag} */,
  {32'hc209de3a, 32'h426e653c} /* (29, 4, 29) {real, imag} */,
  {32'h420c07fc, 32'hc036ad34} /* (29, 4, 28) {real, imag} */,
  {32'hc26983fa, 32'h41a5379e} /* (29, 4, 27) {real, imag} */,
  {32'h40b52336, 32'h4145bc19} /* (29, 4, 26) {real, imag} */,
  {32'hc0eea136, 32'h3efc1050} /* (29, 4, 25) {real, imag} */,
  {32'hc1431488, 32'h3f5d0a88} /* (29, 4, 24) {real, imag} */,
  {32'hc1821620, 32'hc19be7ae} /* (29, 4, 23) {real, imag} */,
  {32'h402a60fc, 32'hc0b751f0} /* (29, 4, 22) {real, imag} */,
  {32'h3ff7d138, 32'hc0ded278} /* (29, 4, 21) {real, imag} */,
  {32'hc0896b6e, 32'hc1055abe} /* (29, 4, 20) {real, imag} */,
  {32'h4100ccfc, 32'hc1386b56} /* (29, 4, 19) {real, imag} */,
  {32'hc1bb638d, 32'hc0535941} /* (29, 4, 18) {real, imag} */,
  {32'h412dada3, 32'hbf72dfa8} /* (29, 4, 17) {real, imag} */,
  {32'hc0a28a79, 32'hbf975a39} /* (29, 4, 16) {real, imag} */,
  {32'hc1214475, 32'hbf01c6e8} /* (29, 4, 15) {real, imag} */,
  {32'hc09c403e, 32'h407cb684} /* (29, 4, 14) {real, imag} */,
  {32'h40b01119, 32'hc178d3d8} /* (29, 4, 13) {real, imag} */,
  {32'hc12d7468, 32'hc123988c} /* (29, 4, 12) {real, imag} */,
  {32'h4020e28b, 32'h416666ec} /* (29, 4, 11) {real, imag} */,
  {32'hbfe8f344, 32'h411e8616} /* (29, 4, 10) {real, imag} */,
  {32'h40c0acc6, 32'hc17ff297} /* (29, 4, 9) {real, imag} */,
  {32'hc11b468f, 32'hc13e9f39} /* (29, 4, 8) {real, imag} */,
  {32'h410d7a3c, 32'hc1388083} /* (29, 4, 7) {real, imag} */,
  {32'hc04db624, 32'h4147aaed} /* (29, 4, 6) {real, imag} */,
  {32'h3fa7d09a, 32'hc1d82390} /* (29, 4, 5) {real, imag} */,
  {32'h41cd952e, 32'h414ac78e} /* (29, 4, 4) {real, imag} */,
  {32'h40f6001b, 32'hc0b49028} /* (29, 4, 3) {real, imag} */,
  {32'hc212ba78, 32'hc27ea0c2} /* (29, 4, 2) {real, imag} */,
  {32'h43204205, 32'h428c80a3} /* (29, 4, 1) {real, imag} */,
  {32'h4253fc1a, 32'h42071e66} /* (29, 4, 0) {real, imag} */,
  {32'hc2f54d4c, 32'h429403bf} /* (29, 3, 31) {real, imag} */,
  {32'h4285dcc3, 32'hc29d31b6} /* (29, 3, 30) {real, imag} */,
  {32'h401a5a4c, 32'h417a681b} /* (29, 3, 29) {real, imag} */,
  {32'h417d76fd, 32'h41e46c6a} /* (29, 3, 28) {real, imag} */,
  {32'hc0bb6a7c, 32'hc21dc348} /* (29, 3, 27) {real, imag} */,
  {32'hc0b11c4a, 32'h41043564} /* (29, 3, 26) {real, imag} */,
  {32'hc1043f86, 32'h411607ae} /* (29, 3, 25) {real, imag} */,
  {32'hc14bbb9a, 32'hc1b5f5b2} /* (29, 3, 24) {real, imag} */,
  {32'h4112f84d, 32'h3fd7fa70} /* (29, 3, 23) {real, imag} */,
  {32'h40b7213a, 32'hbf4ccad8} /* (29, 3, 22) {real, imag} */,
  {32'hc1ef964a, 32'h3fb34a00} /* (29, 3, 21) {real, imag} */,
  {32'h40acb71a, 32'h41336d6a} /* (29, 3, 20) {real, imag} */,
  {32'hc1335c07, 32'h41061542} /* (29, 3, 19) {real, imag} */,
  {32'hc094c728, 32'hbd994f20} /* (29, 3, 18) {real, imag} */,
  {32'h40007b5c, 32'h40477155} /* (29, 3, 17) {real, imag} */,
  {32'hc039534a, 32'hc058d5d9} /* (29, 3, 16) {real, imag} */,
  {32'h40bcc4aa, 32'hc10420a1} /* (29, 3, 15) {real, imag} */,
  {32'h3fea1162, 32'h40b16024} /* (29, 3, 14) {real, imag} */,
  {32'h40d5aaa8, 32'hc0287e92} /* (29, 3, 13) {real, imag} */,
  {32'h4136dc91, 32'h41813486} /* (29, 3, 12) {real, imag} */,
  {32'hbfd2d808, 32'hbf689cf0} /* (29, 3, 11) {real, imag} */,
  {32'h406a5ab8, 32'hc0c01e90} /* (29, 3, 10) {real, imag} */,
  {32'h40dc5bac, 32'hbf83dc8a} /* (29, 3, 9) {real, imag} */,
  {32'hc08a70d2, 32'hbf0cb730} /* (29, 3, 8) {real, imag} */,
  {32'h41da5811, 32'h409c433c} /* (29, 3, 7) {real, imag} */,
  {32'hc1c935f0, 32'hc1a53013} /* (29, 3, 6) {real, imag} */,
  {32'hbed47b00, 32'h4082952c} /* (29, 3, 5) {real, imag} */,
  {32'hc142324c, 32'h41fb9454} /* (29, 3, 4) {real, imag} */,
  {32'h41803b05, 32'h416188aa} /* (29, 3, 3) {real, imag} */,
  {32'hc045ee4c, 32'hc29b7f9e} /* (29, 3, 2) {real, imag} */,
  {32'h428333fa, 32'h42f13afc} /* (29, 3, 1) {real, imag} */,
  {32'h41039992, 32'hbf912a38} /* (29, 3, 0) {real, imag} */,
  {32'hc435e489, 32'hc1c80b8a} /* (29, 2, 31) {real, imag} */,
  {32'h43ccf7ac, 32'hc3103bce} /* (29, 2, 30) {real, imag} */,
  {32'h40fbede4, 32'hc1550b5a} /* (29, 2, 29) {real, imag} */,
  {32'hc20df8e2, 32'h429fef6e} /* (29, 2, 28) {real, imag} */,
  {32'h424bd6e6, 32'hc1cd27c1} /* (29, 2, 27) {real, imag} */,
  {32'h410ebeba, 32'h411c4232} /* (29, 2, 26) {real, imag} */,
  {32'hc027b968, 32'h41f3f13f} /* (29, 2, 25) {real, imag} */,
  {32'h4219f172, 32'hc1ab32ee} /* (29, 2, 24) {real, imag} */,
  {32'hc0edcd34, 32'hc03a5248} /* (29, 2, 23) {real, imag} */,
  {32'h4122f6ad, 32'h419941f3} /* (29, 2, 22) {real, imag} */,
  {32'h413accce, 32'hc132d43e} /* (29, 2, 21) {real, imag} */,
  {32'hc18e3ab9, 32'h4161cc11} /* (29, 2, 20) {real, imag} */,
  {32'hc03966c4, 32'hc1368f86} /* (29, 2, 19) {real, imag} */,
  {32'h4107b257, 32'hbe742080} /* (29, 2, 18) {real, imag} */,
  {32'hbf9e136e, 32'h40d03fb5} /* (29, 2, 17) {real, imag} */,
  {32'h40d61933, 32'hc0d684e9} /* (29, 2, 16) {real, imag} */,
  {32'hc09ed663, 32'hc0e248c8} /* (29, 2, 15) {real, imag} */,
  {32'h4071c924, 32'h40d8a92f} /* (29, 2, 14) {real, imag} */,
  {32'h4097fee6, 32'hc17c5bf3} /* (29, 2, 13) {real, imag} */,
  {32'h3fe7d760, 32'h412baf6c} /* (29, 2, 12) {real, imag} */,
  {32'h41528e85, 32'h4126298e} /* (29, 2, 11) {real, imag} */,
  {32'hc1801f2f, 32'h418c7bd0} /* (29, 2, 10) {real, imag} */,
  {32'h41698acd, 32'h40a2cc1f} /* (29, 2, 9) {real, imag} */,
  {32'hc0ad2634, 32'h410bf4a1} /* (29, 2, 8) {real, imag} */,
  {32'h4154c7f0, 32'hc11d8360} /* (29, 2, 7) {real, imag} */,
  {32'h3f8e2640, 32'h41725786} /* (29, 2, 6) {real, imag} */,
  {32'h421b7092, 32'h413f1c97} /* (29, 2, 5) {real, imag} */,
  {32'hc263036c, 32'hc175a0d6} /* (29, 2, 4) {real, imag} */,
  {32'hc1bd1c38, 32'hc1a3899d} /* (29, 2, 3) {real, imag} */,
  {32'h4388fdd2, 32'hc29f5e9c} /* (29, 2, 2) {real, imag} */,
  {32'hc3e4ca54, 32'h4303ee06} /* (29, 2, 1) {real, imag} */,
  {32'hc3be597d, 32'hc26894af} /* (29, 2, 0) {real, imag} */,
  {32'h4420b567, 32'hc34716e8} /* (29, 1, 31) {real, imag} */,
  {32'hc38976e2, 32'h40729c18} /* (29, 1, 30) {real, imag} */,
  {32'hc0b4d694, 32'hc186f9a0} /* (29, 1, 29) {real, imag} */,
  {32'h4245a46a, 32'h42800d1f} /* (29, 1, 28) {real, imag} */,
  {32'hc2e9e5bc, 32'h4234c304} /* (29, 1, 27) {real, imag} */,
  {32'hc1966796, 32'h407de660} /* (29, 1, 26) {real, imag} */,
  {32'h3f6d8b00, 32'hc23a28f8} /* (29, 1, 25) {real, imag} */,
  {32'h4060bee0, 32'h41c062bd} /* (29, 1, 24) {real, imag} */,
  {32'h409f221c, 32'hc03c9a68} /* (29, 1, 23) {real, imag} */,
  {32'h4135fd69, 32'hc0eb686f} /* (29, 1, 22) {real, imag} */,
  {32'hc09a43f6, 32'h41b2db66} /* (29, 1, 21) {real, imag} */,
  {32'hc0b5c04e, 32'h40b27d7b} /* (29, 1, 20) {real, imag} */,
  {32'h413f87fc, 32'h4039c239} /* (29, 1, 19) {real, imag} */,
  {32'hc18de0e5, 32'h40b41b40} /* (29, 1, 18) {real, imag} */,
  {32'h3fa3cfd8, 32'h3f8d225c} /* (29, 1, 17) {real, imag} */,
  {32'hc0ea626f, 32'hc110d995} /* (29, 1, 16) {real, imag} */,
  {32'h4068306e, 32'h40309a0e} /* (29, 1, 15) {real, imag} */,
  {32'h410d20a3, 32'hc13c3204} /* (29, 1, 14) {real, imag} */,
  {32'h40637cec, 32'hc0f46b4a} /* (29, 1, 13) {real, imag} */,
  {32'h40a18aee, 32'h409d66f0} /* (29, 1, 12) {real, imag} */,
  {32'h40a2a97c, 32'hc177e64d} /* (29, 1, 11) {real, imag} */,
  {32'hc1d014ec, 32'h3f6fafe0} /* (29, 1, 10) {real, imag} */,
  {32'hc12c2cae, 32'h40d8be7f} /* (29, 1, 9) {real, imag} */,
  {32'hc0d3e927, 32'hc1e2fc62} /* (29, 1, 8) {real, imag} */,
  {32'hc1303fd2, 32'h4100b5bc} /* (29, 1, 7) {real, imag} */,
  {32'hc123bcfc, 32'h4155cc87} /* (29, 1, 6) {real, imag} */,
  {32'hc28d7d19, 32'hc2062d79} /* (29, 1, 5) {real, imag} */,
  {32'h423cf852, 32'h420e7a8a} /* (29, 1, 4) {real, imag} */,
  {32'hc1c6232c, 32'h42449552} /* (29, 1, 3) {real, imag} */,
  {32'hc3c0cccc, 32'hc3e3363a} /* (29, 1, 2) {real, imag} */,
  {32'h446981a4, 32'h43c56bdc} /* (29, 1, 1) {real, imag} */,
  {32'h440e6846, 32'h42b994f4} /* (29, 1, 0) {real, imag} */,
  {32'h438603c2, 32'hc38835c3} /* (29, 0, 31) {real, imag} */,
  {32'hc2c32d0d, 32'h43773eef} /* (29, 0, 30) {real, imag} */,
  {32'hc215baf1, 32'hc18c93e8} /* (29, 0, 29) {real, imag} */,
  {32'h4093818c, 32'h41e15320} /* (29, 0, 28) {real, imag} */,
  {32'hc266f9e6, 32'hc1ea217b} /* (29, 0, 27) {real, imag} */,
  {32'hc0c1a960, 32'hc19ed9b6} /* (29, 0, 26) {real, imag} */,
  {32'hc18267a2, 32'hc2064156} /* (29, 0, 25) {real, imag} */,
  {32'h40bb7ca4, 32'h419cadc1} /* (29, 0, 24) {real, imag} */,
  {32'h3f747f40, 32'h417c8a75} /* (29, 0, 23) {real, imag} */,
  {32'h4161b7ee, 32'h410fcec0} /* (29, 0, 22) {real, imag} */,
  {32'h40b1375c, 32'h412b3296} /* (29, 0, 21) {real, imag} */,
  {32'hbf6ff390, 32'hc0a7ebdb} /* (29, 0, 20) {real, imag} */,
  {32'hc0a7f065, 32'hc104b613} /* (29, 0, 19) {real, imag} */,
  {32'h3fbd8f28, 32'h407e152c} /* (29, 0, 18) {real, imag} */,
  {32'h40a7850e, 32'hc14ebffe} /* (29, 0, 17) {real, imag} */,
  {32'hbf52eae4, 32'h00000000} /* (29, 0, 16) {real, imag} */,
  {32'h40a7850e, 32'h414ebffe} /* (29, 0, 15) {real, imag} */,
  {32'h3fbd8f28, 32'hc07e152c} /* (29, 0, 14) {real, imag} */,
  {32'hc0a7f065, 32'h4104b613} /* (29, 0, 13) {real, imag} */,
  {32'hbf6ff390, 32'h40a7ebdb} /* (29, 0, 12) {real, imag} */,
  {32'h40b1375c, 32'hc12b3296} /* (29, 0, 11) {real, imag} */,
  {32'h4161b7ee, 32'hc10fcec0} /* (29, 0, 10) {real, imag} */,
  {32'h3f747f40, 32'hc17c8a75} /* (29, 0, 9) {real, imag} */,
  {32'h40bb7ca4, 32'hc19cadc1} /* (29, 0, 8) {real, imag} */,
  {32'hc18267a2, 32'h42064156} /* (29, 0, 7) {real, imag} */,
  {32'hc0c1a960, 32'h419ed9b6} /* (29, 0, 6) {real, imag} */,
  {32'hc266f9e6, 32'h41ea217b} /* (29, 0, 5) {real, imag} */,
  {32'h4093818c, 32'hc1e15320} /* (29, 0, 4) {real, imag} */,
  {32'hc215baf1, 32'h418c93e8} /* (29, 0, 3) {real, imag} */,
  {32'hc2c32d0d, 32'hc3773eef} /* (29, 0, 2) {real, imag} */,
  {32'h438603c2, 32'h438835c3} /* (29, 0, 1) {real, imag} */,
  {32'h423d556c, 32'h00000000} /* (29, 0, 0) {real, imag} */,
  {32'h444dec3a, 32'hc3afa2b3} /* (28, 31, 31) {real, imag} */,
  {32'hc3bd1793, 32'h43c9ec43} /* (28, 31, 30) {real, imag} */,
  {32'hc282ece5, 32'h3f0ac020} /* (28, 31, 29) {real, imag} */,
  {32'h4239a870, 32'hc109da7e} /* (28, 31, 28) {real, imag} */,
  {32'hc280a52d, 32'h41edc7c4} /* (28, 31, 27) {real, imag} */,
  {32'hbf6f8a40, 32'h413a8ec6} /* (28, 31, 26) {real, imag} */,
  {32'hc17cf2b4, 32'hc1c4bdc6} /* (28, 31, 25) {real, imag} */,
  {32'h3f91aba8, 32'h41bc0a80} /* (28, 31, 24) {real, imag} */,
  {32'hc03a5e10, 32'h411e695c} /* (28, 31, 23) {real, imag} */,
  {32'hc128a226, 32'hc01808ef} /* (28, 31, 22) {real, imag} */,
  {32'hc11b96d6, 32'hc0fef79c} /* (28, 31, 21) {real, imag} */,
  {32'h409ef4c2, 32'h40853a7b} /* (28, 31, 20) {real, imag} */,
  {32'hbf3e7d64, 32'hc10294c1} /* (28, 31, 19) {real, imag} */,
  {32'h415c89a0, 32'h41a9389a} /* (28, 31, 18) {real, imag} */,
  {32'h40921178, 32'hc1250ee0} /* (28, 31, 17) {real, imag} */,
  {32'h40165326, 32'h40aed598} /* (28, 31, 16) {real, imag} */,
  {32'h3fea361c, 32'hc0bc4fa0} /* (28, 31, 15) {real, imag} */,
  {32'h40434f80, 32'hc040008a} /* (28, 31, 14) {real, imag} */,
  {32'hc1221359, 32'hbe85bf20} /* (28, 31, 13) {real, imag} */,
  {32'h400e97fe, 32'h409e0274} /* (28, 31, 12) {real, imag} */,
  {32'hc16114bc, 32'hc0183bde} /* (28, 31, 11) {real, imag} */,
  {32'hc19a26a2, 32'hc1375566} /* (28, 31, 10) {real, imag} */,
  {32'h3cd21e00, 32'hc13aa354} /* (28, 31, 9) {real, imag} */,
  {32'hc17df928, 32'hc0f519ed} /* (28, 31, 8) {real, imag} */,
  {32'hbf9710c0, 32'h41895d26} /* (28, 31, 7) {real, imag} */,
  {32'hc185e7f1, 32'hc041ae04} /* (28, 31, 6) {real, imag} */,
  {32'hc2dfa512, 32'hc20113ad} /* (28, 31, 5) {real, imag} */,
  {32'h42426a2e, 32'hc2184bf4} /* (28, 31, 4) {real, imag} */,
  {32'h4097c6c0, 32'hc1207c5e} /* (28, 31, 3) {real, imag} */,
  {32'hc3836f90, 32'hc21e4a7b} /* (28, 31, 2) {real, imag} */,
  {32'h440cc812, 32'h433e7672} /* (28, 31, 1) {real, imag} */,
  {32'h43dcc76e, 32'hc2721544} /* (28, 31, 0) {real, imag} */,
  {32'hc3c1e4c5, 32'hc2ca20c0} /* (28, 30, 31) {real, imag} */,
  {32'h4397c4b4, 32'h42f7ff4a} /* (28, 30, 30) {real, imag} */,
  {32'hc18954e4, 32'h3fe781ec} /* (28, 30, 29) {real, imag} */,
  {32'hc2b3813b, 32'h4209fa5c} /* (28, 30, 28) {real, imag} */,
  {32'h4232b837, 32'hc1db6217} /* (28, 30, 27) {real, imag} */,
  {32'hc077b184, 32'h4031178c} /* (28, 30, 26) {real, imag} */,
  {32'hc137df7c, 32'h40e00a9f} /* (28, 30, 25) {real, imag} */,
  {32'h41b9549f, 32'hc1abbf56} /* (28, 30, 24) {real, imag} */,
  {32'h40dd10dc, 32'hc1b51a8e} /* (28, 30, 23) {real, imag} */,
  {32'hc179d68c, 32'h40d814a0} /* (28, 30, 22) {real, imag} */,
  {32'h3f5f00b8, 32'hc0c0afd6} /* (28, 30, 21) {real, imag} */,
  {32'hc1190331, 32'h40bd0ec8} /* (28, 30, 20) {real, imag} */,
  {32'hc07cbe84, 32'hc0c38fe1} /* (28, 30, 19) {real, imag} */,
  {32'h3fd3b17e, 32'hc14b86f1} /* (28, 30, 18) {real, imag} */,
  {32'hc0ae6e97, 32'hc0f86131} /* (28, 30, 17) {real, imag} */,
  {32'h4102a39e, 32'h4073909e} /* (28, 30, 16) {real, imag} */,
  {32'hc0a2ff02, 32'hc177f5b3} /* (28, 30, 15) {real, imag} */,
  {32'h4110b6a0, 32'h4163d349} /* (28, 30, 14) {real, imag} */,
  {32'hc0dd4be1, 32'hc1187722} /* (28, 30, 13) {real, imag} */,
  {32'h40bfd038, 32'h40f62b38} /* (28, 30, 12) {real, imag} */,
  {32'h3e913890, 32'h41f6fb7c} /* (28, 30, 11) {real, imag} */,
  {32'h41b84a46, 32'hc035454a} /* (28, 30, 10) {real, imag} */,
  {32'h408152ed, 32'h40e68edf} /* (28, 30, 9) {real, imag} */,
  {32'h4099aa95, 32'h42248af4} /* (28, 30, 8) {real, imag} */,
  {32'hbfb658fa, 32'hc22c00c3} /* (28, 30, 7) {real, imag} */,
  {32'h41b1fa1a, 32'hc1bfc7c6} /* (28, 30, 6) {real, imag} */,
  {32'h41d91d94, 32'h41e88b18} /* (28, 30, 5) {real, imag} */,
  {32'hc1c85007, 32'hc2aefa3a} /* (28, 30, 4) {real, imag} */,
  {32'hc18fec69, 32'h40f64a62} /* (28, 30, 3) {real, imag} */,
  {32'h43c5513e, 32'h431b8fb2} /* (28, 30, 2) {real, imag} */,
  {32'hc425e041, 32'hc1d1e393} /* (28, 30, 1) {real, imag} */,
  {32'hc3af5eb5, 32'h42999eaa} /* (28, 30, 0) {real, imag} */,
  {32'h4293bb0d, 32'hc3198610} /* (28, 29, 31) {real, imag} */,
  {32'hc17b7dbb, 32'h42c77516} /* (28, 29, 30) {real, imag} */,
  {32'h41e276c6, 32'hc180af85} /* (28, 29, 29) {real, imag} */,
  {32'hc004ecfc, 32'hc22cba7a} /* (28, 29, 28) {real, imag} */,
  {32'h41d510a9, 32'h405698e0} /* (28, 29, 27) {real, imag} */,
  {32'hc256890a, 32'h41a326ad} /* (28, 29, 26) {real, imag} */,
  {32'h418c29a3, 32'hc1054129} /* (28, 29, 25) {real, imag} */,
  {32'h400e7b46, 32'h40de8a86} /* (28, 29, 24) {real, imag} */,
  {32'hc09ac983, 32'hc16a7ee3} /* (28, 29, 23) {real, imag} */,
  {32'hc05abf1e, 32'hc0bb725c} /* (28, 29, 22) {real, imag} */,
  {32'h4157585b, 32'h41786ded} /* (28, 29, 21) {real, imag} */,
  {32'hc0d2c720, 32'h4183d950} /* (28, 29, 20) {real, imag} */,
  {32'hc16eccb0, 32'h41a2567f} /* (28, 29, 19) {real, imag} */,
  {32'hc08e4213, 32'h40121e58} /* (28, 29, 18) {real, imag} */,
  {32'h40e1b17c, 32'hbfc854e0} /* (28, 29, 17) {real, imag} */,
  {32'hc10146e2, 32'hbea6fa20} /* (28, 29, 16) {real, imag} */,
  {32'hc0ac6ec9, 32'h411f7e50} /* (28, 29, 15) {real, imag} */,
  {32'h40706cdc, 32'h413feffc} /* (28, 29, 14) {real, imag} */,
  {32'hc0f32a1b, 32'h40b2d14f} /* (28, 29, 13) {real, imag} */,
  {32'h415013f8, 32'h3fea8bca} /* (28, 29, 12) {real, imag} */,
  {32'hc19f03d1, 32'h3ef5abc0} /* (28, 29, 11) {real, imag} */,
  {32'h41f2ea15, 32'hc2077ad3} /* (28, 29, 10) {real, imag} */,
  {32'h410de770, 32'hc182c896} /* (28, 29, 9) {real, imag} */,
  {32'hc07943ea, 32'h41e9089a} /* (28, 29, 8) {real, imag} */,
  {32'hc17a7386, 32'hc1516e46} /* (28, 29, 7) {real, imag} */,
  {32'h4189f571, 32'h400f7f58} /* (28, 29, 6) {real, imag} */,
  {32'hc1283e50, 32'h41e9021b} /* (28, 29, 5) {real, imag} */,
  {32'h413df34d, 32'hc1ce12ce} /* (28, 29, 4) {real, imag} */,
  {32'hc1a15212, 32'hc0ec96c6} /* (28, 29, 3) {real, imag} */,
  {32'h4295b366, 32'h42bf95c8} /* (28, 29, 2) {real, imag} */,
  {32'hc3130f7f, 32'hc222f434} /* (28, 29, 1) {real, imag} */,
  {32'h41afc724, 32'h41837278} /* (28, 29, 0) {real, imag} */,
  {32'h42e49c41, 32'hc298f1ba} /* (28, 28, 31) {real, imag} */,
  {32'hc267b92e, 32'h42971cfb} /* (28, 28, 30) {real, imag} */,
  {32'h41caaf5d, 32'h42067e75} /* (28, 28, 29) {real, imag} */,
  {32'h423cd1c2, 32'h41d339ac} /* (28, 28, 28) {real, imag} */,
  {32'h40d19af8, 32'h412c549a} /* (28, 28, 27) {real, imag} */,
  {32'hbfbf92e0, 32'hc1ab8bc5} /* (28, 28, 26) {real, imag} */,
  {32'hc189befe, 32'hc0107e14} /* (28, 28, 25) {real, imag} */,
  {32'h3fd705cf, 32'h41042c3c} /* (28, 28, 24) {real, imag} */,
  {32'hc17840ee, 32'h412b2690} /* (28, 28, 23) {real, imag} */,
  {32'hc004ea30, 32'hc0824f41} /* (28, 28, 22) {real, imag} */,
  {32'h405bd804, 32'hc14f20ad} /* (28, 28, 21) {real, imag} */,
  {32'h40821d9c, 32'h419e1e44} /* (28, 28, 20) {real, imag} */,
  {32'h406eec6e, 32'hc0ca7927} /* (28, 28, 19) {real, imag} */,
  {32'hc0bd3b40, 32'hc01d4bc6} /* (28, 28, 18) {real, imag} */,
  {32'hc1214080, 32'hc123fe6d} /* (28, 28, 17) {real, imag} */,
  {32'h4032c1a2, 32'h402b470d} /* (28, 28, 16) {real, imag} */,
  {32'hc03bc62e, 32'hc06235a0} /* (28, 28, 15) {real, imag} */,
  {32'h3f28abe8, 32'hc0889076} /* (28, 28, 14) {real, imag} */,
  {32'hbf7f2968, 32'h400e6de5} /* (28, 28, 13) {real, imag} */,
  {32'h41bb9cca, 32'h413c2635} /* (28, 28, 12) {real, imag} */,
  {32'hc1a36ae0, 32'hc0cdaa93} /* (28, 28, 11) {real, imag} */,
  {32'hc10ad9fd, 32'hc0941e22} /* (28, 28, 10) {real, imag} */,
  {32'hc17eac1b, 32'hc0a930be} /* (28, 28, 9) {real, imag} */,
  {32'hc14a3c29, 32'hc01d77fb} /* (28, 28, 8) {real, imag} */,
  {32'h410cca1c, 32'h412b05ac} /* (28, 28, 7) {real, imag} */,
  {32'h4182e4c3, 32'hc174cc02} /* (28, 28, 6) {real, imag} */,
  {32'hc067cb7f, 32'hc0a72a54} /* (28, 28, 5) {real, imag} */,
  {32'h42013465, 32'h4114d7c5} /* (28, 28, 4) {real, imag} */,
  {32'h40be0f14, 32'h401291f4} /* (28, 28, 3) {real, imag} */,
  {32'hc2885c64, 32'h423a225d} /* (28, 28, 2) {real, imag} */,
  {32'h4282ba56, 32'hc28cc1ba} /* (28, 28, 1) {real, imag} */,
  {32'h420b550a, 32'hc24f361d} /* (28, 28, 0) {real, imag} */,
  {32'hc2942d54, 32'h425087b0} /* (28, 27, 31) {real, imag} */,
  {32'h41dd4471, 32'h41d94585} /* (28, 27, 30) {real, imag} */,
  {32'hc1386856, 32'h41a153dc} /* (28, 27, 29) {real, imag} */,
  {32'h405eccb8, 32'hc1a1b553} /* (28, 27, 28) {real, imag} */,
  {32'h41a1eb24, 32'hc1ce45cd} /* (28, 27, 27) {real, imag} */,
  {32'hc03a380e, 32'hc01d063c} /* (28, 27, 26) {real, imag} */,
  {32'h3fb59c66, 32'hc11f0d35} /* (28, 27, 25) {real, imag} */,
  {32'h3ea79cbc, 32'hc1382bf8} /* (28, 27, 24) {real, imag} */,
  {32'h41147aa6, 32'h4180c0eb} /* (28, 27, 23) {real, imag} */,
  {32'hc0dccc51, 32'h416532ad} /* (28, 27, 22) {real, imag} */,
  {32'hc06c5adc, 32'hc0e8cee0} /* (28, 27, 21) {real, imag} */,
  {32'h40f5ef3b, 32'h40dd6a0a} /* (28, 27, 20) {real, imag} */,
  {32'hc009a5ca, 32'h402fa0cc} /* (28, 27, 19) {real, imag} */,
  {32'hc0751552, 32'hc08ff4c6} /* (28, 27, 18) {real, imag} */,
  {32'hc0185527, 32'hc10e20b4} /* (28, 27, 17) {real, imag} */,
  {32'hbfe690c3, 32'h40b02633} /* (28, 27, 16) {real, imag} */,
  {32'hbf9b95e8, 32'h41831d68} /* (28, 27, 15) {real, imag} */,
  {32'hbffada94, 32'hc118b7c9} /* (28, 27, 14) {real, imag} */,
  {32'hc1169420, 32'hbfdc67a0} /* (28, 27, 13) {real, imag} */,
  {32'h3eaa8f78, 32'h3fc27362} /* (28, 27, 12) {real, imag} */,
  {32'h412e30f6, 32'h414c6f27} /* (28, 27, 11) {real, imag} */,
  {32'h4111e984, 32'hbfecf340} /* (28, 27, 10) {real, imag} */,
  {32'h4104279e, 32'hc0b016d9} /* (28, 27, 9) {real, imag} */,
  {32'h40125730, 32'h4039732f} /* (28, 27, 8) {real, imag} */,
  {32'h4165f15d, 32'hc1a7feae} /* (28, 27, 7) {real, imag} */,
  {32'h414ba2aa, 32'h41a832d4} /* (28, 27, 6) {real, imag} */,
  {32'h4214909c, 32'hc0dd58af} /* (28, 27, 5) {real, imag} */,
  {32'hc19e8c5a, 32'hc088a5c8} /* (28, 27, 4) {real, imag} */,
  {32'h40936b43, 32'h41c181aa} /* (28, 27, 3) {real, imag} */,
  {32'h4185815e, 32'h4107527e} /* (28, 27, 2) {real, imag} */,
  {32'hc2d5b67a, 32'h41bb7554} /* (28, 27, 1) {real, imag} */,
  {32'hc2736a56, 32'h421e2570} /* (28, 27, 0) {real, imag} */,
  {32'hc18b3c59, 32'h4121aa63} /* (28, 26, 31) {real, imag} */,
  {32'h40ca8dbc, 32'h3e851f08} /* (28, 26, 30) {real, imag} */,
  {32'h41127e10, 32'hc0da764b} /* (28, 26, 29) {real, imag} */,
  {32'h40e370ce, 32'hc03416b8} /* (28, 26, 28) {real, imag} */,
  {32'hc08edf2f, 32'h3d7837c0} /* (28, 26, 27) {real, imag} */,
  {32'hc128d14f, 32'hc131d618} /* (28, 26, 26) {real, imag} */,
  {32'h41c33aa0, 32'hc183f672} /* (28, 26, 25) {real, imag} */,
  {32'hbfdaa980, 32'h419d89ba} /* (28, 26, 24) {real, imag} */,
  {32'h412d0edc, 32'h4151388c} /* (28, 26, 23) {real, imag} */,
  {32'hc17e4aae, 32'hc1443ff2} /* (28, 26, 22) {real, imag} */,
  {32'h41864051, 32'h3fd48410} /* (28, 26, 21) {real, imag} */,
  {32'h40b9fe10, 32'h403d548c} /* (28, 26, 20) {real, imag} */,
  {32'hc07cedd8, 32'hc1660a54} /* (28, 26, 19) {real, imag} */,
  {32'hc03b76bc, 32'h406bca14} /* (28, 26, 18) {real, imag} */,
  {32'h4050d53f, 32'hc0a819f4} /* (28, 26, 17) {real, imag} */,
  {32'hc00b5341, 32'h4168dd12} /* (28, 26, 16) {real, imag} */,
  {32'h40fe5a48, 32'hc05d92d4} /* (28, 26, 15) {real, imag} */,
  {32'hc1144c0e, 32'hbfe2ea7a} /* (28, 26, 14) {real, imag} */,
  {32'h408e56cb, 32'h413d70b8} /* (28, 26, 13) {real, imag} */,
  {32'h4124a72c, 32'hc048d146} /* (28, 26, 12) {real, imag} */,
  {32'h3eae24d0, 32'h40744f74} /* (28, 26, 11) {real, imag} */,
  {32'h405d1eb2, 32'hc11a2f64} /* (28, 26, 10) {real, imag} */,
  {32'h3fd4e3c4, 32'h40595322} /* (28, 26, 9) {real, imag} */,
  {32'h40d88c08, 32'hc1aba1e5} /* (28, 26, 8) {real, imag} */,
  {32'h40d3b6f0, 32'hc17d03bc} /* (28, 26, 7) {real, imag} */,
  {32'h412f2d98, 32'h3ff7fc68} /* (28, 26, 6) {real, imag} */,
  {32'hc1b11803, 32'h40d403c1} /* (28, 26, 5) {real, imag} */,
  {32'hc0928b16, 32'h414eb5da} /* (28, 26, 4) {real, imag} */,
  {32'h413c8296, 32'hc125708d} /* (28, 26, 3) {real, imag} */,
  {32'h41a44c66, 32'hc1a62a9c} /* (28, 26, 2) {real, imag} */,
  {32'hc1a51b2e, 32'h3f0f16f0} /* (28, 26, 1) {real, imag} */,
  {32'hc0241964, 32'hc163cbaa} /* (28, 26, 0) {real, imag} */,
  {32'h41f54ef2, 32'hc123ccd3} /* (28, 25, 31) {real, imag} */,
  {32'hc14c56b0, 32'hc0ef60a3} /* (28, 25, 30) {real, imag} */,
  {32'hc18ea72a, 32'hc184f07a} /* (28, 25, 29) {real, imag} */,
  {32'hc06310c4, 32'hc104a790} /* (28, 25, 28) {real, imag} */,
  {32'h40e3469c, 32'h3f9adb18} /* (28, 25, 27) {real, imag} */,
  {32'hc0ef16e4, 32'h4045746b} /* (28, 25, 26) {real, imag} */,
  {32'h416c5cd6, 32'hc135bfe3} /* (28, 25, 25) {real, imag} */,
  {32'hc115c0fa, 32'h418f20e6} /* (28, 25, 24) {real, imag} */,
  {32'hc0c789c4, 32'h40052f2a} /* (28, 25, 23) {real, imag} */,
  {32'hbf7fb334, 32'h40b65b9e} /* (28, 25, 22) {real, imag} */,
  {32'hc03e3264, 32'h41619751} /* (28, 25, 21) {real, imag} */,
  {32'hc0746f60, 32'hbffd9f48} /* (28, 25, 20) {real, imag} */,
  {32'hc165cd5a, 32'hbfe96304} /* (28, 25, 19) {real, imag} */,
  {32'h413d555a, 32'h40f03682} /* (28, 25, 18) {real, imag} */,
  {32'h411ca8a7, 32'h3ed7fce0} /* (28, 25, 17) {real, imag} */,
  {32'hc02af9b4, 32'hc114efc2} /* (28, 25, 16) {real, imag} */,
  {32'hbfe9ef76, 32'h402527be} /* (28, 25, 15) {real, imag} */,
  {32'hc0f0a5b5, 32'hc0af31b5} /* (28, 25, 14) {real, imag} */,
  {32'h4175da1a, 32'hc07ecdee} /* (28, 25, 13) {real, imag} */,
  {32'hc058a26f, 32'h417dacbf} /* (28, 25, 12) {real, imag} */,
  {32'h3f5efc88, 32'hc15c7ef8} /* (28, 25, 11) {real, imag} */,
  {32'hc110217d, 32'h41a2ab31} /* (28, 25, 10) {real, imag} */,
  {32'hc08868c6, 32'h411e684c} /* (28, 25, 9) {real, imag} */,
  {32'hc15caef2, 32'hc0846b15} /* (28, 25, 8) {real, imag} */,
  {32'hc0b5d977, 32'hc1461cc3} /* (28, 25, 7) {real, imag} */,
  {32'hc10809b7, 32'h414cea20} /* (28, 25, 6) {real, imag} */,
  {32'hc1a53250, 32'hc18ad63f} /* (28, 25, 5) {real, imag} */,
  {32'hc0a946a7, 32'h41697dd1} /* (28, 25, 4) {real, imag} */,
  {32'hbf93d1a0, 32'h408f31f1} /* (28, 25, 3) {real, imag} */,
  {32'hc12ab9d3, 32'hc174c624} /* (28, 25, 2) {real, imag} */,
  {32'hc162a2c5, 32'hc0449763} /* (28, 25, 1) {real, imag} */,
  {32'h4222f657, 32'hc07c1c54} /* (28, 25, 0) {real, imag} */,
  {32'hc19f16fe, 32'h41c06398} /* (28, 24, 31) {real, imag} */,
  {32'h40022cd4, 32'h4009635e} /* (28, 24, 30) {real, imag} */,
  {32'h3e15a910, 32'hc18b78fe} /* (28, 24, 29) {real, imag} */,
  {32'h4193f97d, 32'h4181ebd8} /* (28, 24, 28) {real, imag} */,
  {32'h415eb9fe, 32'hc010fe70} /* (28, 24, 27) {real, imag} */,
  {32'h410acda3, 32'h4125ba40} /* (28, 24, 26) {real, imag} */,
  {32'hc09e2ad4, 32'h41d67ca9} /* (28, 24, 25) {real, imag} */,
  {32'h3fd2e5f0, 32'h40b46c7a} /* (28, 24, 24) {real, imag} */,
  {32'hc07db988, 32'hc0d14cc2} /* (28, 24, 23) {real, imag} */,
  {32'h4159a0b2, 32'hc1392e61} /* (28, 24, 22) {real, imag} */,
  {32'h410ad7be, 32'hc09bf843} /* (28, 24, 21) {real, imag} */,
  {32'hc0d29a4c, 32'hc121a934} /* (28, 24, 20) {real, imag} */,
  {32'hc0b697b5, 32'h40898519} /* (28, 24, 19) {real, imag} */,
  {32'h404d34de, 32'hc0e75e9c} /* (28, 24, 18) {real, imag} */,
  {32'h40bd625e, 32'hc0af0488} /* (28, 24, 17) {real, imag} */,
  {32'hbef180fc, 32'h412d6cde} /* (28, 24, 16) {real, imag} */,
  {32'hc1494cd6, 32'hc05bf3aa} /* (28, 24, 15) {real, imag} */,
  {32'h40a6b263, 32'hbfd79c27} /* (28, 24, 14) {real, imag} */,
  {32'h416a423c, 32'h416bf5fe} /* (28, 24, 13) {real, imag} */,
  {32'h3fc14118, 32'h40ddf628} /* (28, 24, 12) {real, imag} */,
  {32'h414581e2, 32'h4086f76a} /* (28, 24, 11) {real, imag} */,
  {32'hbe840640, 32'hc045824e} /* (28, 24, 10) {real, imag} */,
  {32'h40286ea0, 32'h41897cde} /* (28, 24, 9) {real, imag} */,
  {32'hc1030f86, 32'hc0cdaa41} /* (28, 24, 8) {real, imag} */,
  {32'h40234b92, 32'h4126f9ba} /* (28, 24, 7) {real, imag} */,
  {32'h3f2c371c, 32'hbffa7c24} /* (28, 24, 6) {real, imag} */,
  {32'hc1f28792, 32'h40ce4eb0} /* (28, 24, 5) {real, imag} */,
  {32'hc199b2ab, 32'h3ea15aec} /* (28, 24, 4) {real, imag} */,
  {32'h41dca3b4, 32'h41886d6e} /* (28, 24, 3) {real, imag} */,
  {32'h4215138a, 32'hc19dfc39} /* (28, 24, 2) {real, imag} */,
  {32'hc2728c1c, 32'h414b2b93} /* (28, 24, 1) {real, imag} */,
  {32'hc19e7bf5, 32'h41863c77} /* (28, 24, 0) {real, imag} */,
  {32'h412e7387, 32'hbfde6f48} /* (28, 23, 31) {real, imag} */,
  {32'h41ec98a6, 32'h40fadd06} /* (28, 23, 30) {real, imag} */,
  {32'hc0b5698b, 32'h4073ca38} /* (28, 23, 29) {real, imag} */,
  {32'h415b7e9a, 32'h406a473e} /* (28, 23, 28) {real, imag} */,
  {32'hc0a20c90, 32'hc1663c13} /* (28, 23, 27) {real, imag} */,
  {32'hc0f66202, 32'hbfcd4cb6} /* (28, 23, 26) {real, imag} */,
  {32'h40d606be, 32'hc0674f8c} /* (28, 23, 25) {real, imag} */,
  {32'h40bfa574, 32'h4192cbe6} /* (28, 23, 24) {real, imag} */,
  {32'hbf338978, 32'hc097d866} /* (28, 23, 23) {real, imag} */,
  {32'h3ff0f540, 32'hc05af5aa} /* (28, 23, 22) {real, imag} */,
  {32'hc11ce7f6, 32'h411794a5} /* (28, 23, 21) {real, imag} */,
  {32'hbfaf8006, 32'hc075dfb2} /* (28, 23, 20) {real, imag} */,
  {32'h406d1168, 32'h40885f9a} /* (28, 23, 19) {real, imag} */,
  {32'hbff04682, 32'hc1062cf3} /* (28, 23, 18) {real, imag} */,
  {32'h41143200, 32'hc0973744} /* (28, 23, 17) {real, imag} */,
  {32'h41577184, 32'hc14dd3be} /* (28, 23, 16) {real, imag} */,
  {32'hc06fb6fa, 32'h4094fd19} /* (28, 23, 15) {real, imag} */,
  {32'h40d47c06, 32'hc0d93c95} /* (28, 23, 14) {real, imag} */,
  {32'hc165df9b, 32'hc1659258} /* (28, 23, 13) {real, imag} */,
  {32'h40bb1284, 32'h405632d6} /* (28, 23, 12) {real, imag} */,
  {32'hc1bf00f3, 32'h41795fbb} /* (28, 23, 11) {real, imag} */,
  {32'hc08bd5e4, 32'h405bab9c} /* (28, 23, 10) {real, imag} */,
  {32'h40a78eea, 32'hc0fb8fc8} /* (28, 23, 9) {real, imag} */,
  {32'hc078260a, 32'hc1416772} /* (28, 23, 8) {real, imag} */,
  {32'h40ce2565, 32'hc0e9ab3e} /* (28, 23, 7) {real, imag} */,
  {32'hc1149a26, 32'hc1675a9c} /* (28, 23, 6) {real, imag} */,
  {32'hc1369914, 32'h418782b7} /* (28, 23, 5) {real, imag} */,
  {32'h3f210a2c, 32'hc0ce5360} /* (28, 23, 4) {real, imag} */,
  {32'hc09988fe, 32'h4072de1c} /* (28, 23, 3) {real, imag} */,
  {32'h41c342b2, 32'h41fbff59} /* (28, 23, 2) {real, imag} */,
  {32'hc1b2bf8d, 32'hc1e6e5c8} /* (28, 23, 1) {real, imag} */,
  {32'hc1ac50ea, 32'hc160da6f} /* (28, 23, 0) {real, imag} */,
  {32'h408a17ea, 32'hc04a38fb} /* (28, 22, 31) {real, imag} */,
  {32'hc1832239, 32'h3f48a720} /* (28, 22, 30) {real, imag} */,
  {32'hbea24bc0, 32'h40d6acd9} /* (28, 22, 29) {real, imag} */,
  {32'h4150bca4, 32'hc0b2b845} /* (28, 22, 28) {real, imag} */,
  {32'hc170a6ab, 32'h41165dbe} /* (28, 22, 27) {real, imag} */,
  {32'hc0104988, 32'hbeca9fa0} /* (28, 22, 26) {real, imag} */,
  {32'h40976aba, 32'hc0b87c6e} /* (28, 22, 25) {real, imag} */,
  {32'hc1c6edfa, 32'hc0a80a21} /* (28, 22, 24) {real, imag} */,
  {32'h411fa5d4, 32'hc0ee7f0d} /* (28, 22, 23) {real, imag} */,
  {32'hbf84cebc, 32'hc11e74a2} /* (28, 22, 22) {real, imag} */,
  {32'hc102966a, 32'hbf7de54c} /* (28, 22, 21) {real, imag} */,
  {32'h3e639680, 32'h417092d8} /* (28, 22, 20) {real, imag} */,
  {32'h40b7d593, 32'h4087cb1c} /* (28, 22, 19) {real, imag} */,
  {32'hc187b31a, 32'h409a5459} /* (28, 22, 18) {real, imag} */,
  {32'hc02fd18c, 32'h40e11de1} /* (28, 22, 17) {real, imag} */,
  {32'h409000c8, 32'hc08d82e0} /* (28, 22, 16) {real, imag} */,
  {32'h40e80d20, 32'h40c29620} /* (28, 22, 15) {real, imag} */,
  {32'h41699b1a, 32'h40c758ca} /* (28, 22, 14) {real, imag} */,
  {32'hc0cf6344, 32'hc1097bf8} /* (28, 22, 13) {real, imag} */,
  {32'h4020534c, 32'h40f86116} /* (28, 22, 12) {real, imag} */,
  {32'h400d501c, 32'h41866cbb} /* (28, 22, 11) {real, imag} */,
  {32'hc01ce48a, 32'hc112992f} /* (28, 22, 10) {real, imag} */,
  {32'h4101690e, 32'hbf3e9c3e} /* (28, 22, 9) {real, imag} */,
  {32'hc123c06b, 32'h40037fd8} /* (28, 22, 8) {real, imag} */,
  {32'h3eb798e0, 32'h415d496d} /* (28, 22, 7) {real, imag} */,
  {32'h4134f770, 32'hc086a1a8} /* (28, 22, 6) {real, imag} */,
  {32'hc160849e, 32'h40f81126} /* (28, 22, 5) {real, imag} */,
  {32'h4010ffc2, 32'h41359732} /* (28, 22, 4) {real, imag} */,
  {32'hc04bed66, 32'hc07d8934} /* (28, 22, 3) {real, imag} */,
  {32'h4054083f, 32'h41887439} /* (28, 22, 2) {real, imag} */,
  {32'h41206018, 32'hc12e1fc9} /* (28, 22, 1) {real, imag} */,
  {32'h3ffcfb4c, 32'hc146fb89} /* (28, 22, 0) {real, imag} */,
  {32'hc0bc8e69, 32'h4196f4b7} /* (28, 21, 31) {real, imag} */,
  {32'hc11dbfd5, 32'hc1ed76ae} /* (28, 21, 30) {real, imag} */,
  {32'h40dabaf9, 32'hc197473b} /* (28, 21, 29) {real, imag} */,
  {32'hc12b68c8, 32'h4195e4b6} /* (28, 21, 28) {real, imag} */,
  {32'h41c99cfc, 32'hc0658230} /* (28, 21, 27) {real, imag} */,
  {32'hc12449da, 32'hc1b6cd14} /* (28, 21, 26) {real, imag} */,
  {32'hbd3bbb00, 32'h40cc2418} /* (28, 21, 25) {real, imag} */,
  {32'h40b482b0, 32'h413fd110} /* (28, 21, 24) {real, imag} */,
  {32'h41642a99, 32'hc0fc7356} /* (28, 21, 23) {real, imag} */,
  {32'h412021d5, 32'hc123b569} /* (28, 21, 22) {real, imag} */,
  {32'hc0ce6e32, 32'hc12ba89a} /* (28, 21, 21) {real, imag} */,
  {32'hbf53d770, 32'hbf6f0cc0} /* (28, 21, 20) {real, imag} */,
  {32'h4083f9e7, 32'hc06232f8} /* (28, 21, 19) {real, imag} */,
  {32'h418b6103, 32'hbf3f0444} /* (28, 21, 18) {real, imag} */,
  {32'h411f2511, 32'hc0830764} /* (28, 21, 17) {real, imag} */,
  {32'hc0870568, 32'hc0dee0f6} /* (28, 21, 16) {real, imag} */,
  {32'h4039cd71, 32'hbfdcb90c} /* (28, 21, 15) {real, imag} */,
  {32'hc10105b2, 32'h409a19e0} /* (28, 21, 14) {real, imag} */,
  {32'hc0cc8d13, 32'hbfe45ddc} /* (28, 21, 13) {real, imag} */,
  {32'hc19a5bae, 32'h3f47b6d0} /* (28, 21, 12) {real, imag} */,
  {32'h40f0c3a4, 32'hc1240018} /* (28, 21, 11) {real, imag} */,
  {32'h409a2862, 32'hc09e350c} /* (28, 21, 10) {real, imag} */,
  {32'hc0d9b0f4, 32'h4174ea66} /* (28, 21, 9) {real, imag} */,
  {32'h40d7fcaa, 32'hbfda859a} /* (28, 21, 8) {real, imag} */,
  {32'h41067dec, 32'h3f2ecfe0} /* (28, 21, 7) {real, imag} */,
  {32'h416653ef, 32'hc003885c} /* (28, 21, 6) {real, imag} */,
  {32'hc0aa9407, 32'hc19a0495} /* (28, 21, 5) {real, imag} */,
  {32'hc073d62b, 32'hc0818fd1} /* (28, 21, 4) {real, imag} */,
  {32'h4069f634, 32'h3f6e5c8e} /* (28, 21, 3) {real, imag} */,
  {32'h418549c1, 32'h3f08c9d0} /* (28, 21, 2) {real, imag} */,
  {32'hc0e8a1d9, 32'hc064f526} /* (28, 21, 1) {real, imag} */,
  {32'hc188439a, 32'h412abdb3} /* (28, 21, 0) {real, imag} */,
  {32'hc0a21920, 32'hc159fe70} /* (28, 20, 31) {real, imag} */,
  {32'h3eefbf28, 32'h4124a17e} /* (28, 20, 30) {real, imag} */,
  {32'h41307ed0, 32'hc0c84cc3} /* (28, 20, 29) {real, imag} */,
  {32'h40a3df49, 32'hbe3eadc0} /* (28, 20, 28) {real, imag} */,
  {32'hc09331ac, 32'hc10a04b6} /* (28, 20, 27) {real, imag} */,
  {32'h40e1bf44, 32'h3f90e632} /* (28, 20, 26) {real, imag} */,
  {32'hbfb9de94, 32'h415253af} /* (28, 20, 25) {real, imag} */,
  {32'h3fdf4fb0, 32'hc0b6bcd2} /* (28, 20, 24) {real, imag} */,
  {32'hc0f648f0, 32'h41289fe2} /* (28, 20, 23) {real, imag} */,
  {32'h4164d32f, 32'h419ca5da} /* (28, 20, 22) {real, imag} */,
  {32'hc029e5ee, 32'hc120e548} /* (28, 20, 21) {real, imag} */,
  {32'hc1837018, 32'h3f8196e8} /* (28, 20, 20) {real, imag} */,
  {32'h41be8bbf, 32'h409393d8} /* (28, 20, 19) {real, imag} */,
  {32'hc0e4d25e, 32'h41478131} /* (28, 20, 18) {real, imag} */,
  {32'h405f60a0, 32'hbfc55b34} /* (28, 20, 17) {real, imag} */,
  {32'hc136c43d, 32'hc0826191} /* (28, 20, 16) {real, imag} */,
  {32'hc02b66a6, 32'h410622f7} /* (28, 20, 15) {real, imag} */,
  {32'hc1971273, 32'h402d14f3} /* (28, 20, 14) {real, imag} */,
  {32'h40de9f3a, 32'hc0c25b30} /* (28, 20, 13) {real, imag} */,
  {32'hc044dc2f, 32'hc14a3908} /* (28, 20, 12) {real, imag} */,
  {32'hc12f4610, 32'hc1209d9d} /* (28, 20, 11) {real, imag} */,
  {32'h414d3a36, 32'hc038b6b4} /* (28, 20, 10) {real, imag} */,
  {32'h4015f4e6, 32'h4091ce18} /* (28, 20, 9) {real, imag} */,
  {32'h3f3e4140, 32'hc1689164} /* (28, 20, 8) {real, imag} */,
  {32'hc1a009cc, 32'hbd82e100} /* (28, 20, 7) {real, imag} */,
  {32'hc13b795e, 32'h40548769} /* (28, 20, 6) {real, imag} */,
  {32'h403e4863, 32'hc1ce03cc} /* (28, 20, 5) {real, imag} */,
  {32'hc0312e36, 32'hc13d2ac6} /* (28, 20, 4) {real, imag} */,
  {32'hc1e2b6ec, 32'h4131ed29} /* (28, 20, 3) {real, imag} */,
  {32'h3fffe810, 32'h40a970a9} /* (28, 20, 2) {real, imag} */,
  {32'h41cfa8a3, 32'hbfc00996} /* (28, 20, 1) {real, imag} */,
  {32'h407d4b44, 32'h416f620a} /* (28, 20, 0) {real, imag} */,
  {32'h408d3a78, 32'hc1063a06} /* (28, 19, 31) {real, imag} */,
  {32'h405e71e0, 32'h410040d4} /* (28, 19, 30) {real, imag} */,
  {32'h3f1eecd8, 32'hc12b474a} /* (28, 19, 29) {real, imag} */,
  {32'hc0374272, 32'hc09ae311} /* (28, 19, 28) {real, imag} */,
  {32'hc0b77ac0, 32'hc0d1b29d} /* (28, 19, 27) {real, imag} */,
  {32'h3f3a14b0, 32'h40e6befe} /* (28, 19, 26) {real, imag} */,
  {32'h409d9b08, 32'h41a2e6d6} /* (28, 19, 25) {real, imag} */,
  {32'h41387566, 32'hc086c0f0} /* (28, 19, 24) {real, imag} */,
  {32'hc097e621, 32'hc092536a} /* (28, 19, 23) {real, imag} */,
  {32'hc1563aca, 32'h4102af7e} /* (28, 19, 22) {real, imag} */,
  {32'hbfd082fa, 32'h41215a0a} /* (28, 19, 21) {real, imag} */,
  {32'h412dba6f, 32'hc0baad72} /* (28, 19, 20) {real, imag} */,
  {32'h411e1d8f, 32'hc133b659} /* (28, 19, 19) {real, imag} */,
  {32'h40d59864, 32'hbfeb6f02} /* (28, 19, 18) {real, imag} */,
  {32'hc1157eda, 32'h4129ff9a} /* (28, 19, 17) {real, imag} */,
  {32'h4069ca40, 32'hc146c9fa} /* (28, 19, 16) {real, imag} */,
  {32'h40db3344, 32'hc0b55246} /* (28, 19, 15) {real, imag} */,
  {32'h416613ae, 32'hc0e28aca} /* (28, 19, 14) {real, imag} */,
  {32'h416bb879, 32'hc093f7f5} /* (28, 19, 13) {real, imag} */,
  {32'hc09f0147, 32'hc04d2f90} /* (28, 19, 12) {real, imag} */,
  {32'hc108f832, 32'h4149641b} /* (28, 19, 11) {real, imag} */,
  {32'hbf79578c, 32'h4193229c} /* (28, 19, 10) {real, imag} */,
  {32'hc08a5a5c, 32'hbfb49414} /* (28, 19, 9) {real, imag} */,
  {32'hc0b2aa70, 32'hbf18a0c4} /* (28, 19, 8) {real, imag} */,
  {32'h4024e457, 32'hc1116ccd} /* (28, 19, 7) {real, imag} */,
  {32'hc05ab0fe, 32'h415108c0} /* (28, 19, 6) {real, imag} */,
  {32'h41c1c11e, 32'hc08ac749} /* (28, 19, 5) {real, imag} */,
  {32'hbf323af9, 32'h40d6ca14} /* (28, 19, 4) {real, imag} */,
  {32'h4122bed2, 32'h4090b919} /* (28, 19, 3) {real, imag} */,
  {32'hbf8ed94e, 32'h408f3965} /* (28, 19, 2) {real, imag} */,
  {32'hc11f1ae9, 32'hc00f2fd2} /* (28, 19, 1) {real, imag} */,
  {32'h41118098, 32'h4131f4a3} /* (28, 19, 0) {real, imag} */,
  {32'h405c2658, 32'h3fab087c} /* (28, 18, 31) {real, imag} */,
  {32'hc1118f1e, 32'hc1ba58fb} /* (28, 18, 30) {real, imag} */,
  {32'h3fa28614, 32'h408f1b03} /* (28, 18, 29) {real, imag} */,
  {32'hc0d18b4f, 32'h410e4f0e} /* (28, 18, 28) {real, imag} */,
  {32'hc10f9c2a, 32'hc0b20a0b} /* (28, 18, 27) {real, imag} */,
  {32'hc1017e8d, 32'hc1166dd2} /* (28, 18, 26) {real, imag} */,
  {32'h3fb732b8, 32'h40f91b1c} /* (28, 18, 25) {real, imag} */,
  {32'hc0871a18, 32'h41290686} /* (28, 18, 24) {real, imag} */,
  {32'h3ff39b58, 32'hc1d57fb4} /* (28, 18, 23) {real, imag} */,
  {32'h417e18b4, 32'hc072dca6} /* (28, 18, 22) {real, imag} */,
  {32'hc0c86722, 32'hc0448dbe} /* (28, 18, 21) {real, imag} */,
  {32'h419f44db, 32'h406ac9f2} /* (28, 18, 20) {real, imag} */,
  {32'hc05098f6, 32'hbfe5ad98} /* (28, 18, 19) {real, imag} */,
  {32'h41511c71, 32'hc022535d} /* (28, 18, 18) {real, imag} */,
  {32'h40162df0, 32'h3f7dbd04} /* (28, 18, 17) {real, imag} */,
  {32'hc0e06173, 32'h410287bc} /* (28, 18, 16) {real, imag} */,
  {32'hc101735f, 32'hc125ebb0} /* (28, 18, 15) {real, imag} */,
  {32'h40a64842, 32'hbfe80748} /* (28, 18, 14) {real, imag} */,
  {32'hc013fd5c, 32'hc0ccec14} /* (28, 18, 13) {real, imag} */,
  {32'h3f85d6ab, 32'h40b04824} /* (28, 18, 12) {real, imag} */,
  {32'hc03fc7a3, 32'hc1275896} /* (28, 18, 11) {real, imag} */,
  {32'hc046ca6b, 32'hc0d07bf6} /* (28, 18, 10) {real, imag} */,
  {32'hc0af2148, 32'h41136113} /* (28, 18, 9) {real, imag} */,
  {32'h407cd028, 32'hc0a5f1c1} /* (28, 18, 8) {real, imag} */,
  {32'h40ce1ce9, 32'h409b572c} /* (28, 18, 7) {real, imag} */,
  {32'hc12a1c5b, 32'h4173b9bf} /* (28, 18, 6) {real, imag} */,
  {32'h41836424, 32'h40798898} /* (28, 18, 5) {real, imag} */,
  {32'h406e56ad, 32'h41860f6a} /* (28, 18, 4) {real, imag} */,
  {32'hc09584cd, 32'hc0c5b62a} /* (28, 18, 3) {real, imag} */,
  {32'h411b33b2, 32'hc13ba2b4} /* (28, 18, 2) {real, imag} */,
  {32'hc136aadc, 32'h41099395} /* (28, 18, 1) {real, imag} */,
  {32'h406381dc, 32'h3ff8e32c} /* (28, 18, 0) {real, imag} */,
  {32'h408908d2, 32'hc00da668} /* (28, 17, 31) {real, imag} */,
  {32'hc1074bc4, 32'h40f547c6} /* (28, 17, 30) {real, imag} */,
  {32'h4094472c, 32'h40ae3736} /* (28, 17, 29) {real, imag} */,
  {32'hc15104ca, 32'hc0a36437} /* (28, 17, 28) {real, imag} */,
  {32'hbf10eef0, 32'h410c0ca0} /* (28, 17, 27) {real, imag} */,
  {32'hc09bd671, 32'hc19a731e} /* (28, 17, 26) {real, imag} */,
  {32'h414959c3, 32'hc0a22f77} /* (28, 17, 25) {real, imag} */,
  {32'h417b4853, 32'h410018c5} /* (28, 17, 24) {real, imag} */,
  {32'hc0b1b805, 32'h409ad822} /* (28, 17, 23) {real, imag} */,
  {32'hc108d1dc, 32'hc0b73272} /* (28, 17, 22) {real, imag} */,
  {32'hc11b3bf7, 32'h4194a21c} /* (28, 17, 21) {real, imag} */,
  {32'hc13da522, 32'h40b0127e} /* (28, 17, 20) {real, imag} */,
  {32'hc18522dd, 32'hc0e1e2f0} /* (28, 17, 19) {real, imag} */,
  {32'hc0cb0ac8, 32'h410626a3} /* (28, 17, 18) {real, imag} */,
  {32'h4067165e, 32'hc0c4fd14} /* (28, 17, 17) {real, imag} */,
  {32'h409b76cf, 32'h4099b4ee} /* (28, 17, 16) {real, imag} */,
  {32'h3f983244, 32'h3f3886e8} /* (28, 17, 15) {real, imag} */,
  {32'hc098aa4a, 32'h3f4cf570} /* (28, 17, 14) {real, imag} */,
  {32'h412caf2e, 32'hbf938580} /* (28, 17, 13) {real, imag} */,
  {32'h410937a7, 32'hbff97b1a} /* (28, 17, 12) {real, imag} */,
  {32'h412f8660, 32'h40a91fad} /* (28, 17, 11) {real, imag} */,
  {32'hbfd0c22c, 32'hc0f0c642} /* (28, 17, 10) {real, imag} */,
  {32'h3fd179da, 32'hc0087cd8} /* (28, 17, 9) {real, imag} */,
  {32'h40b4c0a0, 32'h3f59a21c} /* (28, 17, 8) {real, imag} */,
  {32'hc1022c66, 32'h3e77f2a0} /* (28, 17, 7) {real, imag} */,
  {32'hc109d54a, 32'hc054e458} /* (28, 17, 6) {real, imag} */,
  {32'h4010aa27, 32'hc0b47747} /* (28, 17, 5) {real, imag} */,
  {32'h408a2911, 32'h4051ed2a} /* (28, 17, 4) {real, imag} */,
  {32'h41454c12, 32'hc05c7b18} /* (28, 17, 3) {real, imag} */,
  {32'hc157db43, 32'hc0905df3} /* (28, 17, 2) {real, imag} */,
  {32'h40491b52, 32'h3fca728c} /* (28, 17, 1) {real, imag} */,
  {32'hc12ad55c, 32'h40d64d9d} /* (28, 17, 0) {real, imag} */,
  {32'hbef60160, 32'h4113fac9} /* (28, 16, 31) {real, imag} */,
  {32'hc11abf5c, 32'hbf7e3586} /* (28, 16, 30) {real, imag} */,
  {32'h4123fd33, 32'hc0a48845} /* (28, 16, 29) {real, imag} */,
  {32'h40a00579, 32'h409cd382} /* (28, 16, 28) {real, imag} */,
  {32'h3fc9b8f0, 32'hc10e7545} /* (28, 16, 27) {real, imag} */,
  {32'h408912be, 32'hc100fcd6} /* (28, 16, 26) {real, imag} */,
  {32'h3ffef057, 32'hbf953c70} /* (28, 16, 25) {real, imag} */,
  {32'h3f961dda, 32'hc11e1836} /* (28, 16, 24) {real, imag} */,
  {32'hc1827b7f, 32'hc0f02b0f} /* (28, 16, 23) {real, imag} */,
  {32'h41b3d4e0, 32'h40b05d22} /* (28, 16, 22) {real, imag} */,
  {32'h4011a196, 32'h4074239c} /* (28, 16, 21) {real, imag} */,
  {32'h4097510a, 32'h40c404c9} /* (28, 16, 20) {real, imag} */,
  {32'h40adc39d, 32'h401ebd9a} /* (28, 16, 19) {real, imag} */,
  {32'hc059b85a, 32'hc07cebc6} /* (28, 16, 18) {real, imag} */,
  {32'hc02b466c, 32'hbfc99ec8} /* (28, 16, 17) {real, imag} */,
  {32'h41043b32, 32'h00000000} /* (28, 16, 16) {real, imag} */,
  {32'hc02b466c, 32'h3fc99ec8} /* (28, 16, 15) {real, imag} */,
  {32'hc059b85a, 32'h407cebc6} /* (28, 16, 14) {real, imag} */,
  {32'h40adc39d, 32'hc01ebd9a} /* (28, 16, 13) {real, imag} */,
  {32'h4097510a, 32'hc0c404c9} /* (28, 16, 12) {real, imag} */,
  {32'h4011a196, 32'hc074239c} /* (28, 16, 11) {real, imag} */,
  {32'h41b3d4e0, 32'hc0b05d22} /* (28, 16, 10) {real, imag} */,
  {32'hc1827b7f, 32'h40f02b0f} /* (28, 16, 9) {real, imag} */,
  {32'h3f961dda, 32'h411e1836} /* (28, 16, 8) {real, imag} */,
  {32'h3ffef057, 32'h3f953c70} /* (28, 16, 7) {real, imag} */,
  {32'h408912be, 32'h4100fcd6} /* (28, 16, 6) {real, imag} */,
  {32'h3fc9b8f0, 32'h410e7545} /* (28, 16, 5) {real, imag} */,
  {32'h40a00579, 32'hc09cd382} /* (28, 16, 4) {real, imag} */,
  {32'h4123fd33, 32'h40a48845} /* (28, 16, 3) {real, imag} */,
  {32'hc11abf5c, 32'h3f7e3586} /* (28, 16, 2) {real, imag} */,
  {32'hbef60160, 32'hc113fac9} /* (28, 16, 1) {real, imag} */,
  {32'hc130b84b, 32'h00000000} /* (28, 16, 0) {real, imag} */,
  {32'h40491b52, 32'hbfca728c} /* (28, 15, 31) {real, imag} */,
  {32'hc157db43, 32'h40905df3} /* (28, 15, 30) {real, imag} */,
  {32'h41454c12, 32'h405c7b18} /* (28, 15, 29) {real, imag} */,
  {32'h408a2911, 32'hc051ed2a} /* (28, 15, 28) {real, imag} */,
  {32'h4010aa27, 32'h40b47747} /* (28, 15, 27) {real, imag} */,
  {32'hc109d54a, 32'h4054e458} /* (28, 15, 26) {real, imag} */,
  {32'hc1022c66, 32'hbe77f2a0} /* (28, 15, 25) {real, imag} */,
  {32'h40b4c0a0, 32'hbf59a21c} /* (28, 15, 24) {real, imag} */,
  {32'h3fd179da, 32'h40087cd8} /* (28, 15, 23) {real, imag} */,
  {32'hbfd0c22c, 32'h40f0c642} /* (28, 15, 22) {real, imag} */,
  {32'h412f8660, 32'hc0a91fad} /* (28, 15, 21) {real, imag} */,
  {32'h410937a7, 32'h3ff97b1a} /* (28, 15, 20) {real, imag} */,
  {32'h412caf2e, 32'h3f938580} /* (28, 15, 19) {real, imag} */,
  {32'hc098aa4a, 32'hbf4cf570} /* (28, 15, 18) {real, imag} */,
  {32'h3f983244, 32'hbf3886e8} /* (28, 15, 17) {real, imag} */,
  {32'h409b76cf, 32'hc099b4ee} /* (28, 15, 16) {real, imag} */,
  {32'h4067165e, 32'h40c4fd14} /* (28, 15, 15) {real, imag} */,
  {32'hc0cb0ac8, 32'hc10626a3} /* (28, 15, 14) {real, imag} */,
  {32'hc18522dd, 32'h40e1e2f0} /* (28, 15, 13) {real, imag} */,
  {32'hc13da522, 32'hc0b0127e} /* (28, 15, 12) {real, imag} */,
  {32'hc11b3bf7, 32'hc194a21c} /* (28, 15, 11) {real, imag} */,
  {32'hc108d1dc, 32'h40b73272} /* (28, 15, 10) {real, imag} */,
  {32'hc0b1b805, 32'hc09ad822} /* (28, 15, 9) {real, imag} */,
  {32'h417b4853, 32'hc10018c5} /* (28, 15, 8) {real, imag} */,
  {32'h414959c3, 32'h40a22f77} /* (28, 15, 7) {real, imag} */,
  {32'hc09bd671, 32'h419a731e} /* (28, 15, 6) {real, imag} */,
  {32'hbf10eef0, 32'hc10c0ca0} /* (28, 15, 5) {real, imag} */,
  {32'hc15104ca, 32'h40a36437} /* (28, 15, 4) {real, imag} */,
  {32'h4094472c, 32'hc0ae3736} /* (28, 15, 3) {real, imag} */,
  {32'hc1074bc4, 32'hc0f547c6} /* (28, 15, 2) {real, imag} */,
  {32'h408908d2, 32'h400da668} /* (28, 15, 1) {real, imag} */,
  {32'hc12ad55c, 32'hc0d64d9d} /* (28, 15, 0) {real, imag} */,
  {32'hc136aadc, 32'hc1099395} /* (28, 14, 31) {real, imag} */,
  {32'h411b33b2, 32'h413ba2b4} /* (28, 14, 30) {real, imag} */,
  {32'hc09584cd, 32'h40c5b62a} /* (28, 14, 29) {real, imag} */,
  {32'h406e56ad, 32'hc1860f6a} /* (28, 14, 28) {real, imag} */,
  {32'h41836424, 32'hc0798898} /* (28, 14, 27) {real, imag} */,
  {32'hc12a1c5b, 32'hc173b9bf} /* (28, 14, 26) {real, imag} */,
  {32'h40ce1ce9, 32'hc09b572c} /* (28, 14, 25) {real, imag} */,
  {32'h407cd028, 32'h40a5f1c1} /* (28, 14, 24) {real, imag} */,
  {32'hc0af2148, 32'hc1136113} /* (28, 14, 23) {real, imag} */,
  {32'hc046ca6b, 32'h40d07bf6} /* (28, 14, 22) {real, imag} */,
  {32'hc03fc7a3, 32'h41275896} /* (28, 14, 21) {real, imag} */,
  {32'h3f85d6ab, 32'hc0b04824} /* (28, 14, 20) {real, imag} */,
  {32'hc013fd5c, 32'h40ccec14} /* (28, 14, 19) {real, imag} */,
  {32'h40a64842, 32'h3fe80748} /* (28, 14, 18) {real, imag} */,
  {32'hc101735f, 32'h4125ebb0} /* (28, 14, 17) {real, imag} */,
  {32'hc0e06173, 32'hc10287bc} /* (28, 14, 16) {real, imag} */,
  {32'h40162df0, 32'hbf7dbd04} /* (28, 14, 15) {real, imag} */,
  {32'h41511c71, 32'h4022535d} /* (28, 14, 14) {real, imag} */,
  {32'hc05098f6, 32'h3fe5ad98} /* (28, 14, 13) {real, imag} */,
  {32'h419f44db, 32'hc06ac9f2} /* (28, 14, 12) {real, imag} */,
  {32'hc0c86722, 32'h40448dbe} /* (28, 14, 11) {real, imag} */,
  {32'h417e18b4, 32'h4072dca6} /* (28, 14, 10) {real, imag} */,
  {32'h3ff39b58, 32'h41d57fb4} /* (28, 14, 9) {real, imag} */,
  {32'hc0871a18, 32'hc1290686} /* (28, 14, 8) {real, imag} */,
  {32'h3fb732b8, 32'hc0f91b1c} /* (28, 14, 7) {real, imag} */,
  {32'hc1017e8d, 32'h41166dd2} /* (28, 14, 6) {real, imag} */,
  {32'hc10f9c2a, 32'h40b20a0b} /* (28, 14, 5) {real, imag} */,
  {32'hc0d18b4f, 32'hc10e4f0e} /* (28, 14, 4) {real, imag} */,
  {32'h3fa28614, 32'hc08f1b03} /* (28, 14, 3) {real, imag} */,
  {32'hc1118f1e, 32'h41ba58fb} /* (28, 14, 2) {real, imag} */,
  {32'h405c2658, 32'hbfab087c} /* (28, 14, 1) {real, imag} */,
  {32'h406381dc, 32'hbff8e32c} /* (28, 14, 0) {real, imag} */,
  {32'hc11f1ae9, 32'h400f2fd2} /* (28, 13, 31) {real, imag} */,
  {32'hbf8ed94e, 32'hc08f3965} /* (28, 13, 30) {real, imag} */,
  {32'h4122bed2, 32'hc090b919} /* (28, 13, 29) {real, imag} */,
  {32'hbf323af9, 32'hc0d6ca14} /* (28, 13, 28) {real, imag} */,
  {32'h41c1c11e, 32'h408ac749} /* (28, 13, 27) {real, imag} */,
  {32'hc05ab0fe, 32'hc15108c0} /* (28, 13, 26) {real, imag} */,
  {32'h4024e457, 32'h41116ccd} /* (28, 13, 25) {real, imag} */,
  {32'hc0b2aa70, 32'h3f18a0c4} /* (28, 13, 24) {real, imag} */,
  {32'hc08a5a5c, 32'h3fb49414} /* (28, 13, 23) {real, imag} */,
  {32'hbf79578c, 32'hc193229c} /* (28, 13, 22) {real, imag} */,
  {32'hc108f832, 32'hc149641b} /* (28, 13, 21) {real, imag} */,
  {32'hc09f0147, 32'h404d2f90} /* (28, 13, 20) {real, imag} */,
  {32'h416bb879, 32'h4093f7f5} /* (28, 13, 19) {real, imag} */,
  {32'h416613ae, 32'h40e28aca} /* (28, 13, 18) {real, imag} */,
  {32'h40db3344, 32'h40b55246} /* (28, 13, 17) {real, imag} */,
  {32'h4069ca40, 32'h4146c9fa} /* (28, 13, 16) {real, imag} */,
  {32'hc1157eda, 32'hc129ff9a} /* (28, 13, 15) {real, imag} */,
  {32'h40d59864, 32'h3feb6f02} /* (28, 13, 14) {real, imag} */,
  {32'h411e1d8f, 32'h4133b659} /* (28, 13, 13) {real, imag} */,
  {32'h412dba6f, 32'h40baad72} /* (28, 13, 12) {real, imag} */,
  {32'hbfd082fa, 32'hc1215a0a} /* (28, 13, 11) {real, imag} */,
  {32'hc1563aca, 32'hc102af7e} /* (28, 13, 10) {real, imag} */,
  {32'hc097e621, 32'h4092536a} /* (28, 13, 9) {real, imag} */,
  {32'h41387566, 32'h4086c0f0} /* (28, 13, 8) {real, imag} */,
  {32'h409d9b08, 32'hc1a2e6d6} /* (28, 13, 7) {real, imag} */,
  {32'h3f3a14b0, 32'hc0e6befe} /* (28, 13, 6) {real, imag} */,
  {32'hc0b77ac0, 32'h40d1b29d} /* (28, 13, 5) {real, imag} */,
  {32'hc0374272, 32'h409ae311} /* (28, 13, 4) {real, imag} */,
  {32'h3f1eecd8, 32'h412b474a} /* (28, 13, 3) {real, imag} */,
  {32'h405e71e0, 32'hc10040d4} /* (28, 13, 2) {real, imag} */,
  {32'h408d3a78, 32'h41063a06} /* (28, 13, 1) {real, imag} */,
  {32'h41118098, 32'hc131f4a3} /* (28, 13, 0) {real, imag} */,
  {32'h41cfa8a3, 32'h3fc00996} /* (28, 12, 31) {real, imag} */,
  {32'h3fffe810, 32'hc0a970a9} /* (28, 12, 30) {real, imag} */,
  {32'hc1e2b6ec, 32'hc131ed29} /* (28, 12, 29) {real, imag} */,
  {32'hc0312e36, 32'h413d2ac6} /* (28, 12, 28) {real, imag} */,
  {32'h403e4863, 32'h41ce03cc} /* (28, 12, 27) {real, imag} */,
  {32'hc13b795e, 32'hc0548769} /* (28, 12, 26) {real, imag} */,
  {32'hc1a009cc, 32'h3d82e100} /* (28, 12, 25) {real, imag} */,
  {32'h3f3e4140, 32'h41689164} /* (28, 12, 24) {real, imag} */,
  {32'h4015f4e6, 32'hc091ce18} /* (28, 12, 23) {real, imag} */,
  {32'h414d3a36, 32'h4038b6b4} /* (28, 12, 22) {real, imag} */,
  {32'hc12f4610, 32'h41209d9d} /* (28, 12, 21) {real, imag} */,
  {32'hc044dc2f, 32'h414a3908} /* (28, 12, 20) {real, imag} */,
  {32'h40de9f3a, 32'h40c25b30} /* (28, 12, 19) {real, imag} */,
  {32'hc1971273, 32'hc02d14f3} /* (28, 12, 18) {real, imag} */,
  {32'hc02b66a6, 32'hc10622f7} /* (28, 12, 17) {real, imag} */,
  {32'hc136c43d, 32'h40826191} /* (28, 12, 16) {real, imag} */,
  {32'h405f60a0, 32'h3fc55b34} /* (28, 12, 15) {real, imag} */,
  {32'hc0e4d25e, 32'hc1478131} /* (28, 12, 14) {real, imag} */,
  {32'h41be8bbf, 32'hc09393d8} /* (28, 12, 13) {real, imag} */,
  {32'hc1837018, 32'hbf8196e8} /* (28, 12, 12) {real, imag} */,
  {32'hc029e5ee, 32'h4120e548} /* (28, 12, 11) {real, imag} */,
  {32'h4164d32f, 32'hc19ca5da} /* (28, 12, 10) {real, imag} */,
  {32'hc0f648f0, 32'hc1289fe2} /* (28, 12, 9) {real, imag} */,
  {32'h3fdf4fb0, 32'h40b6bcd2} /* (28, 12, 8) {real, imag} */,
  {32'hbfb9de94, 32'hc15253af} /* (28, 12, 7) {real, imag} */,
  {32'h40e1bf44, 32'hbf90e632} /* (28, 12, 6) {real, imag} */,
  {32'hc09331ac, 32'h410a04b6} /* (28, 12, 5) {real, imag} */,
  {32'h40a3df49, 32'h3e3eadc0} /* (28, 12, 4) {real, imag} */,
  {32'h41307ed0, 32'h40c84cc3} /* (28, 12, 3) {real, imag} */,
  {32'h3eefbf28, 32'hc124a17e} /* (28, 12, 2) {real, imag} */,
  {32'hc0a21920, 32'h4159fe70} /* (28, 12, 1) {real, imag} */,
  {32'h407d4b44, 32'hc16f620a} /* (28, 12, 0) {real, imag} */,
  {32'hc0e8a1d9, 32'h4064f526} /* (28, 11, 31) {real, imag} */,
  {32'h418549c1, 32'hbf08c9d0} /* (28, 11, 30) {real, imag} */,
  {32'h4069f634, 32'hbf6e5c8e} /* (28, 11, 29) {real, imag} */,
  {32'hc073d62b, 32'h40818fd1} /* (28, 11, 28) {real, imag} */,
  {32'hc0aa9407, 32'h419a0495} /* (28, 11, 27) {real, imag} */,
  {32'h416653ef, 32'h4003885c} /* (28, 11, 26) {real, imag} */,
  {32'h41067dec, 32'hbf2ecfe0} /* (28, 11, 25) {real, imag} */,
  {32'h40d7fcaa, 32'h3fda859a} /* (28, 11, 24) {real, imag} */,
  {32'hc0d9b0f4, 32'hc174ea66} /* (28, 11, 23) {real, imag} */,
  {32'h409a2862, 32'h409e350c} /* (28, 11, 22) {real, imag} */,
  {32'h40f0c3a4, 32'h41240018} /* (28, 11, 21) {real, imag} */,
  {32'hc19a5bae, 32'hbf47b6d0} /* (28, 11, 20) {real, imag} */,
  {32'hc0cc8d13, 32'h3fe45ddc} /* (28, 11, 19) {real, imag} */,
  {32'hc10105b2, 32'hc09a19e0} /* (28, 11, 18) {real, imag} */,
  {32'h4039cd71, 32'h3fdcb90c} /* (28, 11, 17) {real, imag} */,
  {32'hc0870568, 32'h40dee0f6} /* (28, 11, 16) {real, imag} */,
  {32'h411f2511, 32'h40830764} /* (28, 11, 15) {real, imag} */,
  {32'h418b6103, 32'h3f3f0444} /* (28, 11, 14) {real, imag} */,
  {32'h4083f9e7, 32'h406232f8} /* (28, 11, 13) {real, imag} */,
  {32'hbf53d770, 32'h3f6f0cc0} /* (28, 11, 12) {real, imag} */,
  {32'hc0ce6e32, 32'h412ba89a} /* (28, 11, 11) {real, imag} */,
  {32'h412021d5, 32'h4123b569} /* (28, 11, 10) {real, imag} */,
  {32'h41642a99, 32'h40fc7356} /* (28, 11, 9) {real, imag} */,
  {32'h40b482b0, 32'hc13fd110} /* (28, 11, 8) {real, imag} */,
  {32'hbd3bbb00, 32'hc0cc2418} /* (28, 11, 7) {real, imag} */,
  {32'hc12449da, 32'h41b6cd14} /* (28, 11, 6) {real, imag} */,
  {32'h41c99cfc, 32'h40658230} /* (28, 11, 5) {real, imag} */,
  {32'hc12b68c8, 32'hc195e4b6} /* (28, 11, 4) {real, imag} */,
  {32'h40dabaf9, 32'h4197473b} /* (28, 11, 3) {real, imag} */,
  {32'hc11dbfd5, 32'h41ed76ae} /* (28, 11, 2) {real, imag} */,
  {32'hc0bc8e69, 32'hc196f4b7} /* (28, 11, 1) {real, imag} */,
  {32'hc188439a, 32'hc12abdb3} /* (28, 11, 0) {real, imag} */,
  {32'h41206018, 32'h412e1fc9} /* (28, 10, 31) {real, imag} */,
  {32'h4054083f, 32'hc1887439} /* (28, 10, 30) {real, imag} */,
  {32'hc04bed66, 32'h407d8934} /* (28, 10, 29) {real, imag} */,
  {32'h4010ffc2, 32'hc1359732} /* (28, 10, 28) {real, imag} */,
  {32'hc160849e, 32'hc0f81126} /* (28, 10, 27) {real, imag} */,
  {32'h4134f770, 32'h4086a1a8} /* (28, 10, 26) {real, imag} */,
  {32'h3eb798e0, 32'hc15d496d} /* (28, 10, 25) {real, imag} */,
  {32'hc123c06b, 32'hc0037fd8} /* (28, 10, 24) {real, imag} */,
  {32'h4101690e, 32'h3f3e9c3e} /* (28, 10, 23) {real, imag} */,
  {32'hc01ce48a, 32'h4112992f} /* (28, 10, 22) {real, imag} */,
  {32'h400d501c, 32'hc1866cbb} /* (28, 10, 21) {real, imag} */,
  {32'h4020534c, 32'hc0f86116} /* (28, 10, 20) {real, imag} */,
  {32'hc0cf6344, 32'h41097bf8} /* (28, 10, 19) {real, imag} */,
  {32'h41699b1a, 32'hc0c758ca} /* (28, 10, 18) {real, imag} */,
  {32'h40e80d20, 32'hc0c29620} /* (28, 10, 17) {real, imag} */,
  {32'h409000c8, 32'h408d82e0} /* (28, 10, 16) {real, imag} */,
  {32'hc02fd18c, 32'hc0e11de1} /* (28, 10, 15) {real, imag} */,
  {32'hc187b31a, 32'hc09a5459} /* (28, 10, 14) {real, imag} */,
  {32'h40b7d593, 32'hc087cb1c} /* (28, 10, 13) {real, imag} */,
  {32'h3e639680, 32'hc17092d8} /* (28, 10, 12) {real, imag} */,
  {32'hc102966a, 32'h3f7de54c} /* (28, 10, 11) {real, imag} */,
  {32'hbf84cebc, 32'h411e74a2} /* (28, 10, 10) {real, imag} */,
  {32'h411fa5d4, 32'h40ee7f0d} /* (28, 10, 9) {real, imag} */,
  {32'hc1c6edfa, 32'h40a80a21} /* (28, 10, 8) {real, imag} */,
  {32'h40976aba, 32'h40b87c6e} /* (28, 10, 7) {real, imag} */,
  {32'hc0104988, 32'h3eca9fa0} /* (28, 10, 6) {real, imag} */,
  {32'hc170a6ab, 32'hc1165dbe} /* (28, 10, 5) {real, imag} */,
  {32'h4150bca4, 32'h40b2b845} /* (28, 10, 4) {real, imag} */,
  {32'hbea24bc0, 32'hc0d6acd9} /* (28, 10, 3) {real, imag} */,
  {32'hc1832239, 32'hbf48a720} /* (28, 10, 2) {real, imag} */,
  {32'h408a17ea, 32'h404a38fb} /* (28, 10, 1) {real, imag} */,
  {32'h3ffcfb4c, 32'h4146fb89} /* (28, 10, 0) {real, imag} */,
  {32'hc1b2bf8d, 32'h41e6e5c8} /* (28, 9, 31) {real, imag} */,
  {32'h41c342b2, 32'hc1fbff59} /* (28, 9, 30) {real, imag} */,
  {32'hc09988fe, 32'hc072de1c} /* (28, 9, 29) {real, imag} */,
  {32'h3f210a2c, 32'h40ce5360} /* (28, 9, 28) {real, imag} */,
  {32'hc1369914, 32'hc18782b7} /* (28, 9, 27) {real, imag} */,
  {32'hc1149a26, 32'h41675a9c} /* (28, 9, 26) {real, imag} */,
  {32'h40ce2565, 32'h40e9ab3e} /* (28, 9, 25) {real, imag} */,
  {32'hc078260a, 32'h41416772} /* (28, 9, 24) {real, imag} */,
  {32'h40a78eea, 32'h40fb8fc8} /* (28, 9, 23) {real, imag} */,
  {32'hc08bd5e4, 32'hc05bab9c} /* (28, 9, 22) {real, imag} */,
  {32'hc1bf00f3, 32'hc1795fbb} /* (28, 9, 21) {real, imag} */,
  {32'h40bb1284, 32'hc05632d6} /* (28, 9, 20) {real, imag} */,
  {32'hc165df9b, 32'h41659258} /* (28, 9, 19) {real, imag} */,
  {32'h40d47c06, 32'h40d93c95} /* (28, 9, 18) {real, imag} */,
  {32'hc06fb6fa, 32'hc094fd19} /* (28, 9, 17) {real, imag} */,
  {32'h41577184, 32'h414dd3be} /* (28, 9, 16) {real, imag} */,
  {32'h41143200, 32'h40973744} /* (28, 9, 15) {real, imag} */,
  {32'hbff04682, 32'h41062cf3} /* (28, 9, 14) {real, imag} */,
  {32'h406d1168, 32'hc0885f9a} /* (28, 9, 13) {real, imag} */,
  {32'hbfaf8006, 32'h4075dfb2} /* (28, 9, 12) {real, imag} */,
  {32'hc11ce7f6, 32'hc11794a5} /* (28, 9, 11) {real, imag} */,
  {32'h3ff0f540, 32'h405af5aa} /* (28, 9, 10) {real, imag} */,
  {32'hbf338978, 32'h4097d866} /* (28, 9, 9) {real, imag} */,
  {32'h40bfa574, 32'hc192cbe6} /* (28, 9, 8) {real, imag} */,
  {32'h40d606be, 32'h40674f8c} /* (28, 9, 7) {real, imag} */,
  {32'hc0f66202, 32'h3fcd4cb6} /* (28, 9, 6) {real, imag} */,
  {32'hc0a20c90, 32'h41663c13} /* (28, 9, 5) {real, imag} */,
  {32'h415b7e9a, 32'hc06a473e} /* (28, 9, 4) {real, imag} */,
  {32'hc0b5698b, 32'hc073ca38} /* (28, 9, 3) {real, imag} */,
  {32'h41ec98a6, 32'hc0fadd06} /* (28, 9, 2) {real, imag} */,
  {32'h412e7387, 32'h3fde6f48} /* (28, 9, 1) {real, imag} */,
  {32'hc1ac50ea, 32'h4160da6f} /* (28, 9, 0) {real, imag} */,
  {32'hc2728c1c, 32'hc14b2b93} /* (28, 8, 31) {real, imag} */,
  {32'h4215138a, 32'h419dfc39} /* (28, 8, 30) {real, imag} */,
  {32'h41dca3b4, 32'hc1886d6e} /* (28, 8, 29) {real, imag} */,
  {32'hc199b2ab, 32'hbea15aec} /* (28, 8, 28) {real, imag} */,
  {32'hc1f28792, 32'hc0ce4eb0} /* (28, 8, 27) {real, imag} */,
  {32'h3f2c371c, 32'h3ffa7c24} /* (28, 8, 26) {real, imag} */,
  {32'h40234b92, 32'hc126f9ba} /* (28, 8, 25) {real, imag} */,
  {32'hc1030f86, 32'h40cdaa41} /* (28, 8, 24) {real, imag} */,
  {32'h40286ea0, 32'hc1897cde} /* (28, 8, 23) {real, imag} */,
  {32'hbe840640, 32'h4045824e} /* (28, 8, 22) {real, imag} */,
  {32'h414581e2, 32'hc086f76a} /* (28, 8, 21) {real, imag} */,
  {32'h3fc14118, 32'hc0ddf628} /* (28, 8, 20) {real, imag} */,
  {32'h416a423c, 32'hc16bf5fe} /* (28, 8, 19) {real, imag} */,
  {32'h40a6b263, 32'h3fd79c27} /* (28, 8, 18) {real, imag} */,
  {32'hc1494cd6, 32'h405bf3aa} /* (28, 8, 17) {real, imag} */,
  {32'hbef180fc, 32'hc12d6cde} /* (28, 8, 16) {real, imag} */,
  {32'h40bd625e, 32'h40af0488} /* (28, 8, 15) {real, imag} */,
  {32'h404d34de, 32'h40e75e9c} /* (28, 8, 14) {real, imag} */,
  {32'hc0b697b5, 32'hc0898519} /* (28, 8, 13) {real, imag} */,
  {32'hc0d29a4c, 32'h4121a934} /* (28, 8, 12) {real, imag} */,
  {32'h410ad7be, 32'h409bf843} /* (28, 8, 11) {real, imag} */,
  {32'h4159a0b2, 32'h41392e61} /* (28, 8, 10) {real, imag} */,
  {32'hc07db988, 32'h40d14cc2} /* (28, 8, 9) {real, imag} */,
  {32'h3fd2e5f0, 32'hc0b46c7a} /* (28, 8, 8) {real, imag} */,
  {32'hc09e2ad4, 32'hc1d67ca9} /* (28, 8, 7) {real, imag} */,
  {32'h410acda3, 32'hc125ba40} /* (28, 8, 6) {real, imag} */,
  {32'h415eb9fe, 32'h4010fe70} /* (28, 8, 5) {real, imag} */,
  {32'h4193f97d, 32'hc181ebd8} /* (28, 8, 4) {real, imag} */,
  {32'h3e15a910, 32'h418b78fe} /* (28, 8, 3) {real, imag} */,
  {32'h40022cd4, 32'hc009635e} /* (28, 8, 2) {real, imag} */,
  {32'hc19f16fe, 32'hc1c06398} /* (28, 8, 1) {real, imag} */,
  {32'hc19e7bf5, 32'hc1863c77} /* (28, 8, 0) {real, imag} */,
  {32'hc162a2c5, 32'h40449763} /* (28, 7, 31) {real, imag} */,
  {32'hc12ab9d3, 32'h4174c624} /* (28, 7, 30) {real, imag} */,
  {32'hbf93d1a0, 32'hc08f31f1} /* (28, 7, 29) {real, imag} */,
  {32'hc0a946a7, 32'hc1697dd1} /* (28, 7, 28) {real, imag} */,
  {32'hc1a53250, 32'h418ad63f} /* (28, 7, 27) {real, imag} */,
  {32'hc10809b7, 32'hc14cea20} /* (28, 7, 26) {real, imag} */,
  {32'hc0b5d977, 32'h41461cc3} /* (28, 7, 25) {real, imag} */,
  {32'hc15caef2, 32'h40846b15} /* (28, 7, 24) {real, imag} */,
  {32'hc08868c6, 32'hc11e684c} /* (28, 7, 23) {real, imag} */,
  {32'hc110217d, 32'hc1a2ab31} /* (28, 7, 22) {real, imag} */,
  {32'h3f5efc88, 32'h415c7ef8} /* (28, 7, 21) {real, imag} */,
  {32'hc058a26f, 32'hc17dacbf} /* (28, 7, 20) {real, imag} */,
  {32'h4175da1a, 32'h407ecdee} /* (28, 7, 19) {real, imag} */,
  {32'hc0f0a5b5, 32'h40af31b5} /* (28, 7, 18) {real, imag} */,
  {32'hbfe9ef76, 32'hc02527be} /* (28, 7, 17) {real, imag} */,
  {32'hc02af9b4, 32'h4114efc2} /* (28, 7, 16) {real, imag} */,
  {32'h411ca8a7, 32'hbed7fce0} /* (28, 7, 15) {real, imag} */,
  {32'h413d555a, 32'hc0f03682} /* (28, 7, 14) {real, imag} */,
  {32'hc165cd5a, 32'h3fe96304} /* (28, 7, 13) {real, imag} */,
  {32'hc0746f60, 32'h3ffd9f48} /* (28, 7, 12) {real, imag} */,
  {32'hc03e3264, 32'hc1619751} /* (28, 7, 11) {real, imag} */,
  {32'hbf7fb334, 32'hc0b65b9e} /* (28, 7, 10) {real, imag} */,
  {32'hc0c789c4, 32'hc0052f2a} /* (28, 7, 9) {real, imag} */,
  {32'hc115c0fa, 32'hc18f20e6} /* (28, 7, 8) {real, imag} */,
  {32'h416c5cd6, 32'h4135bfe3} /* (28, 7, 7) {real, imag} */,
  {32'hc0ef16e4, 32'hc045746b} /* (28, 7, 6) {real, imag} */,
  {32'h40e3469c, 32'hbf9adb18} /* (28, 7, 5) {real, imag} */,
  {32'hc06310c4, 32'h4104a790} /* (28, 7, 4) {real, imag} */,
  {32'hc18ea72a, 32'h4184f07a} /* (28, 7, 3) {real, imag} */,
  {32'hc14c56b0, 32'h40ef60a3} /* (28, 7, 2) {real, imag} */,
  {32'h41f54ef2, 32'h4123ccd3} /* (28, 7, 1) {real, imag} */,
  {32'h4222f657, 32'h407c1c54} /* (28, 7, 0) {real, imag} */,
  {32'hc1a51b2e, 32'hbf0f16f0} /* (28, 6, 31) {real, imag} */,
  {32'h41a44c66, 32'h41a62a9c} /* (28, 6, 30) {real, imag} */,
  {32'h413c8296, 32'h4125708d} /* (28, 6, 29) {real, imag} */,
  {32'hc0928b16, 32'hc14eb5da} /* (28, 6, 28) {real, imag} */,
  {32'hc1b11803, 32'hc0d403c1} /* (28, 6, 27) {real, imag} */,
  {32'h412f2d98, 32'hbff7fc68} /* (28, 6, 26) {real, imag} */,
  {32'h40d3b6f0, 32'h417d03bc} /* (28, 6, 25) {real, imag} */,
  {32'h40d88c08, 32'h41aba1e5} /* (28, 6, 24) {real, imag} */,
  {32'h3fd4e3c4, 32'hc0595322} /* (28, 6, 23) {real, imag} */,
  {32'h405d1eb2, 32'h411a2f64} /* (28, 6, 22) {real, imag} */,
  {32'h3eae24d0, 32'hc0744f74} /* (28, 6, 21) {real, imag} */,
  {32'h4124a72c, 32'h4048d146} /* (28, 6, 20) {real, imag} */,
  {32'h408e56cb, 32'hc13d70b8} /* (28, 6, 19) {real, imag} */,
  {32'hc1144c0e, 32'h3fe2ea7a} /* (28, 6, 18) {real, imag} */,
  {32'h40fe5a48, 32'h405d92d4} /* (28, 6, 17) {real, imag} */,
  {32'hc00b5341, 32'hc168dd12} /* (28, 6, 16) {real, imag} */,
  {32'h4050d53f, 32'h40a819f4} /* (28, 6, 15) {real, imag} */,
  {32'hc03b76bc, 32'hc06bca14} /* (28, 6, 14) {real, imag} */,
  {32'hc07cedd8, 32'h41660a54} /* (28, 6, 13) {real, imag} */,
  {32'h40b9fe10, 32'hc03d548c} /* (28, 6, 12) {real, imag} */,
  {32'h41864051, 32'hbfd48410} /* (28, 6, 11) {real, imag} */,
  {32'hc17e4aae, 32'h41443ff2} /* (28, 6, 10) {real, imag} */,
  {32'h412d0edc, 32'hc151388c} /* (28, 6, 9) {real, imag} */,
  {32'hbfdaa980, 32'hc19d89ba} /* (28, 6, 8) {real, imag} */,
  {32'h41c33aa0, 32'h4183f672} /* (28, 6, 7) {real, imag} */,
  {32'hc128d14f, 32'h4131d618} /* (28, 6, 6) {real, imag} */,
  {32'hc08edf2f, 32'hbd7837c0} /* (28, 6, 5) {real, imag} */,
  {32'h40e370ce, 32'h403416b8} /* (28, 6, 4) {real, imag} */,
  {32'h41127e10, 32'h40da764b} /* (28, 6, 3) {real, imag} */,
  {32'h40ca8dbc, 32'hbe851f08} /* (28, 6, 2) {real, imag} */,
  {32'hc18b3c59, 32'hc121aa63} /* (28, 6, 1) {real, imag} */,
  {32'hc0241964, 32'h4163cbaa} /* (28, 6, 0) {real, imag} */,
  {32'hc2d5b67a, 32'hc1bb7554} /* (28, 5, 31) {real, imag} */,
  {32'h4185815e, 32'hc107527e} /* (28, 5, 30) {real, imag} */,
  {32'h40936b43, 32'hc1c181aa} /* (28, 5, 29) {real, imag} */,
  {32'hc19e8c5a, 32'h4088a5c8} /* (28, 5, 28) {real, imag} */,
  {32'h4214909c, 32'h40dd58af} /* (28, 5, 27) {real, imag} */,
  {32'h414ba2aa, 32'hc1a832d4} /* (28, 5, 26) {real, imag} */,
  {32'h4165f15d, 32'h41a7feae} /* (28, 5, 25) {real, imag} */,
  {32'h40125730, 32'hc039732f} /* (28, 5, 24) {real, imag} */,
  {32'h4104279e, 32'h40b016d9} /* (28, 5, 23) {real, imag} */,
  {32'h4111e984, 32'h3fecf340} /* (28, 5, 22) {real, imag} */,
  {32'h412e30f6, 32'hc14c6f27} /* (28, 5, 21) {real, imag} */,
  {32'h3eaa8f78, 32'hbfc27362} /* (28, 5, 20) {real, imag} */,
  {32'hc1169420, 32'h3fdc67a0} /* (28, 5, 19) {real, imag} */,
  {32'hbffada94, 32'h4118b7c9} /* (28, 5, 18) {real, imag} */,
  {32'hbf9b95e8, 32'hc1831d68} /* (28, 5, 17) {real, imag} */,
  {32'hbfe690c3, 32'hc0b02633} /* (28, 5, 16) {real, imag} */,
  {32'hc0185527, 32'h410e20b4} /* (28, 5, 15) {real, imag} */,
  {32'hc0751552, 32'h408ff4c6} /* (28, 5, 14) {real, imag} */,
  {32'hc009a5ca, 32'hc02fa0cc} /* (28, 5, 13) {real, imag} */,
  {32'h40f5ef3b, 32'hc0dd6a0a} /* (28, 5, 12) {real, imag} */,
  {32'hc06c5adc, 32'h40e8cee0} /* (28, 5, 11) {real, imag} */,
  {32'hc0dccc51, 32'hc16532ad} /* (28, 5, 10) {real, imag} */,
  {32'h41147aa6, 32'hc180c0eb} /* (28, 5, 9) {real, imag} */,
  {32'h3ea79cbc, 32'h41382bf8} /* (28, 5, 8) {real, imag} */,
  {32'h3fb59c66, 32'h411f0d35} /* (28, 5, 7) {real, imag} */,
  {32'hc03a380e, 32'h401d063c} /* (28, 5, 6) {real, imag} */,
  {32'h41a1eb24, 32'h41ce45cd} /* (28, 5, 5) {real, imag} */,
  {32'h405eccb8, 32'h41a1b553} /* (28, 5, 4) {real, imag} */,
  {32'hc1386856, 32'hc1a153dc} /* (28, 5, 3) {real, imag} */,
  {32'h41dd4471, 32'hc1d94585} /* (28, 5, 2) {real, imag} */,
  {32'hc2942d54, 32'hc25087b0} /* (28, 5, 1) {real, imag} */,
  {32'hc2736a56, 32'hc21e2570} /* (28, 5, 0) {real, imag} */,
  {32'h4282ba56, 32'h428cc1ba} /* (28, 4, 31) {real, imag} */,
  {32'hc2885c64, 32'hc23a225d} /* (28, 4, 30) {real, imag} */,
  {32'h40be0f14, 32'hc01291f4} /* (28, 4, 29) {real, imag} */,
  {32'h42013465, 32'hc114d7c5} /* (28, 4, 28) {real, imag} */,
  {32'hc067cb7f, 32'h40a72a54} /* (28, 4, 27) {real, imag} */,
  {32'h4182e4c3, 32'h4174cc02} /* (28, 4, 26) {real, imag} */,
  {32'h410cca1c, 32'hc12b05ac} /* (28, 4, 25) {real, imag} */,
  {32'hc14a3c29, 32'h401d77fb} /* (28, 4, 24) {real, imag} */,
  {32'hc17eac1b, 32'h40a930be} /* (28, 4, 23) {real, imag} */,
  {32'hc10ad9fd, 32'h40941e22} /* (28, 4, 22) {real, imag} */,
  {32'hc1a36ae0, 32'h40cdaa93} /* (28, 4, 21) {real, imag} */,
  {32'h41bb9cca, 32'hc13c2635} /* (28, 4, 20) {real, imag} */,
  {32'hbf7f2968, 32'hc00e6de5} /* (28, 4, 19) {real, imag} */,
  {32'h3f28abe8, 32'h40889076} /* (28, 4, 18) {real, imag} */,
  {32'hc03bc62e, 32'h406235a0} /* (28, 4, 17) {real, imag} */,
  {32'h4032c1a2, 32'hc02b470d} /* (28, 4, 16) {real, imag} */,
  {32'hc1214080, 32'h4123fe6d} /* (28, 4, 15) {real, imag} */,
  {32'hc0bd3b40, 32'h401d4bc6} /* (28, 4, 14) {real, imag} */,
  {32'h406eec6e, 32'h40ca7927} /* (28, 4, 13) {real, imag} */,
  {32'h40821d9c, 32'hc19e1e44} /* (28, 4, 12) {real, imag} */,
  {32'h405bd804, 32'h414f20ad} /* (28, 4, 11) {real, imag} */,
  {32'hc004ea30, 32'h40824f41} /* (28, 4, 10) {real, imag} */,
  {32'hc17840ee, 32'hc12b2690} /* (28, 4, 9) {real, imag} */,
  {32'h3fd705cf, 32'hc1042c3c} /* (28, 4, 8) {real, imag} */,
  {32'hc189befe, 32'h40107e14} /* (28, 4, 7) {real, imag} */,
  {32'hbfbf92e0, 32'h41ab8bc5} /* (28, 4, 6) {real, imag} */,
  {32'h40d19af8, 32'hc12c549a} /* (28, 4, 5) {real, imag} */,
  {32'h423cd1c2, 32'hc1d339ac} /* (28, 4, 4) {real, imag} */,
  {32'h41caaf5d, 32'hc2067e75} /* (28, 4, 3) {real, imag} */,
  {32'hc267b92e, 32'hc2971cfb} /* (28, 4, 2) {real, imag} */,
  {32'h42e49c41, 32'h4298f1ba} /* (28, 4, 1) {real, imag} */,
  {32'h420b550a, 32'h424f361d} /* (28, 4, 0) {real, imag} */,
  {32'hc3130f7f, 32'h4222f434} /* (28, 3, 31) {real, imag} */,
  {32'h4295b366, 32'hc2bf95c8} /* (28, 3, 30) {real, imag} */,
  {32'hc1a15212, 32'h40ec96c6} /* (28, 3, 29) {real, imag} */,
  {32'h413df34d, 32'h41ce12ce} /* (28, 3, 28) {real, imag} */,
  {32'hc1283e50, 32'hc1e9021b} /* (28, 3, 27) {real, imag} */,
  {32'h4189f571, 32'hc00f7f58} /* (28, 3, 26) {real, imag} */,
  {32'hc17a7386, 32'h41516e46} /* (28, 3, 25) {real, imag} */,
  {32'hc07943ea, 32'hc1e9089a} /* (28, 3, 24) {real, imag} */,
  {32'h410de770, 32'h4182c896} /* (28, 3, 23) {real, imag} */,
  {32'h41f2ea15, 32'h42077ad3} /* (28, 3, 22) {real, imag} */,
  {32'hc19f03d1, 32'hbef5abc0} /* (28, 3, 21) {real, imag} */,
  {32'h415013f8, 32'hbfea8bca} /* (28, 3, 20) {real, imag} */,
  {32'hc0f32a1b, 32'hc0b2d14f} /* (28, 3, 19) {real, imag} */,
  {32'h40706cdc, 32'hc13feffc} /* (28, 3, 18) {real, imag} */,
  {32'hc0ac6ec9, 32'hc11f7e50} /* (28, 3, 17) {real, imag} */,
  {32'hc10146e2, 32'h3ea6fa20} /* (28, 3, 16) {real, imag} */,
  {32'h40e1b17c, 32'h3fc854e0} /* (28, 3, 15) {real, imag} */,
  {32'hc08e4213, 32'hc0121e58} /* (28, 3, 14) {real, imag} */,
  {32'hc16eccb0, 32'hc1a2567f} /* (28, 3, 13) {real, imag} */,
  {32'hc0d2c720, 32'hc183d950} /* (28, 3, 12) {real, imag} */,
  {32'h4157585b, 32'hc1786ded} /* (28, 3, 11) {real, imag} */,
  {32'hc05abf1e, 32'h40bb725c} /* (28, 3, 10) {real, imag} */,
  {32'hc09ac983, 32'h416a7ee3} /* (28, 3, 9) {real, imag} */,
  {32'h400e7b46, 32'hc0de8a86} /* (28, 3, 8) {real, imag} */,
  {32'h418c29a3, 32'h41054129} /* (28, 3, 7) {real, imag} */,
  {32'hc256890a, 32'hc1a326ad} /* (28, 3, 6) {real, imag} */,
  {32'h41d510a9, 32'hc05698e0} /* (28, 3, 5) {real, imag} */,
  {32'hc004ecfc, 32'h422cba7a} /* (28, 3, 4) {real, imag} */,
  {32'h41e276c6, 32'h4180af85} /* (28, 3, 3) {real, imag} */,
  {32'hc17b7dbb, 32'hc2c77516} /* (28, 3, 2) {real, imag} */,
  {32'h4293bb0d, 32'h43198610} /* (28, 3, 1) {real, imag} */,
  {32'h41afc724, 32'hc1837278} /* (28, 3, 0) {real, imag} */,
  {32'hc425e041, 32'h41d1e393} /* (28, 2, 31) {real, imag} */,
  {32'h43c5513e, 32'hc31b8fb2} /* (28, 2, 30) {real, imag} */,
  {32'hc18fec69, 32'hc0f64a62} /* (28, 2, 29) {real, imag} */,
  {32'hc1c85007, 32'h42aefa3a} /* (28, 2, 28) {real, imag} */,
  {32'h41d91d94, 32'hc1e88b18} /* (28, 2, 27) {real, imag} */,
  {32'h41b1fa1a, 32'h41bfc7c6} /* (28, 2, 26) {real, imag} */,
  {32'hbfb658fa, 32'h422c00c3} /* (28, 2, 25) {real, imag} */,
  {32'h4099aa95, 32'hc2248af4} /* (28, 2, 24) {real, imag} */,
  {32'h408152ed, 32'hc0e68edf} /* (28, 2, 23) {real, imag} */,
  {32'h41b84a46, 32'h4035454a} /* (28, 2, 22) {real, imag} */,
  {32'h3e913890, 32'hc1f6fb7c} /* (28, 2, 21) {real, imag} */,
  {32'h40bfd038, 32'hc0f62b38} /* (28, 2, 20) {real, imag} */,
  {32'hc0dd4be1, 32'h41187722} /* (28, 2, 19) {real, imag} */,
  {32'h4110b6a0, 32'hc163d349} /* (28, 2, 18) {real, imag} */,
  {32'hc0a2ff02, 32'h4177f5b3} /* (28, 2, 17) {real, imag} */,
  {32'h4102a39e, 32'hc073909e} /* (28, 2, 16) {real, imag} */,
  {32'hc0ae6e97, 32'h40f86131} /* (28, 2, 15) {real, imag} */,
  {32'h3fd3b17e, 32'h414b86f1} /* (28, 2, 14) {real, imag} */,
  {32'hc07cbe84, 32'h40c38fe1} /* (28, 2, 13) {real, imag} */,
  {32'hc1190331, 32'hc0bd0ec8} /* (28, 2, 12) {real, imag} */,
  {32'h3f5f00b8, 32'h40c0afd6} /* (28, 2, 11) {real, imag} */,
  {32'hc179d68c, 32'hc0d814a0} /* (28, 2, 10) {real, imag} */,
  {32'h40dd10dc, 32'h41b51a8e} /* (28, 2, 9) {real, imag} */,
  {32'h41b9549f, 32'h41abbf56} /* (28, 2, 8) {real, imag} */,
  {32'hc137df7c, 32'hc0e00a9f} /* (28, 2, 7) {real, imag} */,
  {32'hc077b184, 32'hc031178c} /* (28, 2, 6) {real, imag} */,
  {32'h4232b837, 32'h41db6217} /* (28, 2, 5) {real, imag} */,
  {32'hc2b3813b, 32'hc209fa5c} /* (28, 2, 4) {real, imag} */,
  {32'hc18954e4, 32'hbfe781ec} /* (28, 2, 3) {real, imag} */,
  {32'h4397c4b4, 32'hc2f7ff4a} /* (28, 2, 2) {real, imag} */,
  {32'hc3c1e4c5, 32'h42ca20c0} /* (28, 2, 1) {real, imag} */,
  {32'hc3af5eb5, 32'hc2999eaa} /* (28, 2, 0) {real, imag} */,
  {32'h440cc812, 32'hc33e7672} /* (28, 1, 31) {real, imag} */,
  {32'hc3836f90, 32'h421e4a7b} /* (28, 1, 30) {real, imag} */,
  {32'h4097c6c0, 32'h41207c5e} /* (28, 1, 29) {real, imag} */,
  {32'h42426a2e, 32'h42184bf4} /* (28, 1, 28) {real, imag} */,
  {32'hc2dfa512, 32'h420113ad} /* (28, 1, 27) {real, imag} */,
  {32'hc185e7f1, 32'h4041ae04} /* (28, 1, 26) {real, imag} */,
  {32'hbf9710c0, 32'hc1895d26} /* (28, 1, 25) {real, imag} */,
  {32'hc17df928, 32'h40f519ed} /* (28, 1, 24) {real, imag} */,
  {32'h3cd21e00, 32'h413aa354} /* (28, 1, 23) {real, imag} */,
  {32'hc19a26a2, 32'h41375566} /* (28, 1, 22) {real, imag} */,
  {32'hc16114bc, 32'h40183bde} /* (28, 1, 21) {real, imag} */,
  {32'h400e97fe, 32'hc09e0274} /* (28, 1, 20) {real, imag} */,
  {32'hc1221359, 32'h3e85bf20} /* (28, 1, 19) {real, imag} */,
  {32'h40434f80, 32'h4040008a} /* (28, 1, 18) {real, imag} */,
  {32'h3fea361c, 32'h40bc4fa0} /* (28, 1, 17) {real, imag} */,
  {32'h40165326, 32'hc0aed598} /* (28, 1, 16) {real, imag} */,
  {32'h40921178, 32'h41250ee0} /* (28, 1, 15) {real, imag} */,
  {32'h415c89a0, 32'hc1a9389a} /* (28, 1, 14) {real, imag} */,
  {32'hbf3e7d64, 32'h410294c1} /* (28, 1, 13) {real, imag} */,
  {32'h409ef4c2, 32'hc0853a7b} /* (28, 1, 12) {real, imag} */,
  {32'hc11b96d6, 32'h40fef79c} /* (28, 1, 11) {real, imag} */,
  {32'hc128a226, 32'h401808ef} /* (28, 1, 10) {real, imag} */,
  {32'hc03a5e10, 32'hc11e695c} /* (28, 1, 9) {real, imag} */,
  {32'h3f91aba8, 32'hc1bc0a80} /* (28, 1, 8) {real, imag} */,
  {32'hc17cf2b4, 32'h41c4bdc6} /* (28, 1, 7) {real, imag} */,
  {32'hbf6f8a40, 32'hc13a8ec6} /* (28, 1, 6) {real, imag} */,
  {32'hc280a52d, 32'hc1edc7c4} /* (28, 1, 5) {real, imag} */,
  {32'h4239a870, 32'h4109da7e} /* (28, 1, 4) {real, imag} */,
  {32'hc282ece5, 32'hbf0ac020} /* (28, 1, 3) {real, imag} */,
  {32'hc3bd1793, 32'hc3c9ec43} /* (28, 1, 2) {real, imag} */,
  {32'h444dec3a, 32'h43afa2b3} /* (28, 1, 1) {real, imag} */,
  {32'h43dcc76e, 32'h42721544} /* (28, 1, 0) {real, imag} */,
  {32'h43191d40, 32'hc3337a0d} /* (28, 0, 31) {real, imag} */,
  {32'hc2ee5408, 32'h435d99ac} /* (28, 0, 30) {real, imag} */,
  {32'hc125f894, 32'hc1bc5b31} /* (28, 0, 29) {real, imag} */,
  {32'hc042034c, 32'h417f8618} /* (28, 0, 28) {real, imag} */,
  {32'hc29a31d0, 32'h4151935a} /* (28, 0, 27) {real, imag} */,
  {32'hc044d628, 32'hc106606f} /* (28, 0, 26) {real, imag} */,
  {32'h40ea5be4, 32'hc22a1411} /* (28, 0, 25) {real, imag} */,
  {32'h416591a7, 32'h40ae1464} /* (28, 0, 24) {real, imag} */,
  {32'h403def34, 32'hc10677e0} /* (28, 0, 23) {real, imag} */,
  {32'h3e853cf0, 32'hc01a6088} /* (28, 0, 22) {real, imag} */,
  {32'hc1693342, 32'h41655b4c} /* (28, 0, 21) {real, imag} */,
  {32'h41223e35, 32'hc181a746} /* (28, 0, 20) {real, imag} */,
  {32'hc0ebddfa, 32'hc122b86e} /* (28, 0, 19) {real, imag} */,
  {32'hbfc73d10, 32'hc0fae38b} /* (28, 0, 18) {real, imag} */,
  {32'hc0a57334, 32'h40d1bd7f} /* (28, 0, 17) {real, imag} */,
  {32'hc0cf6430, 32'h00000000} /* (28, 0, 16) {real, imag} */,
  {32'hc0a57334, 32'hc0d1bd7f} /* (28, 0, 15) {real, imag} */,
  {32'hbfc73d10, 32'h40fae38b} /* (28, 0, 14) {real, imag} */,
  {32'hc0ebddfa, 32'h4122b86e} /* (28, 0, 13) {real, imag} */,
  {32'h41223e35, 32'h4181a746} /* (28, 0, 12) {real, imag} */,
  {32'hc1693342, 32'hc1655b4c} /* (28, 0, 11) {real, imag} */,
  {32'h3e853cf0, 32'h401a6088} /* (28, 0, 10) {real, imag} */,
  {32'h403def34, 32'h410677e0} /* (28, 0, 9) {real, imag} */,
  {32'h416591a7, 32'hc0ae1464} /* (28, 0, 8) {real, imag} */,
  {32'h40ea5be4, 32'h422a1411} /* (28, 0, 7) {real, imag} */,
  {32'hc044d628, 32'h4106606f} /* (28, 0, 6) {real, imag} */,
  {32'hc29a31d0, 32'hc151935a} /* (28, 0, 5) {real, imag} */,
  {32'hc042034c, 32'hc17f8618} /* (28, 0, 4) {real, imag} */,
  {32'hc125f894, 32'h41bc5b31} /* (28, 0, 3) {real, imag} */,
  {32'hc2ee5408, 32'hc35d99ac} /* (28, 0, 2) {real, imag} */,
  {32'h43191d40, 32'h43337a0d} /* (28, 0, 1) {real, imag} */,
  {32'hc2e78278, 32'h00000000} /* (28, 0, 0) {real, imag} */,
  {32'h43d0e7c2, 32'hc3324765} /* (27, 31, 31) {real, imag} */,
  {32'hc38eb0ba, 32'h438aeec8} /* (27, 31, 30) {real, imag} */,
  {32'hc242ca0c, 32'h411fcc40} /* (27, 31, 29) {real, imag} */,
  {32'h41f7485f, 32'hc19830e3} /* (27, 31, 28) {real, imag} */,
  {32'hc2628a12, 32'h41e1ba4d} /* (27, 31, 27) {real, imag} */,
  {32'hc0c6a3e6, 32'h4141f8f7} /* (27, 31, 26) {real, imag} */,
  {32'hc19960fd, 32'hc10c7ef0} /* (27, 31, 25) {real, imag} */,
  {32'hc15b6946, 32'h41fc1033} /* (27, 31, 24) {real, imag} */,
  {32'hc1b191f8, 32'h41574fff} /* (27, 31, 23) {real, imag} */,
  {32'hbf044ed0, 32'hc1b2fc27} /* (27, 31, 22) {real, imag} */,
  {32'hc18df652, 32'h414de1ac} /* (27, 31, 21) {real, imag} */,
  {32'hc13213de, 32'hbfeb1ff4} /* (27, 31, 20) {real, imag} */,
  {32'h418823dd, 32'h3f90da8c} /* (27, 31, 19) {real, imag} */,
  {32'h4153acdd, 32'h4171b2f5} /* (27, 31, 18) {real, imag} */,
  {32'hc11017c2, 32'hc16fa48c} /* (27, 31, 17) {real, imag} */,
  {32'hc084dd01, 32'h4085ad3f} /* (27, 31, 16) {real, imag} */,
  {32'hbf14e0e8, 32'hc08538c1} /* (27, 31, 15) {real, imag} */,
  {32'h413bf42a, 32'hc0f50aae} /* (27, 31, 14) {real, imag} */,
  {32'h3fbe4c1e, 32'h41857a26} /* (27, 31, 13) {real, imag} */,
  {32'hc044237e, 32'hc1ad64e8} /* (27, 31, 12) {real, imag} */,
  {32'hc2016acc, 32'hc11163da} /* (27, 31, 11) {real, imag} */,
  {32'hc051c792, 32'h4090aebb} /* (27, 31, 10) {real, imag} */,
  {32'hc0f35c0a, 32'h419dab4e} /* (27, 31, 9) {real, imag} */,
  {32'h3fbb9ab8, 32'hc13ad6a3} /* (27, 31, 8) {real, imag} */,
  {32'h4119fb76, 32'hc1357ac6} /* (27, 31, 7) {real, imag} */,
  {32'hc125eea1, 32'h418ea87b} /* (27, 31, 6) {real, imag} */,
  {32'hc2c9c86f, 32'hc0f4bf50} /* (27, 31, 5) {real, imag} */,
  {32'h41418f7f, 32'hc1ed56af} /* (27, 31, 4) {real, imag} */,
  {32'h40c1b018, 32'hc0c5ff42} /* (27, 31, 3) {real, imag} */,
  {32'hc32180c4, 32'hc2862957} /* (27, 31, 2) {real, imag} */,
  {32'h439803d0, 32'h42fc004e} /* (27, 31, 1) {real, imag} */,
  {32'h4303ac36, 32'h40997190} /* (27, 31, 0) {real, imag} */,
  {32'hc38244db, 32'hc2eb4504} /* (27, 30, 31) {real, imag} */,
  {32'h438100c2, 32'h42d63fb4} /* (27, 30, 30) {real, imag} */,
  {32'h400c2e84, 32'h416fbccf} /* (27, 30, 29) {real, imag} */,
  {32'hc288be87, 32'h425c77a4} /* (27, 30, 28) {real, imag} */,
  {32'h41dc2f2b, 32'hc214c5a7} /* (27, 30, 27) {real, imag} */,
  {32'hbfa4b296, 32'h40867122} /* (27, 30, 26) {real, imag} */,
  {32'hc1047546, 32'h405c2ea0} /* (27, 30, 25) {real, imag} */,
  {32'h419939e4, 32'hc1be9ff9} /* (27, 30, 24) {real, imag} */,
  {32'h40b30e99, 32'hbf979090} /* (27, 30, 23) {real, imag} */,
  {32'hc126da20, 32'h4187c0b5} /* (27, 30, 22) {real, imag} */,
  {32'hc12115d8, 32'hc1b18e1e} /* (27, 30, 21) {real, imag} */,
  {32'hc166fa1c, 32'hc099587e} /* (27, 30, 20) {real, imag} */,
  {32'h3f7ffe46, 32'h413d37d2} /* (27, 30, 19) {real, imag} */,
  {32'h409c1d65, 32'h3f905c88} /* (27, 30, 18) {real, imag} */,
  {32'h3f802f60, 32'hbdcaf2e0} /* (27, 30, 17) {real, imag} */,
  {32'hc108eb1d, 32'h3f8bdd5c} /* (27, 30, 16) {real, imag} */,
  {32'h4180a813, 32'hc0fd52f0} /* (27, 30, 15) {real, imag} */,
  {32'h41231dcf, 32'h4110e1da} /* (27, 30, 14) {real, imag} */,
  {32'hc0378b54, 32'h401c10a8} /* (27, 30, 13) {real, imag} */,
  {32'h411c30e8, 32'hc0c9bfb0} /* (27, 30, 12) {real, imag} */,
  {32'h3feadc14, 32'h40d81515} /* (27, 30, 11) {real, imag} */,
  {32'hc1001b4f, 32'h4137e102} /* (27, 30, 10) {real, imag} */,
  {32'h416cfb96, 32'hc033add3} /* (27, 30, 9) {real, imag} */,
  {32'h4162d8ce, 32'h419d7c5a} /* (27, 30, 8) {real, imag} */,
  {32'hbfde9688, 32'hc2018f7b} /* (27, 30, 7) {real, imag} */,
  {32'h4104fa0c, 32'h40e894fb} /* (27, 30, 6) {real, imag} */,
  {32'h420615a2, 32'h422dbd5b} /* (27, 30, 5) {real, imag} */,
  {32'hc19e34d9, 32'hc2a75e12} /* (27, 30, 4) {real, imag} */,
  {32'hc1b458b2, 32'hbf9d2510} /* (27, 30, 3) {real, imag} */,
  {32'h439da3ec, 32'h42e59e92} /* (27, 30, 2) {real, imag} */,
  {32'hc3db2dce, 32'hc23d744f} /* (27, 30, 1) {real, imag} */,
  {32'hc34e7eff, 32'h42d9d8f0} /* (27, 30, 0) {real, imag} */,
  {32'h425c4ef9, 32'hc2e695fb} /* (27, 29, 31) {real, imag} */,
  {32'hbfc388a0, 32'h42a5c636} /* (27, 29, 30) {real, imag} */,
  {32'hc069513e, 32'hc107f9b4} /* (27, 29, 29) {real, imag} */,
  {32'hbfc35610, 32'hc1f63c0a} /* (27, 29, 28) {real, imag} */,
  {32'h41233c8c, 32'hc032b51a} /* (27, 29, 27) {real, imag} */,
  {32'hc1ecf93a, 32'h40a967a6} /* (27, 29, 26) {real, imag} */,
  {32'h40abba19, 32'hc14cc0e3} /* (27, 29, 25) {real, imag} */,
  {32'hc135d000, 32'hbdeec340} /* (27, 29, 24) {real, imag} */,
  {32'h4149c73a, 32'hc19171e1} /* (27, 29, 23) {real, imag} */,
  {32'hc1495b6c, 32'h41188ab9} /* (27, 29, 22) {real, imag} */,
  {32'h41526b56, 32'h40691f9e} /* (27, 29, 21) {real, imag} */,
  {32'h3faebc9c, 32'h41d8b63c} /* (27, 29, 20) {real, imag} */,
  {32'h401c88a8, 32'hc017533e} /* (27, 29, 19) {real, imag} */,
  {32'hc094ea3a, 32'hc08d50fe} /* (27, 29, 18) {real, imag} */,
  {32'h4013461c, 32'hc063caee} /* (27, 29, 17) {real, imag} */,
  {32'h40ad2138, 32'h411748c6} /* (27, 29, 16) {real, imag} */,
  {32'hc10ebf6e, 32'h41466ba6} /* (27, 29, 15) {real, imag} */,
  {32'h3fa4de4a, 32'h3f5cf09c} /* (27, 29, 14) {real, imag} */,
  {32'hbfc90cee, 32'hc0fecc16} /* (27, 29, 13) {real, imag} */,
  {32'hc0ad0f9e, 32'h41c00362} /* (27, 29, 12) {real, imag} */,
  {32'hc0095674, 32'hc12c2759} /* (27, 29, 11) {real, imag} */,
  {32'h419c31b4, 32'hc1530580} /* (27, 29, 10) {real, imag} */,
  {32'h414b6aba, 32'hc1303d49} /* (27, 29, 9) {real, imag} */,
  {32'hc1dd36f2, 32'h41760dec} /* (27, 29, 8) {real, imag} */,
  {32'h4170100a, 32'hc0a21a1b} /* (27, 29, 7) {real, imag} */,
  {32'h412fb106, 32'hc1b50600} /* (27, 29, 6) {real, imag} */,
  {32'hc191d7a0, 32'h41a10e02} /* (27, 29, 5) {real, imag} */,
  {32'h41be1560, 32'hc1803889} /* (27, 29, 4) {real, imag} */,
  {32'hc15e59b8, 32'hc030fc20} /* (27, 29, 3) {real, imag} */,
  {32'h429e489b, 32'h428c9735} /* (27, 29, 2) {real, imag} */,
  {32'hc2d3fafa, 32'hc1bd7322} /* (27, 29, 1) {real, imag} */,
  {32'h425e5ea8, 32'hc11ca644} /* (27, 29, 0) {real, imag} */,
  {32'h42b881f6, 32'hc2aadb38} /* (27, 28, 31) {real, imag} */,
  {32'hc24a82ad, 32'h4294c728} /* (27, 28, 30) {real, imag} */,
  {32'h41b2c8af, 32'h40a42fba} /* (27, 28, 29) {real, imag} */,
  {32'h4258aefe, 32'h40d24ab0} /* (27, 28, 28) {real, imag} */,
  {32'hc020e50c, 32'h41c530cf} /* (27, 28, 27) {real, imag} */,
  {32'hc149695b, 32'hbf310b48} /* (27, 28, 26) {real, imag} */,
  {32'h40ef767e, 32'hc1301302} /* (27, 28, 25) {real, imag} */,
  {32'hc13351e2, 32'hc0f245e2} /* (27, 28, 24) {real, imag} */,
  {32'h40263342, 32'h411a8b7e} /* (27, 28, 23) {real, imag} */,
  {32'hc0c30bf0, 32'hc100a57e} /* (27, 28, 22) {real, imag} */,
  {32'hc1adde9c, 32'hc125efe1} /* (27, 28, 21) {real, imag} */,
  {32'hbfd2a578, 32'h412e5a12} /* (27, 28, 20) {real, imag} */,
  {32'h40be8789, 32'hc1324175} /* (27, 28, 19) {real, imag} */,
  {32'hc144270c, 32'hc0ce4517} /* (27, 28, 18) {real, imag} */,
  {32'hc08d67d3, 32'hc09d99a1} /* (27, 28, 17) {real, imag} */,
  {32'h3fdf4456, 32'h4080512e} /* (27, 28, 16) {real, imag} */,
  {32'h408cd94e, 32'h401bc627} /* (27, 28, 15) {real, imag} */,
  {32'hbe5947c0, 32'h40e7ec8a} /* (27, 28, 14) {real, imag} */,
  {32'hc0456931, 32'hc13cbc25} /* (27, 28, 13) {real, imag} */,
  {32'h4080a630, 32'h3fc8b968} /* (27, 28, 12) {real, imag} */,
  {32'hc181b231, 32'hc10bb5a0} /* (27, 28, 11) {real, imag} */,
  {32'h41ee405b, 32'h410c89a5} /* (27, 28, 10) {real, imag} */,
  {32'hc06c8c0b, 32'hc113aad8} /* (27, 28, 9) {real, imag} */,
  {32'h40cdb023, 32'h40185976} /* (27, 28, 8) {real, imag} */,
  {32'hc17703d0, 32'h413294b3} /* (27, 28, 7) {real, imag} */,
  {32'hbf8aef70, 32'hc1da1ab0} /* (27, 28, 6) {real, imag} */,
  {32'h413a01b6, 32'h40d1a504} /* (27, 28, 5) {real, imag} */,
  {32'h3fce1194, 32'h40f2622f} /* (27, 28, 4) {real, imag} */,
  {32'h405e9a15, 32'h41831010} /* (27, 28, 3) {real, imag} */,
  {32'hc255cf0f, 32'h425ed96c} /* (27, 28, 2) {real, imag} */,
  {32'h41a732f9, 32'hc21a1c8a} /* (27, 28, 1) {real, imag} */,
  {32'h40697564, 32'hc0e1ba87} /* (27, 28, 0) {real, imag} */,
  {32'hc25a1798, 32'h420e8ee7} /* (27, 27, 31) {real, imag} */,
  {32'h419fb4a0, 32'h412efa44} /* (27, 27, 30) {real, imag} */,
  {32'hbf4c2f50, 32'h41c7fc55} /* (27, 27, 29) {real, imag} */,
  {32'h4144d278, 32'hc0e2403d} /* (27, 27, 28) {real, imag} */,
  {32'h41cd1ee8, 32'hc10f1eb2} /* (27, 27, 27) {real, imag} */,
  {32'h4138836a, 32'hc104c585} /* (27, 27, 26) {real, imag} */,
  {32'hc1655151, 32'h3fd06f30} /* (27, 27, 25) {real, imag} */,
  {32'hbffe3914, 32'hc072bafd} /* (27, 27, 24) {real, imag} */,
  {32'h404aa73a, 32'h413fe0e8} /* (27, 27, 23) {real, imag} */,
  {32'h41597fe0, 32'hc00e5348} /* (27, 27, 22) {real, imag} */,
  {32'hc1416ad7, 32'h41181a95} /* (27, 27, 21) {real, imag} */,
  {32'hc06847af, 32'h418ca2c5} /* (27, 27, 20) {real, imag} */,
  {32'h403deddc, 32'hc07d825c} /* (27, 27, 19) {real, imag} */,
  {32'hc0e28b64, 32'hc0ba13d0} /* (27, 27, 18) {real, imag} */,
  {32'hc0fd9e44, 32'hc10e523d} /* (27, 27, 17) {real, imag} */,
  {32'h3ff26c78, 32'h3f765758} /* (27, 27, 16) {real, imag} */,
  {32'hc098dda3, 32'hc0367f37} /* (27, 27, 15) {real, imag} */,
  {32'h40f2a8cc, 32'h41798082} /* (27, 27, 14) {real, imag} */,
  {32'hc1a55147, 32'hc0887ca9} /* (27, 27, 13) {real, imag} */,
  {32'h4134bb18, 32'h41956e16} /* (27, 27, 12) {real, imag} */,
  {32'hc039d608, 32'h4096789c} /* (27, 27, 11) {real, imag} */,
  {32'hc027b7aa, 32'h4110f9b8} /* (27, 27, 10) {real, imag} */,
  {32'hbee62460, 32'hc193db7a} /* (27, 27, 9) {real, imag} */,
  {32'hc0b2a3d4, 32'hc1aa7853} /* (27, 27, 8) {real, imag} */,
  {32'h40c886c4, 32'hc03fbf6a} /* (27, 27, 7) {real, imag} */,
  {32'hbfe7b4c8, 32'h3fc0e1a8} /* (27, 27, 6) {real, imag} */,
  {32'h41c9df62, 32'h4194b7b2} /* (27, 27, 5) {real, imag} */,
  {32'hc14237e1, 32'hc2024c48} /* (27, 27, 4) {real, imag} */,
  {32'h40a67210, 32'h40d30ea5} /* (27, 27, 3) {real, imag} */,
  {32'h421b5eb8, 32'h418bbabe} /* (27, 27, 2) {real, imag} */,
  {32'hc29fef84, 32'h420af04b} /* (27, 27, 1) {real, imag} */,
  {32'hc28feb59, 32'h4148c32b} /* (27, 27, 0) {real, imag} */,
  {32'hc02dfe14, 32'h41a57130} /* (27, 26, 31) {real, imag} */,
  {32'h41d0a624, 32'h40d23582} /* (27, 26, 30) {real, imag} */,
  {32'hbfbc99b0, 32'h413bc695} /* (27, 26, 29) {real, imag} */,
  {32'hc0b70dd0, 32'hbc581700} /* (27, 26, 28) {real, imag} */,
  {32'h40ad7e68, 32'hbf16f7c8} /* (27, 26, 27) {real, imag} */,
  {32'h3e8d50f0, 32'hc0af6564} /* (27, 26, 26) {real, imag} */,
  {32'h41200e0c, 32'h409209d7} /* (27, 26, 25) {real, imag} */,
  {32'hc1cfe459, 32'hc0fff674} /* (27, 26, 24) {real, imag} */,
  {32'hbf466a14, 32'h4026e71a} /* (27, 26, 23) {real, imag} */,
  {32'hc196a01e, 32'hc0cb4284} /* (27, 26, 22) {real, imag} */,
  {32'hc09a86a8, 32'hc0cf2ee0} /* (27, 26, 21) {real, imag} */,
  {32'hc044c442, 32'h4125c871} /* (27, 26, 20) {real, imag} */,
  {32'h40bd97ee, 32'hc088c70e} /* (27, 26, 19) {real, imag} */,
  {32'hc0fe628b, 32'h412a3c5b} /* (27, 26, 18) {real, imag} */,
  {32'hc096725e, 32'h41834f5e} /* (27, 26, 17) {real, imag} */,
  {32'hc0801044, 32'hc1269c66} /* (27, 26, 16) {real, imag} */,
  {32'h3e9a4610, 32'hc0a894ec} /* (27, 26, 15) {real, imag} */,
  {32'h412ac7ee, 32'h3ec2f100} /* (27, 26, 14) {real, imag} */,
  {32'hc0855830, 32'h41323663} /* (27, 26, 13) {real, imag} */,
  {32'hc1064031, 32'h4140714a} /* (27, 26, 12) {real, imag} */,
  {32'h40e3a359, 32'hc14ee442} /* (27, 26, 11) {real, imag} */,
  {32'h40fed69b, 32'h3e36ce20} /* (27, 26, 10) {real, imag} */,
  {32'hc008924e, 32'h40a9088c} /* (27, 26, 9) {real, imag} */,
  {32'hc11ed2bc, 32'h40ce50cd} /* (27, 26, 8) {real, imag} */,
  {32'hc0c6cf9a, 32'hc0c8b9d2} /* (27, 26, 7) {real, imag} */,
  {32'h4142f739, 32'h41ae63fe} /* (27, 26, 6) {real, imag} */,
  {32'h418388ae, 32'h3ed6be50} /* (27, 26, 5) {real, imag} */,
  {32'h406a3b5c, 32'hc063e24e} /* (27, 26, 4) {real, imag} */,
  {32'h4179c22e, 32'h4108c7c0} /* (27, 26, 3) {real, imag} */,
  {32'hc0987bb3, 32'hc01b9a10} /* (27, 26, 2) {real, imag} */,
  {32'hc19d2f18, 32'h40021646} /* (27, 26, 1) {real, imag} */,
  {32'h40b5af1c, 32'h41be8495} /* (27, 26, 0) {real, imag} */,
  {32'h41cde80b, 32'hc13e775e} /* (27, 25, 31) {real, imag} */,
  {32'hc100fd82, 32'hc135baad} /* (27, 25, 30) {real, imag} */,
  {32'h41884e1e, 32'h4000a54a} /* (27, 25, 29) {real, imag} */,
  {32'h41492ff8, 32'h3fcd6d6e} /* (27, 25, 28) {real, imag} */,
  {32'hc08a9d38, 32'h40df83dc} /* (27, 25, 27) {real, imag} */,
  {32'h416ad942, 32'hc087d093} /* (27, 25, 26) {real, imag} */,
  {32'h4042be7e, 32'hbf29c564} /* (27, 25, 25) {real, imag} */,
  {32'hc0f48170, 32'h41256cbc} /* (27, 25, 24) {real, imag} */,
  {32'h416edafe, 32'hc0b98fa0} /* (27, 25, 23) {real, imag} */,
  {32'h40883331, 32'hc167915d} /* (27, 25, 22) {real, imag} */,
  {32'hc184fb42, 32'h414b0d4d} /* (27, 25, 21) {real, imag} */,
  {32'h40a1d508, 32'hc0433947} /* (27, 25, 20) {real, imag} */,
  {32'hc03f72a4, 32'h40f728e0} /* (27, 25, 19) {real, imag} */,
  {32'h411a993a, 32'hc01ab95e} /* (27, 25, 18) {real, imag} */,
  {32'h40aeffb7, 32'h40e0b5f2} /* (27, 25, 17) {real, imag} */,
  {32'h418b3f1e, 32'hc100ab4d} /* (27, 25, 16) {real, imag} */,
  {32'hc12712ad, 32'h410b232f} /* (27, 25, 15) {real, imag} */,
  {32'hc0eea909, 32'h409c1046} /* (27, 25, 14) {real, imag} */,
  {32'h4145b795, 32'hc0f2fd00} /* (27, 25, 13) {real, imag} */,
  {32'hc1229f3d, 32'h3ff93b08} /* (27, 25, 12) {real, imag} */,
  {32'h41ea6e13, 32'hc0b75baa} /* (27, 25, 11) {real, imag} */,
  {32'h41b37304, 32'h4126109f} /* (27, 25, 10) {real, imag} */,
  {32'h40116ea4, 32'hc1787966} /* (27, 25, 9) {real, imag} */,
  {32'hc0c59762, 32'hc10510f9} /* (27, 25, 8) {real, imag} */,
  {32'h3e8f2600, 32'hc1a52522} /* (27, 25, 7) {real, imag} */,
  {32'h41199720, 32'hc006b660} /* (27, 25, 6) {real, imag} */,
  {32'hc171542f, 32'h3f34f114} /* (27, 25, 5) {real, imag} */,
  {32'hc1809cec, 32'h4194cf23} /* (27, 25, 4) {real, imag} */,
  {32'h40a54207, 32'hbfe918a5} /* (27, 25, 3) {real, imag} */,
  {32'hc0663b04, 32'h41a7f2e8} /* (27, 25, 2) {real, imag} */,
  {32'hc096fd6c, 32'hc1a6946b} /* (27, 25, 1) {real, imag} */,
  {32'h41a10288, 32'h415520ba} /* (27, 25, 0) {real, imag} */,
  {32'hc1ce83cc, 32'h416deb44} /* (27, 24, 31) {real, imag} */,
  {32'h40d01873, 32'hbff79b60} /* (27, 24, 30) {real, imag} */,
  {32'h3f115460, 32'hc125c898} /* (27, 24, 29) {real, imag} */,
  {32'hc1bd9314, 32'h408971d7} /* (27, 24, 28) {real, imag} */,
  {32'h4116684c, 32'hc19fa76a} /* (27, 24, 27) {real, imag} */,
  {32'hc16254e2, 32'h40f5d222} /* (27, 24, 26) {real, imag} */,
  {32'h41d4cc58, 32'hc14cb8aa} /* (27, 24, 25) {real, imag} */,
  {32'hc10ab63c, 32'hbffdf6e0} /* (27, 24, 24) {real, imag} */,
  {32'hc0e2b0da, 32'hbe2de280} /* (27, 24, 23) {real, imag} */,
  {32'hc0267ba8, 32'h41ad71d9} /* (27, 24, 22) {real, imag} */,
  {32'h418929a5, 32'hc1424e7e} /* (27, 24, 21) {real, imag} */,
  {32'h40be398a, 32'h40c178c4} /* (27, 24, 20) {real, imag} */,
  {32'h402ced20, 32'h3eb13930} /* (27, 24, 19) {real, imag} */,
  {32'hc115a0a0, 32'hc18d1dce} /* (27, 24, 18) {real, imag} */,
  {32'hc14de61a, 32'h401654ba} /* (27, 24, 17) {real, imag} */,
  {32'hbf55a6a0, 32'hbfe0e4e4} /* (27, 24, 16) {real, imag} */,
  {32'h4105f180, 32'hc122f7e2} /* (27, 24, 15) {real, imag} */,
  {32'hc0f27e90, 32'hc07dec6f} /* (27, 24, 14) {real, imag} */,
  {32'hbfd7a99f, 32'hc0a4f782} /* (27, 24, 13) {real, imag} */,
  {32'h419d05d8, 32'h41325e51} /* (27, 24, 12) {real, imag} */,
  {32'h41481968, 32'hc0d29627} /* (27, 24, 11) {real, imag} */,
  {32'hc1876675, 32'h404ccf44} /* (27, 24, 10) {real, imag} */,
  {32'hc1390367, 32'h413e830e} /* (27, 24, 9) {real, imag} */,
  {32'h40a3bfb7, 32'hc14072d8} /* (27, 24, 8) {real, imag} */,
  {32'hc012005e, 32'h414512d8} /* (27, 24, 7) {real, imag} */,
  {32'hc0c8d23e, 32'h3e99a310} /* (27, 24, 6) {real, imag} */,
  {32'hc1abe020, 32'h4148f104} /* (27, 24, 5) {real, imag} */,
  {32'h410f8e1e, 32'h41370c9c} /* (27, 24, 4) {real, imag} */,
  {32'h405ce6f8, 32'h418dd46b} /* (27, 24, 3) {real, imag} */,
  {32'h418709a5, 32'hbe84b248} /* (27, 24, 2) {real, imag} */,
  {32'hc232bee8, 32'h418b7f20} /* (27, 24, 1) {real, imag} */,
  {32'hc19d2840, 32'h41081326} /* (27, 24, 0) {real, imag} */,
  {32'h410d731a, 32'h41cbc9ec} /* (27, 23, 31) {real, imag} */,
  {32'h415fb0f0, 32'h415d2c93} /* (27, 23, 30) {real, imag} */,
  {32'hc1171a36, 32'h4184ea97} /* (27, 23, 29) {real, imag} */,
  {32'h3f52f5f2, 32'hc158fce9} /* (27, 23, 28) {real, imag} */,
  {32'h413e9468, 32'hc1c7569e} /* (27, 23, 27) {real, imag} */,
  {32'hc14d7231, 32'hc181192a} /* (27, 23, 26) {real, imag} */,
  {32'hbee800d0, 32'hc15bdae4} /* (27, 23, 25) {real, imag} */,
  {32'h413d17e1, 32'hbe826b10} /* (27, 23, 24) {real, imag} */,
  {32'h41020308, 32'h413ab4fb} /* (27, 23, 23) {real, imag} */,
  {32'hc1078ed7, 32'h411bf1e8} /* (27, 23, 22) {real, imag} */,
  {32'h40fd792e, 32'hc11b2fc2} /* (27, 23, 21) {real, imag} */,
  {32'h3d2dc9c0, 32'hc0cd9232} /* (27, 23, 20) {real, imag} */,
  {32'h40280d1c, 32'h4106218f} /* (27, 23, 19) {real, imag} */,
  {32'h41876bce, 32'hbf80aef6} /* (27, 23, 18) {real, imag} */,
  {32'hbff36f0c, 32'h408941e4} /* (27, 23, 17) {real, imag} */,
  {32'hc08b0f88, 32'hc1440f96} /* (27, 23, 16) {real, imag} */,
  {32'h40998766, 32'hbfcdf3f8} /* (27, 23, 15) {real, imag} */,
  {32'hc01b5548, 32'h40a5ba98} /* (27, 23, 14) {real, imag} */,
  {32'h40abc49f, 32'h416530a8} /* (27, 23, 13) {real, imag} */,
  {32'h4130fde5, 32'h410ebb2e} /* (27, 23, 12) {real, imag} */,
  {32'h411f7095, 32'hc13837c8} /* (27, 23, 11) {real, imag} */,
  {32'hc0acc7e7, 32'h417ae98a} /* (27, 23, 10) {real, imag} */,
  {32'hc09ffffe, 32'h41594c78} /* (27, 23, 9) {real, imag} */,
  {32'hc13b681f, 32'h4176dccd} /* (27, 23, 8) {real, imag} */,
  {32'h411669b3, 32'hc0f52374} /* (27, 23, 7) {real, imag} */,
  {32'hc1867d48, 32'hc13adc64} /* (27, 23, 6) {real, imag} */,
  {32'hc0cc44fb, 32'hbf75c978} /* (27, 23, 5) {real, imag} */,
  {32'hc16aa86f, 32'hc0da38d2} /* (27, 23, 4) {real, imag} */,
  {32'hbfc91df2, 32'h4081f6a6} /* (27, 23, 3) {real, imag} */,
  {32'h41a7efe4, 32'h40e709a8} /* (27, 23, 2) {real, imag} */,
  {32'hc1c2a1a4, 32'hc18c3b53} /* (27, 23, 1) {real, imag} */,
  {32'hc0cd061c, 32'hc14b7d4a} /* (27, 23, 0) {real, imag} */,
  {32'h419c6399, 32'h3e172d50} /* (27, 22, 31) {real, imag} */,
  {32'hc1c5f5bc, 32'h40551794} /* (27, 22, 30) {real, imag} */,
  {32'hc0ddb25c, 32'hc0dd5135} /* (27, 22, 29) {real, imag} */,
  {32'h415d2c9e, 32'hc19bff3e} /* (27, 22, 28) {real, imag} */,
  {32'h4066c88f, 32'h3f433bca} /* (27, 22, 27) {real, imag} */,
  {32'hc009b1bd, 32'h40d4eb28} /* (27, 22, 26) {real, imag} */,
  {32'h4181cd56, 32'h41a27cf8} /* (27, 22, 25) {real, imag} */,
  {32'h41518eed, 32'hc120a4e4} /* (27, 22, 24) {real, imag} */,
  {32'h3f9e4088, 32'h41221fe0} /* (27, 22, 23) {real, imag} */,
  {32'hc063eb06, 32'h40c74d36} /* (27, 22, 22) {real, imag} */,
  {32'hc08effdb, 32'hbf8cce0e} /* (27, 22, 21) {real, imag} */,
  {32'hc0092b94, 32'hc022aac0} /* (27, 22, 20) {real, imag} */,
  {32'hc0cdbe4c, 32'h41161ae9} /* (27, 22, 19) {real, imag} */,
  {32'h3fae4342, 32'h40a56d52} /* (27, 22, 18) {real, imag} */,
  {32'hc12b0677, 32'hc0f70448} /* (27, 22, 17) {real, imag} */,
  {32'h41205302, 32'h40879754} /* (27, 22, 16) {real, imag} */,
  {32'hc0fdff40, 32'hc16b16ee} /* (27, 22, 15) {real, imag} */,
  {32'hc1004ccd, 32'hc083822a} /* (27, 22, 14) {real, imag} */,
  {32'h3f94931c, 32'h41237553} /* (27, 22, 13) {real, imag} */,
  {32'hbfc7bd32, 32'hc153485e} /* (27, 22, 12) {real, imag} */,
  {32'hc126840c, 32'hc0f69cf0} /* (27, 22, 11) {real, imag} */,
  {32'hc1098f61, 32'h41b08573} /* (27, 22, 10) {real, imag} */,
  {32'h40a89623, 32'hc184a87f} /* (27, 22, 9) {real, imag} */,
  {32'h3f0f5db0, 32'h41246940} /* (27, 22, 8) {real, imag} */,
  {32'hc16fb57a, 32'h41008186} /* (27, 22, 7) {real, imag} */,
  {32'h412888bc, 32'h4122990f} /* (27, 22, 6) {real, imag} */,
  {32'hc117dcc3, 32'h41268340} /* (27, 22, 5) {real, imag} */,
  {32'hc0daede9, 32'h409f6cfd} /* (27, 22, 4) {real, imag} */,
  {32'h408d0f72, 32'hc15940e9} /* (27, 22, 3) {real, imag} */,
  {32'h40ca4acb, 32'h4124678a} /* (27, 22, 2) {real, imag} */,
  {32'hc189b75c, 32'hc16880b5} /* (27, 22, 1) {real, imag} */,
  {32'h408778b5, 32'hc007ef2a} /* (27, 22, 0) {real, imag} */,
  {32'hc0a9e3a4, 32'h419fc7aa} /* (27, 21, 31) {real, imag} */,
  {32'hc09755b1, 32'hc1447bc0} /* (27, 21, 30) {real, imag} */,
  {32'h4121b13e, 32'hc0d36579} /* (27, 21, 29) {real, imag} */,
  {32'hbfa8ca58, 32'h412445a9} /* (27, 21, 28) {real, imag} */,
  {32'hc1a57f29, 32'hc148af01} /* (27, 21, 27) {real, imag} */,
  {32'hc180d48d, 32'hc0bc325e} /* (27, 21, 26) {real, imag} */,
  {32'h40ad90ee, 32'h404a204a} /* (27, 21, 25) {real, imag} */,
  {32'h4038c6ce, 32'hbecad680} /* (27, 21, 24) {real, imag} */,
  {32'h41224d76, 32'hc092147a} /* (27, 21, 23) {real, imag} */,
  {32'h3f8fd1d0, 32'h410aad94} /* (27, 21, 22) {real, imag} */,
  {32'h40dbdbf4, 32'hc05903d5} /* (27, 21, 21) {real, imag} */,
  {32'h41067e8a, 32'hc08a8792} /* (27, 21, 20) {real, imag} */,
  {32'hc1a52468, 32'hc112b7a6} /* (27, 21, 19) {real, imag} */,
  {32'h40b4ed21, 32'h4115d0de} /* (27, 21, 18) {real, imag} */,
  {32'hbe035540, 32'hc0a204b0} /* (27, 21, 17) {real, imag} */,
  {32'hc12b08aa, 32'hc155fdfc} /* (27, 21, 16) {real, imag} */,
  {32'hc10537b9, 32'h4151906f} /* (27, 21, 15) {real, imag} */,
  {32'h40ae2d20, 32'h412ab526} /* (27, 21, 14) {real, imag} */,
  {32'h41026210, 32'hc0824daa} /* (27, 21, 13) {real, imag} */,
  {32'h4118261c, 32'hc149e26c} /* (27, 21, 12) {real, imag} */,
  {32'h410c05bd, 32'hc104c589} /* (27, 21, 11) {real, imag} */,
  {32'h3e74cab0, 32'hc16b50cc} /* (27, 21, 10) {real, imag} */,
  {32'h3feea392, 32'h41048896} /* (27, 21, 9) {real, imag} */,
  {32'hc03fb646, 32'h3da3ccd0} /* (27, 21, 8) {real, imag} */,
  {32'h40b41e2e, 32'h416c93ba} /* (27, 21, 7) {real, imag} */,
  {32'hc0659877, 32'h3ff206f2} /* (27, 21, 6) {real, imag} */,
  {32'hbfb02ef3, 32'hc15ee18c} /* (27, 21, 5) {real, imag} */,
  {32'h3f084b40, 32'hc14fc47e} /* (27, 21, 4) {real, imag} */,
  {32'h4168edf2, 32'h41139a3f} /* (27, 21, 3) {real, imag} */,
  {32'h3fbe9d90, 32'h40bb317e} /* (27, 21, 2) {real, imag} */,
  {32'hc0fde776, 32'h413517f0} /* (27, 21, 1) {real, imag} */,
  {32'hc0c17977, 32'h41312387} /* (27, 21, 0) {real, imag} */,
  {32'hc011d5f4, 32'hc10be7ae} /* (27, 20, 31) {real, imag} */,
  {32'hc13c4246, 32'h408ed098} /* (27, 20, 30) {real, imag} */,
  {32'h412da972, 32'hc0edff76} /* (27, 20, 29) {real, imag} */,
  {32'hc19ac1e2, 32'hbfed672c} /* (27, 20, 28) {real, imag} */,
  {32'h41b6285e, 32'h4145493f} /* (27, 20, 27) {real, imag} */,
  {32'hbf31ab08, 32'h41171c61} /* (27, 20, 26) {real, imag} */,
  {32'hc05f7f08, 32'hbf403350} /* (27, 20, 25) {real, imag} */,
  {32'hc07c5e08, 32'h40b0e956} /* (27, 20, 24) {real, imag} */,
  {32'h40e40f44, 32'h41013058} /* (27, 20, 23) {real, imag} */,
  {32'h4168baa3, 32'hc1080b69} /* (27, 20, 22) {real, imag} */,
  {32'h411a296c, 32'h410abab5} /* (27, 20, 21) {real, imag} */,
  {32'hc081e657, 32'h41489d02} /* (27, 20, 20) {real, imag} */,
  {32'h3ff8e6f4, 32'h405a2499} /* (27, 20, 19) {real, imag} */,
  {32'hc1c65766, 32'h40490880} /* (27, 20, 18) {real, imag} */,
  {32'hbe977a20, 32'hc0861c9c} /* (27, 20, 17) {real, imag} */,
  {32'h3e1d0ff8, 32'hc0608d0d} /* (27, 20, 16) {real, imag} */,
  {32'h408cd60b, 32'hc115634f} /* (27, 20, 15) {real, imag} */,
  {32'hc1074e0c, 32'h3ef6e430} /* (27, 20, 14) {real, imag} */,
  {32'h3fcd6dce, 32'h40cc42d7} /* (27, 20, 13) {real, imag} */,
  {32'hc04da95c, 32'hc18bae9b} /* (27, 20, 12) {real, imag} */,
  {32'h413cba34, 32'h41312f9c} /* (27, 20, 11) {real, imag} */,
  {32'h41972d4c, 32'h40ffa70e} /* (27, 20, 10) {real, imag} */,
  {32'h417a1ee6, 32'h4188e680} /* (27, 20, 9) {real, imag} */,
  {32'hc0e269ae, 32'hc1960bc8} /* (27, 20, 8) {real, imag} */,
  {32'h40ffba5c, 32'h40d56326} /* (27, 20, 7) {real, imag} */,
  {32'hc110f92a, 32'h4188bec2} /* (27, 20, 6) {real, imag} */,
  {32'hc05da597, 32'hc1918175} /* (27, 20, 5) {real, imag} */,
  {32'hc18bb2f2, 32'h4117753b} /* (27, 20, 4) {real, imag} */,
  {32'hc0d670c4, 32'h3f0a6b70} /* (27, 20, 3) {real, imag} */,
  {32'hc11cd02b, 32'h417e1bc4} /* (27, 20, 2) {real, imag} */,
  {32'hbe557330, 32'h3fc036ba} /* (27, 20, 1) {real, imag} */,
  {32'h411361ef, 32'h40c2fb8f} /* (27, 20, 0) {real, imag} */,
  {32'h41064276, 32'hc032e441} /* (27, 19, 31) {real, imag} */,
  {32'hc02bdde8, 32'hc0b06b6e} /* (27, 19, 30) {real, imag} */,
  {32'hc0356b96, 32'h3fe8faf1} /* (27, 19, 29) {real, imag} */,
  {32'hc018aab2, 32'h409d2958} /* (27, 19, 28) {real, imag} */,
  {32'h40fddfa5, 32'hc0c7a856} /* (27, 19, 27) {real, imag} */,
  {32'hc1813305, 32'h407da0e0} /* (27, 19, 26) {real, imag} */,
  {32'h40773c98, 32'hc0110c4e} /* (27, 19, 25) {real, imag} */,
  {32'h3fb8f49d, 32'hc1c0be6e} /* (27, 19, 24) {real, imag} */,
  {32'h40c0cd73, 32'hbfa3b7f0} /* (27, 19, 23) {real, imag} */,
  {32'h411b9e66, 32'h407e4d13} /* (27, 19, 22) {real, imag} */,
  {32'hc0a5734f, 32'hc0e9659a} /* (27, 19, 21) {real, imag} */,
  {32'h41199484, 32'hbfbd785c} /* (27, 19, 20) {real, imag} */,
  {32'h410a1e5c, 32'h4188737e} /* (27, 19, 19) {real, imag} */,
  {32'h40dcb82a, 32'h403719e2} /* (27, 19, 18) {real, imag} */,
  {32'h41043b58, 32'h40b8e938} /* (27, 19, 17) {real, imag} */,
  {32'h401cc122, 32'h40dbd0b1} /* (27, 19, 16) {real, imag} */,
  {32'h3f0774c0, 32'hbedc8a10} /* (27, 19, 15) {real, imag} */,
  {32'hc1583360, 32'h40e9be91} /* (27, 19, 14) {real, imag} */,
  {32'hc0d1e522, 32'h4022e74b} /* (27, 19, 13) {real, imag} */,
  {32'hbff22630, 32'h4085faa2} /* (27, 19, 12) {real, imag} */,
  {32'hc02b8e10, 32'hc0facb24} /* (27, 19, 11) {real, imag} */,
  {32'h4117cafb, 32'hc15797ca} /* (27, 19, 10) {real, imag} */,
  {32'h417f2d3a, 32'hc19924c0} /* (27, 19, 9) {real, imag} */,
  {32'h3f93b004, 32'hc0858018} /* (27, 19, 8) {real, imag} */,
  {32'hc0a3d391, 32'h40cd9c03} /* (27, 19, 7) {real, imag} */,
  {32'hc113c571, 32'hbfda251a} /* (27, 19, 6) {real, imag} */,
  {32'h3ecef4f8, 32'hc08fd09d} /* (27, 19, 5) {real, imag} */,
  {32'h4030d64e, 32'h4122c536} /* (27, 19, 4) {real, imag} */,
  {32'hc121d018, 32'hbf7f2b80} /* (27, 19, 3) {real, imag} */,
  {32'hc04e7bc8, 32'h409a3993} /* (27, 19, 2) {real, imag} */,
  {32'hc10af6b6, 32'h3f102060} /* (27, 19, 1) {real, imag} */,
  {32'hc0dee5a4, 32'h40558886} /* (27, 19, 0) {real, imag} */,
  {32'hc10ee311, 32'h41768990} /* (27, 18, 31) {real, imag} */,
  {32'hc00a0a90, 32'hc18b5d9a} /* (27, 18, 30) {real, imag} */,
  {32'h4193c229, 32'h404324a4} /* (27, 18, 29) {real, imag} */,
  {32'hc14a559e, 32'h416228e5} /* (27, 18, 28) {real, imag} */,
  {32'hc0cf82e6, 32'h40a9b716} /* (27, 18, 27) {real, imag} */,
  {32'hbf01252c, 32'hbdafa3c0} /* (27, 18, 26) {real, imag} */,
  {32'hc071704c, 32'hc02e672c} /* (27, 18, 25) {real, imag} */,
  {32'hc00126e0, 32'hc1aebdf9} /* (27, 18, 24) {real, imag} */,
  {32'hc090af1d, 32'hbd8d4530} /* (27, 18, 23) {real, imag} */,
  {32'hc0c2350a, 32'hc109fc9f} /* (27, 18, 22) {real, imag} */,
  {32'h3f2acc80, 32'h40e24622} /* (27, 18, 21) {real, imag} */,
  {32'hc06a5e24, 32'hc1b36762} /* (27, 18, 20) {real, imag} */,
  {32'hc0891777, 32'h40d2db22} /* (27, 18, 19) {real, imag} */,
  {32'h41025519, 32'hc1141e88} /* (27, 18, 18) {real, imag} */,
  {32'h40d52249, 32'h4120b8dd} /* (27, 18, 17) {real, imag} */,
  {32'hbf4f8fa4, 32'hc07f9f6c} /* (27, 18, 16) {real, imag} */,
  {32'h4032c3fd, 32'hc0dc9c16} /* (27, 18, 15) {real, imag} */,
  {32'h40e1d3d8, 32'h3ff3a24f} /* (27, 18, 14) {real, imag} */,
  {32'h408e9f8d, 32'h3d8812e0} /* (27, 18, 13) {real, imag} */,
  {32'h40ae15e0, 32'h4191e91b} /* (27, 18, 12) {real, imag} */,
  {32'h3fd5ffbc, 32'h40840742} /* (27, 18, 11) {real, imag} */,
  {32'hc1a1104c, 32'h41a40f65} /* (27, 18, 10) {real, imag} */,
  {32'hc0d1663f, 32'h4114efb4} /* (27, 18, 9) {real, imag} */,
  {32'h41112acf, 32'hbfc9619e} /* (27, 18, 8) {real, imag} */,
  {32'h410305a2, 32'h40e48712} /* (27, 18, 7) {real, imag} */,
  {32'hc15e7f45, 32'hc01800a4} /* (27, 18, 6) {real, imag} */,
  {32'h3d09d720, 32'h40ded89d} /* (27, 18, 5) {real, imag} */,
  {32'hc0eda60c, 32'h3fb5b7a8} /* (27, 18, 4) {real, imag} */,
  {32'h40927422, 32'h40277b3b} /* (27, 18, 3) {real, imag} */,
  {32'hc0b08450, 32'hc0f43798} /* (27, 18, 2) {real, imag} */,
  {32'hc1928b0b, 32'h411e58c6} /* (27, 18, 1) {real, imag} */,
  {32'hbe6f9ae0, 32'h41383e98} /* (27, 18, 0) {real, imag} */,
  {32'h40b4d318, 32'h3fe50fac} /* (27, 17, 31) {real, imag} */,
  {32'h4089e59f, 32'h414456e7} /* (27, 17, 30) {real, imag} */,
  {32'hc08c0707, 32'h409cc1ac} /* (27, 17, 29) {real, imag} */,
  {32'hc0253772, 32'h41165f16} /* (27, 17, 28) {real, imag} */,
  {32'h40472588, 32'hc0b042c8} /* (27, 17, 27) {real, imag} */,
  {32'h4099e31a, 32'h4021f763} /* (27, 17, 26) {real, imag} */,
  {32'h4051f98e, 32'hc02e7634} /* (27, 17, 25) {real, imag} */,
  {32'hc05f820a, 32'hc01f9ab3} /* (27, 17, 24) {real, imag} */,
  {32'hc10c098a, 32'hc0deccc6} /* (27, 17, 23) {real, imag} */,
  {32'h40ad94cb, 32'hc03f4b96} /* (27, 17, 22) {real, imag} */,
  {32'h4151b982, 32'hc0503464} /* (27, 17, 21) {real, imag} */,
  {32'hbc02cc00, 32'h40e44f8e} /* (27, 17, 20) {real, imag} */,
  {32'hc0593cf6, 32'hc0806df2} /* (27, 17, 19) {real, imag} */,
  {32'hc0704285, 32'h41b00cb4} /* (27, 17, 18) {real, imag} */,
  {32'h3f816a12, 32'h4149ed56} /* (27, 17, 17) {real, imag} */,
  {32'hc0add904, 32'h4039c482} /* (27, 17, 16) {real, imag} */,
  {32'hc00aff41, 32'hc140f3d8} /* (27, 17, 15) {real, imag} */,
  {32'h40360d2e, 32'h41261f7c} /* (27, 17, 14) {real, imag} */,
  {32'h40c77900, 32'hc0954ebd} /* (27, 17, 13) {real, imag} */,
  {32'hc1488ac1, 32'hc145a090} /* (27, 17, 12) {real, imag} */,
  {32'h3f581940, 32'h414a2758} /* (27, 17, 11) {real, imag} */,
  {32'hbf57ddce, 32'hc1c3271c} /* (27, 17, 10) {real, imag} */,
  {32'h40b11d6d, 32'hbe7e9d00} /* (27, 17, 9) {real, imag} */,
  {32'hbeccc010, 32'hc081902a} /* (27, 17, 8) {real, imag} */,
  {32'h410a0aa6, 32'hc0064ec0} /* (27, 17, 7) {real, imag} */,
  {32'h40e69813, 32'h3fd3dd20} /* (27, 17, 6) {real, imag} */,
  {32'hc145fb9a, 32'h411e791a} /* (27, 17, 5) {real, imag} */,
  {32'h4136a53a, 32'hc061b1aa} /* (27, 17, 4) {real, imag} */,
  {32'h40903185, 32'h41226822} /* (27, 17, 3) {real, imag} */,
  {32'hc159ad6a, 32'h4126d0ba} /* (27, 17, 2) {real, imag} */,
  {32'hc124414e, 32'hc01a3934} /* (27, 17, 1) {real, imag} */,
  {32'hc0a842ad, 32'hc10c4bf7} /* (27, 17, 0) {real, imag} */,
  {32'h3f2e38e4, 32'h411dddea} /* (27, 16, 31) {real, imag} */,
  {32'hc097342c, 32'h40ed45ba} /* (27, 16, 30) {real, imag} */,
  {32'h3fbbdc92, 32'h405c73c0} /* (27, 16, 29) {real, imag} */,
  {32'h40999264, 32'hc09d4dec} /* (27, 16, 28) {real, imag} */,
  {32'hc09c746c, 32'h410b8a02} /* (27, 16, 27) {real, imag} */,
  {32'h400f6aa2, 32'h40b75278} /* (27, 16, 26) {real, imag} */,
  {32'h3c83eb40, 32'hc1297fe4} /* (27, 16, 25) {real, imag} */,
  {32'hbfa1b6d4, 32'h4100af56} /* (27, 16, 24) {real, imag} */,
  {32'hc0359594, 32'h3fa88632} /* (27, 16, 23) {real, imag} */,
  {32'h3f0e2ba0, 32'hbf5a3ebe} /* (27, 16, 22) {real, imag} */,
  {32'h4114c1e3, 32'h3ff32876} /* (27, 16, 21) {real, imag} */,
  {32'h40665a8d, 32'hc13fb4ae} /* (27, 16, 20) {real, imag} */,
  {32'hc140241b, 32'hc194932e} /* (27, 16, 19) {real, imag} */,
  {32'h401f567c, 32'h41330c22} /* (27, 16, 18) {real, imag} */,
  {32'hc0bbacbb, 32'h40c4b335} /* (27, 16, 17) {real, imag} */,
  {32'hbf4f940c, 32'h00000000} /* (27, 16, 16) {real, imag} */,
  {32'hc0bbacbb, 32'hc0c4b335} /* (27, 16, 15) {real, imag} */,
  {32'h401f567c, 32'hc1330c22} /* (27, 16, 14) {real, imag} */,
  {32'hc140241b, 32'h4194932e} /* (27, 16, 13) {real, imag} */,
  {32'h40665a8d, 32'h413fb4ae} /* (27, 16, 12) {real, imag} */,
  {32'h4114c1e3, 32'hbff32876} /* (27, 16, 11) {real, imag} */,
  {32'h3f0e2ba0, 32'h3f5a3ebe} /* (27, 16, 10) {real, imag} */,
  {32'hc0359594, 32'hbfa88632} /* (27, 16, 9) {real, imag} */,
  {32'hbfa1b6d4, 32'hc100af56} /* (27, 16, 8) {real, imag} */,
  {32'h3c83eb40, 32'h41297fe4} /* (27, 16, 7) {real, imag} */,
  {32'h400f6aa2, 32'hc0b75278} /* (27, 16, 6) {real, imag} */,
  {32'hc09c746c, 32'hc10b8a02} /* (27, 16, 5) {real, imag} */,
  {32'h40999264, 32'h409d4dec} /* (27, 16, 4) {real, imag} */,
  {32'h3fbbdc92, 32'hc05c73c0} /* (27, 16, 3) {real, imag} */,
  {32'hc097342c, 32'hc0ed45ba} /* (27, 16, 2) {real, imag} */,
  {32'h3f2e38e4, 32'hc11dddea} /* (27, 16, 1) {real, imag} */,
  {32'hc165da4f, 32'h00000000} /* (27, 16, 0) {real, imag} */,
  {32'hc124414e, 32'h401a3934} /* (27, 15, 31) {real, imag} */,
  {32'hc159ad6a, 32'hc126d0ba} /* (27, 15, 30) {real, imag} */,
  {32'h40903185, 32'hc1226822} /* (27, 15, 29) {real, imag} */,
  {32'h4136a53a, 32'h4061b1aa} /* (27, 15, 28) {real, imag} */,
  {32'hc145fb9a, 32'hc11e791a} /* (27, 15, 27) {real, imag} */,
  {32'h40e69813, 32'hbfd3dd20} /* (27, 15, 26) {real, imag} */,
  {32'h410a0aa6, 32'h40064ec0} /* (27, 15, 25) {real, imag} */,
  {32'hbeccc010, 32'h4081902a} /* (27, 15, 24) {real, imag} */,
  {32'h40b11d6d, 32'h3e7e9d00} /* (27, 15, 23) {real, imag} */,
  {32'hbf57ddce, 32'h41c3271c} /* (27, 15, 22) {real, imag} */,
  {32'h3f581940, 32'hc14a2758} /* (27, 15, 21) {real, imag} */,
  {32'hc1488ac1, 32'h4145a090} /* (27, 15, 20) {real, imag} */,
  {32'h40c77900, 32'h40954ebd} /* (27, 15, 19) {real, imag} */,
  {32'h40360d2e, 32'hc1261f7c} /* (27, 15, 18) {real, imag} */,
  {32'hc00aff41, 32'h4140f3d8} /* (27, 15, 17) {real, imag} */,
  {32'hc0add904, 32'hc039c482} /* (27, 15, 16) {real, imag} */,
  {32'h3f816a12, 32'hc149ed56} /* (27, 15, 15) {real, imag} */,
  {32'hc0704285, 32'hc1b00cb4} /* (27, 15, 14) {real, imag} */,
  {32'hc0593cf6, 32'h40806df2} /* (27, 15, 13) {real, imag} */,
  {32'hbc02cc00, 32'hc0e44f8e} /* (27, 15, 12) {real, imag} */,
  {32'h4151b982, 32'h40503464} /* (27, 15, 11) {real, imag} */,
  {32'h40ad94cb, 32'h403f4b96} /* (27, 15, 10) {real, imag} */,
  {32'hc10c098a, 32'h40deccc6} /* (27, 15, 9) {real, imag} */,
  {32'hc05f820a, 32'h401f9ab3} /* (27, 15, 8) {real, imag} */,
  {32'h4051f98e, 32'h402e7634} /* (27, 15, 7) {real, imag} */,
  {32'h4099e31a, 32'hc021f763} /* (27, 15, 6) {real, imag} */,
  {32'h40472588, 32'h40b042c8} /* (27, 15, 5) {real, imag} */,
  {32'hc0253772, 32'hc1165f16} /* (27, 15, 4) {real, imag} */,
  {32'hc08c0707, 32'hc09cc1ac} /* (27, 15, 3) {real, imag} */,
  {32'h4089e59f, 32'hc14456e7} /* (27, 15, 2) {real, imag} */,
  {32'h40b4d318, 32'hbfe50fac} /* (27, 15, 1) {real, imag} */,
  {32'hc0a842ad, 32'h410c4bf7} /* (27, 15, 0) {real, imag} */,
  {32'hc1928b0b, 32'hc11e58c6} /* (27, 14, 31) {real, imag} */,
  {32'hc0b08450, 32'h40f43798} /* (27, 14, 30) {real, imag} */,
  {32'h40927422, 32'hc0277b3b} /* (27, 14, 29) {real, imag} */,
  {32'hc0eda60c, 32'hbfb5b7a8} /* (27, 14, 28) {real, imag} */,
  {32'h3d09d720, 32'hc0ded89d} /* (27, 14, 27) {real, imag} */,
  {32'hc15e7f45, 32'h401800a4} /* (27, 14, 26) {real, imag} */,
  {32'h410305a2, 32'hc0e48712} /* (27, 14, 25) {real, imag} */,
  {32'h41112acf, 32'h3fc9619e} /* (27, 14, 24) {real, imag} */,
  {32'hc0d1663f, 32'hc114efb4} /* (27, 14, 23) {real, imag} */,
  {32'hc1a1104c, 32'hc1a40f65} /* (27, 14, 22) {real, imag} */,
  {32'h3fd5ffbc, 32'hc0840742} /* (27, 14, 21) {real, imag} */,
  {32'h40ae15e0, 32'hc191e91b} /* (27, 14, 20) {real, imag} */,
  {32'h408e9f8d, 32'hbd8812e0} /* (27, 14, 19) {real, imag} */,
  {32'h40e1d3d8, 32'hbff3a24f} /* (27, 14, 18) {real, imag} */,
  {32'h4032c3fd, 32'h40dc9c16} /* (27, 14, 17) {real, imag} */,
  {32'hbf4f8fa4, 32'h407f9f6c} /* (27, 14, 16) {real, imag} */,
  {32'h40d52249, 32'hc120b8dd} /* (27, 14, 15) {real, imag} */,
  {32'h41025519, 32'h41141e88} /* (27, 14, 14) {real, imag} */,
  {32'hc0891777, 32'hc0d2db22} /* (27, 14, 13) {real, imag} */,
  {32'hc06a5e24, 32'h41b36762} /* (27, 14, 12) {real, imag} */,
  {32'h3f2acc80, 32'hc0e24622} /* (27, 14, 11) {real, imag} */,
  {32'hc0c2350a, 32'h4109fc9f} /* (27, 14, 10) {real, imag} */,
  {32'hc090af1d, 32'h3d8d4530} /* (27, 14, 9) {real, imag} */,
  {32'hc00126e0, 32'h41aebdf9} /* (27, 14, 8) {real, imag} */,
  {32'hc071704c, 32'h402e672c} /* (27, 14, 7) {real, imag} */,
  {32'hbf01252c, 32'h3dafa3c0} /* (27, 14, 6) {real, imag} */,
  {32'hc0cf82e6, 32'hc0a9b716} /* (27, 14, 5) {real, imag} */,
  {32'hc14a559e, 32'hc16228e5} /* (27, 14, 4) {real, imag} */,
  {32'h4193c229, 32'hc04324a4} /* (27, 14, 3) {real, imag} */,
  {32'hc00a0a90, 32'h418b5d9a} /* (27, 14, 2) {real, imag} */,
  {32'hc10ee311, 32'hc1768990} /* (27, 14, 1) {real, imag} */,
  {32'hbe6f9ae0, 32'hc1383e98} /* (27, 14, 0) {real, imag} */,
  {32'hc10af6b6, 32'hbf102060} /* (27, 13, 31) {real, imag} */,
  {32'hc04e7bc8, 32'hc09a3993} /* (27, 13, 30) {real, imag} */,
  {32'hc121d018, 32'h3f7f2b80} /* (27, 13, 29) {real, imag} */,
  {32'h4030d64e, 32'hc122c536} /* (27, 13, 28) {real, imag} */,
  {32'h3ecef4f8, 32'h408fd09d} /* (27, 13, 27) {real, imag} */,
  {32'hc113c571, 32'h3fda251a} /* (27, 13, 26) {real, imag} */,
  {32'hc0a3d391, 32'hc0cd9c03} /* (27, 13, 25) {real, imag} */,
  {32'h3f93b004, 32'h40858018} /* (27, 13, 24) {real, imag} */,
  {32'h417f2d3a, 32'h419924c0} /* (27, 13, 23) {real, imag} */,
  {32'h4117cafb, 32'h415797ca} /* (27, 13, 22) {real, imag} */,
  {32'hc02b8e10, 32'h40facb24} /* (27, 13, 21) {real, imag} */,
  {32'hbff22630, 32'hc085faa2} /* (27, 13, 20) {real, imag} */,
  {32'hc0d1e522, 32'hc022e74b} /* (27, 13, 19) {real, imag} */,
  {32'hc1583360, 32'hc0e9be91} /* (27, 13, 18) {real, imag} */,
  {32'h3f0774c0, 32'h3edc8a10} /* (27, 13, 17) {real, imag} */,
  {32'h401cc122, 32'hc0dbd0b1} /* (27, 13, 16) {real, imag} */,
  {32'h41043b58, 32'hc0b8e938} /* (27, 13, 15) {real, imag} */,
  {32'h40dcb82a, 32'hc03719e2} /* (27, 13, 14) {real, imag} */,
  {32'h410a1e5c, 32'hc188737e} /* (27, 13, 13) {real, imag} */,
  {32'h41199484, 32'h3fbd785c} /* (27, 13, 12) {real, imag} */,
  {32'hc0a5734f, 32'h40e9659a} /* (27, 13, 11) {real, imag} */,
  {32'h411b9e66, 32'hc07e4d13} /* (27, 13, 10) {real, imag} */,
  {32'h40c0cd73, 32'h3fa3b7f0} /* (27, 13, 9) {real, imag} */,
  {32'h3fb8f49d, 32'h41c0be6e} /* (27, 13, 8) {real, imag} */,
  {32'h40773c98, 32'h40110c4e} /* (27, 13, 7) {real, imag} */,
  {32'hc1813305, 32'hc07da0e0} /* (27, 13, 6) {real, imag} */,
  {32'h40fddfa5, 32'h40c7a856} /* (27, 13, 5) {real, imag} */,
  {32'hc018aab2, 32'hc09d2958} /* (27, 13, 4) {real, imag} */,
  {32'hc0356b96, 32'hbfe8faf1} /* (27, 13, 3) {real, imag} */,
  {32'hc02bdde8, 32'h40b06b6e} /* (27, 13, 2) {real, imag} */,
  {32'h41064276, 32'h4032e441} /* (27, 13, 1) {real, imag} */,
  {32'hc0dee5a4, 32'hc0558886} /* (27, 13, 0) {real, imag} */,
  {32'hbe557330, 32'hbfc036ba} /* (27, 12, 31) {real, imag} */,
  {32'hc11cd02b, 32'hc17e1bc4} /* (27, 12, 30) {real, imag} */,
  {32'hc0d670c4, 32'hbf0a6b70} /* (27, 12, 29) {real, imag} */,
  {32'hc18bb2f2, 32'hc117753b} /* (27, 12, 28) {real, imag} */,
  {32'hc05da597, 32'h41918175} /* (27, 12, 27) {real, imag} */,
  {32'hc110f92a, 32'hc188bec2} /* (27, 12, 26) {real, imag} */,
  {32'h40ffba5c, 32'hc0d56326} /* (27, 12, 25) {real, imag} */,
  {32'hc0e269ae, 32'h41960bc8} /* (27, 12, 24) {real, imag} */,
  {32'h417a1ee6, 32'hc188e680} /* (27, 12, 23) {real, imag} */,
  {32'h41972d4c, 32'hc0ffa70e} /* (27, 12, 22) {real, imag} */,
  {32'h413cba34, 32'hc1312f9c} /* (27, 12, 21) {real, imag} */,
  {32'hc04da95c, 32'h418bae9b} /* (27, 12, 20) {real, imag} */,
  {32'h3fcd6dce, 32'hc0cc42d7} /* (27, 12, 19) {real, imag} */,
  {32'hc1074e0c, 32'hbef6e430} /* (27, 12, 18) {real, imag} */,
  {32'h408cd60b, 32'h4115634f} /* (27, 12, 17) {real, imag} */,
  {32'h3e1d0ff8, 32'h40608d0d} /* (27, 12, 16) {real, imag} */,
  {32'hbe977a20, 32'h40861c9c} /* (27, 12, 15) {real, imag} */,
  {32'hc1c65766, 32'hc0490880} /* (27, 12, 14) {real, imag} */,
  {32'h3ff8e6f4, 32'hc05a2499} /* (27, 12, 13) {real, imag} */,
  {32'hc081e657, 32'hc1489d02} /* (27, 12, 12) {real, imag} */,
  {32'h411a296c, 32'hc10abab5} /* (27, 12, 11) {real, imag} */,
  {32'h4168baa3, 32'h41080b69} /* (27, 12, 10) {real, imag} */,
  {32'h40e40f44, 32'hc1013058} /* (27, 12, 9) {real, imag} */,
  {32'hc07c5e08, 32'hc0b0e956} /* (27, 12, 8) {real, imag} */,
  {32'hc05f7f08, 32'h3f403350} /* (27, 12, 7) {real, imag} */,
  {32'hbf31ab08, 32'hc1171c61} /* (27, 12, 6) {real, imag} */,
  {32'h41b6285e, 32'hc145493f} /* (27, 12, 5) {real, imag} */,
  {32'hc19ac1e2, 32'h3fed672c} /* (27, 12, 4) {real, imag} */,
  {32'h412da972, 32'h40edff76} /* (27, 12, 3) {real, imag} */,
  {32'hc13c4246, 32'hc08ed098} /* (27, 12, 2) {real, imag} */,
  {32'hc011d5f4, 32'h410be7ae} /* (27, 12, 1) {real, imag} */,
  {32'h411361ef, 32'hc0c2fb8f} /* (27, 12, 0) {real, imag} */,
  {32'hc0fde776, 32'hc13517f0} /* (27, 11, 31) {real, imag} */,
  {32'h3fbe9d90, 32'hc0bb317e} /* (27, 11, 30) {real, imag} */,
  {32'h4168edf2, 32'hc1139a3f} /* (27, 11, 29) {real, imag} */,
  {32'h3f084b40, 32'h414fc47e} /* (27, 11, 28) {real, imag} */,
  {32'hbfb02ef3, 32'h415ee18c} /* (27, 11, 27) {real, imag} */,
  {32'hc0659877, 32'hbff206f2} /* (27, 11, 26) {real, imag} */,
  {32'h40b41e2e, 32'hc16c93ba} /* (27, 11, 25) {real, imag} */,
  {32'hc03fb646, 32'hbda3ccd0} /* (27, 11, 24) {real, imag} */,
  {32'h3feea392, 32'hc1048896} /* (27, 11, 23) {real, imag} */,
  {32'h3e74cab0, 32'h416b50cc} /* (27, 11, 22) {real, imag} */,
  {32'h410c05bd, 32'h4104c589} /* (27, 11, 21) {real, imag} */,
  {32'h4118261c, 32'h4149e26c} /* (27, 11, 20) {real, imag} */,
  {32'h41026210, 32'h40824daa} /* (27, 11, 19) {real, imag} */,
  {32'h40ae2d20, 32'hc12ab526} /* (27, 11, 18) {real, imag} */,
  {32'hc10537b9, 32'hc151906f} /* (27, 11, 17) {real, imag} */,
  {32'hc12b08aa, 32'h4155fdfc} /* (27, 11, 16) {real, imag} */,
  {32'hbe035540, 32'h40a204b0} /* (27, 11, 15) {real, imag} */,
  {32'h40b4ed21, 32'hc115d0de} /* (27, 11, 14) {real, imag} */,
  {32'hc1a52468, 32'h4112b7a6} /* (27, 11, 13) {real, imag} */,
  {32'h41067e8a, 32'h408a8792} /* (27, 11, 12) {real, imag} */,
  {32'h40dbdbf4, 32'h405903d5} /* (27, 11, 11) {real, imag} */,
  {32'h3f8fd1d0, 32'hc10aad94} /* (27, 11, 10) {real, imag} */,
  {32'h41224d76, 32'h4092147a} /* (27, 11, 9) {real, imag} */,
  {32'h4038c6ce, 32'h3ecad680} /* (27, 11, 8) {real, imag} */,
  {32'h40ad90ee, 32'hc04a204a} /* (27, 11, 7) {real, imag} */,
  {32'hc180d48d, 32'h40bc325e} /* (27, 11, 6) {real, imag} */,
  {32'hc1a57f29, 32'h4148af01} /* (27, 11, 5) {real, imag} */,
  {32'hbfa8ca58, 32'hc12445a9} /* (27, 11, 4) {real, imag} */,
  {32'h4121b13e, 32'h40d36579} /* (27, 11, 3) {real, imag} */,
  {32'hc09755b1, 32'h41447bc0} /* (27, 11, 2) {real, imag} */,
  {32'hc0a9e3a4, 32'hc19fc7aa} /* (27, 11, 1) {real, imag} */,
  {32'hc0c17977, 32'hc1312387} /* (27, 11, 0) {real, imag} */,
  {32'hc189b75c, 32'h416880b5} /* (27, 10, 31) {real, imag} */,
  {32'h40ca4acb, 32'hc124678a} /* (27, 10, 30) {real, imag} */,
  {32'h408d0f72, 32'h415940e9} /* (27, 10, 29) {real, imag} */,
  {32'hc0daede9, 32'hc09f6cfd} /* (27, 10, 28) {real, imag} */,
  {32'hc117dcc3, 32'hc1268340} /* (27, 10, 27) {real, imag} */,
  {32'h412888bc, 32'hc122990f} /* (27, 10, 26) {real, imag} */,
  {32'hc16fb57a, 32'hc1008186} /* (27, 10, 25) {real, imag} */,
  {32'h3f0f5db0, 32'hc1246940} /* (27, 10, 24) {real, imag} */,
  {32'h40a89623, 32'h4184a87f} /* (27, 10, 23) {real, imag} */,
  {32'hc1098f61, 32'hc1b08573} /* (27, 10, 22) {real, imag} */,
  {32'hc126840c, 32'h40f69cf0} /* (27, 10, 21) {real, imag} */,
  {32'hbfc7bd32, 32'h4153485e} /* (27, 10, 20) {real, imag} */,
  {32'h3f94931c, 32'hc1237553} /* (27, 10, 19) {real, imag} */,
  {32'hc1004ccd, 32'h4083822a} /* (27, 10, 18) {real, imag} */,
  {32'hc0fdff40, 32'h416b16ee} /* (27, 10, 17) {real, imag} */,
  {32'h41205302, 32'hc0879754} /* (27, 10, 16) {real, imag} */,
  {32'hc12b0677, 32'h40f70448} /* (27, 10, 15) {real, imag} */,
  {32'h3fae4342, 32'hc0a56d52} /* (27, 10, 14) {real, imag} */,
  {32'hc0cdbe4c, 32'hc1161ae9} /* (27, 10, 13) {real, imag} */,
  {32'hc0092b94, 32'h4022aac0} /* (27, 10, 12) {real, imag} */,
  {32'hc08effdb, 32'h3f8cce0e} /* (27, 10, 11) {real, imag} */,
  {32'hc063eb06, 32'hc0c74d36} /* (27, 10, 10) {real, imag} */,
  {32'h3f9e4088, 32'hc1221fe0} /* (27, 10, 9) {real, imag} */,
  {32'h41518eed, 32'h4120a4e4} /* (27, 10, 8) {real, imag} */,
  {32'h4181cd56, 32'hc1a27cf8} /* (27, 10, 7) {real, imag} */,
  {32'hc009b1bd, 32'hc0d4eb28} /* (27, 10, 6) {real, imag} */,
  {32'h4066c88f, 32'hbf433bca} /* (27, 10, 5) {real, imag} */,
  {32'h415d2c9e, 32'h419bff3e} /* (27, 10, 4) {real, imag} */,
  {32'hc0ddb25c, 32'h40dd5135} /* (27, 10, 3) {real, imag} */,
  {32'hc1c5f5bc, 32'hc0551794} /* (27, 10, 2) {real, imag} */,
  {32'h419c6399, 32'hbe172d50} /* (27, 10, 1) {real, imag} */,
  {32'h408778b5, 32'h4007ef2a} /* (27, 10, 0) {real, imag} */,
  {32'hc1c2a1a4, 32'h418c3b53} /* (27, 9, 31) {real, imag} */,
  {32'h41a7efe4, 32'hc0e709a8} /* (27, 9, 30) {real, imag} */,
  {32'hbfc91df2, 32'hc081f6a6} /* (27, 9, 29) {real, imag} */,
  {32'hc16aa86f, 32'h40da38d2} /* (27, 9, 28) {real, imag} */,
  {32'hc0cc44fb, 32'h3f75c978} /* (27, 9, 27) {real, imag} */,
  {32'hc1867d48, 32'h413adc64} /* (27, 9, 26) {real, imag} */,
  {32'h411669b3, 32'h40f52374} /* (27, 9, 25) {real, imag} */,
  {32'hc13b681f, 32'hc176dccd} /* (27, 9, 24) {real, imag} */,
  {32'hc09ffffe, 32'hc1594c78} /* (27, 9, 23) {real, imag} */,
  {32'hc0acc7e7, 32'hc17ae98a} /* (27, 9, 22) {real, imag} */,
  {32'h411f7095, 32'h413837c8} /* (27, 9, 21) {real, imag} */,
  {32'h4130fde5, 32'hc10ebb2e} /* (27, 9, 20) {real, imag} */,
  {32'h40abc49f, 32'hc16530a8} /* (27, 9, 19) {real, imag} */,
  {32'hc01b5548, 32'hc0a5ba98} /* (27, 9, 18) {real, imag} */,
  {32'h40998766, 32'h3fcdf3f8} /* (27, 9, 17) {real, imag} */,
  {32'hc08b0f88, 32'h41440f96} /* (27, 9, 16) {real, imag} */,
  {32'hbff36f0c, 32'hc08941e4} /* (27, 9, 15) {real, imag} */,
  {32'h41876bce, 32'h3f80aef6} /* (27, 9, 14) {real, imag} */,
  {32'h40280d1c, 32'hc106218f} /* (27, 9, 13) {real, imag} */,
  {32'h3d2dc9c0, 32'h40cd9232} /* (27, 9, 12) {real, imag} */,
  {32'h40fd792e, 32'h411b2fc2} /* (27, 9, 11) {real, imag} */,
  {32'hc1078ed7, 32'hc11bf1e8} /* (27, 9, 10) {real, imag} */,
  {32'h41020308, 32'hc13ab4fb} /* (27, 9, 9) {real, imag} */,
  {32'h413d17e1, 32'h3e826b10} /* (27, 9, 8) {real, imag} */,
  {32'hbee800d0, 32'h415bdae4} /* (27, 9, 7) {real, imag} */,
  {32'hc14d7231, 32'h4181192a} /* (27, 9, 6) {real, imag} */,
  {32'h413e9468, 32'h41c7569e} /* (27, 9, 5) {real, imag} */,
  {32'h3f52f5f2, 32'h4158fce9} /* (27, 9, 4) {real, imag} */,
  {32'hc1171a36, 32'hc184ea97} /* (27, 9, 3) {real, imag} */,
  {32'h415fb0f0, 32'hc15d2c93} /* (27, 9, 2) {real, imag} */,
  {32'h410d731a, 32'hc1cbc9ec} /* (27, 9, 1) {real, imag} */,
  {32'hc0cd061c, 32'h414b7d4a} /* (27, 9, 0) {real, imag} */,
  {32'hc232bee8, 32'hc18b7f20} /* (27, 8, 31) {real, imag} */,
  {32'h418709a5, 32'h3e84b248} /* (27, 8, 30) {real, imag} */,
  {32'h405ce6f8, 32'hc18dd46b} /* (27, 8, 29) {real, imag} */,
  {32'h410f8e1e, 32'hc1370c9c} /* (27, 8, 28) {real, imag} */,
  {32'hc1abe020, 32'hc148f104} /* (27, 8, 27) {real, imag} */,
  {32'hc0c8d23e, 32'hbe99a310} /* (27, 8, 26) {real, imag} */,
  {32'hc012005e, 32'hc14512d8} /* (27, 8, 25) {real, imag} */,
  {32'h40a3bfb7, 32'h414072d8} /* (27, 8, 24) {real, imag} */,
  {32'hc1390367, 32'hc13e830e} /* (27, 8, 23) {real, imag} */,
  {32'hc1876675, 32'hc04ccf44} /* (27, 8, 22) {real, imag} */,
  {32'h41481968, 32'h40d29627} /* (27, 8, 21) {real, imag} */,
  {32'h419d05d8, 32'hc1325e51} /* (27, 8, 20) {real, imag} */,
  {32'hbfd7a99f, 32'h40a4f782} /* (27, 8, 19) {real, imag} */,
  {32'hc0f27e90, 32'h407dec6f} /* (27, 8, 18) {real, imag} */,
  {32'h4105f180, 32'h4122f7e2} /* (27, 8, 17) {real, imag} */,
  {32'hbf55a6a0, 32'h3fe0e4e4} /* (27, 8, 16) {real, imag} */,
  {32'hc14de61a, 32'hc01654ba} /* (27, 8, 15) {real, imag} */,
  {32'hc115a0a0, 32'h418d1dce} /* (27, 8, 14) {real, imag} */,
  {32'h402ced20, 32'hbeb13930} /* (27, 8, 13) {real, imag} */,
  {32'h40be398a, 32'hc0c178c4} /* (27, 8, 12) {real, imag} */,
  {32'h418929a5, 32'h41424e7e} /* (27, 8, 11) {real, imag} */,
  {32'hc0267ba8, 32'hc1ad71d9} /* (27, 8, 10) {real, imag} */,
  {32'hc0e2b0da, 32'h3e2de280} /* (27, 8, 9) {real, imag} */,
  {32'hc10ab63c, 32'h3ffdf6e0} /* (27, 8, 8) {real, imag} */,
  {32'h41d4cc58, 32'h414cb8aa} /* (27, 8, 7) {real, imag} */,
  {32'hc16254e2, 32'hc0f5d222} /* (27, 8, 6) {real, imag} */,
  {32'h4116684c, 32'h419fa76a} /* (27, 8, 5) {real, imag} */,
  {32'hc1bd9314, 32'hc08971d7} /* (27, 8, 4) {real, imag} */,
  {32'h3f115460, 32'h4125c898} /* (27, 8, 3) {real, imag} */,
  {32'h40d01873, 32'h3ff79b60} /* (27, 8, 2) {real, imag} */,
  {32'hc1ce83cc, 32'hc16deb44} /* (27, 8, 1) {real, imag} */,
  {32'hc19d2840, 32'hc1081326} /* (27, 8, 0) {real, imag} */,
  {32'hc096fd6c, 32'h41a6946b} /* (27, 7, 31) {real, imag} */,
  {32'hc0663b04, 32'hc1a7f2e8} /* (27, 7, 30) {real, imag} */,
  {32'h40a54207, 32'h3fe918a5} /* (27, 7, 29) {real, imag} */,
  {32'hc1809cec, 32'hc194cf23} /* (27, 7, 28) {real, imag} */,
  {32'hc171542f, 32'hbf34f114} /* (27, 7, 27) {real, imag} */,
  {32'h41199720, 32'h4006b660} /* (27, 7, 26) {real, imag} */,
  {32'h3e8f2600, 32'h41a52522} /* (27, 7, 25) {real, imag} */,
  {32'hc0c59762, 32'h410510f9} /* (27, 7, 24) {real, imag} */,
  {32'h40116ea4, 32'h41787966} /* (27, 7, 23) {real, imag} */,
  {32'h41b37304, 32'hc126109f} /* (27, 7, 22) {real, imag} */,
  {32'h41ea6e13, 32'h40b75baa} /* (27, 7, 21) {real, imag} */,
  {32'hc1229f3d, 32'hbff93b08} /* (27, 7, 20) {real, imag} */,
  {32'h4145b795, 32'h40f2fd00} /* (27, 7, 19) {real, imag} */,
  {32'hc0eea909, 32'hc09c1046} /* (27, 7, 18) {real, imag} */,
  {32'hc12712ad, 32'hc10b232f} /* (27, 7, 17) {real, imag} */,
  {32'h418b3f1e, 32'h4100ab4d} /* (27, 7, 16) {real, imag} */,
  {32'h40aeffb7, 32'hc0e0b5f2} /* (27, 7, 15) {real, imag} */,
  {32'h411a993a, 32'h401ab95e} /* (27, 7, 14) {real, imag} */,
  {32'hc03f72a4, 32'hc0f728e0} /* (27, 7, 13) {real, imag} */,
  {32'h40a1d508, 32'h40433947} /* (27, 7, 12) {real, imag} */,
  {32'hc184fb42, 32'hc14b0d4d} /* (27, 7, 11) {real, imag} */,
  {32'h40883331, 32'h4167915d} /* (27, 7, 10) {real, imag} */,
  {32'h416edafe, 32'h40b98fa0} /* (27, 7, 9) {real, imag} */,
  {32'hc0f48170, 32'hc1256cbc} /* (27, 7, 8) {real, imag} */,
  {32'h4042be7e, 32'h3f29c564} /* (27, 7, 7) {real, imag} */,
  {32'h416ad942, 32'h4087d093} /* (27, 7, 6) {real, imag} */,
  {32'hc08a9d38, 32'hc0df83dc} /* (27, 7, 5) {real, imag} */,
  {32'h41492ff8, 32'hbfcd6d6e} /* (27, 7, 4) {real, imag} */,
  {32'h41884e1e, 32'hc000a54a} /* (27, 7, 3) {real, imag} */,
  {32'hc100fd82, 32'h4135baad} /* (27, 7, 2) {real, imag} */,
  {32'h41cde80b, 32'h413e775e} /* (27, 7, 1) {real, imag} */,
  {32'h41a10288, 32'hc15520ba} /* (27, 7, 0) {real, imag} */,
  {32'hc19d2f18, 32'hc0021646} /* (27, 6, 31) {real, imag} */,
  {32'hc0987bb3, 32'h401b9a10} /* (27, 6, 30) {real, imag} */,
  {32'h4179c22e, 32'hc108c7c0} /* (27, 6, 29) {real, imag} */,
  {32'h406a3b5c, 32'h4063e24e} /* (27, 6, 28) {real, imag} */,
  {32'h418388ae, 32'hbed6be50} /* (27, 6, 27) {real, imag} */,
  {32'h4142f739, 32'hc1ae63fe} /* (27, 6, 26) {real, imag} */,
  {32'hc0c6cf9a, 32'h40c8b9d2} /* (27, 6, 25) {real, imag} */,
  {32'hc11ed2bc, 32'hc0ce50cd} /* (27, 6, 24) {real, imag} */,
  {32'hc008924e, 32'hc0a9088c} /* (27, 6, 23) {real, imag} */,
  {32'h40fed69b, 32'hbe36ce20} /* (27, 6, 22) {real, imag} */,
  {32'h40e3a359, 32'h414ee442} /* (27, 6, 21) {real, imag} */,
  {32'hc1064031, 32'hc140714a} /* (27, 6, 20) {real, imag} */,
  {32'hc0855830, 32'hc1323663} /* (27, 6, 19) {real, imag} */,
  {32'h412ac7ee, 32'hbec2f100} /* (27, 6, 18) {real, imag} */,
  {32'h3e9a4610, 32'h40a894ec} /* (27, 6, 17) {real, imag} */,
  {32'hc0801044, 32'h41269c66} /* (27, 6, 16) {real, imag} */,
  {32'hc096725e, 32'hc1834f5e} /* (27, 6, 15) {real, imag} */,
  {32'hc0fe628b, 32'hc12a3c5b} /* (27, 6, 14) {real, imag} */,
  {32'h40bd97ee, 32'h4088c70e} /* (27, 6, 13) {real, imag} */,
  {32'hc044c442, 32'hc125c871} /* (27, 6, 12) {real, imag} */,
  {32'hc09a86a8, 32'h40cf2ee0} /* (27, 6, 11) {real, imag} */,
  {32'hc196a01e, 32'h40cb4284} /* (27, 6, 10) {real, imag} */,
  {32'hbf466a14, 32'hc026e71a} /* (27, 6, 9) {real, imag} */,
  {32'hc1cfe459, 32'h40fff674} /* (27, 6, 8) {real, imag} */,
  {32'h41200e0c, 32'hc09209d7} /* (27, 6, 7) {real, imag} */,
  {32'h3e8d50f0, 32'h40af6564} /* (27, 6, 6) {real, imag} */,
  {32'h40ad7e68, 32'h3f16f7c8} /* (27, 6, 5) {real, imag} */,
  {32'hc0b70dd0, 32'h3c581700} /* (27, 6, 4) {real, imag} */,
  {32'hbfbc99b0, 32'hc13bc695} /* (27, 6, 3) {real, imag} */,
  {32'h41d0a624, 32'hc0d23582} /* (27, 6, 2) {real, imag} */,
  {32'hc02dfe14, 32'hc1a57130} /* (27, 6, 1) {real, imag} */,
  {32'h40b5af1c, 32'hc1be8495} /* (27, 6, 0) {real, imag} */,
  {32'hc29fef84, 32'hc20af04b} /* (27, 5, 31) {real, imag} */,
  {32'h421b5eb8, 32'hc18bbabe} /* (27, 5, 30) {real, imag} */,
  {32'h40a67210, 32'hc0d30ea5} /* (27, 5, 29) {real, imag} */,
  {32'hc14237e1, 32'h42024c48} /* (27, 5, 28) {real, imag} */,
  {32'h41c9df62, 32'hc194b7b2} /* (27, 5, 27) {real, imag} */,
  {32'hbfe7b4c8, 32'hbfc0e1a8} /* (27, 5, 26) {real, imag} */,
  {32'h40c886c4, 32'h403fbf6a} /* (27, 5, 25) {real, imag} */,
  {32'hc0b2a3d4, 32'h41aa7853} /* (27, 5, 24) {real, imag} */,
  {32'hbee62460, 32'h4193db7a} /* (27, 5, 23) {real, imag} */,
  {32'hc027b7aa, 32'hc110f9b8} /* (27, 5, 22) {real, imag} */,
  {32'hc039d608, 32'hc096789c} /* (27, 5, 21) {real, imag} */,
  {32'h4134bb18, 32'hc1956e16} /* (27, 5, 20) {real, imag} */,
  {32'hc1a55147, 32'h40887ca9} /* (27, 5, 19) {real, imag} */,
  {32'h40f2a8cc, 32'hc1798082} /* (27, 5, 18) {real, imag} */,
  {32'hc098dda3, 32'h40367f37} /* (27, 5, 17) {real, imag} */,
  {32'h3ff26c78, 32'hbf765758} /* (27, 5, 16) {real, imag} */,
  {32'hc0fd9e44, 32'h410e523d} /* (27, 5, 15) {real, imag} */,
  {32'hc0e28b64, 32'h40ba13d0} /* (27, 5, 14) {real, imag} */,
  {32'h403deddc, 32'h407d825c} /* (27, 5, 13) {real, imag} */,
  {32'hc06847af, 32'hc18ca2c5} /* (27, 5, 12) {real, imag} */,
  {32'hc1416ad7, 32'hc1181a95} /* (27, 5, 11) {real, imag} */,
  {32'h41597fe0, 32'h400e5348} /* (27, 5, 10) {real, imag} */,
  {32'h404aa73a, 32'hc13fe0e8} /* (27, 5, 9) {real, imag} */,
  {32'hbffe3914, 32'h4072bafd} /* (27, 5, 8) {real, imag} */,
  {32'hc1655151, 32'hbfd06f30} /* (27, 5, 7) {real, imag} */,
  {32'h4138836a, 32'h4104c585} /* (27, 5, 6) {real, imag} */,
  {32'h41cd1ee8, 32'h410f1eb2} /* (27, 5, 5) {real, imag} */,
  {32'h4144d278, 32'h40e2403d} /* (27, 5, 4) {real, imag} */,
  {32'hbf4c2f50, 32'hc1c7fc55} /* (27, 5, 3) {real, imag} */,
  {32'h419fb4a0, 32'hc12efa44} /* (27, 5, 2) {real, imag} */,
  {32'hc25a1798, 32'hc20e8ee7} /* (27, 5, 1) {real, imag} */,
  {32'hc28feb59, 32'hc148c32b} /* (27, 5, 0) {real, imag} */,
  {32'h41a732f9, 32'h421a1c8a} /* (27, 4, 31) {real, imag} */,
  {32'hc255cf0f, 32'hc25ed96c} /* (27, 4, 30) {real, imag} */,
  {32'h405e9a15, 32'hc1831010} /* (27, 4, 29) {real, imag} */,
  {32'h3fce1194, 32'hc0f2622f} /* (27, 4, 28) {real, imag} */,
  {32'h413a01b6, 32'hc0d1a504} /* (27, 4, 27) {real, imag} */,
  {32'hbf8aef70, 32'h41da1ab0} /* (27, 4, 26) {real, imag} */,
  {32'hc17703d0, 32'hc13294b3} /* (27, 4, 25) {real, imag} */,
  {32'h40cdb023, 32'hc0185976} /* (27, 4, 24) {real, imag} */,
  {32'hc06c8c0b, 32'h4113aad8} /* (27, 4, 23) {real, imag} */,
  {32'h41ee405b, 32'hc10c89a5} /* (27, 4, 22) {real, imag} */,
  {32'hc181b231, 32'h410bb5a0} /* (27, 4, 21) {real, imag} */,
  {32'h4080a630, 32'hbfc8b968} /* (27, 4, 20) {real, imag} */,
  {32'hc0456931, 32'h413cbc25} /* (27, 4, 19) {real, imag} */,
  {32'hbe5947c0, 32'hc0e7ec8a} /* (27, 4, 18) {real, imag} */,
  {32'h408cd94e, 32'hc01bc627} /* (27, 4, 17) {real, imag} */,
  {32'h3fdf4456, 32'hc080512e} /* (27, 4, 16) {real, imag} */,
  {32'hc08d67d3, 32'h409d99a1} /* (27, 4, 15) {real, imag} */,
  {32'hc144270c, 32'h40ce4517} /* (27, 4, 14) {real, imag} */,
  {32'h40be8789, 32'h41324175} /* (27, 4, 13) {real, imag} */,
  {32'hbfd2a578, 32'hc12e5a12} /* (27, 4, 12) {real, imag} */,
  {32'hc1adde9c, 32'h4125efe1} /* (27, 4, 11) {real, imag} */,
  {32'hc0c30bf0, 32'h4100a57e} /* (27, 4, 10) {real, imag} */,
  {32'h40263342, 32'hc11a8b7e} /* (27, 4, 9) {real, imag} */,
  {32'hc13351e2, 32'h40f245e2} /* (27, 4, 8) {real, imag} */,
  {32'h40ef767e, 32'h41301302} /* (27, 4, 7) {real, imag} */,
  {32'hc149695b, 32'h3f310b48} /* (27, 4, 6) {real, imag} */,
  {32'hc020e50c, 32'hc1c530cf} /* (27, 4, 5) {real, imag} */,
  {32'h4258aefe, 32'hc0d24ab0} /* (27, 4, 4) {real, imag} */,
  {32'h41b2c8af, 32'hc0a42fba} /* (27, 4, 3) {real, imag} */,
  {32'hc24a82ad, 32'hc294c728} /* (27, 4, 2) {real, imag} */,
  {32'h42b881f6, 32'h42aadb38} /* (27, 4, 1) {real, imag} */,
  {32'h40697564, 32'h40e1ba87} /* (27, 4, 0) {real, imag} */,
  {32'hc2d3fafa, 32'h41bd7322} /* (27, 3, 31) {real, imag} */,
  {32'h429e489b, 32'hc28c9735} /* (27, 3, 30) {real, imag} */,
  {32'hc15e59b8, 32'h4030fc20} /* (27, 3, 29) {real, imag} */,
  {32'h41be1560, 32'h41803889} /* (27, 3, 28) {real, imag} */,
  {32'hc191d7a0, 32'hc1a10e02} /* (27, 3, 27) {real, imag} */,
  {32'h412fb106, 32'h41b50600} /* (27, 3, 26) {real, imag} */,
  {32'h4170100a, 32'h40a21a1b} /* (27, 3, 25) {real, imag} */,
  {32'hc1dd36f2, 32'hc1760dec} /* (27, 3, 24) {real, imag} */,
  {32'h414b6aba, 32'h41303d49} /* (27, 3, 23) {real, imag} */,
  {32'h419c31b4, 32'h41530580} /* (27, 3, 22) {real, imag} */,
  {32'hc0095674, 32'h412c2759} /* (27, 3, 21) {real, imag} */,
  {32'hc0ad0f9e, 32'hc1c00362} /* (27, 3, 20) {real, imag} */,
  {32'hbfc90cee, 32'h40fecc16} /* (27, 3, 19) {real, imag} */,
  {32'h3fa4de4a, 32'hbf5cf09c} /* (27, 3, 18) {real, imag} */,
  {32'hc10ebf6e, 32'hc1466ba6} /* (27, 3, 17) {real, imag} */,
  {32'h40ad2138, 32'hc11748c6} /* (27, 3, 16) {real, imag} */,
  {32'h4013461c, 32'h4063caee} /* (27, 3, 15) {real, imag} */,
  {32'hc094ea3a, 32'h408d50fe} /* (27, 3, 14) {real, imag} */,
  {32'h401c88a8, 32'h4017533e} /* (27, 3, 13) {real, imag} */,
  {32'h3faebc9c, 32'hc1d8b63c} /* (27, 3, 12) {real, imag} */,
  {32'h41526b56, 32'hc0691f9e} /* (27, 3, 11) {real, imag} */,
  {32'hc1495b6c, 32'hc1188ab9} /* (27, 3, 10) {real, imag} */,
  {32'h4149c73a, 32'h419171e1} /* (27, 3, 9) {real, imag} */,
  {32'hc135d000, 32'h3deec340} /* (27, 3, 8) {real, imag} */,
  {32'h40abba19, 32'h414cc0e3} /* (27, 3, 7) {real, imag} */,
  {32'hc1ecf93a, 32'hc0a967a6} /* (27, 3, 6) {real, imag} */,
  {32'h41233c8c, 32'h4032b51a} /* (27, 3, 5) {real, imag} */,
  {32'hbfc35610, 32'h41f63c0a} /* (27, 3, 4) {real, imag} */,
  {32'hc069513e, 32'h4107f9b4} /* (27, 3, 3) {real, imag} */,
  {32'hbfc388a0, 32'hc2a5c636} /* (27, 3, 2) {real, imag} */,
  {32'h425c4ef9, 32'h42e695fb} /* (27, 3, 1) {real, imag} */,
  {32'h425e5ea8, 32'h411ca644} /* (27, 3, 0) {real, imag} */,
  {32'hc3db2dce, 32'h423d744f} /* (27, 2, 31) {real, imag} */,
  {32'h439da3ec, 32'hc2e59e92} /* (27, 2, 30) {real, imag} */,
  {32'hc1b458b2, 32'h3f9d2510} /* (27, 2, 29) {real, imag} */,
  {32'hc19e34d9, 32'h42a75e12} /* (27, 2, 28) {real, imag} */,
  {32'h420615a2, 32'hc22dbd5b} /* (27, 2, 27) {real, imag} */,
  {32'h4104fa0c, 32'hc0e894fb} /* (27, 2, 26) {real, imag} */,
  {32'hbfde9688, 32'h42018f7b} /* (27, 2, 25) {real, imag} */,
  {32'h4162d8ce, 32'hc19d7c5a} /* (27, 2, 24) {real, imag} */,
  {32'h416cfb96, 32'h4033add3} /* (27, 2, 23) {real, imag} */,
  {32'hc1001b4f, 32'hc137e102} /* (27, 2, 22) {real, imag} */,
  {32'h3feadc14, 32'hc0d81515} /* (27, 2, 21) {real, imag} */,
  {32'h411c30e8, 32'h40c9bfb0} /* (27, 2, 20) {real, imag} */,
  {32'hc0378b54, 32'hc01c10a8} /* (27, 2, 19) {real, imag} */,
  {32'h41231dcf, 32'hc110e1da} /* (27, 2, 18) {real, imag} */,
  {32'h4180a813, 32'h40fd52f0} /* (27, 2, 17) {real, imag} */,
  {32'hc108eb1d, 32'hbf8bdd5c} /* (27, 2, 16) {real, imag} */,
  {32'h3f802f60, 32'h3dcaf2e0} /* (27, 2, 15) {real, imag} */,
  {32'h409c1d65, 32'hbf905c88} /* (27, 2, 14) {real, imag} */,
  {32'h3f7ffe46, 32'hc13d37d2} /* (27, 2, 13) {real, imag} */,
  {32'hc166fa1c, 32'h4099587e} /* (27, 2, 12) {real, imag} */,
  {32'hc12115d8, 32'h41b18e1e} /* (27, 2, 11) {real, imag} */,
  {32'hc126da20, 32'hc187c0b5} /* (27, 2, 10) {real, imag} */,
  {32'h40b30e99, 32'h3f979090} /* (27, 2, 9) {real, imag} */,
  {32'h419939e4, 32'h41be9ff9} /* (27, 2, 8) {real, imag} */,
  {32'hc1047546, 32'hc05c2ea0} /* (27, 2, 7) {real, imag} */,
  {32'hbfa4b296, 32'hc0867122} /* (27, 2, 6) {real, imag} */,
  {32'h41dc2f2b, 32'h4214c5a7} /* (27, 2, 5) {real, imag} */,
  {32'hc288be87, 32'hc25c77a4} /* (27, 2, 4) {real, imag} */,
  {32'h400c2e84, 32'hc16fbccf} /* (27, 2, 3) {real, imag} */,
  {32'h438100c2, 32'hc2d63fb4} /* (27, 2, 2) {real, imag} */,
  {32'hc38244db, 32'h42eb4504} /* (27, 2, 1) {real, imag} */,
  {32'hc34e7eff, 32'hc2d9d8f0} /* (27, 2, 0) {real, imag} */,
  {32'h439803d0, 32'hc2fc004e} /* (27, 1, 31) {real, imag} */,
  {32'hc32180c4, 32'h42862957} /* (27, 1, 30) {real, imag} */,
  {32'h40c1b018, 32'h40c5ff42} /* (27, 1, 29) {real, imag} */,
  {32'h41418f7f, 32'h41ed56af} /* (27, 1, 28) {real, imag} */,
  {32'hc2c9c86f, 32'h40f4bf50} /* (27, 1, 27) {real, imag} */,
  {32'hc125eea1, 32'hc18ea87b} /* (27, 1, 26) {real, imag} */,
  {32'h4119fb76, 32'h41357ac6} /* (27, 1, 25) {real, imag} */,
  {32'h3fbb9ab8, 32'h413ad6a3} /* (27, 1, 24) {real, imag} */,
  {32'hc0f35c0a, 32'hc19dab4e} /* (27, 1, 23) {real, imag} */,
  {32'hc051c792, 32'hc090aebb} /* (27, 1, 22) {real, imag} */,
  {32'hc2016acc, 32'h411163da} /* (27, 1, 21) {real, imag} */,
  {32'hc044237e, 32'h41ad64e8} /* (27, 1, 20) {real, imag} */,
  {32'h3fbe4c1e, 32'hc1857a26} /* (27, 1, 19) {real, imag} */,
  {32'h413bf42a, 32'h40f50aae} /* (27, 1, 18) {real, imag} */,
  {32'hbf14e0e8, 32'h408538c1} /* (27, 1, 17) {real, imag} */,
  {32'hc084dd01, 32'hc085ad3f} /* (27, 1, 16) {real, imag} */,
  {32'hc11017c2, 32'h416fa48c} /* (27, 1, 15) {real, imag} */,
  {32'h4153acdd, 32'hc171b2f5} /* (27, 1, 14) {real, imag} */,
  {32'h418823dd, 32'hbf90da8c} /* (27, 1, 13) {real, imag} */,
  {32'hc13213de, 32'h3feb1ff4} /* (27, 1, 12) {real, imag} */,
  {32'hc18df652, 32'hc14de1ac} /* (27, 1, 11) {real, imag} */,
  {32'hbf044ed0, 32'h41b2fc27} /* (27, 1, 10) {real, imag} */,
  {32'hc1b191f8, 32'hc1574fff} /* (27, 1, 9) {real, imag} */,
  {32'hc15b6946, 32'hc1fc1033} /* (27, 1, 8) {real, imag} */,
  {32'hc19960fd, 32'h410c7ef0} /* (27, 1, 7) {real, imag} */,
  {32'hc0c6a3e6, 32'hc141f8f7} /* (27, 1, 6) {real, imag} */,
  {32'hc2628a12, 32'hc1e1ba4d} /* (27, 1, 5) {real, imag} */,
  {32'h41f7485f, 32'h419830e3} /* (27, 1, 4) {real, imag} */,
  {32'hc242ca0c, 32'hc11fcc40} /* (27, 1, 3) {real, imag} */,
  {32'hc38eb0ba, 32'hc38aeec8} /* (27, 1, 2) {real, imag} */,
  {32'h43d0e7c2, 32'h43324765} /* (27, 1, 1) {real, imag} */,
  {32'h4303ac36, 32'hc0997190} /* (27, 1, 0) {real, imag} */,
  {32'hc222ca40, 32'h41f603d8} /* (27, 0, 31) {real, imag} */,
  {32'hc29db0b6, 32'h433591de} /* (27, 0, 30) {real, imag} */,
  {32'hc120984c, 32'hc23b3c02} /* (27, 0, 29) {real, imag} */,
  {32'h4202a9ba, 32'h41a85bdc} /* (27, 0, 28) {real, imag} */,
  {32'hc26a827e, 32'h4202a4ca} /* (27, 0, 27) {real, imag} */,
  {32'h41b15af5, 32'h40973e8e} /* (27, 0, 26) {real, imag} */,
  {32'h41978ccf, 32'hc2147a70} /* (27, 0, 25) {real, imag} */,
  {32'hc0b00df0, 32'h421a87bc} /* (27, 0, 24) {real, imag} */,
  {32'hc14ba551, 32'hbfb7a948} /* (27, 0, 23) {real, imag} */,
  {32'hc1493bda, 32'h41558b32} /* (27, 0, 22) {real, imag} */,
  {32'h40472106, 32'h4125794e} /* (27, 0, 21) {real, imag} */,
  {32'h410588f8, 32'h3fd55a2c} /* (27, 0, 20) {real, imag} */,
  {32'h40bbcdfd, 32'hc042d058} /* (27, 0, 19) {real, imag} */,
  {32'h41573f26, 32'h40d5ec14} /* (27, 0, 18) {real, imag} */,
  {32'h40dd1e78, 32'hbfb1b466} /* (27, 0, 17) {real, imag} */,
  {32'hc12fdd7c, 32'h00000000} /* (27, 0, 16) {real, imag} */,
  {32'h40dd1e78, 32'h3fb1b466} /* (27, 0, 15) {real, imag} */,
  {32'h41573f26, 32'hc0d5ec14} /* (27, 0, 14) {real, imag} */,
  {32'h40bbcdfd, 32'h4042d058} /* (27, 0, 13) {real, imag} */,
  {32'h410588f8, 32'hbfd55a2c} /* (27, 0, 12) {real, imag} */,
  {32'h40472106, 32'hc125794e} /* (27, 0, 11) {real, imag} */,
  {32'hc1493bda, 32'hc1558b32} /* (27, 0, 10) {real, imag} */,
  {32'hc14ba551, 32'h3fb7a948} /* (27, 0, 9) {real, imag} */,
  {32'hc0b00df0, 32'hc21a87bc} /* (27, 0, 8) {real, imag} */,
  {32'h41978ccf, 32'h42147a70} /* (27, 0, 7) {real, imag} */,
  {32'h41b15af5, 32'hc0973e8e} /* (27, 0, 6) {real, imag} */,
  {32'hc26a827e, 32'hc202a4ca} /* (27, 0, 5) {real, imag} */,
  {32'h4202a9ba, 32'hc1a85bdc} /* (27, 0, 4) {real, imag} */,
  {32'hc120984c, 32'h423b3c02} /* (27, 0, 3) {real, imag} */,
  {32'hc29db0b6, 32'hc33591de} /* (27, 0, 2) {real, imag} */,
  {32'hc222ca40, 32'hc1f603d8} /* (27, 0, 1) {real, imag} */,
  {32'hc3d271ac, 32'h00000000} /* (27, 0, 0) {real, imag} */,
  {32'hc3910940, 32'h435c801d} /* (26, 31, 31) {real, imag} */,
  {32'hc1fce798, 32'h420169f4} /* (26, 31, 30) {real, imag} */,
  {32'h3e67c600, 32'h41b30c6c} /* (26, 31, 29) {real, imag} */,
  {32'hc192dc72, 32'h4180c656} /* (26, 31, 28) {real, imag} */,
  {32'h3fef3620, 32'hc1247a2e} /* (26, 31, 27) {real, imag} */,
  {32'h416f0c36, 32'h402ae662} /* (26, 31, 26) {real, imag} */,
  {32'h41369168, 32'hc1a6c130} /* (26, 31, 25) {real, imag} */,
  {32'hc12b1098, 32'h419a6005} /* (26, 31, 24) {real, imag} */,
  {32'hc1ae7514, 32'hbf943fe0} /* (26, 31, 23) {real, imag} */,
  {32'hc1dccbee, 32'hbec83278} /* (26, 31, 22) {real, imag} */,
  {32'hc19d1598, 32'hbf832e10} /* (26, 31, 21) {real, imag} */,
  {32'h410907c2, 32'hc14a5faa} /* (26, 31, 20) {real, imag} */,
  {32'h41d95d35, 32'hc0929d18} /* (26, 31, 19) {real, imag} */,
  {32'h407e397a, 32'h40a3ba98} /* (26, 31, 18) {real, imag} */,
  {32'hbde4a4c0, 32'h3f880bcc} /* (26, 31, 17) {real, imag} */,
  {32'hc0ff199a, 32'h3fea115d} /* (26, 31, 16) {real, imag} */,
  {32'h4083bd20, 32'h40fc0667} /* (26, 31, 15) {real, imag} */,
  {32'h41303ef8, 32'hbfb5c9a4} /* (26, 31, 14) {real, imag} */,
  {32'h41850d11, 32'h40be3764} /* (26, 31, 13) {real, imag} */,
  {32'h4139e5a6, 32'hc188db82} /* (26, 31, 12) {real, imag} */,
  {32'hbfe5da08, 32'h41355303} /* (26, 31, 11) {real, imag} */,
  {32'h40013678, 32'hc0a848ee} /* (26, 31, 10) {real, imag} */,
  {32'h410e2b92, 32'hbe7921c0} /* (26, 31, 9) {real, imag} */,
  {32'h41057d44, 32'h408516f1} /* (26, 31, 8) {real, imag} */,
  {32'hc0cce52e, 32'h4128f8e9} /* (26, 31, 7) {real, imag} */,
  {32'hc1d60d2d, 32'h4101b218} /* (26, 31, 6) {real, imag} */,
  {32'hc1947850, 32'h3e416300} /* (26, 31, 5) {real, imag} */,
  {32'hc169817a, 32'hc1941052} /* (26, 31, 4) {real, imag} */,
  {32'h40e986d4, 32'h3fc90a00} /* (26, 31, 3) {real, imag} */,
  {32'h417a1570, 32'hc2d8bf26} /* (26, 31, 2) {real, imag} */,
  {32'hc356de14, 32'hc00695e0} /* (26, 31, 1) {real, imag} */,
  {32'hc3e8fd6c, 32'h42d3370a} /* (26, 31, 0) {real, imag} */,
  {32'h40b59680, 32'hc288b118} /* (26, 30, 31) {real, imag} */,
  {32'h42861f12, 32'h41dc8ee8} /* (26, 30, 30) {real, imag} */,
  {32'hc1f537d2, 32'h4135a3bb} /* (26, 30, 29) {real, imag} */,
  {32'hc1914d0c, 32'h4214c973} /* (26, 30, 28) {real, imag} */,
  {32'hc193011d, 32'hc22263f2} /* (26, 30, 27) {real, imag} */,
  {32'h41609cbe, 32'hc0c3c967} /* (26, 30, 26) {real, imag} */,
  {32'h40cef612, 32'hc1c366d6} /* (26, 30, 25) {real, imag} */,
  {32'hc0945796, 32'hc1a8f5c5} /* (26, 30, 24) {real, imag} */,
  {32'hc194259f, 32'h4152f550} /* (26, 30, 23) {real, imag} */,
  {32'h3edb00b0, 32'hc019b554} /* (26, 30, 22) {real, imag} */,
  {32'h415ede48, 32'hc10115e9} /* (26, 30, 21) {real, imag} */,
  {32'h40b793f8, 32'hc0079494} /* (26, 30, 20) {real, imag} */,
  {32'hc06fe79e, 32'hbff90ac2} /* (26, 30, 19) {real, imag} */,
  {32'hc0826a38, 32'h40eaaffa} /* (26, 30, 18) {real, imag} */,
  {32'hbf6ed506, 32'h40c48894} /* (26, 30, 17) {real, imag} */,
  {32'h401e675e, 32'hc0b9f76d} /* (26, 30, 16) {real, imag} */,
  {32'h411aa0ae, 32'hc0fdfd77} /* (26, 30, 15) {real, imag} */,
  {32'h411b1964, 32'hc140c8cf} /* (26, 30, 14) {real, imag} */,
  {32'hc0f66dda, 32'h3f8b2cb8} /* (26, 30, 13) {real, imag} */,
  {32'hc0f0bd3f, 32'h3ef38940} /* (26, 30, 12) {real, imag} */,
  {32'h40839c7c, 32'hbfbffd80} /* (26, 30, 11) {real, imag} */,
  {32'hc1406eb2, 32'h4036331e} /* (26, 30, 10) {real, imag} */,
  {32'h41e5fcf9, 32'h416ee2d3} /* (26, 30, 9) {real, imag} */,
  {32'h41aafec6, 32'hc128d31d} /* (26, 30, 8) {real, imag} */,
  {32'hc0bffe56, 32'hc221b930} /* (26, 30, 7) {real, imag} */,
  {32'h40b4bb75, 32'hc15f0e50} /* (26, 30, 6) {real, imag} */,
  {32'h41eb715f, 32'h41bef157} /* (26, 30, 5) {real, imag} */,
  {32'hc141df94, 32'hc133531a} /* (26, 30, 4) {real, imag} */,
  {32'hc134a8ec, 32'h40e8e93e} /* (26, 30, 3) {real, imag} */,
  {32'h4262fe10, 32'h427918f2} /* (26, 30, 2) {real, imag} */,
  {32'h41b5c9e0, 32'hc27760bc} /* (26, 30, 1) {real, imag} */,
  {32'h4253d7cc, 32'h428b7808} /* (26, 30, 0) {real, imag} */,
  {32'hc0603680, 32'hc294a578} /* (26, 29, 31) {real, imag} */,
  {32'h41d2df75, 32'h40f5bf94} /* (26, 29, 30) {real, imag} */,
  {32'hc1829350, 32'h3f5002e0} /* (26, 29, 29) {real, imag} */,
  {32'hc0befcea, 32'hc164205d} /* (26, 29, 28) {real, imag} */,
  {32'hc1703418, 32'hc159f036} /* (26, 29, 27) {real, imag} */,
  {32'hc168f290, 32'hc15bf076} /* (26, 29, 26) {real, imag} */,
  {32'hc076243c, 32'hc16a9a5a} /* (26, 29, 25) {real, imag} */,
  {32'hc0eee221, 32'h414d4281} /* (26, 29, 24) {real, imag} */,
  {32'hc08c4b2c, 32'h40fe9390} /* (26, 29, 23) {real, imag} */,
  {32'hc108d650, 32'h4044720a} /* (26, 29, 22) {real, imag} */,
  {32'h40001bc2, 32'h40a36302} /* (26, 29, 21) {real, imag} */,
  {32'h40fe260e, 32'h41172ce0} /* (26, 29, 20) {real, imag} */,
  {32'h41211535, 32'h418d7278} /* (26, 29, 19) {real, imag} */,
  {32'h404c7684, 32'hc18498f4} /* (26, 29, 18) {real, imag} */,
  {32'hc090ab61, 32'h40ce1dc2} /* (26, 29, 17) {real, imag} */,
  {32'h40876e9e, 32'hc10184ef} /* (26, 29, 16) {real, imag} */,
  {32'h419344da, 32'hc0d2d840} /* (26, 29, 15) {real, imag} */,
  {32'hc128e9d6, 32'h419d1ad3} /* (26, 29, 14) {real, imag} */,
  {32'h4143a574, 32'h40cc9c4c} /* (26, 29, 13) {real, imag} */,
  {32'hc137af6a, 32'h4073e51a} /* (26, 29, 12) {real, imag} */,
  {32'h3f1af8c0, 32'hc0a9174a} /* (26, 29, 11) {real, imag} */,
  {32'hc003b432, 32'hc0abd33f} /* (26, 29, 10) {real, imag} */,
  {32'h40c392fb, 32'h411680ba} /* (26, 29, 9) {real, imag} */,
  {32'hc0e0c97e, 32'h413a0988} /* (26, 29, 8) {real, imag} */,
  {32'hc1af19f9, 32'hbf8f2c90} /* (26, 29, 7) {real, imag} */,
  {32'hc1294fdf, 32'hc15d9480} /* (26, 29, 6) {real, imag} */,
  {32'hc016b900, 32'h40f044af} /* (26, 29, 5) {real, imag} */,
  {32'h419f5ad8, 32'hc18a913f} /* (26, 29, 4) {real, imag} */,
  {32'h412bdac1, 32'hc004177e} /* (26, 29, 3) {real, imag} */,
  {32'h42490e17, 32'h415f3e10} /* (26, 29, 2) {real, imag} */,
  {32'hc1d7bc14, 32'hc0917fc8} /* (26, 29, 1) {real, imag} */,
  {32'h429e92db, 32'hc1fd20d5} /* (26, 29, 0) {real, imag} */,
  {32'h41580fc8, 32'hc135c77a} /* (26, 28, 31) {real, imag} */,
  {32'hc1673dec, 32'h4088d008} /* (26, 28, 30) {real, imag} */,
  {32'hc04716f6, 32'h408587e6} /* (26, 28, 29) {real, imag} */,
  {32'h41ae8843, 32'h41e872be} /* (26, 28, 28) {real, imag} */,
  {32'h415aaf09, 32'h3fafaf24} /* (26, 28, 27) {real, imag} */,
  {32'hc1978266, 32'hc11c6e08} /* (26, 28, 26) {real, imag} */,
  {32'hc020d54c, 32'hc14a25f4} /* (26, 28, 25) {real, imag} */,
  {32'h400c760c, 32'h41108507} /* (26, 28, 24) {real, imag} */,
  {32'hc0ba6adf, 32'hc046e62c} /* (26, 28, 23) {real, imag} */,
  {32'h40856319, 32'h40a61476} /* (26, 28, 22) {real, imag} */,
  {32'h41a55f87, 32'hc1192c14} /* (26, 28, 21) {real, imag} */,
  {32'hc13ca03f, 32'h4117b227} /* (26, 28, 20) {real, imag} */,
  {32'h4044e50e, 32'hc1386426} /* (26, 28, 19) {real, imag} */,
  {32'hc1035352, 32'hbfbcd410} /* (26, 28, 18) {real, imag} */,
  {32'hc1750474, 32'h40858686} /* (26, 28, 17) {real, imag} */,
  {32'hc095c904, 32'h3fbce1d4} /* (26, 28, 16) {real, imag} */,
  {32'h40b946b8, 32'h3fc985fc} /* (26, 28, 15) {real, imag} */,
  {32'hc19eec98, 32'h41103573} /* (26, 28, 14) {real, imag} */,
  {32'hbed4757e, 32'h40cb3a8b} /* (26, 28, 13) {real, imag} */,
  {32'h40a03a5c, 32'hc01e0994} /* (26, 28, 12) {real, imag} */,
  {32'hc0a71056, 32'hc1a2e4f0} /* (26, 28, 11) {real, imag} */,
  {32'h41bacb31, 32'hc10cd3cf} /* (26, 28, 10) {real, imag} */,
  {32'hbdbba040, 32'hc10e73ad} /* (26, 28, 9) {real, imag} */,
  {32'h4035ab34, 32'h41327150} /* (26, 28, 8) {real, imag} */,
  {32'hbfbbdcce, 32'hc216858b} /* (26, 28, 7) {real, imag} */,
  {32'hc1c05772, 32'h415577c5} /* (26, 28, 6) {real, imag} */,
  {32'h3f7b8754, 32'hc08909d3} /* (26, 28, 5) {real, imag} */,
  {32'h3f3463f0, 32'h412af775} /* (26, 28, 4) {real, imag} */,
  {32'hc1c4089d, 32'hc022a804} /* (26, 28, 3) {real, imag} */,
  {32'hc135daee, 32'h408d1a58} /* (26, 28, 2) {real, imag} */,
  {32'hc145a5e2, 32'h40069b28} /* (26, 28, 1) {real, imag} */,
  {32'hc1ac42ca, 32'h41fc5812} /* (26, 28, 0) {real, imag} */,
  {32'hc20a3bc1, 32'hc1224b98} /* (26, 27, 31) {real, imag} */,
  {32'hc19275bd, 32'h41367f6a} /* (26, 27, 30) {real, imag} */,
  {32'hc1661926, 32'h41baee14} /* (26, 27, 29) {real, imag} */,
  {32'hc0714a65, 32'h4100f6d3} /* (26, 27, 28) {real, imag} */,
  {32'h4179b22f, 32'hbfb681c0} /* (26, 27, 27) {real, imag} */,
  {32'hc1bb1a1a, 32'hc161ca44} /* (26, 27, 26) {real, imag} */,
  {32'h419a4e22, 32'hc16ad4a6} /* (26, 27, 25) {real, imag} */,
  {32'h41d3f6e6, 32'h40db83d6} /* (26, 27, 24) {real, imag} */,
  {32'h413be2b8, 32'h3f02f2b0} /* (26, 27, 23) {real, imag} */,
  {32'h411af272, 32'hc06562d2} /* (26, 27, 22) {real, imag} */,
  {32'h405e159d, 32'hc18b5dbe} /* (26, 27, 21) {real, imag} */,
  {32'hc0886714, 32'hbf391f70} /* (26, 27, 20) {real, imag} */,
  {32'hc138e9fa, 32'hc1744ae4} /* (26, 27, 19) {real, imag} */,
  {32'hc084cea8, 32'h3ef32e20} /* (26, 27, 18) {real, imag} */,
  {32'hc059c69c, 32'hc00683e4} /* (26, 27, 17) {real, imag} */,
  {32'hc1434b38, 32'h417b725a} /* (26, 27, 16) {real, imag} */,
  {32'h3f95362c, 32'h410950ce} /* (26, 27, 15) {real, imag} */,
  {32'h40db013e, 32'h412715ae} /* (26, 27, 14) {real, imag} */,
  {32'h410ab40e, 32'hc17ecbca} /* (26, 27, 13) {real, imag} */,
  {32'h419e6ae0, 32'hc09c0209} /* (26, 27, 12) {real, imag} */,
  {32'h405bec2a, 32'h414e430a} /* (26, 27, 11) {real, imag} */,
  {32'h416173d6, 32'h3da24080} /* (26, 27, 10) {real, imag} */,
  {32'hc1580ee4, 32'hc158e888} /* (26, 27, 9) {real, imag} */,
  {32'h3ff8d904, 32'h40ab74c9} /* (26, 27, 8) {real, imag} */,
  {32'h3fd23fa2, 32'h41311360} /* (26, 27, 7) {real, imag} */,
  {32'h40867d77, 32'h3f9902e2} /* (26, 27, 6) {real, imag} */,
  {32'hc175a32e, 32'h4122b9dc} /* (26, 27, 5) {real, imag} */,
  {32'hc13bbcf3, 32'hc1ae4bd0} /* (26, 27, 4) {real, imag} */,
  {32'h41d7bcd2, 32'hc004fff4} /* (26, 27, 3) {real, imag} */,
  {32'h418ed5a4, 32'h4124b4dc} /* (26, 27, 2) {real, imag} */,
  {32'hc0594940, 32'h421dd99e} /* (26, 27, 1) {real, imag} */,
  {32'hc2569100, 32'hc1a4f675} /* (26, 27, 0) {real, imag} */,
  {32'hc0c004ec, 32'hc1057943} /* (26, 26, 31) {real, imag} */,
  {32'h410e4984, 32'hc000b062} /* (26, 26, 30) {real, imag} */,
  {32'h41a137d9, 32'h41620997} /* (26, 26, 29) {real, imag} */,
  {32'hc0c36798, 32'h41614baa} /* (26, 26, 28) {real, imag} */,
  {32'h3f9778f8, 32'hc158a6c5} /* (26, 26, 27) {real, imag} */,
  {32'h41908912, 32'h4181811d} /* (26, 26, 26) {real, imag} */,
  {32'h412518f8, 32'hbf93e8c0} /* (26, 26, 25) {real, imag} */,
  {32'h418e19d2, 32'hc1238252} /* (26, 26, 24) {real, imag} */,
  {32'h41a2bcbd, 32'h415876c0} /* (26, 26, 23) {real, imag} */,
  {32'hc09d473b, 32'hbffeb7f8} /* (26, 26, 22) {real, imag} */,
  {32'h4178b646, 32'h40927c61} /* (26, 26, 21) {real, imag} */,
  {32'hc15b3124, 32'hc1531ff6} /* (26, 26, 20) {real, imag} */,
  {32'h414af7d5, 32'h414b920b} /* (26, 26, 19) {real, imag} */,
  {32'h408e04ee, 32'h3e7fcf08} /* (26, 26, 18) {real, imag} */,
  {32'h40c6ad99, 32'hc08c0473} /* (26, 26, 17) {real, imag} */,
  {32'h40d82811, 32'hc0258bd4} /* (26, 26, 16) {real, imag} */,
  {32'hc10e9852, 32'h4155e600} /* (26, 26, 15) {real, imag} */,
  {32'h40401351, 32'hc12ecd0c} /* (26, 26, 14) {real, imag} */,
  {32'hc0ef3dc3, 32'h4136cda9} /* (26, 26, 13) {real, imag} */,
  {32'h4110852e, 32'hc0e04f39} /* (26, 26, 12) {real, imag} */,
  {32'h40aa9500, 32'h4037bd48} /* (26, 26, 11) {real, imag} */,
  {32'h418a8a17, 32'hc11c2d76} /* (26, 26, 10) {real, imag} */,
  {32'h3f62ac38, 32'h403b0c4a} /* (26, 26, 9) {real, imag} */,
  {32'h40e9228a, 32'hc1fcf696} /* (26, 26, 8) {real, imag} */,
  {32'hc155871f, 32'h41497a98} /* (26, 26, 7) {real, imag} */,
  {32'h3ff6b1a8, 32'hc1ad71cd} /* (26, 26, 6) {real, imag} */,
  {32'hbfd9ea4c, 32'hbfb8ed48} /* (26, 26, 5) {real, imag} */,
  {32'h41356916, 32'h416319dd} /* (26, 26, 4) {real, imag} */,
  {32'hc011ce2a, 32'hc09b32d6} /* (26, 26, 3) {real, imag} */,
  {32'hc1af530d, 32'hc017ec3c} /* (26, 26, 2) {real, imag} */,
  {32'hc156d6fe, 32'hc02291d0} /* (26, 26, 1) {real, imag} */,
  {32'h41562ce8, 32'h417b96c0} /* (26, 26, 0) {real, imag} */,
  {32'h42019004, 32'hc1011cea} /* (26, 25, 31) {real, imag} */,
  {32'h4127aad6, 32'hc1a4ae94} /* (26, 25, 30) {real, imag} */,
  {32'h41b61906, 32'h40815854} /* (26, 25, 29) {real, imag} */,
  {32'h41111ffa, 32'h420d3dca} /* (26, 25, 28) {real, imag} */,
  {32'hc1316552, 32'h418c6381} /* (26, 25, 27) {real, imag} */,
  {32'h41a3e214, 32'hc1652827} /* (26, 25, 26) {real, imag} */,
  {32'hc1210d75, 32'h41093c50} /* (26, 25, 25) {real, imag} */,
  {32'h411baaf6, 32'h419c95f7} /* (26, 25, 24) {real, imag} */,
  {32'h41715f48, 32'hc13859de} /* (26, 25, 23) {real, imag} */,
  {32'hc1d5f7ba, 32'h4148deb6} /* (26, 25, 22) {real, imag} */,
  {32'hc0ca93f0, 32'hc180c998} /* (26, 25, 21) {real, imag} */,
  {32'h3f2d3028, 32'h410aeb84} /* (26, 25, 20) {real, imag} */,
  {32'hc0945503, 32'h3fee6d0a} /* (26, 25, 19) {real, imag} */,
  {32'hc18daa64, 32'h3fe6ab3b} /* (26, 25, 18) {real, imag} */,
  {32'h400bc6b4, 32'hbf94ae44} /* (26, 25, 17) {real, imag} */,
  {32'hc1266cd6, 32'h4039db67} /* (26, 25, 16) {real, imag} */,
  {32'hc02c6782, 32'hbf828cae} /* (26, 25, 15) {real, imag} */,
  {32'hc14e3674, 32'hc1104ae8} /* (26, 25, 14) {real, imag} */,
  {32'hc1039bfe, 32'hc1233ede} /* (26, 25, 13) {real, imag} */,
  {32'h41a1a452, 32'hc138a6ea} /* (26, 25, 12) {real, imag} */,
  {32'h3ed97660, 32'h419b5a6c} /* (26, 25, 11) {real, imag} */,
  {32'hbfccaf44, 32'hc1858e57} /* (26, 25, 10) {real, imag} */,
  {32'hc10405ea, 32'hc1893669} /* (26, 25, 9) {real, imag} */,
  {32'h41370ab3, 32'h41dc250c} /* (26, 25, 8) {real, imag} */,
  {32'h3f05bd58, 32'h4043c430} /* (26, 25, 7) {real, imag} */,
  {32'hc042a6e4, 32'hc19a4a94} /* (26, 25, 6) {real, imag} */,
  {32'h417f5eab, 32'hc19a7957} /* (26, 25, 5) {real, imag} */,
  {32'hc0a12fc0, 32'hc0824eb0} /* (26, 25, 4) {real, imag} */,
  {32'h4065c368, 32'h418bdd00} /* (26, 25, 3) {real, imag} */,
  {32'hc0a568ea, 32'h40be00ce} /* (26, 25, 2) {real, imag} */,
  {32'hc1cd02ca, 32'hc0b1503e} /* (26, 25, 1) {real, imag} */,
  {32'hc19c5b62, 32'hbf809baa} /* (26, 25, 0) {real, imag} */,
  {32'hc06c2ee0, 32'h40954f88} /* (26, 24, 31) {real, imag} */,
  {32'hc199902f, 32'h40b16dec} /* (26, 24, 30) {real, imag} */,
  {32'h41cb5d50, 32'hc1e64b8a} /* (26, 24, 29) {real, imag} */,
  {32'hc1aedd4e, 32'hc16dd199} /* (26, 24, 28) {real, imag} */,
  {32'h414ffc8f, 32'hbe8a0828} /* (26, 24, 27) {real, imag} */,
  {32'h407a1a24, 32'hbefa93c8} /* (26, 24, 26) {real, imag} */,
  {32'h41a85fdd, 32'h404430ba} /* (26, 24, 25) {real, imag} */,
  {32'hc18c4e9a, 32'h418c6f4e} /* (26, 24, 24) {real, imag} */,
  {32'h40aedc9c, 32'hc0e54afa} /* (26, 24, 23) {real, imag} */,
  {32'hc16556d4, 32'h412c036a} /* (26, 24, 22) {real, imag} */,
  {32'h4132fe28, 32'h40dcb0d9} /* (26, 24, 21) {real, imag} */,
  {32'h3f7dd9de, 32'h3fd58734} /* (26, 24, 20) {real, imag} */,
  {32'h411836aa, 32'hc091c576} /* (26, 24, 19) {real, imag} */,
  {32'h404f2a30, 32'hc0b1f37a} /* (26, 24, 18) {real, imag} */,
  {32'h40f442d3, 32'hbfc8c350} /* (26, 24, 17) {real, imag} */,
  {32'h407e6c3e, 32'hc053c554} /* (26, 24, 16) {real, imag} */,
  {32'h3ffd60b4, 32'hc1309f67} /* (26, 24, 15) {real, imag} */,
  {32'hc0a22ae0, 32'hc03c2d25} /* (26, 24, 14) {real, imag} */,
  {32'hc1947d64, 32'h3fcf93d4} /* (26, 24, 13) {real, imag} */,
  {32'h40bfa957, 32'hc132b9f2} /* (26, 24, 12) {real, imag} */,
  {32'h3e445880, 32'h41575176} /* (26, 24, 11) {real, imag} */,
  {32'h3eb970e0, 32'h404515ec} /* (26, 24, 10) {real, imag} */,
  {32'hc0e8adf0, 32'h4103859c} /* (26, 24, 9) {real, imag} */,
  {32'h41f2ee4d, 32'hc0e0e254} /* (26, 24, 8) {real, imag} */,
  {32'h40b7418c, 32'h41115e8f} /* (26, 24, 7) {real, imag} */,
  {32'hc194bf92, 32'hc1a135f8} /* (26, 24, 6) {real, imag} */,
  {32'hc1731677, 32'hc10b9ed2} /* (26, 24, 5) {real, imag} */,
  {32'hbffc5cf0, 32'hc10ba91c} /* (26, 24, 4) {real, imag} */,
  {32'hc0e586c8, 32'h41237e35} /* (26, 24, 3) {real, imag} */,
  {32'h410146c1, 32'h3f593bc4} /* (26, 24, 2) {real, imag} */,
  {32'h3fb4f5b8, 32'h41a0619d} /* (26, 24, 1) {real, imag} */,
  {32'hc0fb99ca, 32'h405622e0} /* (26, 24, 0) {real, imag} */,
  {32'h40f66a80, 32'h4183b103} /* (26, 23, 31) {real, imag} */,
  {32'h411e6240, 32'h4181b1d4} /* (26, 23, 30) {real, imag} */,
  {32'hc0e035e4, 32'h40f38ef4} /* (26, 23, 29) {real, imag} */,
  {32'h3fed7868, 32'hc12ac05d} /* (26, 23, 28) {real, imag} */,
  {32'h415886c1, 32'hc1c96e64} /* (26, 23, 27) {real, imag} */,
  {32'h41618bc8, 32'hc0fcef79} /* (26, 23, 26) {real, imag} */,
  {32'h40935104, 32'hc1491233} /* (26, 23, 25) {real, imag} */,
  {32'h3fb37f60, 32'h41aee746} /* (26, 23, 24) {real, imag} */,
  {32'h3e951d80, 32'hc0a02954} /* (26, 23, 23) {real, imag} */,
  {32'hc042a731, 32'hc05c49b8} /* (26, 23, 22) {real, imag} */,
  {32'h404cd736, 32'hc1571efe} /* (26, 23, 21) {real, imag} */,
  {32'h408249d4, 32'hbfe07770} /* (26, 23, 20) {real, imag} */,
  {32'h3eb09090, 32'hc0b20f2b} /* (26, 23, 19) {real, imag} */,
  {32'hc0995e93, 32'hc0984899} /* (26, 23, 18) {real, imag} */,
  {32'hbdf16f80, 32'h4158731b} /* (26, 23, 17) {real, imag} */,
  {32'h407d3eb4, 32'hc0a5602d} /* (26, 23, 16) {real, imag} */,
  {32'h3f81eb24, 32'h409f4ecd} /* (26, 23, 15) {real, imag} */,
  {32'hbd687780, 32'h3fe918f8} /* (26, 23, 14) {real, imag} */,
  {32'h40e027b4, 32'hbfbd7e40} /* (26, 23, 13) {real, imag} */,
  {32'hc1798553, 32'hc1364fd9} /* (26, 23, 12) {real, imag} */,
  {32'hc13b3944, 32'hbfdf0024} /* (26, 23, 11) {real, imag} */,
  {32'hc0d000e1, 32'hc0c1fcca} /* (26, 23, 10) {real, imag} */,
  {32'hc0aa95a7, 32'hc19e7c0c} /* (26, 23, 9) {real, imag} */,
  {32'h3fc043ca, 32'h40b7dd09} /* (26, 23, 8) {real, imag} */,
  {32'h400853bc, 32'hc0089768} /* (26, 23, 7) {real, imag} */,
  {32'hc0a33e48, 32'h413f418b} /* (26, 23, 6) {real, imag} */,
  {32'h40b887cc, 32'hc06dfe79} /* (26, 23, 5) {real, imag} */,
  {32'hc142b5a2, 32'h408fe7a8} /* (26, 23, 4) {real, imag} */,
  {32'h4127ad28, 32'h4060f3ba} /* (26, 23, 3) {real, imag} */,
  {32'hbffd1028, 32'hc1cdfbde} /* (26, 23, 2) {real, imag} */,
  {32'hc0e4b64f, 32'hc1e4d6a6} /* (26, 23, 1) {real, imag} */,
  {32'h403e6910, 32'hc16234a0} /* (26, 23, 0) {real, imag} */,
  {32'h3ff37ea0, 32'hc0b0a3f2} /* (26, 22, 31) {real, imag} */,
  {32'hc191351a, 32'h3f382150} /* (26, 22, 30) {real, imag} */,
  {32'hc0d56b5a, 32'hc0a3f062} /* (26, 22, 29) {real, imag} */,
  {32'hc081c794, 32'hc0f66728} /* (26, 22, 28) {real, imag} */,
  {32'hbf4cb45c, 32'hc1667a43} /* (26, 22, 27) {real, imag} */,
  {32'h4119c96f, 32'hc184ff1d} /* (26, 22, 26) {real, imag} */,
  {32'h41920d6b, 32'hbf1a1684} /* (26, 22, 25) {real, imag} */,
  {32'h4189e765, 32'hc07944a6} /* (26, 22, 24) {real, imag} */,
  {32'hc17351c7, 32'h41543188} /* (26, 22, 23) {real, imag} */,
  {32'hc150e269, 32'hbfff0b48} /* (26, 22, 22) {real, imag} */,
  {32'hc0476a06, 32'hc1538315} /* (26, 22, 21) {real, imag} */,
  {32'hc0966510, 32'hc0f4c794} /* (26, 22, 20) {real, imag} */,
  {32'hbfb67f98, 32'h41b1b2a9} /* (26, 22, 19) {real, imag} */,
  {32'h41e0c595, 32'hc0b12660} /* (26, 22, 18) {real, imag} */,
  {32'hbf334160, 32'h3fa5b0a4} /* (26, 22, 17) {real, imag} */,
  {32'h4116159a, 32'hc0356529} /* (26, 22, 16) {real, imag} */,
  {32'h410358ba, 32'h3f15447a} /* (26, 22, 15) {real, imag} */,
  {32'hbfc7d13e, 32'hc09ceebe} /* (26, 22, 14) {real, imag} */,
  {32'h4170d5be, 32'hc11826d9} /* (26, 22, 13) {real, imag} */,
  {32'hc11c7097, 32'hbfe64184} /* (26, 22, 12) {real, imag} */,
  {32'h40fa354a, 32'h41173496} /* (26, 22, 11) {real, imag} */,
  {32'h4193a47a, 32'h4153c15d} /* (26, 22, 10) {real, imag} */,
  {32'hc09d1f16, 32'hc1f6c6fc} /* (26, 22, 9) {real, imag} */,
  {32'hc14d5566, 32'h41035672} /* (26, 22, 8) {real, imag} */,
  {32'hc1098e7b, 32'h40e4c5fb} /* (26, 22, 7) {real, imag} */,
  {32'hc187f7a3, 32'h40da04f0} /* (26, 22, 6) {real, imag} */,
  {32'h40eaf63f, 32'h40b891b7} /* (26, 22, 5) {real, imag} */,
  {32'hc0d22fe0, 32'hc0379ad2} /* (26, 22, 4) {real, imag} */,
  {32'h4008df6e, 32'hc1313864} /* (26, 22, 3) {real, imag} */,
  {32'h41366c73, 32'hbf379950} /* (26, 22, 2) {real, imag} */,
  {32'hc0eb6042, 32'hc1155927} /* (26, 22, 1) {real, imag} */,
  {32'h40f14cac, 32'hc0d9a308} /* (26, 22, 0) {real, imag} */,
  {32'hc0a93c00, 32'hc101dd33} /* (26, 21, 31) {real, imag} */,
  {32'h40bcddbe, 32'hbfad04f8} /* (26, 21, 30) {real, imag} */,
  {32'hc1b24d69, 32'hc09889c9} /* (26, 21, 29) {real, imag} */,
  {32'hc05944df, 32'hc1b07906} /* (26, 21, 28) {real, imag} */,
  {32'h3fff6f32, 32'h41798328} /* (26, 21, 27) {real, imag} */,
  {32'hc0127096, 32'hc0ed5f42} /* (26, 21, 26) {real, imag} */,
  {32'hc13a0d38, 32'hbf04f020} /* (26, 21, 25) {real, imag} */,
  {32'hc13e31cf, 32'hc11df5b9} /* (26, 21, 24) {real, imag} */,
  {32'h40a4d760, 32'hc08b940b} /* (26, 21, 23) {real, imag} */,
  {32'hc15a5cca, 32'hbfd39c68} /* (26, 21, 22) {real, imag} */,
  {32'hbff9c260, 32'hc19a1442} /* (26, 21, 21) {real, imag} */,
  {32'h4104884c, 32'h41095928} /* (26, 21, 20) {real, imag} */,
  {32'hc19d9f5a, 32'hc10dd217} /* (26, 21, 19) {real, imag} */,
  {32'h4112566b, 32'hbf4887d4} /* (26, 21, 18) {real, imag} */,
  {32'h409a359a, 32'h410ef6a6} /* (26, 21, 17) {real, imag} */,
  {32'h3ebcc8d8, 32'h415125d2} /* (26, 21, 16) {real, imag} */,
  {32'h412e67c8, 32'hc167d40b} /* (26, 21, 15) {real, imag} */,
  {32'hc1a3239a, 32'h416e5c2d} /* (26, 21, 14) {real, imag} */,
  {32'h40aaf216, 32'h40087f90} /* (26, 21, 13) {real, imag} */,
  {32'hc14735f2, 32'h418ff434} /* (26, 21, 12) {real, imag} */,
  {32'hc017cdd8, 32'h40cf0da7} /* (26, 21, 11) {real, imag} */,
  {32'hc16118dc, 32'h40cfce8c} /* (26, 21, 10) {real, imag} */,
  {32'h402963d4, 32'hc0a05b54} /* (26, 21, 9) {real, imag} */,
  {32'hc145db78, 32'h3fec2614} /* (26, 21, 8) {real, imag} */,
  {32'h41141c1c, 32'hc0502d52} /* (26, 21, 7) {real, imag} */,
  {32'hc15add87, 32'h41d67cd0} /* (26, 21, 6) {real, imag} */,
  {32'hc1559f8f, 32'h40b63809} /* (26, 21, 5) {real, imag} */,
  {32'hbf9cd748, 32'hc1594964} /* (26, 21, 4) {real, imag} */,
  {32'h413e9fb4, 32'h40a824ca} /* (26, 21, 3) {real, imag} */,
  {32'h401b8fa9, 32'hbfc70910} /* (26, 21, 2) {real, imag} */,
  {32'hc0fdd766, 32'h41797d7f} /* (26, 21, 1) {real, imag} */,
  {32'hc19cf981, 32'h4168ead4} /* (26, 21, 0) {real, imag} */,
  {32'hc03005fa, 32'hc067c8e0} /* (26, 20, 31) {real, imag} */,
  {32'h3fa33438, 32'hc09f0cc6} /* (26, 20, 30) {real, imag} */,
  {32'h4004af28, 32'hc18577a6} /* (26, 20, 29) {real, imag} */,
  {32'hc06b1312, 32'hbfaefb1e} /* (26, 20, 28) {real, imag} */,
  {32'h3ff1b10e, 32'hbfd79170} /* (26, 20, 27) {real, imag} */,
  {32'hc19193ea, 32'hc0f72b32} /* (26, 20, 26) {real, imag} */,
  {32'h411cf298, 32'hc0f08f68} /* (26, 20, 25) {real, imag} */,
  {32'h401b7768, 32'h3fd5a208} /* (26, 20, 24) {real, imag} */,
  {32'hc17e8487, 32'h417087a2} /* (26, 20, 23) {real, imag} */,
  {32'hc0895ed2, 32'hc0a76729} /* (26, 20, 22) {real, imag} */,
  {32'h409e5f59, 32'hc065074e} /* (26, 20, 21) {real, imag} */,
  {32'hbf7f40ca, 32'h40bd7112} /* (26, 20, 20) {real, imag} */,
  {32'h408877b3, 32'h409ada38} /* (26, 20, 19) {real, imag} */,
  {32'h4101f634, 32'hc022d0bf} /* (26, 20, 18) {real, imag} */,
  {32'hc043800c, 32'hc10c50be} /* (26, 20, 17) {real, imag} */,
  {32'hc02e036a, 32'h414ca1e7} /* (26, 20, 16) {real, imag} */,
  {32'hc1a20a3a, 32'hc146b939} /* (26, 20, 15) {real, imag} */,
  {32'h4070a5ea, 32'hc059479d} /* (26, 20, 14) {real, imag} */,
  {32'h40c75e6c, 32'hc1752ca6} /* (26, 20, 13) {real, imag} */,
  {32'hc058794e, 32'hbfe8e140} /* (26, 20, 12) {real, imag} */,
  {32'hc14e872e, 32'hc07d3d3c} /* (26, 20, 11) {real, imag} */,
  {32'h3e3c67a0, 32'h40a30ca4} /* (26, 20, 10) {real, imag} */,
  {32'h40952f68, 32'h41b60888} /* (26, 20, 9) {real, imag} */,
  {32'hc191d211, 32'h40edda89} /* (26, 20, 8) {real, imag} */,
  {32'hc0fa6148, 32'hc19210ca} /* (26, 20, 7) {real, imag} */,
  {32'h40126fce, 32'h410fd298} /* (26, 20, 6) {real, imag} */,
  {32'hbfb71670, 32'hc03e3716} /* (26, 20, 5) {real, imag} */,
  {32'hc0aa7129, 32'hc0f24096} /* (26, 20, 4) {real, imag} */,
  {32'h40ae339e, 32'h413b52aa} /* (26, 20, 3) {real, imag} */,
  {32'hbf4c53d0, 32'hc13fb70e} /* (26, 20, 2) {real, imag} */,
  {32'hbf855e90, 32'hc1391d7f} /* (26, 20, 1) {real, imag} */,
  {32'h41a336c3, 32'h41e36d4a} /* (26, 20, 0) {real, imag} */,
  {32'hc005bd0e, 32'hc070c2a4} /* (26, 19, 31) {real, imag} */,
  {32'hc0583bba, 32'hc1080ca9} /* (26, 19, 30) {real, imag} */,
  {32'h4149ae4b, 32'hc0017432} /* (26, 19, 29) {real, imag} */,
  {32'hc11a84e1, 32'hc175018c} /* (26, 19, 28) {real, imag} */,
  {32'hbf451770, 32'h412a72f2} /* (26, 19, 27) {real, imag} */,
  {32'hc15a23b0, 32'h40fd65ea} /* (26, 19, 26) {real, imag} */,
  {32'h411c2a31, 32'h409e92d8} /* (26, 19, 25) {real, imag} */,
  {32'h4151ef5d, 32'h4051f536} /* (26, 19, 24) {real, imag} */,
  {32'hc1011c5f, 32'h3e89d5a0} /* (26, 19, 23) {real, imag} */,
  {32'h413709d4, 32'hbfe5ffb2} /* (26, 19, 22) {real, imag} */,
  {32'h4103ad80, 32'hc130b11e} /* (26, 19, 21) {real, imag} */,
  {32'hc11a8176, 32'hbffa4ec8} /* (26, 19, 20) {real, imag} */,
  {32'hc165feea, 32'h41795524} /* (26, 19, 19) {real, imag} */,
  {32'h40e44d9e, 32'h412800a5} /* (26, 19, 18) {real, imag} */,
  {32'h409383ec, 32'hc02863d4} /* (26, 19, 17) {real, imag} */,
  {32'h402bd8ba, 32'h40258bcd} /* (26, 19, 16) {real, imag} */,
  {32'hc151fb1a, 32'hc01413d5} /* (26, 19, 15) {real, imag} */,
  {32'hc0b96370, 32'hc027344d} /* (26, 19, 14) {real, imag} */,
  {32'hc0cf78b8, 32'hc108d67c} /* (26, 19, 13) {real, imag} */,
  {32'hbfe076a0, 32'hc1873aac} /* (26, 19, 12) {real, imag} */,
  {32'hbee9a530, 32'hc08256db} /* (26, 19, 11) {real, imag} */,
  {32'h41301879, 32'hc193a284} /* (26, 19, 10) {real, imag} */,
  {32'h40793d04, 32'h3e975860} /* (26, 19, 9) {real, imag} */,
  {32'h407b26fb, 32'h41957fb6} /* (26, 19, 8) {real, imag} */,
  {32'h4102169a, 32'hc0ac4182} /* (26, 19, 7) {real, imag} */,
  {32'h4149183e, 32'h3fbecd1e} /* (26, 19, 6) {real, imag} */,
  {32'hc0681048, 32'hc12a3c4f} /* (26, 19, 5) {real, imag} */,
  {32'h40ca08f7, 32'hc0fb802c} /* (26, 19, 4) {real, imag} */,
  {32'hbe507aa0, 32'h3f9f8452} /* (26, 19, 3) {real, imag} */,
  {32'h40a3a817, 32'h400f4338} /* (26, 19, 2) {real, imag} */,
  {32'h3ffefd8c, 32'h4165a5f2} /* (26, 19, 1) {real, imag} */,
  {32'hc0469110, 32'hc09656f6} /* (26, 19, 0) {real, imag} */,
  {32'hc143cb49, 32'hc05ac8d6} /* (26, 18, 31) {real, imag} */,
  {32'h40ca0ec2, 32'h4193cfbe} /* (26, 18, 30) {real, imag} */,
  {32'h4131eb71, 32'hc1472c37} /* (26, 18, 29) {real, imag} */,
  {32'hc12b4235, 32'hc0da2794} /* (26, 18, 28) {real, imag} */,
  {32'h40c42bb2, 32'h4136e976} /* (26, 18, 27) {real, imag} */,
  {32'hc12d0114, 32'hc067e7ec} /* (26, 18, 26) {real, imag} */,
  {32'hc10f1161, 32'h41272c00} /* (26, 18, 25) {real, imag} */,
  {32'hc04208fd, 32'hc0872640} /* (26, 18, 24) {real, imag} */,
  {32'h408ef6a6, 32'hc0e00c2a} /* (26, 18, 23) {real, imag} */,
  {32'hbf653800, 32'h41697c82} /* (26, 18, 22) {real, imag} */,
  {32'hc011098c, 32'h41474949} /* (26, 18, 21) {real, imag} */,
  {32'hc15580c5, 32'h40f173b4} /* (26, 18, 20) {real, imag} */,
  {32'h40c65278, 32'hc09704b2} /* (26, 18, 19) {real, imag} */,
  {32'hc0a8d713, 32'h41882daa} /* (26, 18, 18) {real, imag} */,
  {32'hc128db21, 32'hc0815976} /* (26, 18, 17) {real, imag} */,
  {32'h4098af1f, 32'h40c71ac2} /* (26, 18, 16) {real, imag} */,
  {32'h417145d2, 32'h41722df8} /* (26, 18, 15) {real, imag} */,
  {32'hc0cc740e, 32'hc0478f79} /* (26, 18, 14) {real, imag} */,
  {32'h3feb9ff0, 32'h4072dc74} /* (26, 18, 13) {real, imag} */,
  {32'h40ea8b87, 32'h3fc7c508} /* (26, 18, 12) {real, imag} */,
  {32'h41606ae2, 32'h404c6106} /* (26, 18, 11) {real, imag} */,
  {32'h40d3dd1c, 32'hc072ef80} /* (26, 18, 10) {real, imag} */,
  {32'h4106b58a, 32'hc06ba05c} /* (26, 18, 9) {real, imag} */,
  {32'hc067cada, 32'hc1126c1b} /* (26, 18, 8) {real, imag} */,
  {32'h40782f88, 32'hc0b569c8} /* (26, 18, 7) {real, imag} */,
  {32'h410ed0be, 32'hbefc9568} /* (26, 18, 6) {real, imag} */,
  {32'hc0b65743, 32'h40860ad2} /* (26, 18, 5) {real, imag} */,
  {32'hc10b1bf2, 32'h41035dad} /* (26, 18, 4) {real, imag} */,
  {32'h410ac57c, 32'h40502ac0} /* (26, 18, 3) {real, imag} */,
  {32'h415d557a, 32'hc0dd732d} /* (26, 18, 2) {real, imag} */,
  {32'hc0bf0f6c, 32'h4080fe24} /* (26, 18, 1) {real, imag} */,
  {32'h40f4d8d0, 32'hc163b734} /* (26, 18, 0) {real, imag} */,
  {32'hc05ec7e8, 32'hc00d8f37} /* (26, 17, 31) {real, imag} */,
  {32'hbfb7c612, 32'hbf282a30} /* (26, 17, 30) {real, imag} */,
  {32'h40b1db82, 32'h4093d620} /* (26, 17, 29) {real, imag} */,
  {32'hc0911d3e, 32'h3dd1ad00} /* (26, 17, 28) {real, imag} */,
  {32'h41237628, 32'hc0e4be64} /* (26, 17, 27) {real, imag} */,
  {32'hbea43bd4, 32'hc15a4351} /* (26, 17, 26) {real, imag} */,
  {32'h40b73414, 32'hbfb59324} /* (26, 17, 25) {real, imag} */,
  {32'hc1156468, 32'h409e94a9} /* (26, 17, 24) {real, imag} */,
  {32'hc097db80, 32'h4006d8fa} /* (26, 17, 23) {real, imag} */,
  {32'hc1237d38, 32'hc17aee83} /* (26, 17, 22) {real, imag} */,
  {32'h40eab226, 32'h417fba3a} /* (26, 17, 21) {real, imag} */,
  {32'hc12396bc, 32'hc0884e6a} /* (26, 17, 20) {real, imag} */,
  {32'hbf950dae, 32'h40438a91} /* (26, 17, 19) {real, imag} */,
  {32'hbf3c803c, 32'hc141f766} /* (26, 17, 18) {real, imag} */,
  {32'hc0e20a90, 32'hc0ed94f8} /* (26, 17, 17) {real, imag} */,
  {32'h408f8928, 32'h3efaf228} /* (26, 17, 16) {real, imag} */,
  {32'h411716d6, 32'h405ed3e0} /* (26, 17, 15) {real, imag} */,
  {32'h3fa0c60a, 32'h410fc3c4} /* (26, 17, 14) {real, imag} */,
  {32'hc1379f5a, 32'hc08cf49a} /* (26, 17, 13) {real, imag} */,
  {32'h40d626b0, 32'hbe8d8ec8} /* (26, 17, 12) {real, imag} */,
  {32'h408fc810, 32'h40afdcae} /* (26, 17, 11) {real, imag} */,
  {32'hbd907780, 32'hc17743cf} /* (26, 17, 10) {real, imag} */,
  {32'hc0c090db, 32'h411c79b2} /* (26, 17, 9) {real, imag} */,
  {32'hc0bdaafa, 32'hc0f08194} /* (26, 17, 8) {real, imag} */,
  {32'hc01ed18a, 32'h40005a88} /* (26, 17, 7) {real, imag} */,
  {32'h410c5cf3, 32'hc0e03ef3} /* (26, 17, 6) {real, imag} */,
  {32'hc10133ac, 32'h3f8fbfe0} /* (26, 17, 5) {real, imag} */,
  {32'h40cf4178, 32'h41398e5c} /* (26, 17, 4) {real, imag} */,
  {32'hc08abd77, 32'hbba10300} /* (26, 17, 3) {real, imag} */,
  {32'hc0b7f41a, 32'hc082a19f} /* (26, 17, 2) {real, imag} */,
  {32'hc1618874, 32'h411424c0} /* (26, 17, 1) {real, imag} */,
  {32'hc0739cd6, 32'hbf8a1d90} /* (26, 17, 0) {real, imag} */,
  {32'h3faf9696, 32'hc0f62ab7} /* (26, 16, 31) {real, imag} */,
  {32'h40a2568c, 32'hc073ffa2} /* (26, 16, 30) {real, imag} */,
  {32'h3da718a0, 32'hc0c9c2d9} /* (26, 16, 29) {real, imag} */,
  {32'h4033067c, 32'hc0d0a902} /* (26, 16, 28) {real, imag} */,
  {32'hc0a9a95c, 32'hc0fce2b2} /* (26, 16, 27) {real, imag} */,
  {32'hc0e8ac0c, 32'hbeb3d5ee} /* (26, 16, 26) {real, imag} */,
  {32'hbfc9f16e, 32'hbfb9f718} /* (26, 16, 25) {real, imag} */,
  {32'hc0e2eb82, 32'h41148576} /* (26, 16, 24) {real, imag} */,
  {32'h40fb631d, 32'h3f1f1e38} /* (26, 16, 23) {real, imag} */,
  {32'h3f7cf498, 32'hc023e0ac} /* (26, 16, 22) {real, imag} */,
  {32'h40e35c66, 32'hbfd84a12} /* (26, 16, 21) {real, imag} */,
  {32'hc0cc3f01, 32'hc107aa71} /* (26, 16, 20) {real, imag} */,
  {32'hbe1ac210, 32'h40c5c16c} /* (26, 16, 19) {real, imag} */,
  {32'h401bbbd6, 32'hc1246c62} /* (26, 16, 18) {real, imag} */,
  {32'h40da3487, 32'hc04d0cea} /* (26, 16, 17) {real, imag} */,
  {32'h3f16db44, 32'h00000000} /* (26, 16, 16) {real, imag} */,
  {32'h40da3487, 32'h404d0cea} /* (26, 16, 15) {real, imag} */,
  {32'h401bbbd6, 32'h41246c62} /* (26, 16, 14) {real, imag} */,
  {32'hbe1ac210, 32'hc0c5c16c} /* (26, 16, 13) {real, imag} */,
  {32'hc0cc3f01, 32'h4107aa71} /* (26, 16, 12) {real, imag} */,
  {32'h40e35c66, 32'h3fd84a12} /* (26, 16, 11) {real, imag} */,
  {32'h3f7cf498, 32'h4023e0ac} /* (26, 16, 10) {real, imag} */,
  {32'h40fb631d, 32'hbf1f1e38} /* (26, 16, 9) {real, imag} */,
  {32'hc0e2eb82, 32'hc1148576} /* (26, 16, 8) {real, imag} */,
  {32'hbfc9f16e, 32'h3fb9f718} /* (26, 16, 7) {real, imag} */,
  {32'hc0e8ac0c, 32'h3eb3d5ee} /* (26, 16, 6) {real, imag} */,
  {32'hc0a9a95c, 32'h40fce2b2} /* (26, 16, 5) {real, imag} */,
  {32'h4033067c, 32'h40d0a902} /* (26, 16, 4) {real, imag} */,
  {32'h3da718a0, 32'h40c9c2d9} /* (26, 16, 3) {real, imag} */,
  {32'h40a2568c, 32'h4073ffa2} /* (26, 16, 2) {real, imag} */,
  {32'h3faf9696, 32'h40f62ab7} /* (26, 16, 1) {real, imag} */,
  {32'h40bdbece, 32'h00000000} /* (26, 16, 0) {real, imag} */,
  {32'hc1618874, 32'hc11424c0} /* (26, 15, 31) {real, imag} */,
  {32'hc0b7f41a, 32'h4082a19f} /* (26, 15, 30) {real, imag} */,
  {32'hc08abd77, 32'h3ba10300} /* (26, 15, 29) {real, imag} */,
  {32'h40cf4178, 32'hc1398e5c} /* (26, 15, 28) {real, imag} */,
  {32'hc10133ac, 32'hbf8fbfe0} /* (26, 15, 27) {real, imag} */,
  {32'h410c5cf3, 32'h40e03ef3} /* (26, 15, 26) {real, imag} */,
  {32'hc01ed18a, 32'hc0005a88} /* (26, 15, 25) {real, imag} */,
  {32'hc0bdaafa, 32'h40f08194} /* (26, 15, 24) {real, imag} */,
  {32'hc0c090db, 32'hc11c79b2} /* (26, 15, 23) {real, imag} */,
  {32'hbd907780, 32'h417743cf} /* (26, 15, 22) {real, imag} */,
  {32'h408fc810, 32'hc0afdcae} /* (26, 15, 21) {real, imag} */,
  {32'h40d626b0, 32'h3e8d8ec8} /* (26, 15, 20) {real, imag} */,
  {32'hc1379f5a, 32'h408cf49a} /* (26, 15, 19) {real, imag} */,
  {32'h3fa0c60a, 32'hc10fc3c4} /* (26, 15, 18) {real, imag} */,
  {32'h411716d6, 32'hc05ed3e0} /* (26, 15, 17) {real, imag} */,
  {32'h408f8928, 32'hbefaf228} /* (26, 15, 16) {real, imag} */,
  {32'hc0e20a90, 32'h40ed94f8} /* (26, 15, 15) {real, imag} */,
  {32'hbf3c803c, 32'h4141f766} /* (26, 15, 14) {real, imag} */,
  {32'hbf950dae, 32'hc0438a91} /* (26, 15, 13) {real, imag} */,
  {32'hc12396bc, 32'h40884e6a} /* (26, 15, 12) {real, imag} */,
  {32'h40eab226, 32'hc17fba3a} /* (26, 15, 11) {real, imag} */,
  {32'hc1237d38, 32'h417aee83} /* (26, 15, 10) {real, imag} */,
  {32'hc097db80, 32'hc006d8fa} /* (26, 15, 9) {real, imag} */,
  {32'hc1156468, 32'hc09e94a9} /* (26, 15, 8) {real, imag} */,
  {32'h40b73414, 32'h3fb59324} /* (26, 15, 7) {real, imag} */,
  {32'hbea43bd4, 32'h415a4351} /* (26, 15, 6) {real, imag} */,
  {32'h41237628, 32'h40e4be64} /* (26, 15, 5) {real, imag} */,
  {32'hc0911d3e, 32'hbdd1ad00} /* (26, 15, 4) {real, imag} */,
  {32'h40b1db82, 32'hc093d620} /* (26, 15, 3) {real, imag} */,
  {32'hbfb7c612, 32'h3f282a30} /* (26, 15, 2) {real, imag} */,
  {32'hc05ec7e8, 32'h400d8f37} /* (26, 15, 1) {real, imag} */,
  {32'hc0739cd6, 32'h3f8a1d90} /* (26, 15, 0) {real, imag} */,
  {32'hc0bf0f6c, 32'hc080fe24} /* (26, 14, 31) {real, imag} */,
  {32'h415d557a, 32'h40dd732d} /* (26, 14, 30) {real, imag} */,
  {32'h410ac57c, 32'hc0502ac0} /* (26, 14, 29) {real, imag} */,
  {32'hc10b1bf2, 32'hc1035dad} /* (26, 14, 28) {real, imag} */,
  {32'hc0b65743, 32'hc0860ad2} /* (26, 14, 27) {real, imag} */,
  {32'h410ed0be, 32'h3efc9568} /* (26, 14, 26) {real, imag} */,
  {32'h40782f88, 32'h40b569c8} /* (26, 14, 25) {real, imag} */,
  {32'hc067cada, 32'h41126c1b} /* (26, 14, 24) {real, imag} */,
  {32'h4106b58a, 32'h406ba05c} /* (26, 14, 23) {real, imag} */,
  {32'h40d3dd1c, 32'h4072ef80} /* (26, 14, 22) {real, imag} */,
  {32'h41606ae2, 32'hc04c6106} /* (26, 14, 21) {real, imag} */,
  {32'h40ea8b87, 32'hbfc7c508} /* (26, 14, 20) {real, imag} */,
  {32'h3feb9ff0, 32'hc072dc74} /* (26, 14, 19) {real, imag} */,
  {32'hc0cc740e, 32'h40478f79} /* (26, 14, 18) {real, imag} */,
  {32'h417145d2, 32'hc1722df8} /* (26, 14, 17) {real, imag} */,
  {32'h4098af1f, 32'hc0c71ac2} /* (26, 14, 16) {real, imag} */,
  {32'hc128db21, 32'h40815976} /* (26, 14, 15) {real, imag} */,
  {32'hc0a8d713, 32'hc1882daa} /* (26, 14, 14) {real, imag} */,
  {32'h40c65278, 32'h409704b2} /* (26, 14, 13) {real, imag} */,
  {32'hc15580c5, 32'hc0f173b4} /* (26, 14, 12) {real, imag} */,
  {32'hc011098c, 32'hc1474949} /* (26, 14, 11) {real, imag} */,
  {32'hbf653800, 32'hc1697c82} /* (26, 14, 10) {real, imag} */,
  {32'h408ef6a6, 32'h40e00c2a} /* (26, 14, 9) {real, imag} */,
  {32'hc04208fd, 32'h40872640} /* (26, 14, 8) {real, imag} */,
  {32'hc10f1161, 32'hc1272c00} /* (26, 14, 7) {real, imag} */,
  {32'hc12d0114, 32'h4067e7ec} /* (26, 14, 6) {real, imag} */,
  {32'h40c42bb2, 32'hc136e976} /* (26, 14, 5) {real, imag} */,
  {32'hc12b4235, 32'h40da2794} /* (26, 14, 4) {real, imag} */,
  {32'h4131eb71, 32'h41472c37} /* (26, 14, 3) {real, imag} */,
  {32'h40ca0ec2, 32'hc193cfbe} /* (26, 14, 2) {real, imag} */,
  {32'hc143cb49, 32'h405ac8d6} /* (26, 14, 1) {real, imag} */,
  {32'h40f4d8d0, 32'h4163b734} /* (26, 14, 0) {real, imag} */,
  {32'h3ffefd8c, 32'hc165a5f2} /* (26, 13, 31) {real, imag} */,
  {32'h40a3a817, 32'hc00f4338} /* (26, 13, 30) {real, imag} */,
  {32'hbe507aa0, 32'hbf9f8452} /* (26, 13, 29) {real, imag} */,
  {32'h40ca08f7, 32'h40fb802c} /* (26, 13, 28) {real, imag} */,
  {32'hc0681048, 32'h412a3c4f} /* (26, 13, 27) {real, imag} */,
  {32'h4149183e, 32'hbfbecd1e} /* (26, 13, 26) {real, imag} */,
  {32'h4102169a, 32'h40ac4182} /* (26, 13, 25) {real, imag} */,
  {32'h407b26fb, 32'hc1957fb6} /* (26, 13, 24) {real, imag} */,
  {32'h40793d04, 32'hbe975860} /* (26, 13, 23) {real, imag} */,
  {32'h41301879, 32'h4193a284} /* (26, 13, 22) {real, imag} */,
  {32'hbee9a530, 32'h408256db} /* (26, 13, 21) {real, imag} */,
  {32'hbfe076a0, 32'h41873aac} /* (26, 13, 20) {real, imag} */,
  {32'hc0cf78b8, 32'h4108d67c} /* (26, 13, 19) {real, imag} */,
  {32'hc0b96370, 32'h4027344d} /* (26, 13, 18) {real, imag} */,
  {32'hc151fb1a, 32'h401413d5} /* (26, 13, 17) {real, imag} */,
  {32'h402bd8ba, 32'hc0258bcd} /* (26, 13, 16) {real, imag} */,
  {32'h409383ec, 32'h402863d4} /* (26, 13, 15) {real, imag} */,
  {32'h40e44d9e, 32'hc12800a5} /* (26, 13, 14) {real, imag} */,
  {32'hc165feea, 32'hc1795524} /* (26, 13, 13) {real, imag} */,
  {32'hc11a8176, 32'h3ffa4ec8} /* (26, 13, 12) {real, imag} */,
  {32'h4103ad80, 32'h4130b11e} /* (26, 13, 11) {real, imag} */,
  {32'h413709d4, 32'h3fe5ffb2} /* (26, 13, 10) {real, imag} */,
  {32'hc1011c5f, 32'hbe89d5a0} /* (26, 13, 9) {real, imag} */,
  {32'h4151ef5d, 32'hc051f536} /* (26, 13, 8) {real, imag} */,
  {32'h411c2a31, 32'hc09e92d8} /* (26, 13, 7) {real, imag} */,
  {32'hc15a23b0, 32'hc0fd65ea} /* (26, 13, 6) {real, imag} */,
  {32'hbf451770, 32'hc12a72f2} /* (26, 13, 5) {real, imag} */,
  {32'hc11a84e1, 32'h4175018c} /* (26, 13, 4) {real, imag} */,
  {32'h4149ae4b, 32'h40017432} /* (26, 13, 3) {real, imag} */,
  {32'hc0583bba, 32'h41080ca9} /* (26, 13, 2) {real, imag} */,
  {32'hc005bd0e, 32'h4070c2a4} /* (26, 13, 1) {real, imag} */,
  {32'hc0469110, 32'h409656f6} /* (26, 13, 0) {real, imag} */,
  {32'hbf855e90, 32'h41391d7f} /* (26, 12, 31) {real, imag} */,
  {32'hbf4c53d0, 32'h413fb70e} /* (26, 12, 30) {real, imag} */,
  {32'h40ae339e, 32'hc13b52aa} /* (26, 12, 29) {real, imag} */,
  {32'hc0aa7129, 32'h40f24096} /* (26, 12, 28) {real, imag} */,
  {32'hbfb71670, 32'h403e3716} /* (26, 12, 27) {real, imag} */,
  {32'h40126fce, 32'hc10fd298} /* (26, 12, 26) {real, imag} */,
  {32'hc0fa6148, 32'h419210ca} /* (26, 12, 25) {real, imag} */,
  {32'hc191d211, 32'hc0edda89} /* (26, 12, 24) {real, imag} */,
  {32'h40952f68, 32'hc1b60888} /* (26, 12, 23) {real, imag} */,
  {32'h3e3c67a0, 32'hc0a30ca4} /* (26, 12, 22) {real, imag} */,
  {32'hc14e872e, 32'h407d3d3c} /* (26, 12, 21) {real, imag} */,
  {32'hc058794e, 32'h3fe8e140} /* (26, 12, 20) {real, imag} */,
  {32'h40c75e6c, 32'h41752ca6} /* (26, 12, 19) {real, imag} */,
  {32'h4070a5ea, 32'h4059479d} /* (26, 12, 18) {real, imag} */,
  {32'hc1a20a3a, 32'h4146b939} /* (26, 12, 17) {real, imag} */,
  {32'hc02e036a, 32'hc14ca1e7} /* (26, 12, 16) {real, imag} */,
  {32'hc043800c, 32'h410c50be} /* (26, 12, 15) {real, imag} */,
  {32'h4101f634, 32'h4022d0bf} /* (26, 12, 14) {real, imag} */,
  {32'h408877b3, 32'hc09ada38} /* (26, 12, 13) {real, imag} */,
  {32'hbf7f40ca, 32'hc0bd7112} /* (26, 12, 12) {real, imag} */,
  {32'h409e5f59, 32'h4065074e} /* (26, 12, 11) {real, imag} */,
  {32'hc0895ed2, 32'h40a76729} /* (26, 12, 10) {real, imag} */,
  {32'hc17e8487, 32'hc17087a2} /* (26, 12, 9) {real, imag} */,
  {32'h401b7768, 32'hbfd5a208} /* (26, 12, 8) {real, imag} */,
  {32'h411cf298, 32'h40f08f68} /* (26, 12, 7) {real, imag} */,
  {32'hc19193ea, 32'h40f72b32} /* (26, 12, 6) {real, imag} */,
  {32'h3ff1b10e, 32'h3fd79170} /* (26, 12, 5) {real, imag} */,
  {32'hc06b1312, 32'h3faefb1e} /* (26, 12, 4) {real, imag} */,
  {32'h4004af28, 32'h418577a6} /* (26, 12, 3) {real, imag} */,
  {32'h3fa33438, 32'h409f0cc6} /* (26, 12, 2) {real, imag} */,
  {32'hc03005fa, 32'h4067c8e0} /* (26, 12, 1) {real, imag} */,
  {32'h41a336c3, 32'hc1e36d4a} /* (26, 12, 0) {real, imag} */,
  {32'hc0fdd766, 32'hc1797d7f} /* (26, 11, 31) {real, imag} */,
  {32'h401b8fa9, 32'h3fc70910} /* (26, 11, 30) {real, imag} */,
  {32'h413e9fb4, 32'hc0a824ca} /* (26, 11, 29) {real, imag} */,
  {32'hbf9cd748, 32'h41594964} /* (26, 11, 28) {real, imag} */,
  {32'hc1559f8f, 32'hc0b63809} /* (26, 11, 27) {real, imag} */,
  {32'hc15add87, 32'hc1d67cd0} /* (26, 11, 26) {real, imag} */,
  {32'h41141c1c, 32'h40502d52} /* (26, 11, 25) {real, imag} */,
  {32'hc145db78, 32'hbfec2614} /* (26, 11, 24) {real, imag} */,
  {32'h402963d4, 32'h40a05b54} /* (26, 11, 23) {real, imag} */,
  {32'hc16118dc, 32'hc0cfce8c} /* (26, 11, 22) {real, imag} */,
  {32'hc017cdd8, 32'hc0cf0da7} /* (26, 11, 21) {real, imag} */,
  {32'hc14735f2, 32'hc18ff434} /* (26, 11, 20) {real, imag} */,
  {32'h40aaf216, 32'hc0087f90} /* (26, 11, 19) {real, imag} */,
  {32'hc1a3239a, 32'hc16e5c2d} /* (26, 11, 18) {real, imag} */,
  {32'h412e67c8, 32'h4167d40b} /* (26, 11, 17) {real, imag} */,
  {32'h3ebcc8d8, 32'hc15125d2} /* (26, 11, 16) {real, imag} */,
  {32'h409a359a, 32'hc10ef6a6} /* (26, 11, 15) {real, imag} */,
  {32'h4112566b, 32'h3f4887d4} /* (26, 11, 14) {real, imag} */,
  {32'hc19d9f5a, 32'h410dd217} /* (26, 11, 13) {real, imag} */,
  {32'h4104884c, 32'hc1095928} /* (26, 11, 12) {real, imag} */,
  {32'hbff9c260, 32'h419a1442} /* (26, 11, 11) {real, imag} */,
  {32'hc15a5cca, 32'h3fd39c68} /* (26, 11, 10) {real, imag} */,
  {32'h40a4d760, 32'h408b940b} /* (26, 11, 9) {real, imag} */,
  {32'hc13e31cf, 32'h411df5b9} /* (26, 11, 8) {real, imag} */,
  {32'hc13a0d38, 32'h3f04f020} /* (26, 11, 7) {real, imag} */,
  {32'hc0127096, 32'h40ed5f42} /* (26, 11, 6) {real, imag} */,
  {32'h3fff6f32, 32'hc1798328} /* (26, 11, 5) {real, imag} */,
  {32'hc05944df, 32'h41b07906} /* (26, 11, 4) {real, imag} */,
  {32'hc1b24d69, 32'h409889c9} /* (26, 11, 3) {real, imag} */,
  {32'h40bcddbe, 32'h3fad04f8} /* (26, 11, 2) {real, imag} */,
  {32'hc0a93c00, 32'h4101dd33} /* (26, 11, 1) {real, imag} */,
  {32'hc19cf981, 32'hc168ead4} /* (26, 11, 0) {real, imag} */,
  {32'hc0eb6042, 32'h41155927} /* (26, 10, 31) {real, imag} */,
  {32'h41366c73, 32'h3f379950} /* (26, 10, 30) {real, imag} */,
  {32'h4008df6e, 32'h41313864} /* (26, 10, 29) {real, imag} */,
  {32'hc0d22fe0, 32'h40379ad2} /* (26, 10, 28) {real, imag} */,
  {32'h40eaf63f, 32'hc0b891b7} /* (26, 10, 27) {real, imag} */,
  {32'hc187f7a3, 32'hc0da04f0} /* (26, 10, 26) {real, imag} */,
  {32'hc1098e7b, 32'hc0e4c5fb} /* (26, 10, 25) {real, imag} */,
  {32'hc14d5566, 32'hc1035672} /* (26, 10, 24) {real, imag} */,
  {32'hc09d1f16, 32'h41f6c6fc} /* (26, 10, 23) {real, imag} */,
  {32'h4193a47a, 32'hc153c15d} /* (26, 10, 22) {real, imag} */,
  {32'h40fa354a, 32'hc1173496} /* (26, 10, 21) {real, imag} */,
  {32'hc11c7097, 32'h3fe64184} /* (26, 10, 20) {real, imag} */,
  {32'h4170d5be, 32'h411826d9} /* (26, 10, 19) {real, imag} */,
  {32'hbfc7d13e, 32'h409ceebe} /* (26, 10, 18) {real, imag} */,
  {32'h410358ba, 32'hbf15447a} /* (26, 10, 17) {real, imag} */,
  {32'h4116159a, 32'h40356529} /* (26, 10, 16) {real, imag} */,
  {32'hbf334160, 32'hbfa5b0a4} /* (26, 10, 15) {real, imag} */,
  {32'h41e0c595, 32'h40b12660} /* (26, 10, 14) {real, imag} */,
  {32'hbfb67f98, 32'hc1b1b2a9} /* (26, 10, 13) {real, imag} */,
  {32'hc0966510, 32'h40f4c794} /* (26, 10, 12) {real, imag} */,
  {32'hc0476a06, 32'h41538315} /* (26, 10, 11) {real, imag} */,
  {32'hc150e269, 32'h3fff0b48} /* (26, 10, 10) {real, imag} */,
  {32'hc17351c7, 32'hc1543188} /* (26, 10, 9) {real, imag} */,
  {32'h4189e765, 32'h407944a6} /* (26, 10, 8) {real, imag} */,
  {32'h41920d6b, 32'h3f1a1684} /* (26, 10, 7) {real, imag} */,
  {32'h4119c96f, 32'h4184ff1d} /* (26, 10, 6) {real, imag} */,
  {32'hbf4cb45c, 32'h41667a43} /* (26, 10, 5) {real, imag} */,
  {32'hc081c794, 32'h40f66728} /* (26, 10, 4) {real, imag} */,
  {32'hc0d56b5a, 32'h40a3f062} /* (26, 10, 3) {real, imag} */,
  {32'hc191351a, 32'hbf382150} /* (26, 10, 2) {real, imag} */,
  {32'h3ff37ea0, 32'h40b0a3f2} /* (26, 10, 1) {real, imag} */,
  {32'h40f14cac, 32'h40d9a308} /* (26, 10, 0) {real, imag} */,
  {32'hc0e4b64f, 32'h41e4d6a6} /* (26, 9, 31) {real, imag} */,
  {32'hbffd1028, 32'h41cdfbde} /* (26, 9, 30) {real, imag} */,
  {32'h4127ad28, 32'hc060f3ba} /* (26, 9, 29) {real, imag} */,
  {32'hc142b5a2, 32'hc08fe7a8} /* (26, 9, 28) {real, imag} */,
  {32'h40b887cc, 32'h406dfe79} /* (26, 9, 27) {real, imag} */,
  {32'hc0a33e48, 32'hc13f418b} /* (26, 9, 26) {real, imag} */,
  {32'h400853bc, 32'h40089768} /* (26, 9, 25) {real, imag} */,
  {32'h3fc043ca, 32'hc0b7dd09} /* (26, 9, 24) {real, imag} */,
  {32'hc0aa95a7, 32'h419e7c0c} /* (26, 9, 23) {real, imag} */,
  {32'hc0d000e1, 32'h40c1fcca} /* (26, 9, 22) {real, imag} */,
  {32'hc13b3944, 32'h3fdf0024} /* (26, 9, 21) {real, imag} */,
  {32'hc1798553, 32'h41364fd9} /* (26, 9, 20) {real, imag} */,
  {32'h40e027b4, 32'h3fbd7e40} /* (26, 9, 19) {real, imag} */,
  {32'hbd687780, 32'hbfe918f8} /* (26, 9, 18) {real, imag} */,
  {32'h3f81eb24, 32'hc09f4ecd} /* (26, 9, 17) {real, imag} */,
  {32'h407d3eb4, 32'h40a5602d} /* (26, 9, 16) {real, imag} */,
  {32'hbdf16f80, 32'hc158731b} /* (26, 9, 15) {real, imag} */,
  {32'hc0995e93, 32'h40984899} /* (26, 9, 14) {real, imag} */,
  {32'h3eb09090, 32'h40b20f2b} /* (26, 9, 13) {real, imag} */,
  {32'h408249d4, 32'h3fe07770} /* (26, 9, 12) {real, imag} */,
  {32'h404cd736, 32'h41571efe} /* (26, 9, 11) {real, imag} */,
  {32'hc042a731, 32'h405c49b8} /* (26, 9, 10) {real, imag} */,
  {32'h3e951d80, 32'h40a02954} /* (26, 9, 9) {real, imag} */,
  {32'h3fb37f60, 32'hc1aee746} /* (26, 9, 8) {real, imag} */,
  {32'h40935104, 32'h41491233} /* (26, 9, 7) {real, imag} */,
  {32'h41618bc8, 32'h40fcef79} /* (26, 9, 6) {real, imag} */,
  {32'h415886c1, 32'h41c96e64} /* (26, 9, 5) {real, imag} */,
  {32'h3fed7868, 32'h412ac05d} /* (26, 9, 4) {real, imag} */,
  {32'hc0e035e4, 32'hc0f38ef4} /* (26, 9, 3) {real, imag} */,
  {32'h411e6240, 32'hc181b1d4} /* (26, 9, 2) {real, imag} */,
  {32'h40f66a80, 32'hc183b103} /* (26, 9, 1) {real, imag} */,
  {32'h403e6910, 32'h416234a0} /* (26, 9, 0) {real, imag} */,
  {32'h3fb4f5b8, 32'hc1a0619d} /* (26, 8, 31) {real, imag} */,
  {32'h410146c1, 32'hbf593bc4} /* (26, 8, 30) {real, imag} */,
  {32'hc0e586c8, 32'hc1237e35} /* (26, 8, 29) {real, imag} */,
  {32'hbffc5cf0, 32'h410ba91c} /* (26, 8, 28) {real, imag} */,
  {32'hc1731677, 32'h410b9ed2} /* (26, 8, 27) {real, imag} */,
  {32'hc194bf92, 32'h41a135f8} /* (26, 8, 26) {real, imag} */,
  {32'h40b7418c, 32'hc1115e8f} /* (26, 8, 25) {real, imag} */,
  {32'h41f2ee4d, 32'h40e0e254} /* (26, 8, 24) {real, imag} */,
  {32'hc0e8adf0, 32'hc103859c} /* (26, 8, 23) {real, imag} */,
  {32'h3eb970e0, 32'hc04515ec} /* (26, 8, 22) {real, imag} */,
  {32'h3e445880, 32'hc1575176} /* (26, 8, 21) {real, imag} */,
  {32'h40bfa957, 32'h4132b9f2} /* (26, 8, 20) {real, imag} */,
  {32'hc1947d64, 32'hbfcf93d4} /* (26, 8, 19) {real, imag} */,
  {32'hc0a22ae0, 32'h403c2d25} /* (26, 8, 18) {real, imag} */,
  {32'h3ffd60b4, 32'h41309f67} /* (26, 8, 17) {real, imag} */,
  {32'h407e6c3e, 32'h4053c554} /* (26, 8, 16) {real, imag} */,
  {32'h40f442d3, 32'h3fc8c350} /* (26, 8, 15) {real, imag} */,
  {32'h404f2a30, 32'h40b1f37a} /* (26, 8, 14) {real, imag} */,
  {32'h411836aa, 32'h4091c576} /* (26, 8, 13) {real, imag} */,
  {32'h3f7dd9de, 32'hbfd58734} /* (26, 8, 12) {real, imag} */,
  {32'h4132fe28, 32'hc0dcb0d9} /* (26, 8, 11) {real, imag} */,
  {32'hc16556d4, 32'hc12c036a} /* (26, 8, 10) {real, imag} */,
  {32'h40aedc9c, 32'h40e54afa} /* (26, 8, 9) {real, imag} */,
  {32'hc18c4e9a, 32'hc18c6f4e} /* (26, 8, 8) {real, imag} */,
  {32'h41a85fdd, 32'hc04430ba} /* (26, 8, 7) {real, imag} */,
  {32'h407a1a24, 32'h3efa93c8} /* (26, 8, 6) {real, imag} */,
  {32'h414ffc8f, 32'h3e8a0828} /* (26, 8, 5) {real, imag} */,
  {32'hc1aedd4e, 32'h416dd199} /* (26, 8, 4) {real, imag} */,
  {32'h41cb5d50, 32'h41e64b8a} /* (26, 8, 3) {real, imag} */,
  {32'hc199902f, 32'hc0b16dec} /* (26, 8, 2) {real, imag} */,
  {32'hc06c2ee0, 32'hc0954f88} /* (26, 8, 1) {real, imag} */,
  {32'hc0fb99ca, 32'hc05622e0} /* (26, 8, 0) {real, imag} */,
  {32'hc1cd02ca, 32'h40b1503e} /* (26, 7, 31) {real, imag} */,
  {32'hc0a568ea, 32'hc0be00ce} /* (26, 7, 30) {real, imag} */,
  {32'h4065c368, 32'hc18bdd00} /* (26, 7, 29) {real, imag} */,
  {32'hc0a12fc0, 32'h40824eb0} /* (26, 7, 28) {real, imag} */,
  {32'h417f5eab, 32'h419a7957} /* (26, 7, 27) {real, imag} */,
  {32'hc042a6e4, 32'h419a4a94} /* (26, 7, 26) {real, imag} */,
  {32'h3f05bd58, 32'hc043c430} /* (26, 7, 25) {real, imag} */,
  {32'h41370ab3, 32'hc1dc250c} /* (26, 7, 24) {real, imag} */,
  {32'hc10405ea, 32'h41893669} /* (26, 7, 23) {real, imag} */,
  {32'hbfccaf44, 32'h41858e57} /* (26, 7, 22) {real, imag} */,
  {32'h3ed97660, 32'hc19b5a6c} /* (26, 7, 21) {real, imag} */,
  {32'h41a1a452, 32'h4138a6ea} /* (26, 7, 20) {real, imag} */,
  {32'hc1039bfe, 32'h41233ede} /* (26, 7, 19) {real, imag} */,
  {32'hc14e3674, 32'h41104ae8} /* (26, 7, 18) {real, imag} */,
  {32'hc02c6782, 32'h3f828cae} /* (26, 7, 17) {real, imag} */,
  {32'hc1266cd6, 32'hc039db67} /* (26, 7, 16) {real, imag} */,
  {32'h400bc6b4, 32'h3f94ae44} /* (26, 7, 15) {real, imag} */,
  {32'hc18daa64, 32'hbfe6ab3b} /* (26, 7, 14) {real, imag} */,
  {32'hc0945503, 32'hbfee6d0a} /* (26, 7, 13) {real, imag} */,
  {32'h3f2d3028, 32'hc10aeb84} /* (26, 7, 12) {real, imag} */,
  {32'hc0ca93f0, 32'h4180c998} /* (26, 7, 11) {real, imag} */,
  {32'hc1d5f7ba, 32'hc148deb6} /* (26, 7, 10) {real, imag} */,
  {32'h41715f48, 32'h413859de} /* (26, 7, 9) {real, imag} */,
  {32'h411baaf6, 32'hc19c95f7} /* (26, 7, 8) {real, imag} */,
  {32'hc1210d75, 32'hc1093c50} /* (26, 7, 7) {real, imag} */,
  {32'h41a3e214, 32'h41652827} /* (26, 7, 6) {real, imag} */,
  {32'hc1316552, 32'hc18c6381} /* (26, 7, 5) {real, imag} */,
  {32'h41111ffa, 32'hc20d3dca} /* (26, 7, 4) {real, imag} */,
  {32'h41b61906, 32'hc0815854} /* (26, 7, 3) {real, imag} */,
  {32'h4127aad6, 32'h41a4ae94} /* (26, 7, 2) {real, imag} */,
  {32'h42019004, 32'h41011cea} /* (26, 7, 1) {real, imag} */,
  {32'hc19c5b62, 32'h3f809baa} /* (26, 7, 0) {real, imag} */,
  {32'hc156d6fe, 32'h402291d0} /* (26, 6, 31) {real, imag} */,
  {32'hc1af530d, 32'h4017ec3c} /* (26, 6, 30) {real, imag} */,
  {32'hc011ce2a, 32'h409b32d6} /* (26, 6, 29) {real, imag} */,
  {32'h41356916, 32'hc16319dd} /* (26, 6, 28) {real, imag} */,
  {32'hbfd9ea4c, 32'h3fb8ed48} /* (26, 6, 27) {real, imag} */,
  {32'h3ff6b1a8, 32'h41ad71cd} /* (26, 6, 26) {real, imag} */,
  {32'hc155871f, 32'hc1497a98} /* (26, 6, 25) {real, imag} */,
  {32'h40e9228a, 32'h41fcf696} /* (26, 6, 24) {real, imag} */,
  {32'h3f62ac38, 32'hc03b0c4a} /* (26, 6, 23) {real, imag} */,
  {32'h418a8a17, 32'h411c2d76} /* (26, 6, 22) {real, imag} */,
  {32'h40aa9500, 32'hc037bd48} /* (26, 6, 21) {real, imag} */,
  {32'h4110852e, 32'h40e04f39} /* (26, 6, 20) {real, imag} */,
  {32'hc0ef3dc3, 32'hc136cda9} /* (26, 6, 19) {real, imag} */,
  {32'h40401351, 32'h412ecd0c} /* (26, 6, 18) {real, imag} */,
  {32'hc10e9852, 32'hc155e600} /* (26, 6, 17) {real, imag} */,
  {32'h40d82811, 32'h40258bd4} /* (26, 6, 16) {real, imag} */,
  {32'h40c6ad99, 32'h408c0473} /* (26, 6, 15) {real, imag} */,
  {32'h408e04ee, 32'hbe7fcf08} /* (26, 6, 14) {real, imag} */,
  {32'h414af7d5, 32'hc14b920b} /* (26, 6, 13) {real, imag} */,
  {32'hc15b3124, 32'h41531ff6} /* (26, 6, 12) {real, imag} */,
  {32'h4178b646, 32'hc0927c61} /* (26, 6, 11) {real, imag} */,
  {32'hc09d473b, 32'h3ffeb7f8} /* (26, 6, 10) {real, imag} */,
  {32'h41a2bcbd, 32'hc15876c0} /* (26, 6, 9) {real, imag} */,
  {32'h418e19d2, 32'h41238252} /* (26, 6, 8) {real, imag} */,
  {32'h412518f8, 32'h3f93e8c0} /* (26, 6, 7) {real, imag} */,
  {32'h41908912, 32'hc181811d} /* (26, 6, 6) {real, imag} */,
  {32'h3f9778f8, 32'h4158a6c5} /* (26, 6, 5) {real, imag} */,
  {32'hc0c36798, 32'hc1614baa} /* (26, 6, 4) {real, imag} */,
  {32'h41a137d9, 32'hc1620997} /* (26, 6, 3) {real, imag} */,
  {32'h410e4984, 32'h4000b062} /* (26, 6, 2) {real, imag} */,
  {32'hc0c004ec, 32'h41057943} /* (26, 6, 1) {real, imag} */,
  {32'h41562ce8, 32'hc17b96c0} /* (26, 6, 0) {real, imag} */,
  {32'hc0594940, 32'hc21dd99e} /* (26, 5, 31) {real, imag} */,
  {32'h418ed5a4, 32'hc124b4dc} /* (26, 5, 30) {real, imag} */,
  {32'h41d7bcd2, 32'h4004fff4} /* (26, 5, 29) {real, imag} */,
  {32'hc13bbcf3, 32'h41ae4bd0} /* (26, 5, 28) {real, imag} */,
  {32'hc175a32e, 32'hc122b9dc} /* (26, 5, 27) {real, imag} */,
  {32'h40867d77, 32'hbf9902e2} /* (26, 5, 26) {real, imag} */,
  {32'h3fd23fa2, 32'hc1311360} /* (26, 5, 25) {real, imag} */,
  {32'h3ff8d904, 32'hc0ab74c9} /* (26, 5, 24) {real, imag} */,
  {32'hc1580ee4, 32'h4158e888} /* (26, 5, 23) {real, imag} */,
  {32'h416173d6, 32'hbda24080} /* (26, 5, 22) {real, imag} */,
  {32'h405bec2a, 32'hc14e430a} /* (26, 5, 21) {real, imag} */,
  {32'h419e6ae0, 32'h409c0209} /* (26, 5, 20) {real, imag} */,
  {32'h410ab40e, 32'h417ecbca} /* (26, 5, 19) {real, imag} */,
  {32'h40db013e, 32'hc12715ae} /* (26, 5, 18) {real, imag} */,
  {32'h3f95362c, 32'hc10950ce} /* (26, 5, 17) {real, imag} */,
  {32'hc1434b38, 32'hc17b725a} /* (26, 5, 16) {real, imag} */,
  {32'hc059c69c, 32'h400683e4} /* (26, 5, 15) {real, imag} */,
  {32'hc084cea8, 32'hbef32e20} /* (26, 5, 14) {real, imag} */,
  {32'hc138e9fa, 32'h41744ae4} /* (26, 5, 13) {real, imag} */,
  {32'hc0886714, 32'h3f391f70} /* (26, 5, 12) {real, imag} */,
  {32'h405e159d, 32'h418b5dbe} /* (26, 5, 11) {real, imag} */,
  {32'h411af272, 32'h406562d2} /* (26, 5, 10) {real, imag} */,
  {32'h413be2b8, 32'hbf02f2b0} /* (26, 5, 9) {real, imag} */,
  {32'h41d3f6e6, 32'hc0db83d6} /* (26, 5, 8) {real, imag} */,
  {32'h419a4e22, 32'h416ad4a6} /* (26, 5, 7) {real, imag} */,
  {32'hc1bb1a1a, 32'h4161ca44} /* (26, 5, 6) {real, imag} */,
  {32'h4179b22f, 32'h3fb681c0} /* (26, 5, 5) {real, imag} */,
  {32'hc0714a65, 32'hc100f6d3} /* (26, 5, 4) {real, imag} */,
  {32'hc1661926, 32'hc1baee14} /* (26, 5, 3) {real, imag} */,
  {32'hc19275bd, 32'hc1367f6a} /* (26, 5, 2) {real, imag} */,
  {32'hc20a3bc1, 32'h41224b98} /* (26, 5, 1) {real, imag} */,
  {32'hc2569100, 32'h41a4f675} /* (26, 5, 0) {real, imag} */,
  {32'hc145a5e2, 32'hc0069b28} /* (26, 4, 31) {real, imag} */,
  {32'hc135daee, 32'hc08d1a58} /* (26, 4, 30) {real, imag} */,
  {32'hc1c4089d, 32'h4022a804} /* (26, 4, 29) {real, imag} */,
  {32'h3f3463f0, 32'hc12af775} /* (26, 4, 28) {real, imag} */,
  {32'h3f7b8754, 32'h408909d3} /* (26, 4, 27) {real, imag} */,
  {32'hc1c05772, 32'hc15577c5} /* (26, 4, 26) {real, imag} */,
  {32'hbfbbdcce, 32'h4216858b} /* (26, 4, 25) {real, imag} */,
  {32'h4035ab34, 32'hc1327150} /* (26, 4, 24) {real, imag} */,
  {32'hbdbba040, 32'h410e73ad} /* (26, 4, 23) {real, imag} */,
  {32'h41bacb31, 32'h410cd3cf} /* (26, 4, 22) {real, imag} */,
  {32'hc0a71056, 32'h41a2e4f0} /* (26, 4, 21) {real, imag} */,
  {32'h40a03a5c, 32'h401e0994} /* (26, 4, 20) {real, imag} */,
  {32'hbed4757e, 32'hc0cb3a8b} /* (26, 4, 19) {real, imag} */,
  {32'hc19eec98, 32'hc1103573} /* (26, 4, 18) {real, imag} */,
  {32'h40b946b8, 32'hbfc985fc} /* (26, 4, 17) {real, imag} */,
  {32'hc095c904, 32'hbfbce1d4} /* (26, 4, 16) {real, imag} */,
  {32'hc1750474, 32'hc0858686} /* (26, 4, 15) {real, imag} */,
  {32'hc1035352, 32'h3fbcd410} /* (26, 4, 14) {real, imag} */,
  {32'h4044e50e, 32'h41386426} /* (26, 4, 13) {real, imag} */,
  {32'hc13ca03f, 32'hc117b227} /* (26, 4, 12) {real, imag} */,
  {32'h41a55f87, 32'h41192c14} /* (26, 4, 11) {real, imag} */,
  {32'h40856319, 32'hc0a61476} /* (26, 4, 10) {real, imag} */,
  {32'hc0ba6adf, 32'h4046e62c} /* (26, 4, 9) {real, imag} */,
  {32'h400c760c, 32'hc1108507} /* (26, 4, 8) {real, imag} */,
  {32'hc020d54c, 32'h414a25f4} /* (26, 4, 7) {real, imag} */,
  {32'hc1978266, 32'h411c6e08} /* (26, 4, 6) {real, imag} */,
  {32'h415aaf09, 32'hbfafaf24} /* (26, 4, 5) {real, imag} */,
  {32'h41ae8843, 32'hc1e872be} /* (26, 4, 4) {real, imag} */,
  {32'hc04716f6, 32'hc08587e6} /* (26, 4, 3) {real, imag} */,
  {32'hc1673dec, 32'hc088d008} /* (26, 4, 2) {real, imag} */,
  {32'h41580fc8, 32'h4135c77a} /* (26, 4, 1) {real, imag} */,
  {32'hc1ac42ca, 32'hc1fc5812} /* (26, 4, 0) {real, imag} */,
  {32'hc1d7bc14, 32'h40917fc8} /* (26, 3, 31) {real, imag} */,
  {32'h42490e17, 32'hc15f3e10} /* (26, 3, 30) {real, imag} */,
  {32'h412bdac1, 32'h4004177e} /* (26, 3, 29) {real, imag} */,
  {32'h419f5ad8, 32'h418a913f} /* (26, 3, 28) {real, imag} */,
  {32'hc016b900, 32'hc0f044af} /* (26, 3, 27) {real, imag} */,
  {32'hc1294fdf, 32'h415d9480} /* (26, 3, 26) {real, imag} */,
  {32'hc1af19f9, 32'h3f8f2c90} /* (26, 3, 25) {real, imag} */,
  {32'hc0e0c97e, 32'hc13a0988} /* (26, 3, 24) {real, imag} */,
  {32'h40c392fb, 32'hc11680ba} /* (26, 3, 23) {real, imag} */,
  {32'hc003b432, 32'h40abd33f} /* (26, 3, 22) {real, imag} */,
  {32'h3f1af8c0, 32'h40a9174a} /* (26, 3, 21) {real, imag} */,
  {32'hc137af6a, 32'hc073e51a} /* (26, 3, 20) {real, imag} */,
  {32'h4143a574, 32'hc0cc9c4c} /* (26, 3, 19) {real, imag} */,
  {32'hc128e9d6, 32'hc19d1ad3} /* (26, 3, 18) {real, imag} */,
  {32'h419344da, 32'h40d2d840} /* (26, 3, 17) {real, imag} */,
  {32'h40876e9e, 32'h410184ef} /* (26, 3, 16) {real, imag} */,
  {32'hc090ab61, 32'hc0ce1dc2} /* (26, 3, 15) {real, imag} */,
  {32'h404c7684, 32'h418498f4} /* (26, 3, 14) {real, imag} */,
  {32'h41211535, 32'hc18d7278} /* (26, 3, 13) {real, imag} */,
  {32'h40fe260e, 32'hc1172ce0} /* (26, 3, 12) {real, imag} */,
  {32'h40001bc2, 32'hc0a36302} /* (26, 3, 11) {real, imag} */,
  {32'hc108d650, 32'hc044720a} /* (26, 3, 10) {real, imag} */,
  {32'hc08c4b2c, 32'hc0fe9390} /* (26, 3, 9) {real, imag} */,
  {32'hc0eee221, 32'hc14d4281} /* (26, 3, 8) {real, imag} */,
  {32'hc076243c, 32'h416a9a5a} /* (26, 3, 7) {real, imag} */,
  {32'hc168f290, 32'h415bf076} /* (26, 3, 6) {real, imag} */,
  {32'hc1703418, 32'h4159f036} /* (26, 3, 5) {real, imag} */,
  {32'hc0befcea, 32'h4164205d} /* (26, 3, 4) {real, imag} */,
  {32'hc1829350, 32'hbf5002e0} /* (26, 3, 3) {real, imag} */,
  {32'h41d2df75, 32'hc0f5bf94} /* (26, 3, 2) {real, imag} */,
  {32'hc0603680, 32'h4294a578} /* (26, 3, 1) {real, imag} */,
  {32'h429e92db, 32'h41fd20d5} /* (26, 3, 0) {real, imag} */,
  {32'h41b5c9e0, 32'h427760bc} /* (26, 2, 31) {real, imag} */,
  {32'h4262fe10, 32'hc27918f2} /* (26, 2, 30) {real, imag} */,
  {32'hc134a8ec, 32'hc0e8e93e} /* (26, 2, 29) {real, imag} */,
  {32'hc141df94, 32'h4133531a} /* (26, 2, 28) {real, imag} */,
  {32'h41eb715f, 32'hc1bef157} /* (26, 2, 27) {real, imag} */,
  {32'h40b4bb75, 32'h415f0e50} /* (26, 2, 26) {real, imag} */,
  {32'hc0bffe56, 32'h4221b930} /* (26, 2, 25) {real, imag} */,
  {32'h41aafec6, 32'h4128d31d} /* (26, 2, 24) {real, imag} */,
  {32'h41e5fcf9, 32'hc16ee2d3} /* (26, 2, 23) {real, imag} */,
  {32'hc1406eb2, 32'hc036331e} /* (26, 2, 22) {real, imag} */,
  {32'h40839c7c, 32'h3fbffd80} /* (26, 2, 21) {real, imag} */,
  {32'hc0f0bd3f, 32'hbef38940} /* (26, 2, 20) {real, imag} */,
  {32'hc0f66dda, 32'hbf8b2cb8} /* (26, 2, 19) {real, imag} */,
  {32'h411b1964, 32'h4140c8cf} /* (26, 2, 18) {real, imag} */,
  {32'h411aa0ae, 32'h40fdfd77} /* (26, 2, 17) {real, imag} */,
  {32'h401e675e, 32'h40b9f76d} /* (26, 2, 16) {real, imag} */,
  {32'hbf6ed506, 32'hc0c48894} /* (26, 2, 15) {real, imag} */,
  {32'hc0826a38, 32'hc0eaaffa} /* (26, 2, 14) {real, imag} */,
  {32'hc06fe79e, 32'h3ff90ac2} /* (26, 2, 13) {real, imag} */,
  {32'h40b793f8, 32'h40079494} /* (26, 2, 12) {real, imag} */,
  {32'h415ede48, 32'h410115e9} /* (26, 2, 11) {real, imag} */,
  {32'h3edb00b0, 32'h4019b554} /* (26, 2, 10) {real, imag} */,
  {32'hc194259f, 32'hc152f550} /* (26, 2, 9) {real, imag} */,
  {32'hc0945796, 32'h41a8f5c5} /* (26, 2, 8) {real, imag} */,
  {32'h40cef612, 32'h41c366d6} /* (26, 2, 7) {real, imag} */,
  {32'h41609cbe, 32'h40c3c967} /* (26, 2, 6) {real, imag} */,
  {32'hc193011d, 32'h422263f2} /* (26, 2, 5) {real, imag} */,
  {32'hc1914d0c, 32'hc214c973} /* (26, 2, 4) {real, imag} */,
  {32'hc1f537d2, 32'hc135a3bb} /* (26, 2, 3) {real, imag} */,
  {32'h42861f12, 32'hc1dc8ee8} /* (26, 2, 2) {real, imag} */,
  {32'h40b59680, 32'h4288b118} /* (26, 2, 1) {real, imag} */,
  {32'h4253d7cc, 32'hc28b7808} /* (26, 2, 0) {real, imag} */,
  {32'hc356de14, 32'h400695e0} /* (26, 1, 31) {real, imag} */,
  {32'h417a1570, 32'h42d8bf26} /* (26, 1, 30) {real, imag} */,
  {32'h40e986d4, 32'hbfc90a00} /* (26, 1, 29) {real, imag} */,
  {32'hc169817a, 32'h41941052} /* (26, 1, 28) {real, imag} */,
  {32'hc1947850, 32'hbe416300} /* (26, 1, 27) {real, imag} */,
  {32'hc1d60d2d, 32'hc101b218} /* (26, 1, 26) {real, imag} */,
  {32'hc0cce52e, 32'hc128f8e9} /* (26, 1, 25) {real, imag} */,
  {32'h41057d44, 32'hc08516f1} /* (26, 1, 24) {real, imag} */,
  {32'h410e2b92, 32'h3e7921c0} /* (26, 1, 23) {real, imag} */,
  {32'h40013678, 32'h40a848ee} /* (26, 1, 22) {real, imag} */,
  {32'hbfe5da08, 32'hc1355303} /* (26, 1, 21) {real, imag} */,
  {32'h4139e5a6, 32'h4188db82} /* (26, 1, 20) {real, imag} */,
  {32'h41850d11, 32'hc0be3764} /* (26, 1, 19) {real, imag} */,
  {32'h41303ef8, 32'h3fb5c9a4} /* (26, 1, 18) {real, imag} */,
  {32'h4083bd20, 32'hc0fc0667} /* (26, 1, 17) {real, imag} */,
  {32'hc0ff199a, 32'hbfea115d} /* (26, 1, 16) {real, imag} */,
  {32'hbde4a4c0, 32'hbf880bcc} /* (26, 1, 15) {real, imag} */,
  {32'h407e397a, 32'hc0a3ba98} /* (26, 1, 14) {real, imag} */,
  {32'h41d95d35, 32'h40929d18} /* (26, 1, 13) {real, imag} */,
  {32'h410907c2, 32'h414a5faa} /* (26, 1, 12) {real, imag} */,
  {32'hc19d1598, 32'h3f832e10} /* (26, 1, 11) {real, imag} */,
  {32'hc1dccbee, 32'h3ec83278} /* (26, 1, 10) {real, imag} */,
  {32'hc1ae7514, 32'h3f943fe0} /* (26, 1, 9) {real, imag} */,
  {32'hc12b1098, 32'hc19a6005} /* (26, 1, 8) {real, imag} */,
  {32'h41369168, 32'h41a6c130} /* (26, 1, 7) {real, imag} */,
  {32'h416f0c36, 32'hc02ae662} /* (26, 1, 6) {real, imag} */,
  {32'h3fef3620, 32'h41247a2e} /* (26, 1, 5) {real, imag} */,
  {32'hc192dc72, 32'hc180c656} /* (26, 1, 4) {real, imag} */,
  {32'h3e67c600, 32'hc1b30c6c} /* (26, 1, 3) {real, imag} */,
  {32'hc1fce798, 32'hc20169f4} /* (26, 1, 2) {real, imag} */,
  {32'hc3910940, 32'hc35c801d} /* (26, 1, 1) {real, imag} */,
  {32'hc3e8fd6c, 32'hc2d3370a} /* (26, 1, 0) {real, imag} */,
  {32'hc3d295f2, 32'h43aab656} /* (26, 0, 31) {real, imag} */,
  {32'hc1af3b58, 32'h42a48ee9} /* (26, 0, 30) {real, imag} */,
  {32'h416f01e6, 32'hc230bae8} /* (26, 0, 29) {real, imag} */,
  {32'h4221e952, 32'hc13e3a2c} /* (26, 0, 28) {real, imag} */,
  {32'hc0404dc0, 32'h40f4e91e} /* (26, 0, 27) {real, imag} */,
  {32'h41a8150f, 32'hc08dcab4} /* (26, 0, 26) {real, imag} */,
  {32'h411e15f6, 32'hc102dc65} /* (26, 0, 25) {real, imag} */,
  {32'h4098ebc2, 32'hc1db92e7} /* (26, 0, 24) {real, imag} */,
  {32'hc19a73f1, 32'hc071062f} /* (26, 0, 23) {real, imag} */,
  {32'hc13f310c, 32'h4150c886} /* (26, 0, 22) {real, imag} */,
  {32'hc0488daa, 32'h41a3c9df} /* (26, 0, 21) {real, imag} */,
  {32'hbef053d0, 32'hc1251f12} /* (26, 0, 20) {real, imag} */,
  {32'hc0e46985, 32'hc032e116} /* (26, 0, 19) {real, imag} */,
  {32'h40999450, 32'h40915b58} /* (26, 0, 18) {real, imag} */,
  {32'h4091214c, 32'h3fd5a837} /* (26, 0, 17) {real, imag} */,
  {32'h41bfb9f6, 32'h00000000} /* (26, 0, 16) {real, imag} */,
  {32'h4091214c, 32'hbfd5a837} /* (26, 0, 15) {real, imag} */,
  {32'h40999450, 32'hc0915b58} /* (26, 0, 14) {real, imag} */,
  {32'hc0e46985, 32'h4032e116} /* (26, 0, 13) {real, imag} */,
  {32'hbef053d0, 32'h41251f12} /* (26, 0, 12) {real, imag} */,
  {32'hc0488daa, 32'hc1a3c9df} /* (26, 0, 11) {real, imag} */,
  {32'hc13f310c, 32'hc150c886} /* (26, 0, 10) {real, imag} */,
  {32'hc19a73f1, 32'h4071062f} /* (26, 0, 9) {real, imag} */,
  {32'h4098ebc2, 32'h41db92e7} /* (26, 0, 8) {real, imag} */,
  {32'h411e15f6, 32'h4102dc65} /* (26, 0, 7) {real, imag} */,
  {32'h41a8150f, 32'h408dcab4} /* (26, 0, 6) {real, imag} */,
  {32'hc0404dc0, 32'hc0f4e91e} /* (26, 0, 5) {real, imag} */,
  {32'h4221e952, 32'h413e3a2c} /* (26, 0, 4) {real, imag} */,
  {32'h416f01e6, 32'h4230bae8} /* (26, 0, 3) {real, imag} */,
  {32'hc1af3b58, 32'hc2a48ee9} /* (26, 0, 2) {real, imag} */,
  {32'hc3d295f2, 32'hc3aab656} /* (26, 0, 1) {real, imag} */,
  {32'hc46c0ae3, 32'h00000000} /* (26, 0, 0) {real, imag} */,
  {32'hc4924069, 32'h442ea98b} /* (25, 31, 31) {real, imag} */,
  {32'h438543ce, 32'hc38875b1} /* (25, 31, 30) {real, imag} */,
  {32'h421710a7, 32'h3fa5f380} /* (25, 31, 29) {real, imag} */,
  {32'hc00a35c0, 32'h42753126} /* (25, 31, 28) {real, imag} */,
  {32'h42405e16, 32'hc2357b70} /* (25, 31, 27) {real, imag} */,
  {32'h416f6cb3, 32'hc17e8b53} /* (25, 31, 26) {real, imag} */,
  {32'hc081714b, 32'hc0348370} /* (25, 31, 25) {real, imag} */,
  {32'h4103e51f, 32'hc1fb5807} /* (25, 31, 24) {real, imag} */,
  {32'h410b0e3d, 32'h410b89ba} /* (25, 31, 23) {real, imag} */,
  {32'h40b89066, 32'hbfabb4a8} /* (25, 31, 22) {real, imag} */,
  {32'h41442a38, 32'hc1c83c00} /* (25, 31, 21) {real, imag} */,
  {32'hbfb74e4e, 32'hbfe4efcc} /* (25, 31, 20) {real, imag} */,
  {32'h40d69b90, 32'h40ea93da} /* (25, 31, 19) {real, imag} */,
  {32'hc13aaa8d, 32'hc170d1e0} /* (25, 31, 18) {real, imag} */,
  {32'hc123ad74, 32'h416b3d5f} /* (25, 31, 17) {real, imag} */,
  {32'h401de935, 32'hc12cee39} /* (25, 31, 16) {real, imag} */,
  {32'hc05d30c6, 32'hc09e5d68} /* (25, 31, 15) {real, imag} */,
  {32'h40ce2313, 32'h4187981c} /* (25, 31, 14) {real, imag} */,
  {32'hc0bbd3fd, 32'h3f673428} /* (25, 31, 13) {real, imag} */,
  {32'h414f9a2e, 32'h40755af7} /* (25, 31, 12) {real, imag} */,
  {32'h41c12222, 32'h41721ba8} /* (25, 31, 11) {real, imag} */,
  {32'hbfe8b750, 32'h4187fb38} /* (25, 31, 10) {real, imag} */,
  {32'h400856a9, 32'hc172155e} /* (25, 31, 9) {real, imag} */,
  {32'h3fee04f0, 32'h3fbb3408} /* (25, 31, 8) {real, imag} */,
  {32'hc180ef26, 32'hc1283732} /* (25, 31, 7) {real, imag} */,
  {32'hc1b494fb, 32'h40abd18c} /* (25, 31, 6) {real, imag} */,
  {32'h42878014, 32'h414e00d6} /* (25, 31, 5) {real, imag} */,
  {32'hc223353e, 32'h41c8d99e} /* (25, 31, 4) {real, imag} */,
  {32'h41d217c5, 32'h41afe7c8} /* (25, 31, 3) {real, imag} */,
  {32'h433c3442, 32'hc2dfe528} /* (25, 31, 2) {real, imag} */,
  {32'hc4464ef4, 32'hc3323f18} /* (25, 31, 1) {real, imag} */,
  {32'hc493f352, 32'h433fcf31} /* (25, 31, 0) {real, imag} */,
  {32'h43b1396f, 32'hc18b3d40} /* (25, 30, 31) {real, imag} */,
  {32'hc32b65b9, 32'hc2135d2d} /* (25, 30, 30) {real, imag} */,
  {32'hc19386fb, 32'h40f806b4} /* (25, 30, 29) {real, imag} */,
  {32'h42430485, 32'h404e70f4} /* (25, 30, 28) {real, imag} */,
  {32'hc28778e3, 32'h420769b3} /* (25, 30, 27) {real, imag} */,
  {32'hc0a2a9fe, 32'h4143250d} /* (25, 30, 26) {real, imag} */,
  {32'h41ea4924, 32'hc169d390} /* (25, 30, 25) {real, imag} */,
  {32'hc187854d, 32'h40d87b6e} /* (25, 30, 24) {real, imag} */,
  {32'hbfab8274, 32'h416cc5f6} /* (25, 30, 23) {real, imag} */,
  {32'h415f2f14, 32'hc1060087} /* (25, 30, 22) {real, imag} */,
  {32'hc0da26df, 32'h41eec50f} /* (25, 30, 21) {real, imag} */,
  {32'hbfb3a4a8, 32'h4195536b} /* (25, 30, 20) {real, imag} */,
  {32'h4109a426, 32'hbf97197c} /* (25, 30, 19) {real, imag} */,
  {32'hbfe7cd48, 32'hc1503225} /* (25, 30, 18) {real, imag} */,
  {32'h40e0c574, 32'hc09a5ed1} /* (25, 30, 17) {real, imag} */,
  {32'hc0ea1156, 32'hc0cd9fe1} /* (25, 30, 16) {real, imag} */,
  {32'hc0d48374, 32'h414ddffa} /* (25, 30, 15) {real, imag} */,
  {32'hc0a3d4f4, 32'hc0f016c0} /* (25, 30, 14) {real, imag} */,
  {32'h3f2437cc, 32'hbff024f4} /* (25, 30, 13) {real, imag} */,
  {32'hbe8bf2b0, 32'h40f39ca0} /* (25, 30, 12) {real, imag} */,
  {32'hc037db4a, 32'h4116d028} /* (25, 30, 11) {real, imag} */,
  {32'h40f07241, 32'h41c87158} /* (25, 30, 10) {real, imag} */,
  {32'h410fe85f, 32'hbf223f38} /* (25, 30, 9) {real, imag} */,
  {32'hc14ca1ad, 32'hc2022582} /* (25, 30, 8) {real, imag} */,
  {32'hbbaf1800, 32'hc1f92af4} /* (25, 30, 7) {real, imag} */,
  {32'h40c8d3e0, 32'hbf4123f0} /* (25, 30, 6) {real, imag} */,
  {32'h3f98c7f0, 32'h4152c160} /* (25, 30, 5) {real, imag} */,
  {32'h4200646f, 32'h421d9bb9} /* (25, 30, 4) {real, imag} */,
  {32'h41cb205e, 32'h41e52d8e} /* (25, 30, 3) {real, imag} */,
  {32'hc38b0d3a, 32'hc24b1585} /* (25, 30, 2) {real, imag} */,
  {32'h44124ac2, 32'hc2974649} /* (25, 30, 1) {real, imag} */,
  {32'h43af9197, 32'hc1a1350c} /* (25, 30, 0) {real, imag} */,
  {32'hc2b703a1, 32'h423c75bf} /* (25, 29, 31) {real, imag} */,
  {32'h40c3a557, 32'hc2bcd155} /* (25, 29, 30) {real, imag} */,
  {32'hc00c1486, 32'h418dcfcd} /* (25, 29, 29) {real, imag} */,
  {32'h41c5d2e2, 32'h40a516c8} /* (25, 29, 28) {real, imag} */,
  {32'hc1d2fc5e, 32'h4175dcd8} /* (25, 29, 27) {real, imag} */,
  {32'hc03549d8, 32'hc18e9266} /* (25, 29, 26) {real, imag} */,
  {32'hc0c2ff4c, 32'hbf8d42be} /* (25, 29, 25) {real, imag} */,
  {32'hc13b0c1e, 32'h4104cd56} /* (25, 29, 24) {real, imag} */,
  {32'hc0083f66, 32'h40ea6a4a} /* (25, 29, 23) {real, imag} */,
  {32'hbfea2caa, 32'hc03e7304} /* (25, 29, 22) {real, imag} */,
  {32'hc18a8f00, 32'h40529ac4} /* (25, 29, 21) {real, imag} */,
  {32'h4148094d, 32'h40a5df7a} /* (25, 29, 20) {real, imag} */,
  {32'h403f0a54, 32'hc103a276} /* (25, 29, 19) {real, imag} */,
  {32'hc16609ca, 32'h405111b2} /* (25, 29, 18) {real, imag} */,
  {32'h4061958c, 32'hc026a4b7} /* (25, 29, 17) {real, imag} */,
  {32'hc0d9fbd5, 32'hc0cecdf1} /* (25, 29, 16) {real, imag} */,
  {32'h3e0c44b8, 32'h40b46f5d} /* (25, 29, 15) {real, imag} */,
  {32'h41191012, 32'hc0b9eeae} /* (25, 29, 14) {real, imag} */,
  {32'h4148745a, 32'h40afd396} /* (25, 29, 13) {real, imag} */,
  {32'hc03f1ab9, 32'hc12ed7a0} /* (25, 29, 12) {real, imag} */,
  {32'hbf8d6c22, 32'hc0c910e0} /* (25, 29, 11) {real, imag} */,
  {32'hc08e16be, 32'hc0e9ba4a} /* (25, 29, 10) {real, imag} */,
  {32'h407369b4, 32'h41692c34} /* (25, 29, 9) {real, imag} */,
  {32'h415e588d, 32'hc1db916c} /* (25, 29, 8) {real, imag} */,
  {32'h40c9f958, 32'hc109e0fa} /* (25, 29, 7) {real, imag} */,
  {32'hbf2b5230, 32'hc0d4ba12} /* (25, 29, 6) {real, imag} */,
  {32'h416abea8, 32'h401821e8} /* (25, 29, 5) {real, imag} */,
  {32'hc1ce4370, 32'h41a08bd4} /* (25, 29, 4) {real, imag} */,
  {32'h41addf9e, 32'hc1580e26} /* (25, 29, 3) {real, imag} */,
  {32'hc123e0a8, 32'hc26bde3d} /* (25, 29, 2) {real, imag} */,
  {32'h428d6642, 32'h429f3f28} /* (25, 29, 1) {real, imag} */,
  {32'h429cc1ef, 32'hc19c36dc} /* (25, 29, 0) {real, imag} */,
  {32'hc2e053b4, 32'h4181c330} /* (25, 28, 31) {real, imag} */,
  {32'h4264ec3e, 32'hc24350b5} /* (25, 28, 30) {real, imag} */,
  {32'hc0a4025c, 32'h407dc67a} /* (25, 28, 29) {real, imag} */,
  {32'h4111834b, 32'h427eae9b} /* (25, 28, 28) {real, imag} */,
  {32'h4116da0c, 32'hbe118b80} /* (25, 28, 27) {real, imag} */,
  {32'hc1cd1b52, 32'hc1d36dd4} /* (25, 28, 26) {real, imag} */,
  {32'hc1b7d815, 32'hc11fd46d} /* (25, 28, 25) {real, imag} */,
  {32'h417b6267, 32'hc1f982f6} /* (25, 28, 24) {real, imag} */,
  {32'hc0f4b68c, 32'hc13c036e} /* (25, 28, 23) {real, imag} */,
  {32'h40180685, 32'h409312d3} /* (25, 28, 22) {real, imag} */,
  {32'h412afa78, 32'hc1ae7fa2} /* (25, 28, 21) {real, imag} */,
  {32'h40251f20, 32'h3f5f4f30} /* (25, 28, 20) {real, imag} */,
  {32'h410253f6, 32'hc0e1c37c} /* (25, 28, 19) {real, imag} */,
  {32'h3ff3a3e0, 32'h407f2100} /* (25, 28, 18) {real, imag} */,
  {32'hc0b41313, 32'h3fabce2c} /* (25, 28, 17) {real, imag} */,
  {32'hbefc99fe, 32'hc0bab18a} /* (25, 28, 16) {real, imag} */,
  {32'h3fc5be7c, 32'hc0e8a313} /* (25, 28, 15) {real, imag} */,
  {32'h418e9bee, 32'h4093e7d0} /* (25, 28, 14) {real, imag} */,
  {32'hc0e53144, 32'hc1067ab2} /* (25, 28, 13) {real, imag} */,
  {32'h3fe96b78, 32'h3ec33560} /* (25, 28, 12) {real, imag} */,
  {32'h40e2c443, 32'hc1853101} /* (25, 28, 11) {real, imag} */,
  {32'hc13a97a6, 32'h40acdbc0} /* (25, 28, 10) {real, imag} */,
  {32'hc090bfea, 32'h40e6ab51} /* (25, 28, 9) {real, imag} */,
  {32'h3f10c830, 32'hc068e8d0} /* (25, 28, 8) {real, imag} */,
  {32'h410a4d82, 32'hc11e4403} /* (25, 28, 7) {real, imag} */,
  {32'hc078bcd8, 32'h41d79b3c} /* (25, 28, 6) {real, imag} */,
  {32'h40c167df, 32'h3ecb2e10} /* (25, 28, 5) {real, imag} */,
  {32'hc209d772, 32'h421a93f5} /* (25, 28, 4) {real, imag} */,
  {32'hc19e76c3, 32'h40f55a6e} /* (25, 28, 3) {real, imag} */,
  {32'h422bde28, 32'hc292508d} /* (25, 28, 2) {real, imag} */,
  {32'hc20b4cb0, 32'h428ba980} /* (25, 28, 1) {real, imag} */,
  {32'hc24a60d6, 32'h42174fad} /* (25, 28, 0) {real, imag} */,
  {32'h42388489, 32'hc29edf1e} /* (25, 27, 31) {real, imag} */,
  {32'hc20556c6, 32'h4228ec60} /* (25, 27, 30) {real, imag} */,
  {32'h3f711870, 32'h4202c8a4} /* (25, 27, 29) {real, imag} */,
  {32'hc1381486, 32'hc1595528} /* (25, 27, 28) {real, imag} */,
  {32'h41e5cf84, 32'h41176e91} /* (25, 27, 27) {real, imag} */,
  {32'hc040d3c8, 32'hc09cdadc} /* (25, 27, 26) {real, imag} */,
  {32'h4117b582, 32'hc1027211} /* (25, 27, 25) {real, imag} */,
  {32'hc028b09c, 32'h40038a04} /* (25, 27, 24) {real, imag} */,
  {32'hc18dab18, 32'h413fb2b6} /* (25, 27, 23) {real, imag} */,
  {32'h3fde39b0, 32'h416d6cd6} /* (25, 27, 22) {real, imag} */,
  {32'hc04ce098, 32'h41b890b6} /* (25, 27, 21) {real, imag} */,
  {32'h3f9fd11a, 32'hc0ff99e8} /* (25, 27, 20) {real, imag} */,
  {32'hbe169f78, 32'hc0dbadc2} /* (25, 27, 19) {real, imag} */,
  {32'h40a8aa02, 32'hc1004d78} /* (25, 27, 18) {real, imag} */,
  {32'hc058e84e, 32'hc1493f97} /* (25, 27, 17) {real, imag} */,
  {32'h3fcf91ec, 32'hbf0a0bb8} /* (25, 27, 16) {real, imag} */,
  {32'hc1669352, 32'h400d9da0} /* (25, 27, 15) {real, imag} */,
  {32'hc0205594, 32'hc156eca8} /* (25, 27, 14) {real, imag} */,
  {32'h4135ffe8, 32'hc04797a1} /* (25, 27, 13) {real, imag} */,
  {32'h4164da6b, 32'hc0975e26} /* (25, 27, 12) {real, imag} */,
  {32'hc171087e, 32'h3f3e75d8} /* (25, 27, 11) {real, imag} */,
  {32'h40ac70bd, 32'hc0d3b53e} /* (25, 27, 10) {real, imag} */,
  {32'hc0886c84, 32'h4109edc8} /* (25, 27, 9) {real, imag} */,
  {32'hc0a08e68, 32'hc1477fd0} /* (25, 27, 8) {real, imag} */,
  {32'h419d87ad, 32'h416c0be0} /* (25, 27, 7) {real, imag} */,
  {32'h41ba2781, 32'h414dc8c2} /* (25, 27, 6) {real, imag} */,
  {32'hc223f762, 32'hc0ee848c} /* (25, 27, 5) {real, imag} */,
  {32'h40941bb5, 32'hc17b89ec} /* (25, 27, 4) {real, imag} */,
  {32'h41391df4, 32'h40e3ff62} /* (25, 27, 3) {real, imag} */,
  {32'hc2079cda, 32'h41d87950} /* (25, 27, 2) {real, imag} */,
  {32'h42a8f802, 32'h4184a4e4} /* (25, 27, 1) {real, imag} */,
  {32'h4209b2dc, 32'hc24b057a} /* (25, 27, 0) {real, imag} */,
  {32'hc09640a1, 32'hc0b98f75} /* (25, 26, 31) {real, imag} */,
  {32'h41c32d6e, 32'h4084b04c} /* (25, 26, 30) {real, imag} */,
  {32'h40a5fac4, 32'h40880ab0} /* (25, 26, 29) {real, imag} */,
  {32'h40c9778e, 32'h41bc6d8d} /* (25, 26, 28) {real, imag} */,
  {32'h4094659c, 32'h3f39a474} /* (25, 26, 27) {real, imag} */,
  {32'h415f8948, 32'h413474fc} /* (25, 26, 26) {real, imag} */,
  {32'hc196d020, 32'h40da20bc} /* (25, 26, 25) {real, imag} */,
  {32'h4188e4c9, 32'hc10a2690} /* (25, 26, 24) {real, imag} */,
  {32'h4115293a, 32'hbfd1856e} /* (25, 26, 23) {real, imag} */,
  {32'h418a54e5, 32'hc0ccf76c} /* (25, 26, 22) {real, imag} */,
  {32'hc0d28e72, 32'h403eab44} /* (25, 26, 21) {real, imag} */,
  {32'hbf489ac8, 32'hbfa0caa0} /* (25, 26, 20) {real, imag} */,
  {32'h4158a848, 32'h40f042f2} /* (25, 26, 19) {real, imag} */,
  {32'hc0d180a6, 32'hc06e0796} /* (25, 26, 18) {real, imag} */,
  {32'hbe800178, 32'hc14e1e4e} /* (25, 26, 17) {real, imag} */,
  {32'h417b1526, 32'hbef9ddf0} /* (25, 26, 16) {real, imag} */,
  {32'h409b5be2, 32'h40029d40} /* (25, 26, 15) {real, imag} */,
  {32'hc0e17fd8, 32'hbf117988} /* (25, 26, 14) {real, imag} */,
  {32'hc0d25501, 32'h40a4ee69} /* (25, 26, 13) {real, imag} */,
  {32'h4126afd0, 32'h4033dab0} /* (25, 26, 12) {real, imag} */,
  {32'h40951cbb, 32'h40a12a8a} /* (25, 26, 11) {real, imag} */,
  {32'h40a5008c, 32'hc13060ff} /* (25, 26, 10) {real, imag} */,
  {32'h40e7204d, 32'hc1841b3f} /* (25, 26, 9) {real, imag} */,
  {32'h4094aca2, 32'h40a33576} /* (25, 26, 8) {real, imag} */,
  {32'hc0a6f290, 32'hc1183f23} /* (25, 26, 7) {real, imag} */,
  {32'hc0a827f4, 32'hc1f9ee26} /* (25, 26, 6) {real, imag} */,
  {32'hc0aad513, 32'h4141be39} /* (25, 26, 5) {real, imag} */,
  {32'h41c482ea, 32'h41bcf13c} /* (25, 26, 4) {real, imag} */,
  {32'hc0f522e7, 32'hc07e53f2} /* (25, 26, 3) {real, imag} */,
  {32'hc1789a47, 32'hc16784f3} /* (25, 26, 2) {real, imag} */,
  {32'h412161d2, 32'h41495ee7} /* (25, 26, 1) {real, imag} */,
  {32'h4009d972, 32'hbf520d00} /* (25, 26, 0) {real, imag} */,
  {32'hc1d708f7, 32'h41a0f6b1} /* (25, 25, 31) {real, imag} */,
  {32'h400180a4, 32'hc1d14108} /* (25, 25, 30) {real, imag} */,
  {32'h40fe936a, 32'hc1d584cc} /* (25, 25, 29) {real, imag} */,
  {32'h41a2fe4c, 32'h41b202f3} /* (25, 25, 28) {real, imag} */,
  {32'hc18c5bf6, 32'hc1528bfe} /* (25, 25, 27) {real, imag} */,
  {32'hc145a902, 32'h3ea7a840} /* (25, 25, 26) {real, imag} */,
  {32'h40522f0c, 32'h4140a940} /* (25, 25, 25) {real, imag} */,
  {32'h409f565b, 32'hc0f4d1f4} /* (25, 25, 24) {real, imag} */,
  {32'hc09ce534, 32'h41350910} /* (25, 25, 23) {real, imag} */,
  {32'hc1b2401c, 32'h41568c1b} /* (25, 25, 22) {real, imag} */,
  {32'h40de08b8, 32'h41376f92} /* (25, 25, 21) {real, imag} */,
  {32'hc091ff30, 32'hc15ac813} /* (25, 25, 20) {real, imag} */,
  {32'h4184969e, 32'hc12c9750} /* (25, 25, 19) {real, imag} */,
  {32'hbf20a488, 32'h404e5f6d} /* (25, 25, 18) {real, imag} */,
  {32'hc0d4377c, 32'hc0d2e07a} /* (25, 25, 17) {real, imag} */,
  {32'hc02d7ade, 32'hbfe27d44} /* (25, 25, 16) {real, imag} */,
  {32'h4052ab41, 32'hc12081d8} /* (25, 25, 15) {real, imag} */,
  {32'h40b43fe1, 32'h40f45803} /* (25, 25, 14) {real, imag} */,
  {32'hc15da76d, 32'h41715148} /* (25, 25, 13) {real, imag} */,
  {32'hbe9a2168, 32'hc06cdbb9} /* (25, 25, 12) {real, imag} */,
  {32'hc0662472, 32'h4172fa71} /* (25, 25, 11) {real, imag} */,
  {32'hc14378fe, 32'hc0823dcc} /* (25, 25, 10) {real, imag} */,
  {32'h40d87688, 32'hc12d5b1f} /* (25, 25, 9) {real, imag} */,
  {32'h4030ec86, 32'h42049174} /* (25, 25, 8) {real, imag} */,
  {32'h40d82542, 32'h41327b17} /* (25, 25, 7) {real, imag} */,
  {32'hc1184002, 32'h412415e0} /* (25, 25, 6) {real, imag} */,
  {32'h3f69e68c, 32'hc0b4e45e} /* (25, 25, 5) {real, imag} */,
  {32'hc11fbb24, 32'hc0c8adcc} /* (25, 25, 4) {real, imag} */,
  {32'hc07e4b14, 32'h41b347a6} /* (25, 25, 3) {real, imag} */,
  {32'h40af3e3c, 32'h40faa3a0} /* (25, 25, 2) {real, imag} */,
  {32'hc18ad48b, 32'h41354daa} /* (25, 25, 1) {real, imag} */,
  {32'hc203d5fe, 32'h4029c4ca} /* (25, 25, 0) {real, imag} */,
  {32'h4233094d, 32'hc14f4c7a} /* (25, 24, 31) {real, imag} */,
  {32'hc1f39902, 32'h41083a64} /* (25, 24, 30) {real, imag} */,
  {32'hc1dff362, 32'hc11297d6} /* (25, 24, 29) {real, imag} */,
  {32'hc0f5d92a, 32'hc1ee730f} /* (25, 24, 28) {real, imag} */,
  {32'hbf9c7080, 32'hbff5b8fc} /* (25, 24, 27) {real, imag} */,
  {32'hc1754518, 32'h40c2cf94} /* (25, 24, 26) {real, imag} */,
  {32'hc02d0482, 32'h414e6344} /* (25, 24, 25) {real, imag} */,
  {32'hc0ae9970, 32'h41989e30} /* (25, 24, 24) {real, imag} */,
  {32'h409e7b40, 32'hc01a89b4} /* (25, 24, 23) {real, imag} */,
  {32'h411aab6a, 32'hc0698a8a} /* (25, 24, 22) {real, imag} */,
  {32'h413d8652, 32'h4129b408} /* (25, 24, 21) {real, imag} */,
  {32'hc14d2d90, 32'hc1343660} /* (25, 24, 20) {real, imag} */,
  {32'h3fc591d8, 32'h419cc25b} /* (25, 24, 19) {real, imag} */,
  {32'h405383a8, 32'h418d106b} /* (25, 24, 18) {real, imag} */,
  {32'h40fd077a, 32'hc177d72c} /* (25, 24, 17) {real, imag} */,
  {32'h4129fbac, 32'h410bc557} /* (25, 24, 16) {real, imag} */,
  {32'hc0995df7, 32'h401e6d7a} /* (25, 24, 15) {real, imag} */,
  {32'hc156d18a, 32'hc0a4b51e} /* (25, 24, 14) {real, imag} */,
  {32'hc0f4286e, 32'hc1000618} /* (25, 24, 13) {real, imag} */,
  {32'h3edfb9a8, 32'hc10a896a} /* (25, 24, 12) {real, imag} */,
  {32'hc04136c6, 32'h4114641c} /* (25, 24, 11) {real, imag} */,
  {32'h40b8494c, 32'h40717172} /* (25, 24, 10) {real, imag} */,
  {32'h419a0ad0, 32'h418a2d84} /* (25, 24, 9) {real, imag} */,
  {32'h40e836ea, 32'h3f901770} /* (25, 24, 8) {real, imag} */,
  {32'h41a9f621, 32'h40667b06} /* (25, 24, 7) {real, imag} */,
  {32'hbe54f1a0, 32'h3fcc1ee8} /* (25, 24, 6) {real, imag} */,
  {32'hc1733594, 32'hbfa57604} /* (25, 24, 5) {real, imag} */,
  {32'hc04f6da0, 32'h3fc94e4c} /* (25, 24, 4) {real, imag} */,
  {32'h4192d514, 32'hc04f0906} /* (25, 24, 3) {real, imag} */,
  {32'hc1970cdf, 32'hc118abe0} /* (25, 24, 2) {real, imag} */,
  {32'h4249ab45, 32'hc15213d0} /* (25, 24, 1) {real, imag} */,
  {32'h417df5fa, 32'hc07e68ee} /* (25, 24, 0) {real, imag} */,
  {32'hc0d33190, 32'h4183e02d} /* (25, 23, 31) {real, imag} */,
  {32'h4053a19e, 32'h4111e0a8} /* (25, 23, 30) {real, imag} */,
  {32'h3fdddd02, 32'h41bc249c} /* (25, 23, 29) {real, imag} */,
  {32'hc112c907, 32'h4150214c} /* (25, 23, 28) {real, imag} */,
  {32'hc029d784, 32'hc1913a2c} /* (25, 23, 27) {real, imag} */,
  {32'h41aac6b4, 32'hc037de98} /* (25, 23, 26) {real, imag} */,
  {32'hc0742fda, 32'h412caaec} /* (25, 23, 25) {real, imag} */,
  {32'h4142affe, 32'h40f2ef23} /* (25, 23, 24) {real, imag} */,
  {32'hc0c0a2df, 32'hbfcfef68} /* (25, 23, 23) {real, imag} */,
  {32'hc1063128, 32'h402739f4} /* (25, 23, 22) {real, imag} */,
  {32'hc081ad3c, 32'hc16e45a4} /* (25, 23, 21) {real, imag} */,
  {32'hc0f9a1a6, 32'hc03b3bba} /* (25, 23, 20) {real, imag} */,
  {32'hc15747d5, 32'hc0cb3a78} /* (25, 23, 19) {real, imag} */,
  {32'h4112ffa8, 32'h3f7facc4} /* (25, 23, 18) {real, imag} */,
  {32'hc0ad79e2, 32'h40ea9c48} /* (25, 23, 17) {real, imag} */,
  {32'h3fb790d9, 32'hbf1ef7a8} /* (25, 23, 16) {real, imag} */,
  {32'hc0e928b7, 32'hc17f7810} /* (25, 23, 15) {real, imag} */,
  {32'hc0abb44e, 32'hbf455a28} /* (25, 23, 14) {real, imag} */,
  {32'h40d10ebc, 32'hc104d225} /* (25, 23, 13) {real, imag} */,
  {32'h4157b1c0, 32'hc1076b61} /* (25, 23, 12) {real, imag} */,
  {32'h4157b435, 32'hbfc9b99e} /* (25, 23, 11) {real, imag} */,
  {32'hc0e33bbe, 32'h3fc171ec} /* (25, 23, 10) {real, imag} */,
  {32'h413dbab7, 32'hc15bd3b3} /* (25, 23, 9) {real, imag} */,
  {32'h4122a3cc, 32'h3f292728} /* (25, 23, 8) {real, imag} */,
  {32'h3fc4f110, 32'h41012b9a} /* (25, 23, 7) {real, imag} */,
  {32'hc1b18670, 32'h40f9ba44} /* (25, 23, 6) {real, imag} */,
  {32'h41a550b6, 32'hc1317aed} /* (25, 23, 5) {real, imag} */,
  {32'hc104af65, 32'h40ada943} /* (25, 23, 4) {real, imag} */,
  {32'h416bdb40, 32'hc0a20095} /* (25, 23, 3) {real, imag} */,
  {32'hc0a81d80, 32'hc09aaea2} /* (25, 23, 2) {real, imag} */,
  {32'h4169b67c, 32'h41126a5e} /* (25, 23, 1) {real, imag} */,
  {32'hc1a0a077, 32'h4080c449} /* (25, 23, 0) {real, imag} */,
  {32'h4068e4d0, 32'h41b1cc26} /* (25, 22, 31) {real, imag} */,
  {32'hc1831662, 32'h405efbe2} /* (25, 22, 30) {real, imag} */,
  {32'h4143f4f0, 32'hc14022e4} /* (25, 22, 29) {real, imag} */,
  {32'h403c37fb, 32'h418996aa} /* (25, 22, 28) {real, imag} */,
  {32'hc1034ea6, 32'hc19342b2} /* (25, 22, 27) {real, imag} */,
  {32'h40e7ffde, 32'h405b69ea} /* (25, 22, 26) {real, imag} */,
  {32'h410bb1b5, 32'h3ffc65c4} /* (25, 22, 25) {real, imag} */,
  {32'h412c89a0, 32'h40c682a1} /* (25, 22, 24) {real, imag} */,
  {32'h4132273e, 32'hc0afc0b5} /* (25, 22, 23) {real, imag} */,
  {32'hc03a60c6, 32'hc09c273f} /* (25, 22, 22) {real, imag} */,
  {32'h3e8399f8, 32'h41221763} /* (25, 22, 21) {real, imag} */,
  {32'hc150a59a, 32'h418bc40f} /* (25, 22, 20) {real, imag} */,
  {32'h3ffc87ec, 32'h41acf721} /* (25, 22, 19) {real, imag} */,
  {32'hc11451c1, 32'hc12d13b5} /* (25, 22, 18) {real, imag} */,
  {32'hbeb85f72, 32'h409e581e} /* (25, 22, 17) {real, imag} */,
  {32'hc09873c9, 32'hc11087e1} /* (25, 22, 16) {real, imag} */,
  {32'h40a9db15, 32'hc110168c} /* (25, 22, 15) {real, imag} */,
  {32'h4156773b, 32'hc171ac66} /* (25, 22, 14) {real, imag} */,
  {32'h4065bfd2, 32'hc04f5b94} /* (25, 22, 13) {real, imag} */,
  {32'h3fb418e0, 32'h3eb33c70} /* (25, 22, 12) {real, imag} */,
  {32'hbfacd130, 32'h3fe014a0} /* (25, 22, 11) {real, imag} */,
  {32'h4164a091, 32'hc16f449a} /* (25, 22, 10) {real, imag} */,
  {32'h418d794f, 32'h4165bb35} /* (25, 22, 9) {real, imag} */,
  {32'hc1bd6904, 32'h4008373d} /* (25, 22, 8) {real, imag} */,
  {32'h413d357a, 32'hc05f23e2} /* (25, 22, 7) {real, imag} */,
  {32'hc12ca2f7, 32'h411d6012} /* (25, 22, 6) {real, imag} */,
  {32'h4112f74a, 32'h412b7c2d} /* (25, 22, 5) {real, imag} */,
  {32'hc0accca0, 32'h40b00e5c} /* (25, 22, 4) {real, imag} */,
  {32'hc0e21b00, 32'h41031b2d} /* (25, 22, 3) {real, imag} */,
  {32'h413ece1c, 32'hc1b3439e} /* (25, 22, 2) {real, imag} */,
  {32'hbfbefed0, 32'h414b8bde} /* (25, 22, 1) {real, imag} */,
  {32'h41122290, 32'h40a91a48} /* (25, 22, 0) {real, imag} */,
  {32'h414c079a, 32'hc105b702} /* (25, 21, 31) {real, imag} */,
  {32'hc069898a, 32'h4192a943} /* (25, 21, 30) {real, imag} */,
  {32'h40df8e7d, 32'h4117befa} /* (25, 21, 29) {real, imag} */,
  {32'h40cd3f70, 32'hc1aa1eb6} /* (25, 21, 28) {real, imag} */,
  {32'h40b966d0, 32'hc0108cf2} /* (25, 21, 27) {real, imag} */,
  {32'hc00b932a, 32'h4128040f} /* (25, 21, 26) {real, imag} */,
  {32'hc0fc8673, 32'h3ec45fa0} /* (25, 21, 25) {real, imag} */,
  {32'h40e483ee, 32'hc0aa05ba} /* (25, 21, 24) {real, imag} */,
  {32'hc10e420a, 32'h40b5bd45} /* (25, 21, 23) {real, imag} */,
  {32'hc10d809c, 32'hbfb01eb8} /* (25, 21, 22) {real, imag} */,
  {32'h41aafa01, 32'hc0cc6831} /* (25, 21, 21) {real, imag} */,
  {32'h41320440, 32'h3f97d278} /* (25, 21, 20) {real, imag} */,
  {32'hc0e0986c, 32'h40b6cf51} /* (25, 21, 19) {real, imag} */,
  {32'h404f0028, 32'h40f4c5d4} /* (25, 21, 18) {real, imag} */,
  {32'hc0d182a8, 32'h3f9758b4} /* (25, 21, 17) {real, imag} */,
  {32'h3f8b2e0c, 32'h407a8964} /* (25, 21, 16) {real, imag} */,
  {32'hbfeb65e4, 32'h4062fe4a} /* (25, 21, 15) {real, imag} */,
  {32'h40a37ab6, 32'hc1788787} /* (25, 21, 14) {real, imag} */,
  {32'h40f6fae2, 32'h40edea47} /* (25, 21, 13) {real, imag} */,
  {32'h3f3c1a70, 32'h3feb1292} /* (25, 21, 12) {real, imag} */,
  {32'hc1725a01, 32'hbeb2cb30} /* (25, 21, 11) {real, imag} */,
  {32'hc12073df, 32'hc19aa84a} /* (25, 21, 10) {real, imag} */,
  {32'hc0b51fde, 32'h3fba5b38} /* (25, 21, 9) {real, imag} */,
  {32'h417d159b, 32'hc16bdcee} /* (25, 21, 8) {real, imag} */,
  {32'h4119293c, 32'hbd9ff450} /* (25, 21, 7) {real, imag} */,
  {32'hc06742dd, 32'hc09c8d6b} /* (25, 21, 6) {real, imag} */,
  {32'hc16f310f, 32'h40c0eec4} /* (25, 21, 5) {real, imag} */,
  {32'h3f922b7c, 32'h3f3a48a0} /* (25, 21, 4) {real, imag} */,
  {32'h4145181c, 32'h40b7cff4} /* (25, 21, 3) {real, imag} */,
  {32'hc0f1983e, 32'h41c1dd03} /* (25, 21, 2) {real, imag} */,
  {32'h419d9d56, 32'hc0cf2a3a} /* (25, 21, 1) {real, imag} */,
  {32'hbfaaafa8, 32'hc199c7ce} /* (25, 21, 0) {real, imag} */,
  {32'h412b1cef, 32'hbfda24b2} /* (25, 20, 31) {real, imag} */,
  {32'h418c0c6e, 32'hc0222958} /* (25, 20, 30) {real, imag} */,
  {32'hc0ad9835, 32'h40acce55} /* (25, 20, 29) {real, imag} */,
  {32'hc08998f7, 32'hc12d6d65} /* (25, 20, 28) {real, imag} */,
  {32'hc188a032, 32'hc02e0780} /* (25, 20, 27) {real, imag} */,
  {32'hc0d0c6fa, 32'hbfe5dc40} /* (25, 20, 26) {real, imag} */,
  {32'h40246c70, 32'h3ffd2e80} /* (25, 20, 25) {real, imag} */,
  {32'hc167e9c6, 32'hc127a1c8} /* (25, 20, 24) {real, imag} */,
  {32'hc11d7e38, 32'h419e1bb4} /* (25, 20, 23) {real, imag} */,
  {32'h3e31d5a0, 32'h40ca8346} /* (25, 20, 22) {real, imag} */,
  {32'hc0efda4e, 32'hc0ee98b6} /* (25, 20, 21) {real, imag} */,
  {32'h417449a3, 32'hc0570608} /* (25, 20, 20) {real, imag} */,
  {32'hc1278d47, 32'h413105ef} /* (25, 20, 19) {real, imag} */,
  {32'h412ffccd, 32'h3fc191f4} /* (25, 20, 18) {real, imag} */,
  {32'h41575087, 32'hc1a1c4cc} /* (25, 20, 17) {real, imag} */,
  {32'hc06da0d9, 32'hc14c3502} /* (25, 20, 16) {real, imag} */,
  {32'h4114f071, 32'hc12bf2d4} /* (25, 20, 15) {real, imag} */,
  {32'h3f1f7fb8, 32'h40f06742} /* (25, 20, 14) {real, imag} */,
  {32'h4189b32d, 32'h3fbcb7fc} /* (25, 20, 13) {real, imag} */,
  {32'hc10067a2, 32'h405f0a12} /* (25, 20, 12) {real, imag} */,
  {32'hc143b987, 32'hc0d0aeb2} /* (25, 20, 11) {real, imag} */,
  {32'h412b4d47, 32'hc0a9c37c} /* (25, 20, 10) {real, imag} */,
  {32'h419ea32f, 32'hc0eeff41} /* (25, 20, 9) {real, imag} */,
  {32'h418af56f, 32'h4005e7b9} /* (25, 20, 8) {real, imag} */,
  {32'h41060159, 32'hc09f15c4} /* (25, 20, 7) {real, imag} */,
  {32'h40bac52a, 32'hc14254f3} /* (25, 20, 6) {real, imag} */,
  {32'h419b422c, 32'h40a0b1bf} /* (25, 20, 5) {real, imag} */,
  {32'h3ea73450, 32'h41517c7a} /* (25, 20, 4) {real, imag} */,
  {32'hc187dcf2, 32'h41364248} /* (25, 20, 3) {real, imag} */,
  {32'hc0ab25fe, 32'hc0a8e3ac} /* (25, 20, 2) {real, imag} */,
  {32'hc0b9d765, 32'h4027b078} /* (25, 20, 1) {real, imag} */,
  {32'h41090201, 32'h40c060c6} /* (25, 20, 0) {real, imag} */,
  {32'hc1950b53, 32'hc117c71a} /* (25, 19, 31) {real, imag} */,
  {32'hc0e6c07d, 32'hc1022e14} /* (25, 19, 30) {real, imag} */,
  {32'h40df3386, 32'hc120a616} /* (25, 19, 29) {real, imag} */,
  {32'hc0c6f82a, 32'hc03db487} /* (25, 19, 28) {real, imag} */,
  {32'hc0c4ddbb, 32'hc14521b4} /* (25, 19, 27) {real, imag} */,
  {32'h3f9342eb, 32'hc0d92c34} /* (25, 19, 26) {real, imag} */,
  {32'h40f28d39, 32'hc117c3c9} /* (25, 19, 25) {real, imag} */,
  {32'h4114ef65, 32'h3fb87d64} /* (25, 19, 24) {real, imag} */,
  {32'hc0f044ca, 32'hc0ce8fd1} /* (25, 19, 23) {real, imag} */,
  {32'h3f36d9e0, 32'hc0e70eec} /* (25, 19, 22) {real, imag} */,
  {32'hc115ba59, 32'h40a81f8c} /* (25, 19, 21) {real, imag} */,
  {32'h40c69097, 32'hc15cefdc} /* (25, 19, 20) {real, imag} */,
  {32'hc06135a6, 32'h4060d2df} /* (25, 19, 19) {real, imag} */,
  {32'h41a3cc90, 32'h402040ac} /* (25, 19, 18) {real, imag} */,
  {32'hbff62f48, 32'hc05feff9} /* (25, 19, 17) {real, imag} */,
  {32'hc1862a87, 32'h40c5ccb6} /* (25, 19, 16) {real, imag} */,
  {32'h412e70ed, 32'h40007f52} /* (25, 19, 15) {real, imag} */,
  {32'h40e20a0a, 32'h4148ad99} /* (25, 19, 14) {real, imag} */,
  {32'h3ede60c0, 32'hc0220898} /* (25, 19, 13) {real, imag} */,
  {32'hc045d75c, 32'h4147b3c2} /* (25, 19, 12) {real, imag} */,
  {32'hc1615d7d, 32'hc1972ed8} /* (25, 19, 11) {real, imag} */,
  {32'h40b87ae3, 32'hc193ad19} /* (25, 19, 10) {real, imag} */,
  {32'hc1368fe2, 32'h40c45710} /* (25, 19, 9) {real, imag} */,
  {32'hbdd22040, 32'hbf9771c0} /* (25, 19, 8) {real, imag} */,
  {32'hc1600281, 32'h3fe37da9} /* (25, 19, 7) {real, imag} */,
  {32'h4112cef3, 32'hc13e07ea} /* (25, 19, 6) {real, imag} */,
  {32'h406c640a, 32'h40c67d6e} /* (25, 19, 5) {real, imag} */,
  {32'hbe540c20, 32'hc088cfa4} /* (25, 19, 4) {real, imag} */,
  {32'h4063864f, 32'h416eccf5} /* (25, 19, 3) {real, imag} */,
  {32'h3fdc20b4, 32'h41410978} /* (25, 19, 2) {real, imag} */,
  {32'hc12eb6ef, 32'h3ff98054} /* (25, 19, 1) {real, imag} */,
  {32'hc0b62b90, 32'h4127397e} /* (25, 19, 0) {real, imag} */,
  {32'hc0518b5f, 32'hc1932681} /* (25, 18, 31) {real, imag} */,
  {32'h4160ff0a, 32'h4105905a} /* (25, 18, 30) {real, imag} */,
  {32'hc03f135b, 32'hc0ad08d8} /* (25, 18, 29) {real, imag} */,
  {32'hc031aace, 32'hc12e7b2e} /* (25, 18, 28) {real, imag} */,
  {32'h4185f016, 32'hc06469fe} /* (25, 18, 27) {real, imag} */,
  {32'h41679860, 32'hc0dab92f} /* (25, 18, 26) {real, imag} */,
  {32'hc122a343, 32'h3edd65c2} /* (25, 18, 25) {real, imag} */,
  {32'h417aadd8, 32'hbff3837c} /* (25, 18, 24) {real, imag} */,
  {32'h413d7af6, 32'hc0ce879d} /* (25, 18, 23) {real, imag} */,
  {32'h40e200aa, 32'hc13bd6ed} /* (25, 18, 22) {real, imag} */,
  {32'h408cc244, 32'hc0748534} /* (25, 18, 21) {real, imag} */,
  {32'h4046891a, 32'h412afca9} /* (25, 18, 20) {real, imag} */,
  {32'h40c187b2, 32'h413a611e} /* (25, 18, 19) {real, imag} */,
  {32'h4040642c, 32'h3fb51e48} /* (25, 18, 18) {real, imag} */,
  {32'h3ec677e0, 32'hbe9b29fc} /* (25, 18, 17) {real, imag} */,
  {32'h401c77f0, 32'hbec5eee0} /* (25, 18, 16) {real, imag} */,
  {32'h40450272, 32'h40a390cf} /* (25, 18, 15) {real, imag} */,
  {32'h40991a0a, 32'hc0efd804} /* (25, 18, 14) {real, imag} */,
  {32'hc1612b79, 32'h40a6d64b} /* (25, 18, 13) {real, imag} */,
  {32'hc182d1d0, 32'hc0c29d54} /* (25, 18, 12) {real, imag} */,
  {32'h40dc8888, 32'hc05d2e98} /* (25, 18, 11) {real, imag} */,
  {32'h417673a9, 32'h4070cfa2} /* (25, 18, 10) {real, imag} */,
  {32'hc17e280a, 32'h41aa4a28} /* (25, 18, 9) {real, imag} */,
  {32'hc11d24a9, 32'hc1468f3e} /* (25, 18, 8) {real, imag} */,
  {32'hc1fbcbc4, 32'hc120a711} /* (25, 18, 7) {real, imag} */,
  {32'hbff5f708, 32'h40d4fdcb} /* (25, 18, 6) {real, imag} */,
  {32'h40deb84c, 32'hc12122a4} /* (25, 18, 5) {real, imag} */,
  {32'h4182ba72, 32'h41267177} /* (25, 18, 4) {real, imag} */,
  {32'hc0d8397a, 32'hc0df44ce} /* (25, 18, 3) {real, imag} */,
  {32'hbe984c38, 32'hc05bd707} /* (25, 18, 2) {real, imag} */,
  {32'h4066c5ee, 32'hc1adf588} /* (25, 18, 1) {real, imag} */,
  {32'hc0c35684, 32'hc1b02eb2} /* (25, 18, 0) {real, imag} */,
  {32'hc0c6f8d6, 32'h3fdd3a00} /* (25, 17, 31) {real, imag} */,
  {32'hbff15749, 32'hc1a20e93} /* (25, 17, 30) {real, imag} */,
  {32'hbf33ccf4, 32'h40ab5640} /* (25, 17, 29) {real, imag} */,
  {32'hc0a72e3e, 32'hc00c06ba} /* (25, 17, 28) {real, imag} */,
  {32'hc08f430e, 32'h414f686c} /* (25, 17, 27) {real, imag} */,
  {32'hc00613d7, 32'hc0ae916a} /* (25, 17, 26) {real, imag} */,
  {32'h40b3e910, 32'h40e0b1c0} /* (25, 17, 25) {real, imag} */,
  {32'h41459995, 32'hc0b41c65} /* (25, 17, 24) {real, imag} */,
  {32'h3f457f8c, 32'h40dc8569} /* (25, 17, 23) {real, imag} */,
  {32'h41001151, 32'h403f5674} /* (25, 17, 22) {real, imag} */,
  {32'hc139e1aa, 32'h410c63d8} /* (25, 17, 21) {real, imag} */,
  {32'h405552f0, 32'h40fea7fc} /* (25, 17, 20) {real, imag} */,
  {32'hbfed5b72, 32'hc10fb30b} /* (25, 17, 19) {real, imag} */,
  {32'h416e9a46, 32'h41414abc} /* (25, 17, 18) {real, imag} */,
  {32'h40aa1482, 32'h3f8abe26} /* (25, 17, 17) {real, imag} */,
  {32'h3fb264dc, 32'h409d6b44} /* (25, 17, 16) {real, imag} */,
  {32'hc116ac7a, 32'hc114fbde} /* (25, 17, 15) {real, imag} */,
  {32'hc115c3e4, 32'hc0db70d0} /* (25, 17, 14) {real, imag} */,
  {32'h408d0f65, 32'hc071b0c5} /* (25, 17, 13) {real, imag} */,
  {32'h40d75a82, 32'h40a0c56e} /* (25, 17, 12) {real, imag} */,
  {32'h40bfd4cc, 32'hc0d38299} /* (25, 17, 11) {real, imag} */,
  {32'h408e87f4, 32'h41a37046} /* (25, 17, 10) {real, imag} */,
  {32'h40eb9aa3, 32'hc050f03b} /* (25, 17, 9) {real, imag} */,
  {32'h3f832d3a, 32'hbf827390} /* (25, 17, 8) {real, imag} */,
  {32'hc0c0d2e0, 32'h41b47ef0} /* (25, 17, 7) {real, imag} */,
  {32'h4093d434, 32'hc0875b0d} /* (25, 17, 6) {real, imag} */,
  {32'hc0e740f8, 32'h3f97c9d0} /* (25, 17, 5) {real, imag} */,
  {32'h3f3e7a24, 32'h3f5a9a2e} /* (25, 17, 4) {real, imag} */,
  {32'hbd6a9f40, 32'hc0593240} /* (25, 17, 3) {real, imag} */,
  {32'hbf88695c, 32'hc0b499cd} /* (25, 17, 2) {real, imag} */,
  {32'hc1181c16, 32'h4160ad96} /* (25, 17, 1) {real, imag} */,
  {32'h4184a911, 32'hbff7fe70} /* (25, 17, 0) {real, imag} */,
  {32'h40af8c82, 32'h40b7c0fa} /* (25, 16, 31) {real, imag} */,
  {32'h4082b66c, 32'hbf75b7d4} /* (25, 16, 30) {real, imag} */,
  {32'hc0c54254, 32'hbf749246} /* (25, 16, 29) {real, imag} */,
  {32'h40aad96e, 32'h41287ee1} /* (25, 16, 28) {real, imag} */,
  {32'h403fbe34, 32'h403c30e2} /* (25, 16, 27) {real, imag} */,
  {32'h41235f08, 32'h4103eb6c} /* (25, 16, 26) {real, imag} */,
  {32'hc0ae39b8, 32'hc0cb99ce} /* (25, 16, 25) {real, imag} */,
  {32'hc0c6da56, 32'h3fefcd16} /* (25, 16, 24) {real, imag} */,
  {32'hc15f2bba, 32'hbf6dff00} /* (25, 16, 23) {real, imag} */,
  {32'hc02b4bee, 32'hc09ad0b5} /* (25, 16, 22) {real, imag} */,
  {32'hbfa6ddd2, 32'h40e29ec8} /* (25, 16, 21) {real, imag} */,
  {32'h3f003798, 32'h41670a12} /* (25, 16, 20) {real, imag} */,
  {32'hc115297a, 32'h3e79b650} /* (25, 16, 19) {real, imag} */,
  {32'hc081a8fe, 32'h3f03c3e7} /* (25, 16, 18) {real, imag} */,
  {32'hc0467dd8, 32'hc0ccec62} /* (25, 16, 17) {real, imag} */,
  {32'h3f3443c8, 32'h00000000} /* (25, 16, 16) {real, imag} */,
  {32'hc0467dd8, 32'h40ccec62} /* (25, 16, 15) {real, imag} */,
  {32'hc081a8fe, 32'hbf03c3e7} /* (25, 16, 14) {real, imag} */,
  {32'hc115297a, 32'hbe79b650} /* (25, 16, 13) {real, imag} */,
  {32'h3f003798, 32'hc1670a12} /* (25, 16, 12) {real, imag} */,
  {32'hbfa6ddd2, 32'hc0e29ec8} /* (25, 16, 11) {real, imag} */,
  {32'hc02b4bee, 32'h409ad0b5} /* (25, 16, 10) {real, imag} */,
  {32'hc15f2bba, 32'h3f6dff00} /* (25, 16, 9) {real, imag} */,
  {32'hc0c6da56, 32'hbfefcd16} /* (25, 16, 8) {real, imag} */,
  {32'hc0ae39b8, 32'h40cb99ce} /* (25, 16, 7) {real, imag} */,
  {32'h41235f08, 32'hc103eb6c} /* (25, 16, 6) {real, imag} */,
  {32'h403fbe34, 32'hc03c30e2} /* (25, 16, 5) {real, imag} */,
  {32'h40aad96e, 32'hc1287ee1} /* (25, 16, 4) {real, imag} */,
  {32'hc0c54254, 32'h3f749246} /* (25, 16, 3) {real, imag} */,
  {32'h4082b66c, 32'h3f75b7d4} /* (25, 16, 2) {real, imag} */,
  {32'h40af8c82, 32'hc0b7c0fa} /* (25, 16, 1) {real, imag} */,
  {32'h41564851, 32'h00000000} /* (25, 16, 0) {real, imag} */,
  {32'hc1181c16, 32'hc160ad96} /* (25, 15, 31) {real, imag} */,
  {32'hbf88695c, 32'h40b499cd} /* (25, 15, 30) {real, imag} */,
  {32'hbd6a9f40, 32'h40593240} /* (25, 15, 29) {real, imag} */,
  {32'h3f3e7a24, 32'hbf5a9a2e} /* (25, 15, 28) {real, imag} */,
  {32'hc0e740f8, 32'hbf97c9d0} /* (25, 15, 27) {real, imag} */,
  {32'h4093d434, 32'h40875b0d} /* (25, 15, 26) {real, imag} */,
  {32'hc0c0d2e0, 32'hc1b47ef0} /* (25, 15, 25) {real, imag} */,
  {32'h3f832d3a, 32'h3f827390} /* (25, 15, 24) {real, imag} */,
  {32'h40eb9aa3, 32'h4050f03b} /* (25, 15, 23) {real, imag} */,
  {32'h408e87f4, 32'hc1a37046} /* (25, 15, 22) {real, imag} */,
  {32'h40bfd4cc, 32'h40d38299} /* (25, 15, 21) {real, imag} */,
  {32'h40d75a82, 32'hc0a0c56e} /* (25, 15, 20) {real, imag} */,
  {32'h408d0f65, 32'h4071b0c5} /* (25, 15, 19) {real, imag} */,
  {32'hc115c3e4, 32'h40db70d0} /* (25, 15, 18) {real, imag} */,
  {32'hc116ac7a, 32'h4114fbde} /* (25, 15, 17) {real, imag} */,
  {32'h3fb264dc, 32'hc09d6b44} /* (25, 15, 16) {real, imag} */,
  {32'h40aa1482, 32'hbf8abe26} /* (25, 15, 15) {real, imag} */,
  {32'h416e9a46, 32'hc1414abc} /* (25, 15, 14) {real, imag} */,
  {32'hbfed5b72, 32'h410fb30b} /* (25, 15, 13) {real, imag} */,
  {32'h405552f0, 32'hc0fea7fc} /* (25, 15, 12) {real, imag} */,
  {32'hc139e1aa, 32'hc10c63d8} /* (25, 15, 11) {real, imag} */,
  {32'h41001151, 32'hc03f5674} /* (25, 15, 10) {real, imag} */,
  {32'h3f457f8c, 32'hc0dc8569} /* (25, 15, 9) {real, imag} */,
  {32'h41459995, 32'h40b41c65} /* (25, 15, 8) {real, imag} */,
  {32'h40b3e910, 32'hc0e0b1c0} /* (25, 15, 7) {real, imag} */,
  {32'hc00613d7, 32'h40ae916a} /* (25, 15, 6) {real, imag} */,
  {32'hc08f430e, 32'hc14f686c} /* (25, 15, 5) {real, imag} */,
  {32'hc0a72e3e, 32'h400c06ba} /* (25, 15, 4) {real, imag} */,
  {32'hbf33ccf4, 32'hc0ab5640} /* (25, 15, 3) {real, imag} */,
  {32'hbff15749, 32'h41a20e93} /* (25, 15, 2) {real, imag} */,
  {32'hc0c6f8d6, 32'hbfdd3a00} /* (25, 15, 1) {real, imag} */,
  {32'h4184a911, 32'h3ff7fe70} /* (25, 15, 0) {real, imag} */,
  {32'h4066c5ee, 32'h41adf588} /* (25, 14, 31) {real, imag} */,
  {32'hbe984c38, 32'h405bd707} /* (25, 14, 30) {real, imag} */,
  {32'hc0d8397a, 32'h40df44ce} /* (25, 14, 29) {real, imag} */,
  {32'h4182ba72, 32'hc1267177} /* (25, 14, 28) {real, imag} */,
  {32'h40deb84c, 32'h412122a4} /* (25, 14, 27) {real, imag} */,
  {32'hbff5f708, 32'hc0d4fdcb} /* (25, 14, 26) {real, imag} */,
  {32'hc1fbcbc4, 32'h4120a711} /* (25, 14, 25) {real, imag} */,
  {32'hc11d24a9, 32'h41468f3e} /* (25, 14, 24) {real, imag} */,
  {32'hc17e280a, 32'hc1aa4a28} /* (25, 14, 23) {real, imag} */,
  {32'h417673a9, 32'hc070cfa2} /* (25, 14, 22) {real, imag} */,
  {32'h40dc8888, 32'h405d2e98} /* (25, 14, 21) {real, imag} */,
  {32'hc182d1d0, 32'h40c29d54} /* (25, 14, 20) {real, imag} */,
  {32'hc1612b79, 32'hc0a6d64b} /* (25, 14, 19) {real, imag} */,
  {32'h40991a0a, 32'h40efd804} /* (25, 14, 18) {real, imag} */,
  {32'h40450272, 32'hc0a390cf} /* (25, 14, 17) {real, imag} */,
  {32'h401c77f0, 32'h3ec5eee0} /* (25, 14, 16) {real, imag} */,
  {32'h3ec677e0, 32'h3e9b29fc} /* (25, 14, 15) {real, imag} */,
  {32'h4040642c, 32'hbfb51e48} /* (25, 14, 14) {real, imag} */,
  {32'h40c187b2, 32'hc13a611e} /* (25, 14, 13) {real, imag} */,
  {32'h4046891a, 32'hc12afca9} /* (25, 14, 12) {real, imag} */,
  {32'h408cc244, 32'h40748534} /* (25, 14, 11) {real, imag} */,
  {32'h40e200aa, 32'h413bd6ed} /* (25, 14, 10) {real, imag} */,
  {32'h413d7af6, 32'h40ce879d} /* (25, 14, 9) {real, imag} */,
  {32'h417aadd8, 32'h3ff3837c} /* (25, 14, 8) {real, imag} */,
  {32'hc122a343, 32'hbedd65c2} /* (25, 14, 7) {real, imag} */,
  {32'h41679860, 32'h40dab92f} /* (25, 14, 6) {real, imag} */,
  {32'h4185f016, 32'h406469fe} /* (25, 14, 5) {real, imag} */,
  {32'hc031aace, 32'h412e7b2e} /* (25, 14, 4) {real, imag} */,
  {32'hc03f135b, 32'h40ad08d8} /* (25, 14, 3) {real, imag} */,
  {32'h4160ff0a, 32'hc105905a} /* (25, 14, 2) {real, imag} */,
  {32'hc0518b5f, 32'h41932681} /* (25, 14, 1) {real, imag} */,
  {32'hc0c35684, 32'h41b02eb2} /* (25, 14, 0) {real, imag} */,
  {32'hc12eb6ef, 32'hbff98054} /* (25, 13, 31) {real, imag} */,
  {32'h3fdc20b4, 32'hc1410978} /* (25, 13, 30) {real, imag} */,
  {32'h4063864f, 32'hc16eccf5} /* (25, 13, 29) {real, imag} */,
  {32'hbe540c20, 32'h4088cfa4} /* (25, 13, 28) {real, imag} */,
  {32'h406c640a, 32'hc0c67d6e} /* (25, 13, 27) {real, imag} */,
  {32'h4112cef3, 32'h413e07ea} /* (25, 13, 26) {real, imag} */,
  {32'hc1600281, 32'hbfe37da9} /* (25, 13, 25) {real, imag} */,
  {32'hbdd22040, 32'h3f9771c0} /* (25, 13, 24) {real, imag} */,
  {32'hc1368fe2, 32'hc0c45710} /* (25, 13, 23) {real, imag} */,
  {32'h40b87ae3, 32'h4193ad19} /* (25, 13, 22) {real, imag} */,
  {32'hc1615d7d, 32'h41972ed8} /* (25, 13, 21) {real, imag} */,
  {32'hc045d75c, 32'hc147b3c2} /* (25, 13, 20) {real, imag} */,
  {32'h3ede60c0, 32'h40220898} /* (25, 13, 19) {real, imag} */,
  {32'h40e20a0a, 32'hc148ad99} /* (25, 13, 18) {real, imag} */,
  {32'h412e70ed, 32'hc0007f52} /* (25, 13, 17) {real, imag} */,
  {32'hc1862a87, 32'hc0c5ccb6} /* (25, 13, 16) {real, imag} */,
  {32'hbff62f48, 32'h405feff9} /* (25, 13, 15) {real, imag} */,
  {32'h41a3cc90, 32'hc02040ac} /* (25, 13, 14) {real, imag} */,
  {32'hc06135a6, 32'hc060d2df} /* (25, 13, 13) {real, imag} */,
  {32'h40c69097, 32'h415cefdc} /* (25, 13, 12) {real, imag} */,
  {32'hc115ba59, 32'hc0a81f8c} /* (25, 13, 11) {real, imag} */,
  {32'h3f36d9e0, 32'h40e70eec} /* (25, 13, 10) {real, imag} */,
  {32'hc0f044ca, 32'h40ce8fd1} /* (25, 13, 9) {real, imag} */,
  {32'h4114ef65, 32'hbfb87d64} /* (25, 13, 8) {real, imag} */,
  {32'h40f28d39, 32'h4117c3c9} /* (25, 13, 7) {real, imag} */,
  {32'h3f9342eb, 32'h40d92c34} /* (25, 13, 6) {real, imag} */,
  {32'hc0c4ddbb, 32'h414521b4} /* (25, 13, 5) {real, imag} */,
  {32'hc0c6f82a, 32'h403db487} /* (25, 13, 4) {real, imag} */,
  {32'h40df3386, 32'h4120a616} /* (25, 13, 3) {real, imag} */,
  {32'hc0e6c07d, 32'h41022e14} /* (25, 13, 2) {real, imag} */,
  {32'hc1950b53, 32'h4117c71a} /* (25, 13, 1) {real, imag} */,
  {32'hc0b62b90, 32'hc127397e} /* (25, 13, 0) {real, imag} */,
  {32'hc0b9d765, 32'hc027b078} /* (25, 12, 31) {real, imag} */,
  {32'hc0ab25fe, 32'h40a8e3ac} /* (25, 12, 30) {real, imag} */,
  {32'hc187dcf2, 32'hc1364248} /* (25, 12, 29) {real, imag} */,
  {32'h3ea73450, 32'hc1517c7a} /* (25, 12, 28) {real, imag} */,
  {32'h419b422c, 32'hc0a0b1bf} /* (25, 12, 27) {real, imag} */,
  {32'h40bac52a, 32'h414254f3} /* (25, 12, 26) {real, imag} */,
  {32'h41060159, 32'h409f15c4} /* (25, 12, 25) {real, imag} */,
  {32'h418af56f, 32'hc005e7b9} /* (25, 12, 24) {real, imag} */,
  {32'h419ea32f, 32'h40eeff41} /* (25, 12, 23) {real, imag} */,
  {32'h412b4d47, 32'h40a9c37c} /* (25, 12, 22) {real, imag} */,
  {32'hc143b987, 32'h40d0aeb2} /* (25, 12, 21) {real, imag} */,
  {32'hc10067a2, 32'hc05f0a12} /* (25, 12, 20) {real, imag} */,
  {32'h4189b32d, 32'hbfbcb7fc} /* (25, 12, 19) {real, imag} */,
  {32'h3f1f7fb8, 32'hc0f06742} /* (25, 12, 18) {real, imag} */,
  {32'h4114f071, 32'h412bf2d4} /* (25, 12, 17) {real, imag} */,
  {32'hc06da0d9, 32'h414c3502} /* (25, 12, 16) {real, imag} */,
  {32'h41575087, 32'h41a1c4cc} /* (25, 12, 15) {real, imag} */,
  {32'h412ffccd, 32'hbfc191f4} /* (25, 12, 14) {real, imag} */,
  {32'hc1278d47, 32'hc13105ef} /* (25, 12, 13) {real, imag} */,
  {32'h417449a3, 32'h40570608} /* (25, 12, 12) {real, imag} */,
  {32'hc0efda4e, 32'h40ee98b6} /* (25, 12, 11) {real, imag} */,
  {32'h3e31d5a0, 32'hc0ca8346} /* (25, 12, 10) {real, imag} */,
  {32'hc11d7e38, 32'hc19e1bb4} /* (25, 12, 9) {real, imag} */,
  {32'hc167e9c6, 32'h4127a1c8} /* (25, 12, 8) {real, imag} */,
  {32'h40246c70, 32'hbffd2e80} /* (25, 12, 7) {real, imag} */,
  {32'hc0d0c6fa, 32'h3fe5dc40} /* (25, 12, 6) {real, imag} */,
  {32'hc188a032, 32'h402e0780} /* (25, 12, 5) {real, imag} */,
  {32'hc08998f7, 32'h412d6d65} /* (25, 12, 4) {real, imag} */,
  {32'hc0ad9835, 32'hc0acce55} /* (25, 12, 3) {real, imag} */,
  {32'h418c0c6e, 32'h40222958} /* (25, 12, 2) {real, imag} */,
  {32'h412b1cef, 32'h3fda24b2} /* (25, 12, 1) {real, imag} */,
  {32'h41090201, 32'hc0c060c6} /* (25, 12, 0) {real, imag} */,
  {32'h419d9d56, 32'h40cf2a3a} /* (25, 11, 31) {real, imag} */,
  {32'hc0f1983e, 32'hc1c1dd03} /* (25, 11, 30) {real, imag} */,
  {32'h4145181c, 32'hc0b7cff4} /* (25, 11, 29) {real, imag} */,
  {32'h3f922b7c, 32'hbf3a48a0} /* (25, 11, 28) {real, imag} */,
  {32'hc16f310f, 32'hc0c0eec4} /* (25, 11, 27) {real, imag} */,
  {32'hc06742dd, 32'h409c8d6b} /* (25, 11, 26) {real, imag} */,
  {32'h4119293c, 32'h3d9ff450} /* (25, 11, 25) {real, imag} */,
  {32'h417d159b, 32'h416bdcee} /* (25, 11, 24) {real, imag} */,
  {32'hc0b51fde, 32'hbfba5b38} /* (25, 11, 23) {real, imag} */,
  {32'hc12073df, 32'h419aa84a} /* (25, 11, 22) {real, imag} */,
  {32'hc1725a01, 32'h3eb2cb30} /* (25, 11, 21) {real, imag} */,
  {32'h3f3c1a70, 32'hbfeb1292} /* (25, 11, 20) {real, imag} */,
  {32'h40f6fae2, 32'hc0edea47} /* (25, 11, 19) {real, imag} */,
  {32'h40a37ab6, 32'h41788787} /* (25, 11, 18) {real, imag} */,
  {32'hbfeb65e4, 32'hc062fe4a} /* (25, 11, 17) {real, imag} */,
  {32'h3f8b2e0c, 32'hc07a8964} /* (25, 11, 16) {real, imag} */,
  {32'hc0d182a8, 32'hbf9758b4} /* (25, 11, 15) {real, imag} */,
  {32'h404f0028, 32'hc0f4c5d4} /* (25, 11, 14) {real, imag} */,
  {32'hc0e0986c, 32'hc0b6cf51} /* (25, 11, 13) {real, imag} */,
  {32'h41320440, 32'hbf97d278} /* (25, 11, 12) {real, imag} */,
  {32'h41aafa01, 32'h40cc6831} /* (25, 11, 11) {real, imag} */,
  {32'hc10d809c, 32'h3fb01eb8} /* (25, 11, 10) {real, imag} */,
  {32'hc10e420a, 32'hc0b5bd45} /* (25, 11, 9) {real, imag} */,
  {32'h40e483ee, 32'h40aa05ba} /* (25, 11, 8) {real, imag} */,
  {32'hc0fc8673, 32'hbec45fa0} /* (25, 11, 7) {real, imag} */,
  {32'hc00b932a, 32'hc128040f} /* (25, 11, 6) {real, imag} */,
  {32'h40b966d0, 32'h40108cf2} /* (25, 11, 5) {real, imag} */,
  {32'h40cd3f70, 32'h41aa1eb6} /* (25, 11, 4) {real, imag} */,
  {32'h40df8e7d, 32'hc117befa} /* (25, 11, 3) {real, imag} */,
  {32'hc069898a, 32'hc192a943} /* (25, 11, 2) {real, imag} */,
  {32'h414c079a, 32'h4105b702} /* (25, 11, 1) {real, imag} */,
  {32'hbfaaafa8, 32'h4199c7ce} /* (25, 11, 0) {real, imag} */,
  {32'hbfbefed0, 32'hc14b8bde} /* (25, 10, 31) {real, imag} */,
  {32'h413ece1c, 32'h41b3439e} /* (25, 10, 30) {real, imag} */,
  {32'hc0e21b00, 32'hc1031b2d} /* (25, 10, 29) {real, imag} */,
  {32'hc0accca0, 32'hc0b00e5c} /* (25, 10, 28) {real, imag} */,
  {32'h4112f74a, 32'hc12b7c2d} /* (25, 10, 27) {real, imag} */,
  {32'hc12ca2f7, 32'hc11d6012} /* (25, 10, 26) {real, imag} */,
  {32'h413d357a, 32'h405f23e2} /* (25, 10, 25) {real, imag} */,
  {32'hc1bd6904, 32'hc008373d} /* (25, 10, 24) {real, imag} */,
  {32'h418d794f, 32'hc165bb35} /* (25, 10, 23) {real, imag} */,
  {32'h4164a091, 32'h416f449a} /* (25, 10, 22) {real, imag} */,
  {32'hbfacd130, 32'hbfe014a0} /* (25, 10, 21) {real, imag} */,
  {32'h3fb418e0, 32'hbeb33c70} /* (25, 10, 20) {real, imag} */,
  {32'h4065bfd2, 32'h404f5b94} /* (25, 10, 19) {real, imag} */,
  {32'h4156773b, 32'h4171ac66} /* (25, 10, 18) {real, imag} */,
  {32'h40a9db15, 32'h4110168c} /* (25, 10, 17) {real, imag} */,
  {32'hc09873c9, 32'h411087e1} /* (25, 10, 16) {real, imag} */,
  {32'hbeb85f72, 32'hc09e581e} /* (25, 10, 15) {real, imag} */,
  {32'hc11451c1, 32'h412d13b5} /* (25, 10, 14) {real, imag} */,
  {32'h3ffc87ec, 32'hc1acf721} /* (25, 10, 13) {real, imag} */,
  {32'hc150a59a, 32'hc18bc40f} /* (25, 10, 12) {real, imag} */,
  {32'h3e8399f8, 32'hc1221763} /* (25, 10, 11) {real, imag} */,
  {32'hc03a60c6, 32'h409c273f} /* (25, 10, 10) {real, imag} */,
  {32'h4132273e, 32'h40afc0b5} /* (25, 10, 9) {real, imag} */,
  {32'h412c89a0, 32'hc0c682a1} /* (25, 10, 8) {real, imag} */,
  {32'h410bb1b5, 32'hbffc65c4} /* (25, 10, 7) {real, imag} */,
  {32'h40e7ffde, 32'hc05b69ea} /* (25, 10, 6) {real, imag} */,
  {32'hc1034ea6, 32'h419342b2} /* (25, 10, 5) {real, imag} */,
  {32'h403c37fb, 32'hc18996aa} /* (25, 10, 4) {real, imag} */,
  {32'h4143f4f0, 32'h414022e4} /* (25, 10, 3) {real, imag} */,
  {32'hc1831662, 32'hc05efbe2} /* (25, 10, 2) {real, imag} */,
  {32'h4068e4d0, 32'hc1b1cc26} /* (25, 10, 1) {real, imag} */,
  {32'h41122290, 32'hc0a91a48} /* (25, 10, 0) {real, imag} */,
  {32'h4169b67c, 32'hc1126a5e} /* (25, 9, 31) {real, imag} */,
  {32'hc0a81d80, 32'h409aaea2} /* (25, 9, 30) {real, imag} */,
  {32'h416bdb40, 32'h40a20095} /* (25, 9, 29) {real, imag} */,
  {32'hc104af65, 32'hc0ada943} /* (25, 9, 28) {real, imag} */,
  {32'h41a550b6, 32'h41317aed} /* (25, 9, 27) {real, imag} */,
  {32'hc1b18670, 32'hc0f9ba44} /* (25, 9, 26) {real, imag} */,
  {32'h3fc4f110, 32'hc1012b9a} /* (25, 9, 25) {real, imag} */,
  {32'h4122a3cc, 32'hbf292728} /* (25, 9, 24) {real, imag} */,
  {32'h413dbab7, 32'h415bd3b3} /* (25, 9, 23) {real, imag} */,
  {32'hc0e33bbe, 32'hbfc171ec} /* (25, 9, 22) {real, imag} */,
  {32'h4157b435, 32'h3fc9b99e} /* (25, 9, 21) {real, imag} */,
  {32'h4157b1c0, 32'h41076b61} /* (25, 9, 20) {real, imag} */,
  {32'h40d10ebc, 32'h4104d225} /* (25, 9, 19) {real, imag} */,
  {32'hc0abb44e, 32'h3f455a28} /* (25, 9, 18) {real, imag} */,
  {32'hc0e928b7, 32'h417f7810} /* (25, 9, 17) {real, imag} */,
  {32'h3fb790d9, 32'h3f1ef7a8} /* (25, 9, 16) {real, imag} */,
  {32'hc0ad79e2, 32'hc0ea9c48} /* (25, 9, 15) {real, imag} */,
  {32'h4112ffa8, 32'hbf7facc4} /* (25, 9, 14) {real, imag} */,
  {32'hc15747d5, 32'h40cb3a78} /* (25, 9, 13) {real, imag} */,
  {32'hc0f9a1a6, 32'h403b3bba} /* (25, 9, 12) {real, imag} */,
  {32'hc081ad3c, 32'h416e45a4} /* (25, 9, 11) {real, imag} */,
  {32'hc1063128, 32'hc02739f4} /* (25, 9, 10) {real, imag} */,
  {32'hc0c0a2df, 32'h3fcfef68} /* (25, 9, 9) {real, imag} */,
  {32'h4142affe, 32'hc0f2ef23} /* (25, 9, 8) {real, imag} */,
  {32'hc0742fda, 32'hc12caaec} /* (25, 9, 7) {real, imag} */,
  {32'h41aac6b4, 32'h4037de98} /* (25, 9, 6) {real, imag} */,
  {32'hc029d784, 32'h41913a2c} /* (25, 9, 5) {real, imag} */,
  {32'hc112c907, 32'hc150214c} /* (25, 9, 4) {real, imag} */,
  {32'h3fdddd02, 32'hc1bc249c} /* (25, 9, 3) {real, imag} */,
  {32'h4053a19e, 32'hc111e0a8} /* (25, 9, 2) {real, imag} */,
  {32'hc0d33190, 32'hc183e02d} /* (25, 9, 1) {real, imag} */,
  {32'hc1a0a077, 32'hc080c449} /* (25, 9, 0) {real, imag} */,
  {32'h4249ab45, 32'h415213d0} /* (25, 8, 31) {real, imag} */,
  {32'hc1970cdf, 32'h4118abe0} /* (25, 8, 30) {real, imag} */,
  {32'h4192d514, 32'h404f0906} /* (25, 8, 29) {real, imag} */,
  {32'hc04f6da0, 32'hbfc94e4c} /* (25, 8, 28) {real, imag} */,
  {32'hc1733594, 32'h3fa57604} /* (25, 8, 27) {real, imag} */,
  {32'hbe54f1a0, 32'hbfcc1ee8} /* (25, 8, 26) {real, imag} */,
  {32'h41a9f621, 32'hc0667b06} /* (25, 8, 25) {real, imag} */,
  {32'h40e836ea, 32'hbf901770} /* (25, 8, 24) {real, imag} */,
  {32'h419a0ad0, 32'hc18a2d84} /* (25, 8, 23) {real, imag} */,
  {32'h40b8494c, 32'hc0717172} /* (25, 8, 22) {real, imag} */,
  {32'hc04136c6, 32'hc114641c} /* (25, 8, 21) {real, imag} */,
  {32'h3edfb9a8, 32'h410a896a} /* (25, 8, 20) {real, imag} */,
  {32'hc0f4286e, 32'h41000618} /* (25, 8, 19) {real, imag} */,
  {32'hc156d18a, 32'h40a4b51e} /* (25, 8, 18) {real, imag} */,
  {32'hc0995df7, 32'hc01e6d7a} /* (25, 8, 17) {real, imag} */,
  {32'h4129fbac, 32'hc10bc557} /* (25, 8, 16) {real, imag} */,
  {32'h40fd077a, 32'h4177d72c} /* (25, 8, 15) {real, imag} */,
  {32'h405383a8, 32'hc18d106b} /* (25, 8, 14) {real, imag} */,
  {32'h3fc591d8, 32'hc19cc25b} /* (25, 8, 13) {real, imag} */,
  {32'hc14d2d90, 32'h41343660} /* (25, 8, 12) {real, imag} */,
  {32'h413d8652, 32'hc129b408} /* (25, 8, 11) {real, imag} */,
  {32'h411aab6a, 32'h40698a8a} /* (25, 8, 10) {real, imag} */,
  {32'h409e7b40, 32'h401a89b4} /* (25, 8, 9) {real, imag} */,
  {32'hc0ae9970, 32'hc1989e30} /* (25, 8, 8) {real, imag} */,
  {32'hc02d0482, 32'hc14e6344} /* (25, 8, 7) {real, imag} */,
  {32'hc1754518, 32'hc0c2cf94} /* (25, 8, 6) {real, imag} */,
  {32'hbf9c7080, 32'h3ff5b8fc} /* (25, 8, 5) {real, imag} */,
  {32'hc0f5d92a, 32'h41ee730f} /* (25, 8, 4) {real, imag} */,
  {32'hc1dff362, 32'h411297d6} /* (25, 8, 3) {real, imag} */,
  {32'hc1f39902, 32'hc1083a64} /* (25, 8, 2) {real, imag} */,
  {32'h4233094d, 32'h414f4c7a} /* (25, 8, 1) {real, imag} */,
  {32'h417df5fa, 32'h407e68ee} /* (25, 8, 0) {real, imag} */,
  {32'hc18ad48b, 32'hc1354daa} /* (25, 7, 31) {real, imag} */,
  {32'h40af3e3c, 32'hc0faa3a0} /* (25, 7, 30) {real, imag} */,
  {32'hc07e4b14, 32'hc1b347a6} /* (25, 7, 29) {real, imag} */,
  {32'hc11fbb24, 32'h40c8adcc} /* (25, 7, 28) {real, imag} */,
  {32'h3f69e68c, 32'h40b4e45e} /* (25, 7, 27) {real, imag} */,
  {32'hc1184002, 32'hc12415e0} /* (25, 7, 26) {real, imag} */,
  {32'h40d82542, 32'hc1327b17} /* (25, 7, 25) {real, imag} */,
  {32'h4030ec86, 32'hc2049174} /* (25, 7, 24) {real, imag} */,
  {32'h40d87688, 32'h412d5b1f} /* (25, 7, 23) {real, imag} */,
  {32'hc14378fe, 32'h40823dcc} /* (25, 7, 22) {real, imag} */,
  {32'hc0662472, 32'hc172fa71} /* (25, 7, 21) {real, imag} */,
  {32'hbe9a2168, 32'h406cdbb9} /* (25, 7, 20) {real, imag} */,
  {32'hc15da76d, 32'hc1715148} /* (25, 7, 19) {real, imag} */,
  {32'h40b43fe1, 32'hc0f45803} /* (25, 7, 18) {real, imag} */,
  {32'h4052ab41, 32'h412081d8} /* (25, 7, 17) {real, imag} */,
  {32'hc02d7ade, 32'h3fe27d44} /* (25, 7, 16) {real, imag} */,
  {32'hc0d4377c, 32'h40d2e07a} /* (25, 7, 15) {real, imag} */,
  {32'hbf20a488, 32'hc04e5f6d} /* (25, 7, 14) {real, imag} */,
  {32'h4184969e, 32'h412c9750} /* (25, 7, 13) {real, imag} */,
  {32'hc091ff30, 32'h415ac813} /* (25, 7, 12) {real, imag} */,
  {32'h40de08b8, 32'hc1376f92} /* (25, 7, 11) {real, imag} */,
  {32'hc1b2401c, 32'hc1568c1b} /* (25, 7, 10) {real, imag} */,
  {32'hc09ce534, 32'hc1350910} /* (25, 7, 9) {real, imag} */,
  {32'h409f565b, 32'h40f4d1f4} /* (25, 7, 8) {real, imag} */,
  {32'h40522f0c, 32'hc140a940} /* (25, 7, 7) {real, imag} */,
  {32'hc145a902, 32'hbea7a840} /* (25, 7, 6) {real, imag} */,
  {32'hc18c5bf6, 32'h41528bfe} /* (25, 7, 5) {real, imag} */,
  {32'h41a2fe4c, 32'hc1b202f3} /* (25, 7, 4) {real, imag} */,
  {32'h40fe936a, 32'h41d584cc} /* (25, 7, 3) {real, imag} */,
  {32'h400180a4, 32'h41d14108} /* (25, 7, 2) {real, imag} */,
  {32'hc1d708f7, 32'hc1a0f6b1} /* (25, 7, 1) {real, imag} */,
  {32'hc203d5fe, 32'hc029c4ca} /* (25, 7, 0) {real, imag} */,
  {32'h412161d2, 32'hc1495ee7} /* (25, 6, 31) {real, imag} */,
  {32'hc1789a47, 32'h416784f3} /* (25, 6, 30) {real, imag} */,
  {32'hc0f522e7, 32'h407e53f2} /* (25, 6, 29) {real, imag} */,
  {32'h41c482ea, 32'hc1bcf13c} /* (25, 6, 28) {real, imag} */,
  {32'hc0aad513, 32'hc141be39} /* (25, 6, 27) {real, imag} */,
  {32'hc0a827f4, 32'h41f9ee26} /* (25, 6, 26) {real, imag} */,
  {32'hc0a6f290, 32'h41183f23} /* (25, 6, 25) {real, imag} */,
  {32'h4094aca2, 32'hc0a33576} /* (25, 6, 24) {real, imag} */,
  {32'h40e7204d, 32'h41841b3f} /* (25, 6, 23) {real, imag} */,
  {32'h40a5008c, 32'h413060ff} /* (25, 6, 22) {real, imag} */,
  {32'h40951cbb, 32'hc0a12a8a} /* (25, 6, 21) {real, imag} */,
  {32'h4126afd0, 32'hc033dab0} /* (25, 6, 20) {real, imag} */,
  {32'hc0d25501, 32'hc0a4ee69} /* (25, 6, 19) {real, imag} */,
  {32'hc0e17fd8, 32'h3f117988} /* (25, 6, 18) {real, imag} */,
  {32'h409b5be2, 32'hc0029d40} /* (25, 6, 17) {real, imag} */,
  {32'h417b1526, 32'h3ef9ddf0} /* (25, 6, 16) {real, imag} */,
  {32'hbe800178, 32'h414e1e4e} /* (25, 6, 15) {real, imag} */,
  {32'hc0d180a6, 32'h406e0796} /* (25, 6, 14) {real, imag} */,
  {32'h4158a848, 32'hc0f042f2} /* (25, 6, 13) {real, imag} */,
  {32'hbf489ac8, 32'h3fa0caa0} /* (25, 6, 12) {real, imag} */,
  {32'hc0d28e72, 32'hc03eab44} /* (25, 6, 11) {real, imag} */,
  {32'h418a54e5, 32'h40ccf76c} /* (25, 6, 10) {real, imag} */,
  {32'h4115293a, 32'h3fd1856e} /* (25, 6, 9) {real, imag} */,
  {32'h4188e4c9, 32'h410a2690} /* (25, 6, 8) {real, imag} */,
  {32'hc196d020, 32'hc0da20bc} /* (25, 6, 7) {real, imag} */,
  {32'h415f8948, 32'hc13474fc} /* (25, 6, 6) {real, imag} */,
  {32'h4094659c, 32'hbf39a474} /* (25, 6, 5) {real, imag} */,
  {32'h40c9778e, 32'hc1bc6d8d} /* (25, 6, 4) {real, imag} */,
  {32'h40a5fac4, 32'hc0880ab0} /* (25, 6, 3) {real, imag} */,
  {32'h41c32d6e, 32'hc084b04c} /* (25, 6, 2) {real, imag} */,
  {32'hc09640a1, 32'h40b98f75} /* (25, 6, 1) {real, imag} */,
  {32'h4009d972, 32'h3f520d00} /* (25, 6, 0) {real, imag} */,
  {32'h42a8f802, 32'hc184a4e4} /* (25, 5, 31) {real, imag} */,
  {32'hc2079cda, 32'hc1d87950} /* (25, 5, 30) {real, imag} */,
  {32'h41391df4, 32'hc0e3ff62} /* (25, 5, 29) {real, imag} */,
  {32'h40941bb5, 32'h417b89ec} /* (25, 5, 28) {real, imag} */,
  {32'hc223f762, 32'h40ee848c} /* (25, 5, 27) {real, imag} */,
  {32'h41ba2781, 32'hc14dc8c2} /* (25, 5, 26) {real, imag} */,
  {32'h419d87ad, 32'hc16c0be0} /* (25, 5, 25) {real, imag} */,
  {32'hc0a08e68, 32'h41477fd0} /* (25, 5, 24) {real, imag} */,
  {32'hc0886c84, 32'hc109edc8} /* (25, 5, 23) {real, imag} */,
  {32'h40ac70bd, 32'h40d3b53e} /* (25, 5, 22) {real, imag} */,
  {32'hc171087e, 32'hbf3e75d8} /* (25, 5, 21) {real, imag} */,
  {32'h4164da6b, 32'h40975e26} /* (25, 5, 20) {real, imag} */,
  {32'h4135ffe8, 32'h404797a1} /* (25, 5, 19) {real, imag} */,
  {32'hc0205594, 32'h4156eca8} /* (25, 5, 18) {real, imag} */,
  {32'hc1669352, 32'hc00d9da0} /* (25, 5, 17) {real, imag} */,
  {32'h3fcf91ec, 32'h3f0a0bb8} /* (25, 5, 16) {real, imag} */,
  {32'hc058e84e, 32'h41493f97} /* (25, 5, 15) {real, imag} */,
  {32'h40a8aa02, 32'h41004d78} /* (25, 5, 14) {real, imag} */,
  {32'hbe169f78, 32'h40dbadc2} /* (25, 5, 13) {real, imag} */,
  {32'h3f9fd11a, 32'h40ff99e8} /* (25, 5, 12) {real, imag} */,
  {32'hc04ce098, 32'hc1b890b6} /* (25, 5, 11) {real, imag} */,
  {32'h3fde39b0, 32'hc16d6cd6} /* (25, 5, 10) {real, imag} */,
  {32'hc18dab18, 32'hc13fb2b6} /* (25, 5, 9) {real, imag} */,
  {32'hc028b09c, 32'hc0038a04} /* (25, 5, 8) {real, imag} */,
  {32'h4117b582, 32'h41027211} /* (25, 5, 7) {real, imag} */,
  {32'hc040d3c8, 32'h409cdadc} /* (25, 5, 6) {real, imag} */,
  {32'h41e5cf84, 32'hc1176e91} /* (25, 5, 5) {real, imag} */,
  {32'hc1381486, 32'h41595528} /* (25, 5, 4) {real, imag} */,
  {32'h3f711870, 32'hc202c8a4} /* (25, 5, 3) {real, imag} */,
  {32'hc20556c6, 32'hc228ec60} /* (25, 5, 2) {real, imag} */,
  {32'h42388489, 32'h429edf1e} /* (25, 5, 1) {real, imag} */,
  {32'h4209b2dc, 32'h424b057a} /* (25, 5, 0) {real, imag} */,
  {32'hc20b4cb0, 32'hc28ba980} /* (25, 4, 31) {real, imag} */,
  {32'h422bde28, 32'h4292508d} /* (25, 4, 30) {real, imag} */,
  {32'hc19e76c3, 32'hc0f55a6e} /* (25, 4, 29) {real, imag} */,
  {32'hc209d772, 32'hc21a93f5} /* (25, 4, 28) {real, imag} */,
  {32'h40c167df, 32'hbecb2e10} /* (25, 4, 27) {real, imag} */,
  {32'hc078bcd8, 32'hc1d79b3c} /* (25, 4, 26) {real, imag} */,
  {32'h410a4d82, 32'h411e4403} /* (25, 4, 25) {real, imag} */,
  {32'h3f10c830, 32'h4068e8d0} /* (25, 4, 24) {real, imag} */,
  {32'hc090bfea, 32'hc0e6ab51} /* (25, 4, 23) {real, imag} */,
  {32'hc13a97a6, 32'hc0acdbc0} /* (25, 4, 22) {real, imag} */,
  {32'h40e2c443, 32'h41853101} /* (25, 4, 21) {real, imag} */,
  {32'h3fe96b78, 32'hbec33560} /* (25, 4, 20) {real, imag} */,
  {32'hc0e53144, 32'h41067ab2} /* (25, 4, 19) {real, imag} */,
  {32'h418e9bee, 32'hc093e7d0} /* (25, 4, 18) {real, imag} */,
  {32'h3fc5be7c, 32'h40e8a313} /* (25, 4, 17) {real, imag} */,
  {32'hbefc99fe, 32'h40bab18a} /* (25, 4, 16) {real, imag} */,
  {32'hc0b41313, 32'hbfabce2c} /* (25, 4, 15) {real, imag} */,
  {32'h3ff3a3e0, 32'hc07f2100} /* (25, 4, 14) {real, imag} */,
  {32'h410253f6, 32'h40e1c37c} /* (25, 4, 13) {real, imag} */,
  {32'h40251f20, 32'hbf5f4f30} /* (25, 4, 12) {real, imag} */,
  {32'h412afa78, 32'h41ae7fa2} /* (25, 4, 11) {real, imag} */,
  {32'h40180685, 32'hc09312d3} /* (25, 4, 10) {real, imag} */,
  {32'hc0f4b68c, 32'h413c036e} /* (25, 4, 9) {real, imag} */,
  {32'h417b6267, 32'h41f982f6} /* (25, 4, 8) {real, imag} */,
  {32'hc1b7d815, 32'h411fd46d} /* (25, 4, 7) {real, imag} */,
  {32'hc1cd1b52, 32'h41d36dd4} /* (25, 4, 6) {real, imag} */,
  {32'h4116da0c, 32'h3e118b80} /* (25, 4, 5) {real, imag} */,
  {32'h4111834b, 32'hc27eae9b} /* (25, 4, 4) {real, imag} */,
  {32'hc0a4025c, 32'hc07dc67a} /* (25, 4, 3) {real, imag} */,
  {32'h4264ec3e, 32'h424350b5} /* (25, 4, 2) {real, imag} */,
  {32'hc2e053b4, 32'hc181c330} /* (25, 4, 1) {real, imag} */,
  {32'hc24a60d6, 32'hc2174fad} /* (25, 4, 0) {real, imag} */,
  {32'h428d6642, 32'hc29f3f28} /* (25, 3, 31) {real, imag} */,
  {32'hc123e0a8, 32'h426bde3d} /* (25, 3, 30) {real, imag} */,
  {32'h41addf9e, 32'h41580e26} /* (25, 3, 29) {real, imag} */,
  {32'hc1ce4370, 32'hc1a08bd4} /* (25, 3, 28) {real, imag} */,
  {32'h416abea8, 32'hc01821e8} /* (25, 3, 27) {real, imag} */,
  {32'hbf2b5230, 32'h40d4ba12} /* (25, 3, 26) {real, imag} */,
  {32'h40c9f958, 32'h4109e0fa} /* (25, 3, 25) {real, imag} */,
  {32'h415e588d, 32'h41db916c} /* (25, 3, 24) {real, imag} */,
  {32'h407369b4, 32'hc1692c34} /* (25, 3, 23) {real, imag} */,
  {32'hc08e16be, 32'h40e9ba4a} /* (25, 3, 22) {real, imag} */,
  {32'hbf8d6c22, 32'h40c910e0} /* (25, 3, 21) {real, imag} */,
  {32'hc03f1ab9, 32'h412ed7a0} /* (25, 3, 20) {real, imag} */,
  {32'h4148745a, 32'hc0afd396} /* (25, 3, 19) {real, imag} */,
  {32'h41191012, 32'h40b9eeae} /* (25, 3, 18) {real, imag} */,
  {32'h3e0c44b8, 32'hc0b46f5d} /* (25, 3, 17) {real, imag} */,
  {32'hc0d9fbd5, 32'h40cecdf1} /* (25, 3, 16) {real, imag} */,
  {32'h4061958c, 32'h4026a4b7} /* (25, 3, 15) {real, imag} */,
  {32'hc16609ca, 32'hc05111b2} /* (25, 3, 14) {real, imag} */,
  {32'h403f0a54, 32'h4103a276} /* (25, 3, 13) {real, imag} */,
  {32'h4148094d, 32'hc0a5df7a} /* (25, 3, 12) {real, imag} */,
  {32'hc18a8f00, 32'hc0529ac4} /* (25, 3, 11) {real, imag} */,
  {32'hbfea2caa, 32'h403e7304} /* (25, 3, 10) {real, imag} */,
  {32'hc0083f66, 32'hc0ea6a4a} /* (25, 3, 9) {real, imag} */,
  {32'hc13b0c1e, 32'hc104cd56} /* (25, 3, 8) {real, imag} */,
  {32'hc0c2ff4c, 32'h3f8d42be} /* (25, 3, 7) {real, imag} */,
  {32'hc03549d8, 32'h418e9266} /* (25, 3, 6) {real, imag} */,
  {32'hc1d2fc5e, 32'hc175dcd8} /* (25, 3, 5) {real, imag} */,
  {32'h41c5d2e2, 32'hc0a516c8} /* (25, 3, 4) {real, imag} */,
  {32'hc00c1486, 32'hc18dcfcd} /* (25, 3, 3) {real, imag} */,
  {32'h40c3a557, 32'h42bcd155} /* (25, 3, 2) {real, imag} */,
  {32'hc2b703a1, 32'hc23c75bf} /* (25, 3, 1) {real, imag} */,
  {32'h429cc1ef, 32'h419c36dc} /* (25, 3, 0) {real, imag} */,
  {32'h44124ac2, 32'h42974649} /* (25, 2, 31) {real, imag} */,
  {32'hc38b0d3a, 32'h424b1585} /* (25, 2, 30) {real, imag} */,
  {32'h41cb205e, 32'hc1e52d8e} /* (25, 2, 29) {real, imag} */,
  {32'h4200646f, 32'hc21d9bb9} /* (25, 2, 28) {real, imag} */,
  {32'h3f98c7f0, 32'hc152c160} /* (25, 2, 27) {real, imag} */,
  {32'h40c8d3e0, 32'h3f4123f0} /* (25, 2, 26) {real, imag} */,
  {32'hbbaf1800, 32'h41f92af4} /* (25, 2, 25) {real, imag} */,
  {32'hc14ca1ad, 32'h42022582} /* (25, 2, 24) {real, imag} */,
  {32'h410fe85f, 32'h3f223f38} /* (25, 2, 23) {real, imag} */,
  {32'h40f07241, 32'hc1c87158} /* (25, 2, 22) {real, imag} */,
  {32'hc037db4a, 32'hc116d028} /* (25, 2, 21) {real, imag} */,
  {32'hbe8bf2b0, 32'hc0f39ca0} /* (25, 2, 20) {real, imag} */,
  {32'h3f2437cc, 32'h3ff024f4} /* (25, 2, 19) {real, imag} */,
  {32'hc0a3d4f4, 32'h40f016c0} /* (25, 2, 18) {real, imag} */,
  {32'hc0d48374, 32'hc14ddffa} /* (25, 2, 17) {real, imag} */,
  {32'hc0ea1156, 32'h40cd9fe1} /* (25, 2, 16) {real, imag} */,
  {32'h40e0c574, 32'h409a5ed1} /* (25, 2, 15) {real, imag} */,
  {32'hbfe7cd48, 32'h41503225} /* (25, 2, 14) {real, imag} */,
  {32'h4109a426, 32'h3f97197c} /* (25, 2, 13) {real, imag} */,
  {32'hbfb3a4a8, 32'hc195536b} /* (25, 2, 12) {real, imag} */,
  {32'hc0da26df, 32'hc1eec50f} /* (25, 2, 11) {real, imag} */,
  {32'h415f2f14, 32'h41060087} /* (25, 2, 10) {real, imag} */,
  {32'hbfab8274, 32'hc16cc5f6} /* (25, 2, 9) {real, imag} */,
  {32'hc187854d, 32'hc0d87b6e} /* (25, 2, 8) {real, imag} */,
  {32'h41ea4924, 32'h4169d390} /* (25, 2, 7) {real, imag} */,
  {32'hc0a2a9fe, 32'hc143250d} /* (25, 2, 6) {real, imag} */,
  {32'hc28778e3, 32'hc20769b3} /* (25, 2, 5) {real, imag} */,
  {32'h42430485, 32'hc04e70f4} /* (25, 2, 4) {real, imag} */,
  {32'hc19386fb, 32'hc0f806b4} /* (25, 2, 3) {real, imag} */,
  {32'hc32b65b9, 32'h42135d2d} /* (25, 2, 2) {real, imag} */,
  {32'h43b1396f, 32'h418b3d40} /* (25, 2, 1) {real, imag} */,
  {32'h43af9197, 32'h41a1350c} /* (25, 2, 0) {real, imag} */,
  {32'hc4464ef4, 32'h43323f18} /* (25, 1, 31) {real, imag} */,
  {32'h433c3442, 32'h42dfe528} /* (25, 1, 30) {real, imag} */,
  {32'h41d217c5, 32'hc1afe7c8} /* (25, 1, 29) {real, imag} */,
  {32'hc223353e, 32'hc1c8d99e} /* (25, 1, 28) {real, imag} */,
  {32'h42878014, 32'hc14e00d6} /* (25, 1, 27) {real, imag} */,
  {32'hc1b494fb, 32'hc0abd18c} /* (25, 1, 26) {real, imag} */,
  {32'hc180ef26, 32'h41283732} /* (25, 1, 25) {real, imag} */,
  {32'h3fee04f0, 32'hbfbb3408} /* (25, 1, 24) {real, imag} */,
  {32'h400856a9, 32'h4172155e} /* (25, 1, 23) {real, imag} */,
  {32'hbfe8b750, 32'hc187fb38} /* (25, 1, 22) {real, imag} */,
  {32'h41c12222, 32'hc1721ba8} /* (25, 1, 21) {real, imag} */,
  {32'h414f9a2e, 32'hc0755af7} /* (25, 1, 20) {real, imag} */,
  {32'hc0bbd3fd, 32'hbf673428} /* (25, 1, 19) {real, imag} */,
  {32'h40ce2313, 32'hc187981c} /* (25, 1, 18) {real, imag} */,
  {32'hc05d30c6, 32'h409e5d68} /* (25, 1, 17) {real, imag} */,
  {32'h401de935, 32'h412cee39} /* (25, 1, 16) {real, imag} */,
  {32'hc123ad74, 32'hc16b3d5f} /* (25, 1, 15) {real, imag} */,
  {32'hc13aaa8d, 32'h4170d1e0} /* (25, 1, 14) {real, imag} */,
  {32'h40d69b90, 32'hc0ea93da} /* (25, 1, 13) {real, imag} */,
  {32'hbfb74e4e, 32'h3fe4efcc} /* (25, 1, 12) {real, imag} */,
  {32'h41442a38, 32'h41c83c00} /* (25, 1, 11) {real, imag} */,
  {32'h40b89066, 32'h3fabb4a8} /* (25, 1, 10) {real, imag} */,
  {32'h410b0e3d, 32'hc10b89ba} /* (25, 1, 9) {real, imag} */,
  {32'h4103e51f, 32'h41fb5807} /* (25, 1, 8) {real, imag} */,
  {32'hc081714b, 32'h40348370} /* (25, 1, 7) {real, imag} */,
  {32'h416f6cb3, 32'h417e8b53} /* (25, 1, 6) {real, imag} */,
  {32'h42405e16, 32'h42357b70} /* (25, 1, 5) {real, imag} */,
  {32'hc00a35c0, 32'hc2753126} /* (25, 1, 4) {real, imag} */,
  {32'h421710a7, 32'hbfa5f380} /* (25, 1, 3) {real, imag} */,
  {32'h438543ce, 32'h438875b1} /* (25, 1, 2) {real, imag} */,
  {32'hc4924069, 32'hc42ea98b} /* (25, 1, 1) {real, imag} */,
  {32'hc493f352, 32'hc33fcf31} /* (25, 1, 0) {real, imag} */,
  {32'hc463a334, 32'h442d9fb2} /* (25, 0, 31) {real, imag} */,
  {32'h4274f99d, 32'hc233c9a4} /* (25, 0, 30) {real, imag} */,
  {32'h41d1fbc1, 32'hc1d782d7} /* (25, 0, 29) {real, imag} */,
  {32'h41c42766, 32'hc2901663} /* (25, 0, 28) {real, imag} */,
  {32'h42885bc8, 32'hc1213bfc} /* (25, 0, 27) {real, imag} */,
  {32'hc094cec5, 32'h41717d91} /* (25, 0, 26) {real, imag} */,
  {32'hbf10e378, 32'h3de11400} /* (25, 0, 25) {real, imag} */,
  {32'hc1a6ce92, 32'hc25e0c8a} /* (25, 0, 24) {real, imag} */,
  {32'h41384fc4, 32'hc1ae4e71} /* (25, 0, 23) {real, imag} */,
  {32'h3fe3dd04, 32'hbe906d68} /* (25, 0, 22) {real, imag} */,
  {32'h415fcbac, 32'hc0e65d57} /* (25, 0, 21) {real, imag} */,
  {32'hc157e5f8, 32'hc141688c} /* (25, 0, 20) {real, imag} */,
  {32'h4100d74c, 32'h40a12a80} /* (25, 0, 19) {real, imag} */,
  {32'hc0b86dc6, 32'hc1b4cefd} /* (25, 0, 18) {real, imag} */,
  {32'h40a9387c, 32'h3f3ff458} /* (25, 0, 17) {real, imag} */,
  {32'h419c8272, 32'h00000000} /* (25, 0, 16) {real, imag} */,
  {32'h40a9387c, 32'hbf3ff458} /* (25, 0, 15) {real, imag} */,
  {32'hc0b86dc6, 32'h41b4cefd} /* (25, 0, 14) {real, imag} */,
  {32'h4100d74c, 32'hc0a12a80} /* (25, 0, 13) {real, imag} */,
  {32'hc157e5f8, 32'h4141688c} /* (25, 0, 12) {real, imag} */,
  {32'h415fcbac, 32'h40e65d57} /* (25, 0, 11) {real, imag} */,
  {32'h3fe3dd04, 32'h3e906d68} /* (25, 0, 10) {real, imag} */,
  {32'h41384fc4, 32'h41ae4e71} /* (25, 0, 9) {real, imag} */,
  {32'hc1a6ce92, 32'h425e0c8a} /* (25, 0, 8) {real, imag} */,
  {32'hbf10e378, 32'hbde11400} /* (25, 0, 7) {real, imag} */,
  {32'hc094cec5, 32'hc1717d91} /* (25, 0, 6) {real, imag} */,
  {32'h42885bc8, 32'h41213bfc} /* (25, 0, 5) {real, imag} */,
  {32'h41c42766, 32'h42901663} /* (25, 0, 4) {real, imag} */,
  {32'h41d1fbc1, 32'h41d782d7} /* (25, 0, 3) {real, imag} */,
  {32'h4274f99d, 32'h4233c9a4} /* (25, 0, 2) {real, imag} */,
  {32'hc463a334, 32'hc42d9fb2} /* (25, 0, 1) {real, imag} */,
  {32'hc4bbf222, 32'h00000000} /* (25, 0, 0) {real, imag} */,
  {32'hc4da1b49, 32'h447ba9e1} /* (24, 31, 31) {real, imag} */,
  {32'h43d3f596, 32'hc3cc952c} /* (24, 31, 30) {real, imag} */,
  {32'h41acdc58, 32'hc176266a} /* (24, 31, 29) {real, imag} */,
  {32'hc1c8c5bc, 32'h4240efb0} /* (24, 31, 28) {real, imag} */,
  {32'h4286aabc, 32'hc23d260a} /* (24, 31, 27) {real, imag} */,
  {32'h417a6cdc, 32'h3fa01aa8} /* (24, 31, 26) {real, imag} */,
  {32'hc1465812, 32'h416b890a} /* (24, 31, 25) {real, imag} */,
  {32'h41c97c17, 32'hc1d9d703} /* (24, 31, 24) {real, imag} */,
  {32'hbd73f480, 32'hc0fdbbe6} /* (24, 31, 23) {real, imag} */,
  {32'hc0d7a006, 32'h40f6db3a} /* (24, 31, 22) {real, imag} */,
  {32'h40cc3c0d, 32'hc1811cc6} /* (24, 31, 21) {real, imag} */,
  {32'hc05c2fc6, 32'h3f340ca0} /* (24, 31, 20) {real, imag} */,
  {32'hbdbb4ba0, 32'h414efacc} /* (24, 31, 19) {real, imag} */,
  {32'hc0e9c1a8, 32'hc17d4c14} /* (24, 31, 18) {real, imag} */,
  {32'hbebd1c00, 32'h405c9e08} /* (24, 31, 17) {real, imag} */,
  {32'h3f446fc8, 32'h404209b4} /* (24, 31, 16) {real, imag} */,
  {32'h401bd268, 32'hc0dfb4ea} /* (24, 31, 15) {real, imag} */,
  {32'hbfd87bf8, 32'h418aa1f2} /* (24, 31, 14) {real, imag} */,
  {32'h4097426a, 32'h4191c677} /* (24, 31, 13) {real, imag} */,
  {32'hc1a3941a, 32'hc10842c2} /* (24, 31, 12) {real, imag} */,
  {32'h411b3418, 32'h41ce1184} /* (24, 31, 11) {real, imag} */,
  {32'h40ad67a2, 32'h41a21b46} /* (24, 31, 10) {real, imag} */,
  {32'h415fb864, 32'hc09fab2d} /* (24, 31, 9) {real, imag} */,
  {32'h41edf247, 32'h41f56b36} /* (24, 31, 8) {real, imag} */,
  {32'hc1a995b9, 32'hc1971191} /* (24, 31, 7) {real, imag} */,
  {32'hc1e4ff74, 32'h40de3bb6} /* (24, 31, 6) {real, imag} */,
  {32'h42bd1066, 32'h411dc783} /* (24, 31, 5) {real, imag} */,
  {32'hc2b1d835, 32'h418f146e} /* (24, 31, 4) {real, imag} */,
  {32'h423cef3e, 32'h41d067d0} /* (24, 31, 3) {real, imag} */,
  {32'h438a21ab, 32'hc2b55130} /* (24, 31, 2) {real, imag} */,
  {32'hc4977b8b, 32'hc397591a} /* (24, 31, 1) {real, imag} */,
  {32'hc4cea4af, 32'h435bd352} /* (24, 31, 0) {real, imag} */,
  {32'h4403bf18, 32'h420b6cb7} /* (24, 30, 31) {real, imag} */,
  {32'hc384b84e, 32'hc221f5cc} /* (24, 30, 30) {real, imag} */,
  {32'h410689ce, 32'h4224e195} /* (24, 30, 29) {real, imag} */,
  {32'h42b49c5c, 32'hc1a8ef62} /* (24, 30, 28) {real, imag} */,
  {32'hc29e93f2, 32'h421c20fb} /* (24, 30, 27) {real, imag} */,
  {32'h41c85b5a, 32'hbd8a57c0} /* (24, 30, 26) {real, imag} */,
  {32'h417633d0, 32'hc0e0b594} /* (24, 30, 25) {real, imag} */,
  {32'hc18d9b6e, 32'hc0d1e0cf} /* (24, 30, 24) {real, imag} */,
  {32'h40f9165d, 32'hbed1be70} /* (24, 30, 23) {real, imag} */,
  {32'h4121e90f, 32'h418abe24} /* (24, 30, 22) {real, imag} */,
  {32'hc106951e, 32'h418a8943} /* (24, 30, 21) {real, imag} */,
  {32'h411e9f07, 32'hc13eb63c} /* (24, 30, 20) {real, imag} */,
  {32'hc0929db8, 32'h416cd54e} /* (24, 30, 19) {real, imag} */,
  {32'hbfb76e04, 32'h409ec6f6} /* (24, 30, 18) {real, imag} */,
  {32'h40435ade, 32'h40c50d37} /* (24, 30, 17) {real, imag} */,
  {32'hc0b2c55c, 32'hc07b3631} /* (24, 30, 16) {real, imag} */,
  {32'hc0bc473e, 32'hbf3f3598} /* (24, 30, 15) {real, imag} */,
  {32'h3fe81c4a, 32'hc0e1a8ff} /* (24, 30, 14) {real, imag} */,
  {32'hc0b67834, 32'hc124fbdf} /* (24, 30, 13) {real, imag} */,
  {32'hc00870b4, 32'h41743f38} /* (24, 30, 12) {real, imag} */,
  {32'h41e617f8, 32'hc158d9fe} /* (24, 30, 11) {real, imag} */,
  {32'hc11f356f, 32'h41611de0} /* (24, 30, 10) {real, imag} */,
  {32'h418916ba, 32'hc036bbbe} /* (24, 30, 9) {real, imag} */,
  {32'h3ecd80c0, 32'hc21581f2} /* (24, 30, 8) {real, imag} */,
  {32'hc12a64c7, 32'hc12798e2} /* (24, 30, 7) {real, imag} */,
  {32'hc1c1d6bc, 32'hc12976a5} /* (24, 30, 6) {real, imag} */,
  {32'hc1fe4eb0, 32'hc127d3d1} /* (24, 30, 5) {real, imag} */,
  {32'h424c8c7c, 32'h4244b9aa} /* (24, 30, 4) {real, imag} */,
  {32'h42371b66, 32'h41e04c0a} /* (24, 30, 3) {real, imag} */,
  {32'hc3d475c7, 32'hc2c91990} /* (24, 30, 2) {real, imag} */,
  {32'h4461eb34, 32'hc26216af} /* (24, 30, 1) {real, imag} */,
  {32'h43f0ba5e, 32'hc2921bb6} /* (24, 30, 0) {real, imag} */,
  {32'hc2ea3ab7, 32'h42ae5ab6} /* (24, 29, 31) {real, imag} */,
  {32'hc1bd8f3c, 32'hc2fb3b78} /* (24, 29, 30) {real, imag} */,
  {32'h3e641d40, 32'h4072ac48} /* (24, 29, 29) {real, imag} */,
  {32'h42353f41, 32'h419c749e} /* (24, 29, 28) {real, imag} */,
  {32'hc0f4c42d, 32'h41974d74} /* (24, 29, 27) {real, imag} */,
  {32'hc17947b9, 32'hc1fb27a8} /* (24, 29, 26) {real, imag} */,
  {32'hc140b7c2, 32'h3f6a4a60} /* (24, 29, 25) {real, imag} */,
  {32'h404e781c, 32'hc07f605e} /* (24, 29, 24) {real, imag} */,
  {32'h41237a9c, 32'h403111da} /* (24, 29, 23) {real, imag} */,
  {32'h40bfb824, 32'h3e9e5a58} /* (24, 29, 22) {real, imag} */,
  {32'h40f486fe, 32'hbf30a94c} /* (24, 29, 21) {real, imag} */,
  {32'hbfefeac8, 32'h3fa97c70} /* (24, 29, 20) {real, imag} */,
  {32'hc1c7c258, 32'h40757863} /* (24, 29, 19) {real, imag} */,
  {32'hbe8f6978, 32'hc011da00} /* (24, 29, 18) {real, imag} */,
  {32'h3fa1a4e8, 32'h3fc732c0} /* (24, 29, 17) {real, imag} */,
  {32'h40ce5534, 32'h405980f4} /* (24, 29, 16) {real, imag} */,
  {32'hc03d6eac, 32'hc01c51d3} /* (24, 29, 15) {real, imag} */,
  {32'h4119eda7, 32'hc1b70f59} /* (24, 29, 14) {real, imag} */,
  {32'hc00d48ac, 32'h41981ee6} /* (24, 29, 13) {real, imag} */,
  {32'h3fe88362, 32'hc0c514c1} /* (24, 29, 12) {real, imag} */,
  {32'hc08808b6, 32'h418ab045} /* (24, 29, 11) {real, imag} */,
  {32'h40d07c55, 32'hc10b42fe} /* (24, 29, 10) {real, imag} */,
  {32'hc19c1dc0, 32'hc0997d6d} /* (24, 29, 9) {real, imag} */,
  {32'hc11ddd94, 32'hc1abcb94} /* (24, 29, 8) {real, imag} */,
  {32'hc0b0bddc, 32'h415e12ca} /* (24, 29, 7) {real, imag} */,
  {32'hc0b24cc2, 32'hc12762ec} /* (24, 29, 6) {real, imag} */,
  {32'h4219523e, 32'hc109de0d} /* (24, 29, 5) {real, imag} */,
  {32'hc1b0c5a2, 32'h41fcc259} /* (24, 29, 4) {real, imag} */,
  {32'h412e0e67, 32'hc1ee17d9} /* (24, 29, 3) {real, imag} */,
  {32'hc28909d8, 32'hc2aa7b68} /* (24, 29, 2) {real, imag} */,
  {32'h42ee42f4, 32'h42bb5b5c} /* (24, 29, 1) {real, imag} */,
  {32'h42baac1c, 32'hc1332833} /* (24, 29, 0) {real, imag} */,
  {32'hc30f7771, 32'h420d80e7} /* (24, 28, 31) {real, imag} */,
  {32'h42f69f0c, 32'hc24e413e} /* (24, 28, 30) {real, imag} */,
  {32'h41acbf7c, 32'h4144c790} /* (24, 28, 29) {real, imag} */,
  {32'h41d9b7e6, 32'h425d0dee} /* (24, 28, 28) {real, imag} */,
  {32'hc11622e1, 32'hc1adfb16} /* (24, 28, 27) {real, imag} */,
  {32'hc1d12acd, 32'hc05b0574} /* (24, 28, 26) {real, imag} */,
  {32'hc1a91dd4, 32'hc0d561fc} /* (24, 28, 25) {real, imag} */,
  {32'hc09c8886, 32'hc1558dee} /* (24, 28, 24) {real, imag} */,
  {32'h41724d46, 32'hc0bee805} /* (24, 28, 23) {real, imag} */,
  {32'h4138bd7f, 32'h41808031} /* (24, 28, 22) {real, imag} */,
  {32'hc029feda, 32'hc18213d6} /* (24, 28, 21) {real, imag} */,
  {32'hc11711e0, 32'h4116043e} /* (24, 28, 20) {real, imag} */,
  {32'h40c6e964, 32'h41215006} /* (24, 28, 19) {real, imag} */,
  {32'h408160ae, 32'hc1126220} /* (24, 28, 18) {real, imag} */,
  {32'hbdcd8680, 32'h40f6ca73} /* (24, 28, 17) {real, imag} */,
  {32'hc0d567d2, 32'hc03c08e7} /* (24, 28, 16) {real, imag} */,
  {32'h40e572e8, 32'hc1699fd0} /* (24, 28, 15) {real, imag} */,
  {32'h40a72405, 32'h40bc16ea} /* (24, 28, 14) {real, imag} */,
  {32'hc0a60275, 32'h40f022ee} /* (24, 28, 13) {real, imag} */,
  {32'hbfe7ece0, 32'h3fee9530} /* (24, 28, 12) {real, imag} */,
  {32'h412f6748, 32'hc0b77b8e} /* (24, 28, 11) {real, imag} */,
  {32'hc1885499, 32'hc0db455c} /* (24, 28, 10) {real, imag} */,
  {32'h41ac2990, 32'h41613998} /* (24, 28, 9) {real, imag} */,
  {32'h418adde4, 32'hc142ceab} /* (24, 28, 8) {real, imag} */,
  {32'hbff18830, 32'hc03a8748} /* (24, 28, 7) {real, imag} */,
  {32'h41adbcfe, 32'h419a5c43} /* (24, 28, 6) {real, imag} */,
  {32'h414795a8, 32'h416f6cb8} /* (24, 28, 5) {real, imag} */,
  {32'hc263deca, 32'h42123c7d} /* (24, 28, 4) {real, imag} */,
  {32'h3f981108, 32'h41ea39f2} /* (24, 28, 3) {real, imag} */,
  {32'h4292366f, 32'hc2c99c03} /* (24, 28, 2) {real, imag} */,
  {32'hc22f51f3, 32'h42bb7c9e} /* (24, 28, 1) {real, imag} */,
  {32'hc2970c33, 32'h41f776a4} /* (24, 28, 0) {real, imag} */,
  {32'h42543057, 32'hc2a7e872} /* (24, 27, 31) {real, imag} */,
  {32'hc205c5e0, 32'h42314f54} /* (24, 27, 30) {real, imag} */,
  {32'h4164cd44, 32'h411e4582} /* (24, 27, 29) {real, imag} */,
  {32'h4050ba0c, 32'hc20157cc} /* (24, 27, 28) {real, imag} */,
  {32'h3fe7c470, 32'h418a69a6} /* (24, 27, 27) {real, imag} */,
  {32'hc13fe688, 32'h3e59b380} /* (24, 27, 26) {real, imag} */,
  {32'h4141b58c, 32'hc0f56444} /* (24, 27, 25) {real, imag} */,
  {32'h402801d8, 32'h41849e9a} /* (24, 27, 24) {real, imag} */,
  {32'hc18812e2, 32'hc0c1b86e} /* (24, 27, 23) {real, imag} */,
  {32'h410477ec, 32'h40c158ee} /* (24, 27, 22) {real, imag} */,
  {32'h403c3e9b, 32'hc06423d4} /* (24, 27, 21) {real, imag} */,
  {32'h40dbe933, 32'h3fc2e406} /* (24, 27, 20) {real, imag} */,
  {32'hc17b5636, 32'h4138926b} /* (24, 27, 19) {real, imag} */,
  {32'hc0bc3010, 32'h415183d1} /* (24, 27, 18) {real, imag} */,
  {32'hc113444c, 32'h40726188} /* (24, 27, 17) {real, imag} */,
  {32'h40dccb34, 32'hc050c612} /* (24, 27, 16) {real, imag} */,
  {32'hc0ade89a, 32'hbf1ff5e6} /* (24, 27, 15) {real, imag} */,
  {32'hc0c25a2a, 32'hc0829510} /* (24, 27, 14) {real, imag} */,
  {32'h4101c6c8, 32'h411be939} /* (24, 27, 13) {real, imag} */,
  {32'hc04875de, 32'hbfe29874} /* (24, 27, 12) {real, imag} */,
  {32'hc0da5e72, 32'h3f0fa0a0} /* (24, 27, 11) {real, imag} */,
  {32'hc100da3d, 32'hc1223213} /* (24, 27, 10) {real, imag} */,
  {32'h3ffd82fa, 32'hbf780d18} /* (24, 27, 9) {real, imag} */,
  {32'hc0c03cbc, 32'h4114f407} /* (24, 27, 8) {real, imag} */,
  {32'hc1406f0a, 32'h413cb7fe} /* (24, 27, 7) {real, imag} */,
  {32'h41a48003, 32'hbfc5ef68} /* (24, 27, 6) {real, imag} */,
  {32'hc1fcc1ae, 32'hc1b5833a} /* (24, 27, 5) {real, imag} */,
  {32'h40b7cb82, 32'hc03eeb96} /* (24, 27, 4) {real, imag} */,
  {32'h40fc0ebd, 32'h418639f2} /* (24, 27, 3) {real, imag} */,
  {32'hc262499d, 32'hbf620c40} /* (24, 27, 2) {real, imag} */,
  {32'h42e763bc, 32'hc170a48d} /* (24, 27, 1) {real, imag} */,
  {32'h4241438a, 32'hc1f6d6c1} /* (24, 27, 0) {real, imag} */,
  {32'hc1111978, 32'h4089fe5b} /* (24, 26, 31) {real, imag} */,
  {32'h4210c538, 32'h405c70aa} /* (24, 26, 30) {real, imag} */,
  {32'h3f95d6bc, 32'hc0617376} /* (24, 26, 29) {real, imag} */,
  {32'h414c1193, 32'hc137ad74} /* (24, 26, 28) {real, imag} */,
  {32'h41b70c02, 32'hbfe556f8} /* (24, 26, 27) {real, imag} */,
  {32'h3d7d6880, 32'h41d33a36} /* (24, 26, 26) {real, imag} */,
  {32'hc137e425, 32'hc0e13e98} /* (24, 26, 25) {real, imag} */,
  {32'hc106aba6, 32'h41153478} /* (24, 26, 24) {real, imag} */,
  {32'h41bfcafa, 32'h4122c0ca} /* (24, 26, 23) {real, imag} */,
  {32'hc149e764, 32'hc10ac272} /* (24, 26, 22) {real, imag} */,
  {32'hc1b46da8, 32'hbe86fa20} /* (24, 26, 21) {real, imag} */,
  {32'hc0760737, 32'h4194597c} /* (24, 26, 20) {real, imag} */,
  {32'hc10f0e0a, 32'h4009e157} /* (24, 26, 19) {real, imag} */,
  {32'h41188a54, 32'hc0c4a596} /* (24, 26, 18) {real, imag} */,
  {32'h4085609e, 32'h40781e8c} /* (24, 26, 17) {real, imag} */,
  {32'hbe69df00, 32'h3fc71596} /* (24, 26, 16) {real, imag} */,
  {32'h3ddaefb0, 32'hc12713a1} /* (24, 26, 15) {real, imag} */,
  {32'h3fcf319c, 32'h410f6c61} /* (24, 26, 14) {real, imag} */,
  {32'h41b10193, 32'h40f64879} /* (24, 26, 13) {real, imag} */,
  {32'h4169c9fc, 32'h3f8576c0} /* (24, 26, 12) {real, imag} */,
  {32'hc1415463, 32'hc0dd6df0} /* (24, 26, 11) {real, imag} */,
  {32'hc120375e, 32'h40c233b3} /* (24, 26, 10) {real, imag} */,
  {32'hc1546a88, 32'hbe8d88c0} /* (24, 26, 9) {real, imag} */,
  {32'hbf372104, 32'h41b94bda} /* (24, 26, 8) {real, imag} */,
  {32'hc02aef31, 32'hc190c9a1} /* (24, 26, 7) {real, imag} */,
  {32'hc1e5bf77, 32'hc16318a0} /* (24, 26, 6) {real, imag} */,
  {32'hbf91848c, 32'h3f33a7c0} /* (24, 26, 5) {real, imag} */,
  {32'h41a1d446, 32'hc1a9c722} /* (24, 26, 4) {real, imag} */,
  {32'hc1028e68, 32'h41439cf5} /* (24, 26, 3) {real, imag} */,
  {32'hc0e28d1e, 32'hc17450aa} /* (24, 26, 2) {real, imag} */,
  {32'h4127404c, 32'h409de668} /* (24, 26, 1) {real, imag} */,
  {32'hc014d688, 32'h408ee3cc} /* (24, 26, 0) {real, imag} */,
  {32'hc1ce74de, 32'h41f477c7} /* (24, 25, 31) {real, imag} */,
  {32'hbefc3f30, 32'hc203b6c0} /* (24, 25, 30) {real, imag} */,
  {32'hc18363fa, 32'hc1b04c2c} /* (24, 25, 29) {real, imag} */,
  {32'h4104a084, 32'h3fdc8cab} /* (24, 25, 28) {real, imag} */,
  {32'hc115c452, 32'hc154f8c1} /* (24, 25, 27) {real, imag} */,
  {32'h3f3a2f40, 32'h40875817} /* (24, 25, 26) {real, imag} */,
  {32'hc0eb2600, 32'h414de22a} /* (24, 25, 25) {real, imag} */,
  {32'h40fc305a, 32'hc2026b74} /* (24, 25, 24) {real, imag} */,
  {32'h41810876, 32'h3ffa1908} /* (24, 25, 23) {real, imag} */,
  {32'hc136deb8, 32'hc1b31fa9} /* (24, 25, 22) {real, imag} */,
  {32'hc08d0b2b, 32'hc05a5912} /* (24, 25, 21) {real, imag} */,
  {32'h413a12ba, 32'hc11800a2} /* (24, 25, 20) {real, imag} */,
  {32'h4154befa, 32'h3fd5d662} /* (24, 25, 19) {real, imag} */,
  {32'h4191d8fa, 32'hc14aea74} /* (24, 25, 18) {real, imag} */,
  {32'hc0ad6530, 32'hc0f72870} /* (24, 25, 17) {real, imag} */,
  {32'hc09015ad, 32'h40bc8549} /* (24, 25, 16) {real, imag} */,
  {32'h4117384d, 32'h40e73fb3} /* (24, 25, 15) {real, imag} */,
  {32'hc17f155e, 32'hbfada0f4} /* (24, 25, 14) {real, imag} */,
  {32'hc0e54f6c, 32'hc0b39b78} /* (24, 25, 13) {real, imag} */,
  {32'h4010c83f, 32'hc15e7e2c} /* (24, 25, 12) {real, imag} */,
  {32'hc1931e78, 32'h40383abc} /* (24, 25, 11) {real, imag} */,
  {32'hc00f8e96, 32'h4071a820} /* (24, 25, 10) {real, imag} */,
  {32'h41a675bf, 32'hc1315da0} /* (24, 25, 9) {real, imag} */,
  {32'h41268770, 32'hc12b7aa4} /* (24, 25, 8) {real, imag} */,
  {32'h40c7b414, 32'hc15ec1aa} /* (24, 25, 7) {real, imag} */,
  {32'hc0ed6f4d, 32'h41eafd46} /* (24, 25, 6) {real, imag} */,
  {32'hc14289f5, 32'hc0242070} /* (24, 25, 5) {real, imag} */,
  {32'hc180d10b, 32'h4144eefd} /* (24, 25, 4) {real, imag} */,
  {32'hc1231d50, 32'hc0a75ee3} /* (24, 25, 3) {real, imag} */,
  {32'h40826bdc, 32'hc118e15e} /* (24, 25, 2) {real, imag} */,
  {32'hc1f6203b, 32'hbeca1e40} /* (24, 25, 1) {real, imag} */,
  {32'hc1982442, 32'h41270262} /* (24, 25, 0) {real, imag} */,
  {32'h4212f4bd, 32'hc19e7531} /* (24, 24, 31) {real, imag} */,
  {32'hc1f5980a, 32'h41783853} /* (24, 24, 30) {real, imag} */,
  {32'hc1748a33, 32'h4138e8c0} /* (24, 24, 29) {real, imag} */,
  {32'h419a0965, 32'h3f51fdf0} /* (24, 24, 28) {real, imag} */,
  {32'hc19fe7d8, 32'h40ac280d} /* (24, 24, 27) {real, imag} */,
  {32'h416f4b3e, 32'h417f90bd} /* (24, 24, 26) {real, imag} */,
  {32'h3fc15558, 32'h4159cfe2} /* (24, 24, 25) {real, imag} */,
  {32'hc13c57cc, 32'h4135a0d7} /* (24, 24, 24) {real, imag} */,
  {32'hc09808df, 32'hc0f62e16} /* (24, 24, 23) {real, imag} */,
  {32'hc044c118, 32'hc016ab60} /* (24, 24, 22) {real, imag} */,
  {32'h4053779f, 32'hc0b9c296} /* (24, 24, 21) {real, imag} */,
  {32'h412455d0, 32'h40e5f22e} /* (24, 24, 20) {real, imag} */,
  {32'h41034d81, 32'h3fed91fc} /* (24, 24, 19) {real, imag} */,
  {32'hc0220cf6, 32'hc1070902} /* (24, 24, 18) {real, imag} */,
  {32'h408fbca5, 32'hc097b9b1} /* (24, 24, 17) {real, imag} */,
  {32'hbeb01240, 32'h4125a4be} /* (24, 24, 16) {real, imag} */,
  {32'h4021087a, 32'hc01e3d86} /* (24, 24, 15) {real, imag} */,
  {32'h3fbdc57c, 32'hbf527c88} /* (24, 24, 14) {real, imag} */,
  {32'hc096cfd5, 32'hc096372a} /* (24, 24, 13) {real, imag} */,
  {32'h40ed8fe1, 32'hc149a799} /* (24, 24, 12) {real, imag} */,
  {32'h3f6a3504, 32'hc180678e} /* (24, 24, 11) {real, imag} */,
  {32'hbf143b35, 32'hc169c6b8} /* (24, 24, 10) {real, imag} */,
  {32'h3eaa2c7c, 32'hc13f9592} /* (24, 24, 9) {real, imag} */,
  {32'hc0612076, 32'h4166ae6b} /* (24, 24, 8) {real, imag} */,
  {32'h4193ccb2, 32'h41c23c84} /* (24, 24, 7) {real, imag} */,
  {32'h41140d74, 32'h4195afd0} /* (24, 24, 6) {real, imag} */,
  {32'hc17cf1e8, 32'hc146e3bc} /* (24, 24, 5) {real, imag} */,
  {32'h41494199, 32'h40b25374} /* (24, 24, 4) {real, imag} */,
  {32'h408c7710, 32'hc0748fed} /* (24, 24, 3) {real, imag} */,
  {32'hc1cf68e0, 32'h4111f9a2} /* (24, 24, 2) {real, imag} */,
  {32'h423ea0ad, 32'hc1b7e9ca} /* (24, 24, 1) {real, imag} */,
  {32'h403e2992, 32'hc12422e0} /* (24, 24, 0) {real, imag} */,
  {32'hc214bd6a, 32'hbf2fb200} /* (24, 23, 31) {real, imag} */,
  {32'h3c409d00, 32'hc056d3b0} /* (24, 23, 30) {real, imag} */,
  {32'h3d9a5fa0, 32'h419945a3} /* (24, 23, 29) {real, imag} */,
  {32'hc086f494, 32'h40bea6ca} /* (24, 23, 28) {real, imag} */,
  {32'h41181b3f, 32'hc0c78497} /* (24, 23, 27) {real, imag} */,
  {32'h4130991c, 32'hc044bb36} /* (24, 23, 26) {real, imag} */,
  {32'hc17a4be0, 32'hc0ab0c5c} /* (24, 23, 25) {real, imag} */,
  {32'hc0f9c855, 32'hc09f3391} /* (24, 23, 24) {real, imag} */,
  {32'hc0b03e2e, 32'h3f32c678} /* (24, 23, 23) {real, imag} */,
  {32'hc0b1215f, 32'hc172cc30} /* (24, 23, 22) {real, imag} */,
  {32'hc1229b35, 32'h3d1032c0} /* (24, 23, 21) {real, imag} */,
  {32'hc0508558, 32'h4092f3f2} /* (24, 23, 20) {real, imag} */,
  {32'hc0d5b216, 32'h402ae604} /* (24, 23, 19) {real, imag} */,
  {32'hc1315790, 32'hc0f17428} /* (24, 23, 18) {real, imag} */,
  {32'h4035411c, 32'h400f8e60} /* (24, 23, 17) {real, imag} */,
  {32'hc0123430, 32'h4189b418} /* (24, 23, 16) {real, imag} */,
  {32'hc066dbc3, 32'h40fc1b06} /* (24, 23, 15) {real, imag} */,
  {32'hbe7d56c0, 32'hc157e0d0} /* (24, 23, 14) {real, imag} */,
  {32'h412109a5, 32'hc1054a9e} /* (24, 23, 13) {real, imag} */,
  {32'h4048896c, 32'h408274a1} /* (24, 23, 12) {real, imag} */,
  {32'h3f60a6fc, 32'h4129ac20} /* (24, 23, 11) {real, imag} */,
  {32'h40ffd569, 32'h407ebdc9} /* (24, 23, 10) {real, imag} */,
  {32'hc18c6f1b, 32'h40fa9d9c} /* (24, 23, 9) {real, imag} */,
  {32'hc0023e49, 32'hc001099c} /* (24, 23, 8) {real, imag} */,
  {32'hbf9be4ca, 32'h3ffa5898} /* (24, 23, 7) {real, imag} */,
  {32'hc14c16d0, 32'hc05b5f3e} /* (24, 23, 6) {real, imag} */,
  {32'h419e404f, 32'hc1c2193e} /* (24, 23, 5) {real, imag} */,
  {32'h40fb9904, 32'hbf9bc604} /* (24, 23, 4) {real, imag} */,
  {32'h40f5eb89, 32'h415aff92} /* (24, 23, 3) {real, imag} */,
  {32'hc1366cbe, 32'hc19d4058} /* (24, 23, 2) {real, imag} */,
  {32'h406e9c08, 32'h412b8bb6} /* (24, 23, 1) {real, imag} */,
  {32'h3f3079d0, 32'h407e9448} /* (24, 23, 0) {real, imag} */,
  {32'hc112045a, 32'h419c347a} /* (24, 22, 31) {real, imag} */,
  {32'h41128ae3, 32'h40801d62} /* (24, 22, 30) {real, imag} */,
  {32'hc12a3755, 32'h3fc56079} /* (24, 22, 29) {real, imag} */,
  {32'h405e68da, 32'h40f0e17a} /* (24, 22, 28) {real, imag} */,
  {32'h3f4ed038, 32'hc12accb4} /* (24, 22, 27) {real, imag} */,
  {32'hc18d138d, 32'hc1057efa} /* (24, 22, 26) {real, imag} */,
  {32'h413add4a, 32'h40c4a7b2} /* (24, 22, 25) {real, imag} */,
  {32'h4143f3cc, 32'h41989c6b} /* (24, 22, 24) {real, imag} */,
  {32'hc07ddb80, 32'hc08b1a43} /* (24, 22, 23) {real, imag} */,
  {32'hc15ad57f, 32'h4080304a} /* (24, 22, 22) {real, imag} */,
  {32'h40978dae, 32'h412cc08a} /* (24, 22, 21) {real, imag} */,
  {32'hc1039f4d, 32'hc17a25c8} /* (24, 22, 20) {real, imag} */,
  {32'h410ea27a, 32'hc12b0729} /* (24, 22, 19) {real, imag} */,
  {32'h40bb774b, 32'h4170863e} /* (24, 22, 18) {real, imag} */,
  {32'hc0841bec, 32'hc1873266} /* (24, 22, 17) {real, imag} */,
  {32'hc019db70, 32'h4085d796} /* (24, 22, 16) {real, imag} */,
  {32'h409a63ba, 32'h4151e6ac} /* (24, 22, 15) {real, imag} */,
  {32'hc1b2ed17, 32'hbfbeea62} /* (24, 22, 14) {real, imag} */,
  {32'hc11a1510, 32'hbeea5550} /* (24, 22, 13) {real, imag} */,
  {32'hc124e66b, 32'hc10b6dd9} /* (24, 22, 12) {real, imag} */,
  {32'h41340d0a, 32'h41b6ec60} /* (24, 22, 11) {real, imag} */,
  {32'hbee8ca30, 32'hc09f082f} /* (24, 22, 10) {real, imag} */,
  {32'h41801bfe, 32'h4155eefe} /* (24, 22, 9) {real, imag} */,
  {32'hc1443eb8, 32'h40589574} /* (24, 22, 8) {real, imag} */,
  {32'h404d92a8, 32'h40b1b27f} /* (24, 22, 7) {real, imag} */,
  {32'hc07aa384, 32'h418583b0} /* (24, 22, 6) {real, imag} */,
  {32'h4096cd40, 32'hc11e5ace} /* (24, 22, 5) {real, imag} */,
  {32'hc1a4bd3b, 32'h410d3c4a} /* (24, 22, 4) {real, imag} */,
  {32'hc181d08a, 32'h40ceeb42} /* (24, 22, 3) {real, imag} */,
  {32'hbf604be0, 32'hc2182f52} /* (24, 22, 2) {real, imag} */,
  {32'hc1480bb6, 32'h41de4132} /* (24, 22, 1) {real, imag} */,
  {32'hc0d4c971, 32'h419ec9d3} /* (24, 22, 0) {real, imag} */,
  {32'h403858b0, 32'hc184702a} /* (24, 21, 31) {real, imag} */,
  {32'h41924f42, 32'h413c856a} /* (24, 21, 30) {real, imag} */,
  {32'h41d909b0, 32'hc00aa81f} /* (24, 21, 29) {real, imag} */,
  {32'hc010a0b0, 32'hbf31699c} /* (24, 21, 28) {real, imag} */,
  {32'hc0e9af4c, 32'h4091bbc0} /* (24, 21, 27) {real, imag} */,
  {32'hc1611a50, 32'h406e5f47} /* (24, 21, 26) {real, imag} */,
  {32'hbfa0e374, 32'hc1dfc24e} /* (24, 21, 25) {real, imag} */,
  {32'hc0d2021f, 32'h413ea240} /* (24, 21, 24) {real, imag} */,
  {32'h414f2bc4, 32'h41394251} /* (24, 21, 23) {real, imag} */,
  {32'hc0be1c88, 32'hc14bdd49} /* (24, 21, 22) {real, imag} */,
  {32'h4070e3f9, 32'hc025747e} /* (24, 21, 21) {real, imag} */,
  {32'h40b31fa0, 32'h41393168} /* (24, 21, 20) {real, imag} */,
  {32'hbd8c6f00, 32'h4172f065} /* (24, 21, 19) {real, imag} */,
  {32'h413d2ec0, 32'hc0145c36} /* (24, 21, 18) {real, imag} */,
  {32'hc1179c04, 32'hc13384e4} /* (24, 21, 17) {real, imag} */,
  {32'h4181bfa4, 32'hc0f75f83} /* (24, 21, 16) {real, imag} */,
  {32'hc15f703c, 32'h3f1c2f38} /* (24, 21, 15) {real, imag} */,
  {32'h403d91c3, 32'h3fc3caf6} /* (24, 21, 14) {real, imag} */,
  {32'hbfe92e8a, 32'h3ef23de0} /* (24, 21, 13) {real, imag} */,
  {32'h3efc5250, 32'hc0e1488e} /* (24, 21, 12) {real, imag} */,
  {32'h4091b849, 32'hc1c5bf44} /* (24, 21, 11) {real, imag} */,
  {32'h41152c3b, 32'h40a9a86a} /* (24, 21, 10) {real, imag} */,
  {32'hbffcd69b, 32'h40804dc2} /* (24, 21, 9) {real, imag} */,
  {32'h40bb12f7, 32'hc0fca492} /* (24, 21, 8) {real, imag} */,
  {32'h41958501, 32'h415470b2} /* (24, 21, 7) {real, imag} */,
  {32'hbfa8ba10, 32'h41082fd8} /* (24, 21, 6) {real, imag} */,
  {32'h40e54d04, 32'h3fc316dc} /* (24, 21, 5) {real, imag} */,
  {32'hbfb7d342, 32'hbfa48180} /* (24, 21, 4) {real, imag} */,
  {32'hc135840e, 32'hc04b3a98} /* (24, 21, 3) {real, imag} */,
  {32'hc0fe4dd2, 32'h41b0a015} /* (24, 21, 2) {real, imag} */,
  {32'h41cc71ec, 32'hc101c8a6} /* (24, 21, 1) {real, imag} */,
  {32'h40e01e50, 32'hc153983a} /* (24, 21, 0) {real, imag} */,
  {32'h3fba5a0c, 32'hc01db146} /* (24, 20, 31) {real, imag} */,
  {32'hc0c47a34, 32'h3f0b6c00} /* (24, 20, 30) {real, imag} */,
  {32'h3fbb02e1, 32'h40bfb4d6} /* (24, 20, 29) {real, imag} */,
  {32'hbdb24e80, 32'hc15422d8} /* (24, 20, 28) {real, imag} */,
  {32'h3fdaa0f8, 32'h40c704f2} /* (24, 20, 27) {real, imag} */,
  {32'h40c8a023, 32'hc0422a38} /* (24, 20, 26) {real, imag} */,
  {32'h4170bbe9, 32'hc1006952} /* (24, 20, 25) {real, imag} */,
  {32'hc08c6f30, 32'hc0cc0da4} /* (24, 20, 24) {real, imag} */,
  {32'hc10ac9ab, 32'h4140faec} /* (24, 20, 23) {real, imag} */,
  {32'hc19cc2d6, 32'hc00b2156} /* (24, 20, 22) {real, imag} */,
  {32'hc0d47caf, 32'h418ace78} /* (24, 20, 21) {real, imag} */,
  {32'hc06876ca, 32'h40a6e40a} /* (24, 20, 20) {real, imag} */,
  {32'hc009b3e4, 32'hc07b5132} /* (24, 20, 19) {real, imag} */,
  {32'h3fc9a7b6, 32'h40ac6563} /* (24, 20, 18) {real, imag} */,
  {32'h3d235d80, 32'h415ab6dc} /* (24, 20, 17) {real, imag} */,
  {32'h3ffa75b4, 32'hbfe8f5df} /* (24, 20, 16) {real, imag} */,
  {32'h40dc1436, 32'h3f9f7b66} /* (24, 20, 15) {real, imag} */,
  {32'hc09e1ba4, 32'h414c7dd2} /* (24, 20, 14) {real, imag} */,
  {32'h40d75c7d, 32'hc00908de} /* (24, 20, 13) {real, imag} */,
  {32'h41c76918, 32'h40a8039c} /* (24, 20, 12) {real, imag} */,
  {32'hc0ced349, 32'hc028e81e} /* (24, 20, 11) {real, imag} */,
  {32'h3fdffd58, 32'hc15f1668} /* (24, 20, 10) {real, imag} */,
  {32'hc124f667, 32'hbf123bc8} /* (24, 20, 9) {real, imag} */,
  {32'hc14681c4, 32'hc1922c55} /* (24, 20, 8) {real, imag} */,
  {32'hbd8d5e00, 32'h41166a26} /* (24, 20, 7) {real, imag} */,
  {32'h3eaa48b0, 32'hc15fa9d0} /* (24, 20, 6) {real, imag} */,
  {32'hc14780ae, 32'h41ab1b8c} /* (24, 20, 5) {real, imag} */,
  {32'h41264843, 32'h411d08ec} /* (24, 20, 4) {real, imag} */,
  {32'h3f9deb16, 32'h40406e2c} /* (24, 20, 3) {real, imag} */,
  {32'h407a99e0, 32'hc0039e31} /* (24, 20, 2) {real, imag} */,
  {32'hc13fa884, 32'hc135012d} /* (24, 20, 1) {real, imag} */,
  {32'h419b8a8c, 32'hc0f3ea75} /* (24, 20, 0) {real, imag} */,
  {32'hc01b6f24, 32'hc18d3268} /* (24, 19, 31) {real, imag} */,
  {32'h40d499b4, 32'h415eda4a} /* (24, 19, 30) {real, imag} */,
  {32'h40a2bde8, 32'h3f897c98} /* (24, 19, 29) {real, imag} */,
  {32'hc17a2577, 32'h41938afa} /* (24, 19, 28) {real, imag} */,
  {32'h41783d75, 32'h3f24dd90} /* (24, 19, 27) {real, imag} */,
  {32'h414097b6, 32'hc0ad6860} /* (24, 19, 26) {real, imag} */,
  {32'h41112ef1, 32'hc051b588} /* (24, 19, 25) {real, imag} */,
  {32'h40ebb7d3, 32'hc07559b2} /* (24, 19, 24) {real, imag} */,
  {32'h4076a91a, 32'hc12295bb} /* (24, 19, 23) {real, imag} */,
  {32'h409f7ae2, 32'h409a3e78} /* (24, 19, 22) {real, imag} */,
  {32'h40516af3, 32'h40f299a0} /* (24, 19, 21) {real, imag} */,
  {32'h3fafb2de, 32'hc06d7b4b} /* (24, 19, 20) {real, imag} */,
  {32'hc0c61f6b, 32'hbf41e5c0} /* (24, 19, 19) {real, imag} */,
  {32'hc15a21b4, 32'h40f5dd28} /* (24, 19, 18) {real, imag} */,
  {32'hc1364b66, 32'hbfb4bc6c} /* (24, 19, 17) {real, imag} */,
  {32'hc06b5159, 32'hc0eb1194} /* (24, 19, 16) {real, imag} */,
  {32'h411a3447, 32'h41200188} /* (24, 19, 15) {real, imag} */,
  {32'hc05c5277, 32'hbe32f610} /* (24, 19, 14) {real, imag} */,
  {32'h4153f967, 32'hc1168564} /* (24, 19, 13) {real, imag} */,
  {32'hc031b2ec, 32'h4184923c} /* (24, 19, 12) {real, imag} */,
  {32'h40f2e8d2, 32'h40c90523} /* (24, 19, 11) {real, imag} */,
  {32'hc11bed9a, 32'hc13b4c50} /* (24, 19, 10) {real, imag} */,
  {32'hc14973f2, 32'h40cc1806} /* (24, 19, 9) {real, imag} */,
  {32'hc05beb4e, 32'h3feaa68e} /* (24, 19, 8) {real, imag} */,
  {32'hc0b46cef, 32'hc184a811} /* (24, 19, 7) {real, imag} */,
  {32'hc0a9392e, 32'hc15b2eea} /* (24, 19, 6) {real, imag} */,
  {32'hc09dda8e, 32'hc0e72e82} /* (24, 19, 5) {real, imag} */,
  {32'hc11db17d, 32'hc0d94316} /* (24, 19, 4) {real, imag} */,
  {32'h412b4f9f, 32'hc002339c} /* (24, 19, 3) {real, imag} */,
  {32'hc0c41cc4, 32'h412a2aca} /* (24, 19, 2) {real, imag} */,
  {32'hc1895488, 32'hc0c05505} /* (24, 19, 1) {real, imag} */,
  {32'hbfd8b280, 32'h40c8c809} /* (24, 19, 0) {real, imag} */,
  {32'hc01fd9de, 32'hc1183f5e} /* (24, 18, 31) {real, imag} */,
  {32'hc0f7994a, 32'h413bb441} /* (24, 18, 30) {real, imag} */,
  {32'h403159f1, 32'hc006dbae} /* (24, 18, 29) {real, imag} */,
  {32'h3d972f50, 32'hbf1a0cdc} /* (24, 18, 28) {real, imag} */,
  {32'hc120df2b, 32'h4155225e} /* (24, 18, 27) {real, imag} */,
  {32'h40c834e6, 32'h3f90435c} /* (24, 18, 26) {real, imag} */,
  {32'hc186390e, 32'hc00c8741} /* (24, 18, 25) {real, imag} */,
  {32'hc056c781, 32'h4129e3dc} /* (24, 18, 24) {real, imag} */,
  {32'h414095e9, 32'hc13a99ef} /* (24, 18, 23) {real, imag} */,
  {32'hc14afcfd, 32'hc0f8f612} /* (24, 18, 22) {real, imag} */,
  {32'h41214010, 32'hc0d18f34} /* (24, 18, 21) {real, imag} */,
  {32'hc02dbc2f, 32'hbf4881a8} /* (24, 18, 20) {real, imag} */,
  {32'hc09f94f3, 32'hbfacb50c} /* (24, 18, 19) {real, imag} */,
  {32'h3f3497b0, 32'h3f93ca24} /* (24, 18, 18) {real, imag} */,
  {32'hc01486d8, 32'hbfa95fc4} /* (24, 18, 17) {real, imag} */,
  {32'h41243521, 32'h405527f4} /* (24, 18, 16) {real, imag} */,
  {32'hc1063afc, 32'hc0792380} /* (24, 18, 15) {real, imag} */,
  {32'hc0f0f6d8, 32'hc1478d2c} /* (24, 18, 14) {real, imag} */,
  {32'h40c2a475, 32'h40beeb0a} /* (24, 18, 13) {real, imag} */,
  {32'hc0aa265c, 32'h40838755} /* (24, 18, 12) {real, imag} */,
  {32'hc18661a3, 32'h403c3f86} /* (24, 18, 11) {real, imag} */,
  {32'h40b69508, 32'h3fdda50c} /* (24, 18, 10) {real, imag} */,
  {32'h4145852e, 32'hbf9116f8} /* (24, 18, 9) {real, imag} */,
  {32'hc13a5d0a, 32'hc097aa42} /* (24, 18, 8) {real, imag} */,
  {32'h400dc1ee, 32'h3c8531c0} /* (24, 18, 7) {real, imag} */,
  {32'hc0a332c8, 32'hc15106bc} /* (24, 18, 6) {real, imag} */,
  {32'h4036262e, 32'h3fd97088} /* (24, 18, 5) {real, imag} */,
  {32'h4188c6b2, 32'h414e6208} /* (24, 18, 4) {real, imag} */,
  {32'h41621400, 32'hbf913834} /* (24, 18, 3) {real, imag} */,
  {32'hc1a0a493, 32'h40aabf5c} /* (24, 18, 2) {real, imag} */,
  {32'h40bb989f, 32'hc15c8a74} /* (24, 18, 1) {real, imag} */,
  {32'h410356ea, 32'hc07d10e6} /* (24, 18, 0) {real, imag} */,
  {32'hbdaa5e90, 32'hbfa3c850} /* (24, 17, 31) {real, imag} */,
  {32'hc0ac079f, 32'hc0cfe5fd} /* (24, 17, 30) {real, imag} */,
  {32'hc1175e34, 32'hc0bec5bc} /* (24, 17, 29) {real, imag} */,
  {32'h4107c13c, 32'h41028813} /* (24, 17, 28) {real, imag} */,
  {32'h3d2a4100, 32'hbebca7a0} /* (24, 17, 27) {real, imag} */,
  {32'hbf335200, 32'h410b3ba2} /* (24, 17, 26) {real, imag} */,
  {32'hc0b0e526, 32'hc14b15b2} /* (24, 17, 25) {real, imag} */,
  {32'h40d50642, 32'hbfa77960} /* (24, 17, 24) {real, imag} */,
  {32'hc189185a, 32'hc08d4442} /* (24, 17, 23) {real, imag} */,
  {32'hc1036360, 32'h4113a241} /* (24, 17, 22) {real, imag} */,
  {32'h413afad6, 32'hc1846e95} /* (24, 17, 21) {real, imag} */,
  {32'hbf00a88c, 32'h402edbe0} /* (24, 17, 20) {real, imag} */,
  {32'h40d850ce, 32'hbe5e4040} /* (24, 17, 19) {real, imag} */,
  {32'h411200d2, 32'h408dff4b} /* (24, 17, 18) {real, imag} */,
  {32'hc0317624, 32'hc06a5802} /* (24, 17, 17) {real, imag} */,
  {32'hbf707d60, 32'h400e501e} /* (24, 17, 16) {real, imag} */,
  {32'hbfb760b8, 32'h3f5c0a40} /* (24, 17, 15) {real, imag} */,
  {32'hc088a77a, 32'h409425b8} /* (24, 17, 14) {real, imag} */,
  {32'h401eb17f, 32'hc08cd7f0} /* (24, 17, 13) {real, imag} */,
  {32'h3ee3eaa8, 32'hc02c11ad} /* (24, 17, 12) {real, imag} */,
  {32'hc0035fc2, 32'hc0d66a77} /* (24, 17, 11) {real, imag} */,
  {32'hbf0275d0, 32'h40c3c394} /* (24, 17, 10) {real, imag} */,
  {32'h4149335f, 32'h40d70928} /* (24, 17, 9) {real, imag} */,
  {32'h409dee31, 32'h40432bba} /* (24, 17, 8) {real, imag} */,
  {32'h3fbf76d4, 32'hc1948829} /* (24, 17, 7) {real, imag} */,
  {32'h4096b012, 32'hc1243290} /* (24, 17, 6) {real, imag} */,
  {32'hbe9a3fa4, 32'h401df903} /* (24, 17, 5) {real, imag} */,
  {32'hc099ee8c, 32'h3fbc5b47} /* (24, 17, 4) {real, imag} */,
  {32'hc1201314, 32'h4099370c} /* (24, 17, 3) {real, imag} */,
  {32'h4101e38f, 32'hbfbfed4c} /* (24, 17, 2) {real, imag} */,
  {32'hbf8315e7, 32'h3f876098} /* (24, 17, 1) {real, imag} */,
  {32'hc01ac802, 32'h40e1093a} /* (24, 17, 0) {real, imag} */,
  {32'h40d8811a, 32'hbdcf2c60} /* (24, 16, 31) {real, imag} */,
  {32'h407460aa, 32'hc0143ba8} /* (24, 16, 30) {real, imag} */,
  {32'hc0b0b48b, 32'h40532096} /* (24, 16, 29) {real, imag} */,
  {32'h3fc2c97c, 32'h3fba561a} /* (24, 16, 28) {real, imag} */,
  {32'hc0e22ab7, 32'hc0ebadab} /* (24, 16, 27) {real, imag} */,
  {32'h40516367, 32'hc1457bd1} /* (24, 16, 26) {real, imag} */,
  {32'h411c54a8, 32'h408a0896} /* (24, 16, 25) {real, imag} */,
  {32'h40e310f4, 32'h41355262} /* (24, 16, 24) {real, imag} */,
  {32'h3f7d5e40, 32'h41649adc} /* (24, 16, 23) {real, imag} */,
  {32'hc14cf9fb, 32'hc09ce1fe} /* (24, 16, 22) {real, imag} */,
  {32'hbcb1cd00, 32'h40832f6d} /* (24, 16, 21) {real, imag} */,
  {32'h4081ce9a, 32'hc0998052} /* (24, 16, 20) {real, imag} */,
  {32'h405642a4, 32'hc04c8054} /* (24, 16, 19) {real, imag} */,
  {32'hc047aa54, 32'hc0882b0f} /* (24, 16, 18) {real, imag} */,
  {32'hc1007c81, 32'hc0a383f8} /* (24, 16, 17) {real, imag} */,
  {32'hc0aa69bc, 32'h00000000} /* (24, 16, 16) {real, imag} */,
  {32'hc1007c81, 32'h40a383f8} /* (24, 16, 15) {real, imag} */,
  {32'hc047aa54, 32'h40882b0f} /* (24, 16, 14) {real, imag} */,
  {32'h405642a4, 32'h404c8054} /* (24, 16, 13) {real, imag} */,
  {32'h4081ce9a, 32'h40998052} /* (24, 16, 12) {real, imag} */,
  {32'hbcb1cd00, 32'hc0832f6d} /* (24, 16, 11) {real, imag} */,
  {32'hc14cf9fb, 32'h409ce1fe} /* (24, 16, 10) {real, imag} */,
  {32'h3f7d5e40, 32'hc1649adc} /* (24, 16, 9) {real, imag} */,
  {32'h40e310f4, 32'hc1355262} /* (24, 16, 8) {real, imag} */,
  {32'h411c54a8, 32'hc08a0896} /* (24, 16, 7) {real, imag} */,
  {32'h40516367, 32'h41457bd1} /* (24, 16, 6) {real, imag} */,
  {32'hc0e22ab7, 32'h40ebadab} /* (24, 16, 5) {real, imag} */,
  {32'h3fc2c97c, 32'hbfba561a} /* (24, 16, 4) {real, imag} */,
  {32'hc0b0b48b, 32'hc0532096} /* (24, 16, 3) {real, imag} */,
  {32'h407460aa, 32'h40143ba8} /* (24, 16, 2) {real, imag} */,
  {32'h40d8811a, 32'h3dcf2c60} /* (24, 16, 1) {real, imag} */,
  {32'hc02b64c0, 32'h00000000} /* (24, 16, 0) {real, imag} */,
  {32'hbf8315e7, 32'hbf876098} /* (24, 15, 31) {real, imag} */,
  {32'h4101e38f, 32'h3fbfed4c} /* (24, 15, 30) {real, imag} */,
  {32'hc1201314, 32'hc099370c} /* (24, 15, 29) {real, imag} */,
  {32'hc099ee8c, 32'hbfbc5b47} /* (24, 15, 28) {real, imag} */,
  {32'hbe9a3fa4, 32'hc01df903} /* (24, 15, 27) {real, imag} */,
  {32'h4096b012, 32'h41243290} /* (24, 15, 26) {real, imag} */,
  {32'h3fbf76d4, 32'h41948829} /* (24, 15, 25) {real, imag} */,
  {32'h409dee31, 32'hc0432bba} /* (24, 15, 24) {real, imag} */,
  {32'h4149335f, 32'hc0d70928} /* (24, 15, 23) {real, imag} */,
  {32'hbf0275d0, 32'hc0c3c394} /* (24, 15, 22) {real, imag} */,
  {32'hc0035fc2, 32'h40d66a77} /* (24, 15, 21) {real, imag} */,
  {32'h3ee3eaa8, 32'h402c11ad} /* (24, 15, 20) {real, imag} */,
  {32'h401eb17f, 32'h408cd7f0} /* (24, 15, 19) {real, imag} */,
  {32'hc088a77a, 32'hc09425b8} /* (24, 15, 18) {real, imag} */,
  {32'hbfb760b8, 32'hbf5c0a40} /* (24, 15, 17) {real, imag} */,
  {32'hbf707d60, 32'hc00e501e} /* (24, 15, 16) {real, imag} */,
  {32'hc0317624, 32'h406a5802} /* (24, 15, 15) {real, imag} */,
  {32'h411200d2, 32'hc08dff4b} /* (24, 15, 14) {real, imag} */,
  {32'h40d850ce, 32'h3e5e4040} /* (24, 15, 13) {real, imag} */,
  {32'hbf00a88c, 32'hc02edbe0} /* (24, 15, 12) {real, imag} */,
  {32'h413afad6, 32'h41846e95} /* (24, 15, 11) {real, imag} */,
  {32'hc1036360, 32'hc113a241} /* (24, 15, 10) {real, imag} */,
  {32'hc189185a, 32'h408d4442} /* (24, 15, 9) {real, imag} */,
  {32'h40d50642, 32'h3fa77960} /* (24, 15, 8) {real, imag} */,
  {32'hc0b0e526, 32'h414b15b2} /* (24, 15, 7) {real, imag} */,
  {32'hbf335200, 32'hc10b3ba2} /* (24, 15, 6) {real, imag} */,
  {32'h3d2a4100, 32'h3ebca7a0} /* (24, 15, 5) {real, imag} */,
  {32'h4107c13c, 32'hc1028813} /* (24, 15, 4) {real, imag} */,
  {32'hc1175e34, 32'h40bec5bc} /* (24, 15, 3) {real, imag} */,
  {32'hc0ac079f, 32'h40cfe5fd} /* (24, 15, 2) {real, imag} */,
  {32'hbdaa5e90, 32'h3fa3c850} /* (24, 15, 1) {real, imag} */,
  {32'hc01ac802, 32'hc0e1093a} /* (24, 15, 0) {real, imag} */,
  {32'h40bb989f, 32'h415c8a74} /* (24, 14, 31) {real, imag} */,
  {32'hc1a0a493, 32'hc0aabf5c} /* (24, 14, 30) {real, imag} */,
  {32'h41621400, 32'h3f913834} /* (24, 14, 29) {real, imag} */,
  {32'h4188c6b2, 32'hc14e6208} /* (24, 14, 28) {real, imag} */,
  {32'h4036262e, 32'hbfd97088} /* (24, 14, 27) {real, imag} */,
  {32'hc0a332c8, 32'h415106bc} /* (24, 14, 26) {real, imag} */,
  {32'h400dc1ee, 32'hbc8531c0} /* (24, 14, 25) {real, imag} */,
  {32'hc13a5d0a, 32'h4097aa42} /* (24, 14, 24) {real, imag} */,
  {32'h4145852e, 32'h3f9116f8} /* (24, 14, 23) {real, imag} */,
  {32'h40b69508, 32'hbfdda50c} /* (24, 14, 22) {real, imag} */,
  {32'hc18661a3, 32'hc03c3f86} /* (24, 14, 21) {real, imag} */,
  {32'hc0aa265c, 32'hc0838755} /* (24, 14, 20) {real, imag} */,
  {32'h40c2a475, 32'hc0beeb0a} /* (24, 14, 19) {real, imag} */,
  {32'hc0f0f6d8, 32'h41478d2c} /* (24, 14, 18) {real, imag} */,
  {32'hc1063afc, 32'h40792380} /* (24, 14, 17) {real, imag} */,
  {32'h41243521, 32'hc05527f4} /* (24, 14, 16) {real, imag} */,
  {32'hc01486d8, 32'h3fa95fc4} /* (24, 14, 15) {real, imag} */,
  {32'h3f3497b0, 32'hbf93ca24} /* (24, 14, 14) {real, imag} */,
  {32'hc09f94f3, 32'h3facb50c} /* (24, 14, 13) {real, imag} */,
  {32'hc02dbc2f, 32'h3f4881a8} /* (24, 14, 12) {real, imag} */,
  {32'h41214010, 32'h40d18f34} /* (24, 14, 11) {real, imag} */,
  {32'hc14afcfd, 32'h40f8f612} /* (24, 14, 10) {real, imag} */,
  {32'h414095e9, 32'h413a99ef} /* (24, 14, 9) {real, imag} */,
  {32'hc056c781, 32'hc129e3dc} /* (24, 14, 8) {real, imag} */,
  {32'hc186390e, 32'h400c8741} /* (24, 14, 7) {real, imag} */,
  {32'h40c834e6, 32'hbf90435c} /* (24, 14, 6) {real, imag} */,
  {32'hc120df2b, 32'hc155225e} /* (24, 14, 5) {real, imag} */,
  {32'h3d972f50, 32'h3f1a0cdc} /* (24, 14, 4) {real, imag} */,
  {32'h403159f1, 32'h4006dbae} /* (24, 14, 3) {real, imag} */,
  {32'hc0f7994a, 32'hc13bb441} /* (24, 14, 2) {real, imag} */,
  {32'hc01fd9de, 32'h41183f5e} /* (24, 14, 1) {real, imag} */,
  {32'h410356ea, 32'h407d10e6} /* (24, 14, 0) {real, imag} */,
  {32'hc1895488, 32'h40c05505} /* (24, 13, 31) {real, imag} */,
  {32'hc0c41cc4, 32'hc12a2aca} /* (24, 13, 30) {real, imag} */,
  {32'h412b4f9f, 32'h4002339c} /* (24, 13, 29) {real, imag} */,
  {32'hc11db17d, 32'h40d94316} /* (24, 13, 28) {real, imag} */,
  {32'hc09dda8e, 32'h40e72e82} /* (24, 13, 27) {real, imag} */,
  {32'hc0a9392e, 32'h415b2eea} /* (24, 13, 26) {real, imag} */,
  {32'hc0b46cef, 32'h4184a811} /* (24, 13, 25) {real, imag} */,
  {32'hc05beb4e, 32'hbfeaa68e} /* (24, 13, 24) {real, imag} */,
  {32'hc14973f2, 32'hc0cc1806} /* (24, 13, 23) {real, imag} */,
  {32'hc11bed9a, 32'h413b4c50} /* (24, 13, 22) {real, imag} */,
  {32'h40f2e8d2, 32'hc0c90523} /* (24, 13, 21) {real, imag} */,
  {32'hc031b2ec, 32'hc184923c} /* (24, 13, 20) {real, imag} */,
  {32'h4153f967, 32'h41168564} /* (24, 13, 19) {real, imag} */,
  {32'hc05c5277, 32'h3e32f610} /* (24, 13, 18) {real, imag} */,
  {32'h411a3447, 32'hc1200188} /* (24, 13, 17) {real, imag} */,
  {32'hc06b5159, 32'h40eb1194} /* (24, 13, 16) {real, imag} */,
  {32'hc1364b66, 32'h3fb4bc6c} /* (24, 13, 15) {real, imag} */,
  {32'hc15a21b4, 32'hc0f5dd28} /* (24, 13, 14) {real, imag} */,
  {32'hc0c61f6b, 32'h3f41e5c0} /* (24, 13, 13) {real, imag} */,
  {32'h3fafb2de, 32'h406d7b4b} /* (24, 13, 12) {real, imag} */,
  {32'h40516af3, 32'hc0f299a0} /* (24, 13, 11) {real, imag} */,
  {32'h409f7ae2, 32'hc09a3e78} /* (24, 13, 10) {real, imag} */,
  {32'h4076a91a, 32'h412295bb} /* (24, 13, 9) {real, imag} */,
  {32'h40ebb7d3, 32'h407559b2} /* (24, 13, 8) {real, imag} */,
  {32'h41112ef1, 32'h4051b588} /* (24, 13, 7) {real, imag} */,
  {32'h414097b6, 32'h40ad6860} /* (24, 13, 6) {real, imag} */,
  {32'h41783d75, 32'hbf24dd90} /* (24, 13, 5) {real, imag} */,
  {32'hc17a2577, 32'hc1938afa} /* (24, 13, 4) {real, imag} */,
  {32'h40a2bde8, 32'hbf897c98} /* (24, 13, 3) {real, imag} */,
  {32'h40d499b4, 32'hc15eda4a} /* (24, 13, 2) {real, imag} */,
  {32'hc01b6f24, 32'h418d3268} /* (24, 13, 1) {real, imag} */,
  {32'hbfd8b280, 32'hc0c8c809} /* (24, 13, 0) {real, imag} */,
  {32'hc13fa884, 32'h4135012d} /* (24, 12, 31) {real, imag} */,
  {32'h407a99e0, 32'h40039e31} /* (24, 12, 30) {real, imag} */,
  {32'h3f9deb16, 32'hc0406e2c} /* (24, 12, 29) {real, imag} */,
  {32'h41264843, 32'hc11d08ec} /* (24, 12, 28) {real, imag} */,
  {32'hc14780ae, 32'hc1ab1b8c} /* (24, 12, 27) {real, imag} */,
  {32'h3eaa48b0, 32'h415fa9d0} /* (24, 12, 26) {real, imag} */,
  {32'hbd8d5e00, 32'hc1166a26} /* (24, 12, 25) {real, imag} */,
  {32'hc14681c4, 32'h41922c55} /* (24, 12, 24) {real, imag} */,
  {32'hc124f667, 32'h3f123bc8} /* (24, 12, 23) {real, imag} */,
  {32'h3fdffd58, 32'h415f1668} /* (24, 12, 22) {real, imag} */,
  {32'hc0ced349, 32'h4028e81e} /* (24, 12, 21) {real, imag} */,
  {32'h41c76918, 32'hc0a8039c} /* (24, 12, 20) {real, imag} */,
  {32'h40d75c7d, 32'h400908de} /* (24, 12, 19) {real, imag} */,
  {32'hc09e1ba4, 32'hc14c7dd2} /* (24, 12, 18) {real, imag} */,
  {32'h40dc1436, 32'hbf9f7b66} /* (24, 12, 17) {real, imag} */,
  {32'h3ffa75b4, 32'h3fe8f5df} /* (24, 12, 16) {real, imag} */,
  {32'h3d235d80, 32'hc15ab6dc} /* (24, 12, 15) {real, imag} */,
  {32'h3fc9a7b6, 32'hc0ac6563} /* (24, 12, 14) {real, imag} */,
  {32'hc009b3e4, 32'h407b5132} /* (24, 12, 13) {real, imag} */,
  {32'hc06876ca, 32'hc0a6e40a} /* (24, 12, 12) {real, imag} */,
  {32'hc0d47caf, 32'hc18ace78} /* (24, 12, 11) {real, imag} */,
  {32'hc19cc2d6, 32'h400b2156} /* (24, 12, 10) {real, imag} */,
  {32'hc10ac9ab, 32'hc140faec} /* (24, 12, 9) {real, imag} */,
  {32'hc08c6f30, 32'h40cc0da4} /* (24, 12, 8) {real, imag} */,
  {32'h4170bbe9, 32'h41006952} /* (24, 12, 7) {real, imag} */,
  {32'h40c8a023, 32'h40422a38} /* (24, 12, 6) {real, imag} */,
  {32'h3fdaa0f8, 32'hc0c704f2} /* (24, 12, 5) {real, imag} */,
  {32'hbdb24e80, 32'h415422d8} /* (24, 12, 4) {real, imag} */,
  {32'h3fbb02e1, 32'hc0bfb4d6} /* (24, 12, 3) {real, imag} */,
  {32'hc0c47a34, 32'hbf0b6c00} /* (24, 12, 2) {real, imag} */,
  {32'h3fba5a0c, 32'h401db146} /* (24, 12, 1) {real, imag} */,
  {32'h419b8a8c, 32'h40f3ea75} /* (24, 12, 0) {real, imag} */,
  {32'h41cc71ec, 32'h4101c8a6} /* (24, 11, 31) {real, imag} */,
  {32'hc0fe4dd2, 32'hc1b0a015} /* (24, 11, 30) {real, imag} */,
  {32'hc135840e, 32'h404b3a98} /* (24, 11, 29) {real, imag} */,
  {32'hbfb7d342, 32'h3fa48180} /* (24, 11, 28) {real, imag} */,
  {32'h40e54d04, 32'hbfc316dc} /* (24, 11, 27) {real, imag} */,
  {32'hbfa8ba10, 32'hc1082fd8} /* (24, 11, 26) {real, imag} */,
  {32'h41958501, 32'hc15470b2} /* (24, 11, 25) {real, imag} */,
  {32'h40bb12f7, 32'h40fca492} /* (24, 11, 24) {real, imag} */,
  {32'hbffcd69b, 32'hc0804dc2} /* (24, 11, 23) {real, imag} */,
  {32'h41152c3b, 32'hc0a9a86a} /* (24, 11, 22) {real, imag} */,
  {32'h4091b849, 32'h41c5bf44} /* (24, 11, 21) {real, imag} */,
  {32'h3efc5250, 32'h40e1488e} /* (24, 11, 20) {real, imag} */,
  {32'hbfe92e8a, 32'hbef23de0} /* (24, 11, 19) {real, imag} */,
  {32'h403d91c3, 32'hbfc3caf6} /* (24, 11, 18) {real, imag} */,
  {32'hc15f703c, 32'hbf1c2f38} /* (24, 11, 17) {real, imag} */,
  {32'h4181bfa4, 32'h40f75f83} /* (24, 11, 16) {real, imag} */,
  {32'hc1179c04, 32'h413384e4} /* (24, 11, 15) {real, imag} */,
  {32'h413d2ec0, 32'h40145c36} /* (24, 11, 14) {real, imag} */,
  {32'hbd8c6f00, 32'hc172f065} /* (24, 11, 13) {real, imag} */,
  {32'h40b31fa0, 32'hc1393168} /* (24, 11, 12) {real, imag} */,
  {32'h4070e3f9, 32'h4025747e} /* (24, 11, 11) {real, imag} */,
  {32'hc0be1c88, 32'h414bdd49} /* (24, 11, 10) {real, imag} */,
  {32'h414f2bc4, 32'hc1394251} /* (24, 11, 9) {real, imag} */,
  {32'hc0d2021f, 32'hc13ea240} /* (24, 11, 8) {real, imag} */,
  {32'hbfa0e374, 32'h41dfc24e} /* (24, 11, 7) {real, imag} */,
  {32'hc1611a50, 32'hc06e5f47} /* (24, 11, 6) {real, imag} */,
  {32'hc0e9af4c, 32'hc091bbc0} /* (24, 11, 5) {real, imag} */,
  {32'hc010a0b0, 32'h3f31699c} /* (24, 11, 4) {real, imag} */,
  {32'h41d909b0, 32'h400aa81f} /* (24, 11, 3) {real, imag} */,
  {32'h41924f42, 32'hc13c856a} /* (24, 11, 2) {real, imag} */,
  {32'h403858b0, 32'h4184702a} /* (24, 11, 1) {real, imag} */,
  {32'h40e01e50, 32'h4153983a} /* (24, 11, 0) {real, imag} */,
  {32'hc1480bb6, 32'hc1de4132} /* (24, 10, 31) {real, imag} */,
  {32'hbf604be0, 32'h42182f52} /* (24, 10, 30) {real, imag} */,
  {32'hc181d08a, 32'hc0ceeb42} /* (24, 10, 29) {real, imag} */,
  {32'hc1a4bd3b, 32'hc10d3c4a} /* (24, 10, 28) {real, imag} */,
  {32'h4096cd40, 32'h411e5ace} /* (24, 10, 27) {real, imag} */,
  {32'hc07aa384, 32'hc18583b0} /* (24, 10, 26) {real, imag} */,
  {32'h404d92a8, 32'hc0b1b27f} /* (24, 10, 25) {real, imag} */,
  {32'hc1443eb8, 32'hc0589574} /* (24, 10, 24) {real, imag} */,
  {32'h41801bfe, 32'hc155eefe} /* (24, 10, 23) {real, imag} */,
  {32'hbee8ca30, 32'h409f082f} /* (24, 10, 22) {real, imag} */,
  {32'h41340d0a, 32'hc1b6ec60} /* (24, 10, 21) {real, imag} */,
  {32'hc124e66b, 32'h410b6dd9} /* (24, 10, 20) {real, imag} */,
  {32'hc11a1510, 32'h3eea5550} /* (24, 10, 19) {real, imag} */,
  {32'hc1b2ed17, 32'h3fbeea62} /* (24, 10, 18) {real, imag} */,
  {32'h409a63ba, 32'hc151e6ac} /* (24, 10, 17) {real, imag} */,
  {32'hc019db70, 32'hc085d796} /* (24, 10, 16) {real, imag} */,
  {32'hc0841bec, 32'h41873266} /* (24, 10, 15) {real, imag} */,
  {32'h40bb774b, 32'hc170863e} /* (24, 10, 14) {real, imag} */,
  {32'h410ea27a, 32'h412b0729} /* (24, 10, 13) {real, imag} */,
  {32'hc1039f4d, 32'h417a25c8} /* (24, 10, 12) {real, imag} */,
  {32'h40978dae, 32'hc12cc08a} /* (24, 10, 11) {real, imag} */,
  {32'hc15ad57f, 32'hc080304a} /* (24, 10, 10) {real, imag} */,
  {32'hc07ddb80, 32'h408b1a43} /* (24, 10, 9) {real, imag} */,
  {32'h4143f3cc, 32'hc1989c6b} /* (24, 10, 8) {real, imag} */,
  {32'h413add4a, 32'hc0c4a7b2} /* (24, 10, 7) {real, imag} */,
  {32'hc18d138d, 32'h41057efa} /* (24, 10, 6) {real, imag} */,
  {32'h3f4ed038, 32'h412accb4} /* (24, 10, 5) {real, imag} */,
  {32'h405e68da, 32'hc0f0e17a} /* (24, 10, 4) {real, imag} */,
  {32'hc12a3755, 32'hbfc56079} /* (24, 10, 3) {real, imag} */,
  {32'h41128ae3, 32'hc0801d62} /* (24, 10, 2) {real, imag} */,
  {32'hc112045a, 32'hc19c347a} /* (24, 10, 1) {real, imag} */,
  {32'hc0d4c971, 32'hc19ec9d3} /* (24, 10, 0) {real, imag} */,
  {32'h406e9c08, 32'hc12b8bb6} /* (24, 9, 31) {real, imag} */,
  {32'hc1366cbe, 32'h419d4058} /* (24, 9, 30) {real, imag} */,
  {32'h40f5eb89, 32'hc15aff92} /* (24, 9, 29) {real, imag} */,
  {32'h40fb9904, 32'h3f9bc604} /* (24, 9, 28) {real, imag} */,
  {32'h419e404f, 32'h41c2193e} /* (24, 9, 27) {real, imag} */,
  {32'hc14c16d0, 32'h405b5f3e} /* (24, 9, 26) {real, imag} */,
  {32'hbf9be4ca, 32'hbffa5898} /* (24, 9, 25) {real, imag} */,
  {32'hc0023e49, 32'h4001099c} /* (24, 9, 24) {real, imag} */,
  {32'hc18c6f1b, 32'hc0fa9d9c} /* (24, 9, 23) {real, imag} */,
  {32'h40ffd569, 32'hc07ebdc9} /* (24, 9, 22) {real, imag} */,
  {32'h3f60a6fc, 32'hc129ac20} /* (24, 9, 21) {real, imag} */,
  {32'h4048896c, 32'hc08274a1} /* (24, 9, 20) {real, imag} */,
  {32'h412109a5, 32'h41054a9e} /* (24, 9, 19) {real, imag} */,
  {32'hbe7d56c0, 32'h4157e0d0} /* (24, 9, 18) {real, imag} */,
  {32'hc066dbc3, 32'hc0fc1b06} /* (24, 9, 17) {real, imag} */,
  {32'hc0123430, 32'hc189b418} /* (24, 9, 16) {real, imag} */,
  {32'h4035411c, 32'hc00f8e60} /* (24, 9, 15) {real, imag} */,
  {32'hc1315790, 32'h40f17428} /* (24, 9, 14) {real, imag} */,
  {32'hc0d5b216, 32'hc02ae604} /* (24, 9, 13) {real, imag} */,
  {32'hc0508558, 32'hc092f3f2} /* (24, 9, 12) {real, imag} */,
  {32'hc1229b35, 32'hbd1032c0} /* (24, 9, 11) {real, imag} */,
  {32'hc0b1215f, 32'h4172cc30} /* (24, 9, 10) {real, imag} */,
  {32'hc0b03e2e, 32'hbf32c678} /* (24, 9, 9) {real, imag} */,
  {32'hc0f9c855, 32'h409f3391} /* (24, 9, 8) {real, imag} */,
  {32'hc17a4be0, 32'h40ab0c5c} /* (24, 9, 7) {real, imag} */,
  {32'h4130991c, 32'h4044bb36} /* (24, 9, 6) {real, imag} */,
  {32'h41181b3f, 32'h40c78497} /* (24, 9, 5) {real, imag} */,
  {32'hc086f494, 32'hc0bea6ca} /* (24, 9, 4) {real, imag} */,
  {32'h3d9a5fa0, 32'hc19945a3} /* (24, 9, 3) {real, imag} */,
  {32'h3c409d00, 32'h4056d3b0} /* (24, 9, 2) {real, imag} */,
  {32'hc214bd6a, 32'h3f2fb200} /* (24, 9, 1) {real, imag} */,
  {32'h3f3079d0, 32'hc07e9448} /* (24, 9, 0) {real, imag} */,
  {32'h423ea0ad, 32'h41b7e9ca} /* (24, 8, 31) {real, imag} */,
  {32'hc1cf68e0, 32'hc111f9a2} /* (24, 8, 30) {real, imag} */,
  {32'h408c7710, 32'h40748fed} /* (24, 8, 29) {real, imag} */,
  {32'h41494199, 32'hc0b25374} /* (24, 8, 28) {real, imag} */,
  {32'hc17cf1e8, 32'h4146e3bc} /* (24, 8, 27) {real, imag} */,
  {32'h41140d74, 32'hc195afd0} /* (24, 8, 26) {real, imag} */,
  {32'h4193ccb2, 32'hc1c23c84} /* (24, 8, 25) {real, imag} */,
  {32'hc0612076, 32'hc166ae6b} /* (24, 8, 24) {real, imag} */,
  {32'h3eaa2c7c, 32'h413f9592} /* (24, 8, 23) {real, imag} */,
  {32'hbf143b35, 32'h4169c6b8} /* (24, 8, 22) {real, imag} */,
  {32'h3f6a3504, 32'h4180678e} /* (24, 8, 21) {real, imag} */,
  {32'h40ed8fe1, 32'h4149a799} /* (24, 8, 20) {real, imag} */,
  {32'hc096cfd5, 32'h4096372a} /* (24, 8, 19) {real, imag} */,
  {32'h3fbdc57c, 32'h3f527c88} /* (24, 8, 18) {real, imag} */,
  {32'h4021087a, 32'h401e3d86} /* (24, 8, 17) {real, imag} */,
  {32'hbeb01240, 32'hc125a4be} /* (24, 8, 16) {real, imag} */,
  {32'h408fbca5, 32'h4097b9b1} /* (24, 8, 15) {real, imag} */,
  {32'hc0220cf6, 32'h41070902} /* (24, 8, 14) {real, imag} */,
  {32'h41034d81, 32'hbfed91fc} /* (24, 8, 13) {real, imag} */,
  {32'h412455d0, 32'hc0e5f22e} /* (24, 8, 12) {real, imag} */,
  {32'h4053779f, 32'h40b9c296} /* (24, 8, 11) {real, imag} */,
  {32'hc044c118, 32'h4016ab60} /* (24, 8, 10) {real, imag} */,
  {32'hc09808df, 32'h40f62e16} /* (24, 8, 9) {real, imag} */,
  {32'hc13c57cc, 32'hc135a0d7} /* (24, 8, 8) {real, imag} */,
  {32'h3fc15558, 32'hc159cfe2} /* (24, 8, 7) {real, imag} */,
  {32'h416f4b3e, 32'hc17f90bd} /* (24, 8, 6) {real, imag} */,
  {32'hc19fe7d8, 32'hc0ac280d} /* (24, 8, 5) {real, imag} */,
  {32'h419a0965, 32'hbf51fdf0} /* (24, 8, 4) {real, imag} */,
  {32'hc1748a33, 32'hc138e8c0} /* (24, 8, 3) {real, imag} */,
  {32'hc1f5980a, 32'hc1783853} /* (24, 8, 2) {real, imag} */,
  {32'h4212f4bd, 32'h419e7531} /* (24, 8, 1) {real, imag} */,
  {32'h403e2992, 32'h412422e0} /* (24, 8, 0) {real, imag} */,
  {32'hc1f6203b, 32'h3eca1e40} /* (24, 7, 31) {real, imag} */,
  {32'h40826bdc, 32'h4118e15e} /* (24, 7, 30) {real, imag} */,
  {32'hc1231d50, 32'h40a75ee3} /* (24, 7, 29) {real, imag} */,
  {32'hc180d10b, 32'hc144eefd} /* (24, 7, 28) {real, imag} */,
  {32'hc14289f5, 32'h40242070} /* (24, 7, 27) {real, imag} */,
  {32'hc0ed6f4d, 32'hc1eafd46} /* (24, 7, 26) {real, imag} */,
  {32'h40c7b414, 32'h415ec1aa} /* (24, 7, 25) {real, imag} */,
  {32'h41268770, 32'h412b7aa4} /* (24, 7, 24) {real, imag} */,
  {32'h41a675bf, 32'h41315da0} /* (24, 7, 23) {real, imag} */,
  {32'hc00f8e96, 32'hc071a820} /* (24, 7, 22) {real, imag} */,
  {32'hc1931e78, 32'hc0383abc} /* (24, 7, 21) {real, imag} */,
  {32'h4010c83f, 32'h415e7e2c} /* (24, 7, 20) {real, imag} */,
  {32'hc0e54f6c, 32'h40b39b78} /* (24, 7, 19) {real, imag} */,
  {32'hc17f155e, 32'h3fada0f4} /* (24, 7, 18) {real, imag} */,
  {32'h4117384d, 32'hc0e73fb3} /* (24, 7, 17) {real, imag} */,
  {32'hc09015ad, 32'hc0bc8549} /* (24, 7, 16) {real, imag} */,
  {32'hc0ad6530, 32'h40f72870} /* (24, 7, 15) {real, imag} */,
  {32'h4191d8fa, 32'h414aea74} /* (24, 7, 14) {real, imag} */,
  {32'h4154befa, 32'hbfd5d662} /* (24, 7, 13) {real, imag} */,
  {32'h413a12ba, 32'h411800a2} /* (24, 7, 12) {real, imag} */,
  {32'hc08d0b2b, 32'h405a5912} /* (24, 7, 11) {real, imag} */,
  {32'hc136deb8, 32'h41b31fa9} /* (24, 7, 10) {real, imag} */,
  {32'h41810876, 32'hbffa1908} /* (24, 7, 9) {real, imag} */,
  {32'h40fc305a, 32'h42026b74} /* (24, 7, 8) {real, imag} */,
  {32'hc0eb2600, 32'hc14de22a} /* (24, 7, 7) {real, imag} */,
  {32'h3f3a2f40, 32'hc0875817} /* (24, 7, 6) {real, imag} */,
  {32'hc115c452, 32'h4154f8c1} /* (24, 7, 5) {real, imag} */,
  {32'h4104a084, 32'hbfdc8cab} /* (24, 7, 4) {real, imag} */,
  {32'hc18363fa, 32'h41b04c2c} /* (24, 7, 3) {real, imag} */,
  {32'hbefc3f30, 32'h4203b6c0} /* (24, 7, 2) {real, imag} */,
  {32'hc1ce74de, 32'hc1f477c7} /* (24, 7, 1) {real, imag} */,
  {32'hc1982442, 32'hc1270262} /* (24, 7, 0) {real, imag} */,
  {32'h4127404c, 32'hc09de668} /* (24, 6, 31) {real, imag} */,
  {32'hc0e28d1e, 32'h417450aa} /* (24, 6, 30) {real, imag} */,
  {32'hc1028e68, 32'hc1439cf5} /* (24, 6, 29) {real, imag} */,
  {32'h41a1d446, 32'h41a9c722} /* (24, 6, 28) {real, imag} */,
  {32'hbf91848c, 32'hbf33a7c0} /* (24, 6, 27) {real, imag} */,
  {32'hc1e5bf77, 32'h416318a0} /* (24, 6, 26) {real, imag} */,
  {32'hc02aef31, 32'h4190c9a1} /* (24, 6, 25) {real, imag} */,
  {32'hbf372104, 32'hc1b94bda} /* (24, 6, 24) {real, imag} */,
  {32'hc1546a88, 32'h3e8d88c0} /* (24, 6, 23) {real, imag} */,
  {32'hc120375e, 32'hc0c233b3} /* (24, 6, 22) {real, imag} */,
  {32'hc1415463, 32'h40dd6df0} /* (24, 6, 21) {real, imag} */,
  {32'h4169c9fc, 32'hbf8576c0} /* (24, 6, 20) {real, imag} */,
  {32'h41b10193, 32'hc0f64879} /* (24, 6, 19) {real, imag} */,
  {32'h3fcf319c, 32'hc10f6c61} /* (24, 6, 18) {real, imag} */,
  {32'h3ddaefb0, 32'h412713a1} /* (24, 6, 17) {real, imag} */,
  {32'hbe69df00, 32'hbfc71596} /* (24, 6, 16) {real, imag} */,
  {32'h4085609e, 32'hc0781e8c} /* (24, 6, 15) {real, imag} */,
  {32'h41188a54, 32'h40c4a596} /* (24, 6, 14) {real, imag} */,
  {32'hc10f0e0a, 32'hc009e157} /* (24, 6, 13) {real, imag} */,
  {32'hc0760737, 32'hc194597c} /* (24, 6, 12) {real, imag} */,
  {32'hc1b46da8, 32'h3e86fa20} /* (24, 6, 11) {real, imag} */,
  {32'hc149e764, 32'h410ac272} /* (24, 6, 10) {real, imag} */,
  {32'h41bfcafa, 32'hc122c0ca} /* (24, 6, 9) {real, imag} */,
  {32'hc106aba6, 32'hc1153478} /* (24, 6, 8) {real, imag} */,
  {32'hc137e425, 32'h40e13e98} /* (24, 6, 7) {real, imag} */,
  {32'h3d7d6880, 32'hc1d33a36} /* (24, 6, 6) {real, imag} */,
  {32'h41b70c02, 32'h3fe556f8} /* (24, 6, 5) {real, imag} */,
  {32'h414c1193, 32'h4137ad74} /* (24, 6, 4) {real, imag} */,
  {32'h3f95d6bc, 32'h40617376} /* (24, 6, 3) {real, imag} */,
  {32'h4210c538, 32'hc05c70aa} /* (24, 6, 2) {real, imag} */,
  {32'hc1111978, 32'hc089fe5b} /* (24, 6, 1) {real, imag} */,
  {32'hc014d688, 32'hc08ee3cc} /* (24, 6, 0) {real, imag} */,
  {32'h42e763bc, 32'h4170a48d} /* (24, 5, 31) {real, imag} */,
  {32'hc262499d, 32'h3f620c40} /* (24, 5, 30) {real, imag} */,
  {32'h40fc0ebd, 32'hc18639f2} /* (24, 5, 29) {real, imag} */,
  {32'h40b7cb82, 32'h403eeb96} /* (24, 5, 28) {real, imag} */,
  {32'hc1fcc1ae, 32'h41b5833a} /* (24, 5, 27) {real, imag} */,
  {32'h41a48003, 32'h3fc5ef68} /* (24, 5, 26) {real, imag} */,
  {32'hc1406f0a, 32'hc13cb7fe} /* (24, 5, 25) {real, imag} */,
  {32'hc0c03cbc, 32'hc114f407} /* (24, 5, 24) {real, imag} */,
  {32'h3ffd82fa, 32'h3f780d18} /* (24, 5, 23) {real, imag} */,
  {32'hc100da3d, 32'h41223213} /* (24, 5, 22) {real, imag} */,
  {32'hc0da5e72, 32'hbf0fa0a0} /* (24, 5, 21) {real, imag} */,
  {32'hc04875de, 32'h3fe29874} /* (24, 5, 20) {real, imag} */,
  {32'h4101c6c8, 32'hc11be939} /* (24, 5, 19) {real, imag} */,
  {32'hc0c25a2a, 32'h40829510} /* (24, 5, 18) {real, imag} */,
  {32'hc0ade89a, 32'h3f1ff5e6} /* (24, 5, 17) {real, imag} */,
  {32'h40dccb34, 32'h4050c612} /* (24, 5, 16) {real, imag} */,
  {32'hc113444c, 32'hc0726188} /* (24, 5, 15) {real, imag} */,
  {32'hc0bc3010, 32'hc15183d1} /* (24, 5, 14) {real, imag} */,
  {32'hc17b5636, 32'hc138926b} /* (24, 5, 13) {real, imag} */,
  {32'h40dbe933, 32'hbfc2e406} /* (24, 5, 12) {real, imag} */,
  {32'h403c3e9b, 32'h406423d4} /* (24, 5, 11) {real, imag} */,
  {32'h410477ec, 32'hc0c158ee} /* (24, 5, 10) {real, imag} */,
  {32'hc18812e2, 32'h40c1b86e} /* (24, 5, 9) {real, imag} */,
  {32'h402801d8, 32'hc1849e9a} /* (24, 5, 8) {real, imag} */,
  {32'h4141b58c, 32'h40f56444} /* (24, 5, 7) {real, imag} */,
  {32'hc13fe688, 32'hbe59b380} /* (24, 5, 6) {real, imag} */,
  {32'h3fe7c470, 32'hc18a69a6} /* (24, 5, 5) {real, imag} */,
  {32'h4050ba0c, 32'h420157cc} /* (24, 5, 4) {real, imag} */,
  {32'h4164cd44, 32'hc11e4582} /* (24, 5, 3) {real, imag} */,
  {32'hc205c5e0, 32'hc2314f54} /* (24, 5, 2) {real, imag} */,
  {32'h42543057, 32'h42a7e872} /* (24, 5, 1) {real, imag} */,
  {32'h4241438a, 32'h41f6d6c1} /* (24, 5, 0) {real, imag} */,
  {32'hc22f51f3, 32'hc2bb7c9e} /* (24, 4, 31) {real, imag} */,
  {32'h4292366f, 32'h42c99c03} /* (24, 4, 30) {real, imag} */,
  {32'h3f981108, 32'hc1ea39f2} /* (24, 4, 29) {real, imag} */,
  {32'hc263deca, 32'hc2123c7d} /* (24, 4, 28) {real, imag} */,
  {32'h414795a8, 32'hc16f6cb8} /* (24, 4, 27) {real, imag} */,
  {32'h41adbcfe, 32'hc19a5c43} /* (24, 4, 26) {real, imag} */,
  {32'hbff18830, 32'h403a8748} /* (24, 4, 25) {real, imag} */,
  {32'h418adde4, 32'h4142ceab} /* (24, 4, 24) {real, imag} */,
  {32'h41ac2990, 32'hc1613998} /* (24, 4, 23) {real, imag} */,
  {32'hc1885499, 32'h40db455c} /* (24, 4, 22) {real, imag} */,
  {32'h412f6748, 32'h40b77b8e} /* (24, 4, 21) {real, imag} */,
  {32'hbfe7ece0, 32'hbfee9530} /* (24, 4, 20) {real, imag} */,
  {32'hc0a60275, 32'hc0f022ee} /* (24, 4, 19) {real, imag} */,
  {32'h40a72405, 32'hc0bc16ea} /* (24, 4, 18) {real, imag} */,
  {32'h40e572e8, 32'h41699fd0} /* (24, 4, 17) {real, imag} */,
  {32'hc0d567d2, 32'h403c08e7} /* (24, 4, 16) {real, imag} */,
  {32'hbdcd8680, 32'hc0f6ca73} /* (24, 4, 15) {real, imag} */,
  {32'h408160ae, 32'h41126220} /* (24, 4, 14) {real, imag} */,
  {32'h40c6e964, 32'hc1215006} /* (24, 4, 13) {real, imag} */,
  {32'hc11711e0, 32'hc116043e} /* (24, 4, 12) {real, imag} */,
  {32'hc029feda, 32'h418213d6} /* (24, 4, 11) {real, imag} */,
  {32'h4138bd7f, 32'hc1808031} /* (24, 4, 10) {real, imag} */,
  {32'h41724d46, 32'h40bee805} /* (24, 4, 9) {real, imag} */,
  {32'hc09c8886, 32'h41558dee} /* (24, 4, 8) {real, imag} */,
  {32'hc1a91dd4, 32'h40d561fc} /* (24, 4, 7) {real, imag} */,
  {32'hc1d12acd, 32'h405b0574} /* (24, 4, 6) {real, imag} */,
  {32'hc11622e1, 32'h41adfb16} /* (24, 4, 5) {real, imag} */,
  {32'h41d9b7e6, 32'hc25d0dee} /* (24, 4, 4) {real, imag} */,
  {32'h41acbf7c, 32'hc144c790} /* (24, 4, 3) {real, imag} */,
  {32'h42f69f0c, 32'h424e413e} /* (24, 4, 2) {real, imag} */,
  {32'hc30f7771, 32'hc20d80e7} /* (24, 4, 1) {real, imag} */,
  {32'hc2970c33, 32'hc1f776a4} /* (24, 4, 0) {real, imag} */,
  {32'h42ee42f4, 32'hc2bb5b5c} /* (24, 3, 31) {real, imag} */,
  {32'hc28909d8, 32'h42aa7b68} /* (24, 3, 30) {real, imag} */,
  {32'h412e0e67, 32'h41ee17d9} /* (24, 3, 29) {real, imag} */,
  {32'hc1b0c5a2, 32'hc1fcc259} /* (24, 3, 28) {real, imag} */,
  {32'h4219523e, 32'h4109de0d} /* (24, 3, 27) {real, imag} */,
  {32'hc0b24cc2, 32'h412762ec} /* (24, 3, 26) {real, imag} */,
  {32'hc0b0bddc, 32'hc15e12ca} /* (24, 3, 25) {real, imag} */,
  {32'hc11ddd94, 32'h41abcb94} /* (24, 3, 24) {real, imag} */,
  {32'hc19c1dc0, 32'h40997d6d} /* (24, 3, 23) {real, imag} */,
  {32'h40d07c55, 32'h410b42fe} /* (24, 3, 22) {real, imag} */,
  {32'hc08808b6, 32'hc18ab045} /* (24, 3, 21) {real, imag} */,
  {32'h3fe88362, 32'h40c514c1} /* (24, 3, 20) {real, imag} */,
  {32'hc00d48ac, 32'hc1981ee6} /* (24, 3, 19) {real, imag} */,
  {32'h4119eda7, 32'h41b70f59} /* (24, 3, 18) {real, imag} */,
  {32'hc03d6eac, 32'h401c51d3} /* (24, 3, 17) {real, imag} */,
  {32'h40ce5534, 32'hc05980f4} /* (24, 3, 16) {real, imag} */,
  {32'h3fa1a4e8, 32'hbfc732c0} /* (24, 3, 15) {real, imag} */,
  {32'hbe8f6978, 32'h4011da00} /* (24, 3, 14) {real, imag} */,
  {32'hc1c7c258, 32'hc0757863} /* (24, 3, 13) {real, imag} */,
  {32'hbfefeac8, 32'hbfa97c70} /* (24, 3, 12) {real, imag} */,
  {32'h40f486fe, 32'h3f30a94c} /* (24, 3, 11) {real, imag} */,
  {32'h40bfb824, 32'hbe9e5a58} /* (24, 3, 10) {real, imag} */,
  {32'h41237a9c, 32'hc03111da} /* (24, 3, 9) {real, imag} */,
  {32'h404e781c, 32'h407f605e} /* (24, 3, 8) {real, imag} */,
  {32'hc140b7c2, 32'hbf6a4a60} /* (24, 3, 7) {real, imag} */,
  {32'hc17947b9, 32'h41fb27a8} /* (24, 3, 6) {real, imag} */,
  {32'hc0f4c42d, 32'hc1974d74} /* (24, 3, 5) {real, imag} */,
  {32'h42353f41, 32'hc19c749e} /* (24, 3, 4) {real, imag} */,
  {32'h3e641d40, 32'hc072ac48} /* (24, 3, 3) {real, imag} */,
  {32'hc1bd8f3c, 32'h42fb3b78} /* (24, 3, 2) {real, imag} */,
  {32'hc2ea3ab7, 32'hc2ae5ab6} /* (24, 3, 1) {real, imag} */,
  {32'h42baac1c, 32'h41332833} /* (24, 3, 0) {real, imag} */,
  {32'h4461eb34, 32'h426216af} /* (24, 2, 31) {real, imag} */,
  {32'hc3d475c7, 32'h42c91990} /* (24, 2, 30) {real, imag} */,
  {32'h42371b66, 32'hc1e04c0a} /* (24, 2, 29) {real, imag} */,
  {32'h424c8c7c, 32'hc244b9aa} /* (24, 2, 28) {real, imag} */,
  {32'hc1fe4eb0, 32'h4127d3d1} /* (24, 2, 27) {real, imag} */,
  {32'hc1c1d6bc, 32'h412976a5} /* (24, 2, 26) {real, imag} */,
  {32'hc12a64c7, 32'h412798e2} /* (24, 2, 25) {real, imag} */,
  {32'h3ecd80c0, 32'h421581f2} /* (24, 2, 24) {real, imag} */,
  {32'h418916ba, 32'h4036bbbe} /* (24, 2, 23) {real, imag} */,
  {32'hc11f356f, 32'hc1611de0} /* (24, 2, 22) {real, imag} */,
  {32'h41e617f8, 32'h4158d9fe} /* (24, 2, 21) {real, imag} */,
  {32'hc00870b4, 32'hc1743f38} /* (24, 2, 20) {real, imag} */,
  {32'hc0b67834, 32'h4124fbdf} /* (24, 2, 19) {real, imag} */,
  {32'h3fe81c4a, 32'h40e1a8ff} /* (24, 2, 18) {real, imag} */,
  {32'hc0bc473e, 32'h3f3f3598} /* (24, 2, 17) {real, imag} */,
  {32'hc0b2c55c, 32'h407b3631} /* (24, 2, 16) {real, imag} */,
  {32'h40435ade, 32'hc0c50d37} /* (24, 2, 15) {real, imag} */,
  {32'hbfb76e04, 32'hc09ec6f6} /* (24, 2, 14) {real, imag} */,
  {32'hc0929db8, 32'hc16cd54e} /* (24, 2, 13) {real, imag} */,
  {32'h411e9f07, 32'h413eb63c} /* (24, 2, 12) {real, imag} */,
  {32'hc106951e, 32'hc18a8943} /* (24, 2, 11) {real, imag} */,
  {32'h4121e90f, 32'hc18abe24} /* (24, 2, 10) {real, imag} */,
  {32'h40f9165d, 32'h3ed1be70} /* (24, 2, 9) {real, imag} */,
  {32'hc18d9b6e, 32'h40d1e0cf} /* (24, 2, 8) {real, imag} */,
  {32'h417633d0, 32'h40e0b594} /* (24, 2, 7) {real, imag} */,
  {32'h41c85b5a, 32'h3d8a57c0} /* (24, 2, 6) {real, imag} */,
  {32'hc29e93f2, 32'hc21c20fb} /* (24, 2, 5) {real, imag} */,
  {32'h42b49c5c, 32'h41a8ef62} /* (24, 2, 4) {real, imag} */,
  {32'h410689ce, 32'hc224e195} /* (24, 2, 3) {real, imag} */,
  {32'hc384b84e, 32'h4221f5cc} /* (24, 2, 2) {real, imag} */,
  {32'h4403bf18, 32'hc20b6cb7} /* (24, 2, 1) {real, imag} */,
  {32'h43f0ba5e, 32'h42921bb6} /* (24, 2, 0) {real, imag} */,
  {32'hc4977b8b, 32'h4397591a} /* (24, 1, 31) {real, imag} */,
  {32'h438a21ab, 32'h42b55130} /* (24, 1, 30) {real, imag} */,
  {32'h423cef3e, 32'hc1d067d0} /* (24, 1, 29) {real, imag} */,
  {32'hc2b1d835, 32'hc18f146e} /* (24, 1, 28) {real, imag} */,
  {32'h42bd1066, 32'hc11dc783} /* (24, 1, 27) {real, imag} */,
  {32'hc1e4ff74, 32'hc0de3bb6} /* (24, 1, 26) {real, imag} */,
  {32'hc1a995b9, 32'h41971191} /* (24, 1, 25) {real, imag} */,
  {32'h41edf247, 32'hc1f56b36} /* (24, 1, 24) {real, imag} */,
  {32'h415fb864, 32'h409fab2d} /* (24, 1, 23) {real, imag} */,
  {32'h40ad67a2, 32'hc1a21b46} /* (24, 1, 22) {real, imag} */,
  {32'h411b3418, 32'hc1ce1184} /* (24, 1, 21) {real, imag} */,
  {32'hc1a3941a, 32'h410842c2} /* (24, 1, 20) {real, imag} */,
  {32'h4097426a, 32'hc191c677} /* (24, 1, 19) {real, imag} */,
  {32'hbfd87bf8, 32'hc18aa1f2} /* (24, 1, 18) {real, imag} */,
  {32'h401bd268, 32'h40dfb4ea} /* (24, 1, 17) {real, imag} */,
  {32'h3f446fc8, 32'hc04209b4} /* (24, 1, 16) {real, imag} */,
  {32'hbebd1c00, 32'hc05c9e08} /* (24, 1, 15) {real, imag} */,
  {32'hc0e9c1a8, 32'h417d4c14} /* (24, 1, 14) {real, imag} */,
  {32'hbdbb4ba0, 32'hc14efacc} /* (24, 1, 13) {real, imag} */,
  {32'hc05c2fc6, 32'hbf340ca0} /* (24, 1, 12) {real, imag} */,
  {32'h40cc3c0d, 32'h41811cc6} /* (24, 1, 11) {real, imag} */,
  {32'hc0d7a006, 32'hc0f6db3a} /* (24, 1, 10) {real, imag} */,
  {32'hbd73f480, 32'h40fdbbe6} /* (24, 1, 9) {real, imag} */,
  {32'h41c97c17, 32'h41d9d703} /* (24, 1, 8) {real, imag} */,
  {32'hc1465812, 32'hc16b890a} /* (24, 1, 7) {real, imag} */,
  {32'h417a6cdc, 32'hbfa01aa8} /* (24, 1, 6) {real, imag} */,
  {32'h4286aabc, 32'h423d260a} /* (24, 1, 5) {real, imag} */,
  {32'hc1c8c5bc, 32'hc240efb0} /* (24, 1, 4) {real, imag} */,
  {32'h41acdc58, 32'h4176266a} /* (24, 1, 3) {real, imag} */,
  {32'h43d3f596, 32'h43cc952c} /* (24, 1, 2) {real, imag} */,
  {32'hc4da1b49, 32'hc47ba9e1} /* (24, 1, 1) {real, imag} */,
  {32'hc4cea4af, 32'hc35bd352} /* (24, 1, 0) {real, imag} */,
  {32'hc498aeef, 32'h446ece01} /* (24, 0, 31) {real, imag} */,
  {32'h43036024, 32'hc31e667a} /* (24, 0, 30) {real, imag} */,
  {32'h4202c1d0, 32'h41ae93e5} /* (24, 0, 29) {real, imag} */,
  {32'h420c1c00, 32'hc2afa9ed} /* (24, 0, 28) {real, imag} */,
  {32'h425a5078, 32'hc198fd08} /* (24, 0, 27) {real, imag} */,
  {32'h41af62fa, 32'h40315f7c} /* (24, 0, 26) {real, imag} */,
  {32'h41b98a10, 32'h40d82484} /* (24, 0, 25) {real, imag} */,
  {32'h40b77c1e, 32'hc1207ca8} /* (24, 0, 24) {real, imag} */,
  {32'hc1b25277, 32'hc1278586} /* (24, 0, 23) {real, imag} */,
  {32'hc07a43db, 32'hc0fd8f1c} /* (24, 0, 22) {real, imag} */,
  {32'hbf01da88, 32'hbe9a1e60} /* (24, 0, 21) {real, imag} */,
  {32'hc1944378, 32'hc0378edc} /* (24, 0, 20) {real, imag} */,
  {32'hc031880c, 32'h3f9b49fb} /* (24, 0, 19) {real, imag} */,
  {32'h41774a8e, 32'hbfea3550} /* (24, 0, 18) {real, imag} */,
  {32'hc0483e7f, 32'h3f720684} /* (24, 0, 17) {real, imag} */,
  {32'h415e1625, 32'h00000000} /* (24, 0, 16) {real, imag} */,
  {32'hc0483e7f, 32'hbf720684} /* (24, 0, 15) {real, imag} */,
  {32'h41774a8e, 32'h3fea3550} /* (24, 0, 14) {real, imag} */,
  {32'hc031880c, 32'hbf9b49fb} /* (24, 0, 13) {real, imag} */,
  {32'hc1944378, 32'h40378edc} /* (24, 0, 12) {real, imag} */,
  {32'hbf01da88, 32'h3e9a1e60} /* (24, 0, 11) {real, imag} */,
  {32'hc07a43db, 32'h40fd8f1c} /* (24, 0, 10) {real, imag} */,
  {32'hc1b25277, 32'h41278586} /* (24, 0, 9) {real, imag} */,
  {32'h40b77c1e, 32'h41207ca8} /* (24, 0, 8) {real, imag} */,
  {32'h41b98a10, 32'hc0d82484} /* (24, 0, 7) {real, imag} */,
  {32'h41af62fa, 32'hc0315f7c} /* (24, 0, 6) {real, imag} */,
  {32'h425a5078, 32'h4198fd08} /* (24, 0, 5) {real, imag} */,
  {32'h420c1c00, 32'h42afa9ed} /* (24, 0, 4) {real, imag} */,
  {32'h4202c1d0, 32'hc1ae93e5} /* (24, 0, 3) {real, imag} */,
  {32'h43036024, 32'h431e667a} /* (24, 0, 2) {real, imag} */,
  {32'hc498aeef, 32'hc46ece01} /* (24, 0, 1) {real, imag} */,
  {32'hc4f08769, 32'h00000000} /* (24, 0, 0) {real, imag} */,
  {32'hc5068bfc, 32'h4497fdc2} /* (23, 31, 31) {real, imag} */,
  {32'h4403b620, 32'hc3f4792e} /* (23, 31, 30) {real, imag} */,
  {32'h426795ba, 32'hc1917c12} /* (23, 31, 29) {real, imag} */,
  {32'hc2779290, 32'h424e75d0} /* (23, 31, 28) {real, imag} */,
  {32'h4289667e, 32'hc23c3ea8} /* (23, 31, 27) {real, imag} */,
  {32'h41fa9161, 32'h419f313e} /* (23, 31, 26) {real, imag} */,
  {32'hc19b6a79, 32'h41713484} /* (23, 31, 25) {real, imag} */,
  {32'h4188e354, 32'hc1847db0} /* (23, 31, 24) {real, imag} */,
  {32'h41a2d8b8, 32'hc0d60520} /* (23, 31, 23) {real, imag} */,
  {32'h410a7593, 32'h4025abe0} /* (23, 31, 22) {real, imag} */,
  {32'hc0957f2a, 32'hc1c9ef1c} /* (23, 31, 21) {real, imag} */,
  {32'h401276c0, 32'h400b597a} /* (23, 31, 20) {real, imag} */,
  {32'h3fc12f58, 32'h411cd642} /* (23, 31, 19) {real, imag} */,
  {32'hbdfaf530, 32'hc0f11340} /* (23, 31, 18) {real, imag} */,
  {32'h40957fdf, 32'h4045ed62} /* (23, 31, 17) {real, imag} */,
  {32'hbf4096e4, 32'hbfb7c518} /* (23, 31, 16) {real, imag} */,
  {32'h40261db8, 32'h414b530e} /* (23, 31, 15) {real, imag} */,
  {32'hc115d8c3, 32'h4101f154} /* (23, 31, 14) {real, imag} */,
  {32'h3f431cb4, 32'hc0a416b5} /* (23, 31, 13) {real, imag} */,
  {32'hc03680a9, 32'hbfa71c0e} /* (23, 31, 12) {real, imag} */,
  {32'h4154f591, 32'h40e26385} /* (23, 31, 11) {real, imag} */,
  {32'hc135a73e, 32'h3e746030} /* (23, 31, 10) {real, imag} */,
  {32'h410b3e58, 32'h4182ef78} /* (23, 31, 9) {real, imag} */,
  {32'h4164f898, 32'h4198423e} /* (23, 31, 8) {real, imag} */,
  {32'hc188bbaa, 32'hc1b2af03} /* (23, 31, 7) {real, imag} */,
  {32'h41800e6c, 32'hc08ba27f} /* (23, 31, 6) {real, imag} */,
  {32'h43035292, 32'h410a4b87} /* (23, 31, 5) {real, imag} */,
  {32'hc2f497c3, 32'h41bb464a} /* (23, 31, 4) {real, imag} */,
  {32'h423ed4c7, 32'h42117ce6} /* (23, 31, 3) {real, imag} */,
  {32'h43b97e08, 32'hc2c7a4af} /* (23, 31, 2) {real, imag} */,
  {32'hc4bef642, 32'hc3c64375} /* (23, 31, 1) {real, imag} */,
  {32'hc4f7c643, 32'h43749fae} /* (23, 31, 0) {real, imag} */,
  {32'h4423b111, 32'h428030bb} /* (23, 30, 31) {real, imag} */,
  {32'hc3b782d9, 32'hc26039dd} /* (23, 30, 30) {real, imag} */,
  {32'h40b051ae, 32'h4204bbfa} /* (23, 30, 29) {real, imag} */,
  {32'h42bae243, 32'hc26f8566} /* (23, 30, 28) {real, imag} */,
  {32'hc29969ca, 32'h42895e65} /* (23, 30, 27) {real, imag} */,
  {32'hbfdb9b90, 32'hc094fb42} /* (23, 30, 26) {real, imag} */,
  {32'h4192a0e2, 32'hc118f4de} /* (23, 30, 25) {real, imag} */,
  {32'hc1c7eb87, 32'hc1c0f53e} /* (23, 30, 24) {real, imag} */,
  {32'h4134e1ee, 32'hc149d1cb} /* (23, 30, 23) {real, imag} */,
  {32'h407705b6, 32'hc13f5da4} /* (23, 30, 22) {real, imag} */,
  {32'hc128cdde, 32'h4169f938} /* (23, 30, 21) {real, imag} */,
  {32'hc0901495, 32'hc083563e} /* (23, 30, 20) {real, imag} */,
  {32'hc08d3392, 32'h3f436538} /* (23, 30, 19) {real, imag} */,
  {32'hc0ddafee, 32'h3ffc2230} /* (23, 30, 18) {real, imag} */,
  {32'h414d39ba, 32'hc1040d6c} /* (23, 30, 17) {real, imag} */,
  {32'hc10054e7, 32'hc14cd86c} /* (23, 30, 16) {real, imag} */,
  {32'hc116f083, 32'h414a5172} /* (23, 30, 15) {real, imag} */,
  {32'h3f77215d, 32'hbf4684e0} /* (23, 30, 14) {real, imag} */,
  {32'h40e81410, 32'hc10996f8} /* (23, 30, 13) {real, imag} */,
  {32'h40b49ca0, 32'hc1035139} /* (23, 30, 12) {real, imag} */,
  {32'hc0219e03, 32'h3f1d9d76} /* (23, 30, 11) {real, imag} */,
  {32'h404a5c8e, 32'hc10e57a6} /* (23, 30, 10) {real, imag} */,
  {32'hc112a177, 32'hc0ea2e14} /* (23, 30, 9) {real, imag} */,
  {32'hc08e63de, 32'hc1875939} /* (23, 30, 8) {real, imag} */,
  {32'h409d8022, 32'hc0c9aef5} /* (23, 30, 7) {real, imag} */,
  {32'hc14dc896, 32'hc1a648f5} /* (23, 30, 6) {real, imag} */,
  {32'hc26f603e, 32'hc170b745} /* (23, 30, 5) {real, imag} */,
  {32'h4210b104, 32'h42a6d48d} /* (23, 30, 4) {real, imag} */,
  {32'h4205622a, 32'h41fe6136} /* (23, 30, 3) {real, imag} */,
  {32'hc4004dd6, 32'hc318de2e} /* (23, 30, 2) {real, imag} */,
  {32'h448d8d54, 32'hc28929ed} /* (23, 30, 1) {real, imag} */,
  {32'h44136f1d, 32'hc2debdb6} /* (23, 30, 0) {real, imag} */,
  {32'hc2fa0378, 32'h428b5b6e} /* (23, 29, 31) {real, imag} */,
  {32'hc18fba7a, 32'hc314b7e2} /* (23, 29, 30) {real, imag} */,
  {32'hc1098167, 32'h40f2d87c} /* (23, 29, 29) {real, imag} */,
  {32'h4219a45a, 32'h42171346} /* (23, 29, 28) {real, imag} */,
  {32'hc17f5bf6, 32'h4198e7ab} /* (23, 29, 27) {real, imag} */,
  {32'hc1475569, 32'hc1aba4e3} /* (23, 29, 26) {real, imag} */,
  {32'hc135a23a, 32'h41afadc0} /* (23, 29, 25) {real, imag} */,
  {32'hc1060738, 32'hc161a9de} /* (23, 29, 24) {real, imag} */,
  {32'h40047a64, 32'hbe970c38} /* (23, 29, 23) {real, imag} */,
  {32'hc0b28a51, 32'hc0efe7f5} /* (23, 29, 22) {real, imag} */,
  {32'h411452f5, 32'h40dfc04f} /* (23, 29, 21) {real, imag} */,
  {32'hc1860867, 32'h417bb03a} /* (23, 29, 20) {real, imag} */,
  {32'h403bc1ae, 32'hc009c567} /* (23, 29, 19) {real, imag} */,
  {32'h3f6ab118, 32'hc121dce6} /* (23, 29, 18) {real, imag} */,
  {32'h4091f61f, 32'h405af65c} /* (23, 29, 17) {real, imag} */,
  {32'h4189be82, 32'hbf8e9e6c} /* (23, 29, 16) {real, imag} */,
  {32'hc11b4e51, 32'hc07626b0} /* (23, 29, 15) {real, imag} */,
  {32'h40e61327, 32'hc0c2aa06} /* (23, 29, 14) {real, imag} */,
  {32'hc0f5e146, 32'hc12f8656} /* (23, 29, 13) {real, imag} */,
  {32'hc10803fc, 32'h415798a4} /* (23, 29, 12) {real, imag} */,
  {32'h3ff34252, 32'h40dd369b} /* (23, 29, 11) {real, imag} */,
  {32'hc044a30c, 32'h400b2673} /* (23, 29, 10) {real, imag} */,
  {32'hc13a70ab, 32'h4169f307} /* (23, 29, 9) {real, imag} */,
  {32'hc0f842c4, 32'hc1518260} /* (23, 29, 8) {real, imag} */,
  {32'hbed1c5c0, 32'h41f302c2} /* (23, 29, 7) {real, imag} */,
  {32'hc1210dfb, 32'hc0b854ed} /* (23, 29, 6) {real, imag} */,
  {32'h423e318e, 32'hc044c28c} /* (23, 29, 5) {real, imag} */,
  {32'hc21632bb, 32'h41d38c60} /* (23, 29, 4) {real, imag} */,
  {32'hc16b201a, 32'hc122248a} /* (23, 29, 3) {real, imag} */,
  {32'hc284e30c, 32'hc2cca452} /* (23, 29, 2) {real, imag} */,
  {32'h4307fc76, 32'h42aade2e} /* (23, 29, 1) {real, imag} */,
  {32'h42b289dc, 32'hc10fab8d} /* (23, 29, 0) {real, imag} */,
  {32'hc304c3d7, 32'h426f1274} /* (23, 28, 31) {real, imag} */,
  {32'h42ec2057, 32'hc2618a3b} /* (23, 28, 30) {real, imag} */,
  {32'h41702ed0, 32'h41c49130} /* (23, 28, 29) {real, imag} */,
  {32'h4206d6d6, 32'h42265bf0} /* (23, 28, 28) {real, imag} */,
  {32'h410a241c, 32'hc0270af4} /* (23, 28, 27) {real, imag} */,
  {32'hc19cb234, 32'hc0a4a876} /* (23, 28, 26) {real, imag} */,
  {32'hc1c39506, 32'h41049418} /* (23, 28, 25) {real, imag} */,
  {32'h408b4bbe, 32'h414c0111} /* (23, 28, 24) {real, imag} */,
  {32'hc0ef21ae, 32'h412f7851} /* (23, 28, 23) {real, imag} */,
  {32'h40fdbe28, 32'hc10a49f0} /* (23, 28, 22) {real, imag} */,
  {32'hc1621ae0, 32'hc14690a3} /* (23, 28, 21) {real, imag} */,
  {32'hc06f15c8, 32'hbf94386c} /* (23, 28, 20) {real, imag} */,
  {32'hc033f2ec, 32'hc0f2c11e} /* (23, 28, 19) {real, imag} */,
  {32'h3e9399c8, 32'hc15b53d6} /* (23, 28, 18) {real, imag} */,
  {32'h412fde39, 32'h40adc509} /* (23, 28, 17) {real, imag} */,
  {32'hc017fd9a, 32'hc0539c0b} /* (23, 28, 16) {real, imag} */,
  {32'h3f257258, 32'h4134ff53} /* (23, 28, 15) {real, imag} */,
  {32'h3fd6d6cc, 32'hc115c101} /* (23, 28, 14) {real, imag} */,
  {32'h41615fd6, 32'h40cb687f} /* (23, 28, 13) {real, imag} */,
  {32'h410448f0, 32'hc155fba0} /* (23, 28, 12) {real, imag} */,
  {32'h3ec42a58, 32'h410d2907} /* (23, 28, 11) {real, imag} */,
  {32'hc171ffd4, 32'hc1027f1a} /* (23, 28, 10) {real, imag} */,
  {32'hc039c4ba, 32'h3e500048} /* (23, 28, 9) {real, imag} */,
  {32'h424a805e, 32'hc08fce1c} /* (23, 28, 8) {real, imag} */,
  {32'hc14e9410, 32'h400da686} /* (23, 28, 7) {real, imag} */,
  {32'hc0942418, 32'h40ae4926} /* (23, 28, 6) {real, imag} */,
  {32'h41d12176, 32'h41d4c085} /* (23, 28, 5) {real, imag} */,
  {32'hc2433705, 32'h41777f69} /* (23, 28, 4) {real, imag} */,
  {32'h40f356ad, 32'h40457254} /* (23, 28, 3) {real, imag} */,
  {32'h42be3f20, 32'hc2b6ddde} /* (23, 28, 2) {real, imag} */,
  {32'hc24c40d1, 32'h42c23c90} /* (23, 28, 1) {real, imag} */,
  {32'hc29b529e, 32'hc1a18e94} /* (23, 28, 0) {real, imag} */,
  {32'h428039a0, 32'hc2a4d11e} /* (23, 27, 31) {real, imag} */,
  {32'hc17ae3ee, 32'h420f6100} /* (23, 27, 30) {real, imag} */,
  {32'h409f5de4, 32'h4191ecb0} /* (23, 27, 29) {real, imag} */,
  {32'h40f41b86, 32'hc23d769c} /* (23, 27, 28) {real, imag} */,
  {32'h3f1a0680, 32'h41e1f99c} /* (23, 27, 27) {real, imag} */,
  {32'h3eeb3bc0, 32'hc17f234c} /* (23, 27, 26) {real, imag} */,
  {32'h3e1a4540, 32'h3fb70114} /* (23, 27, 25) {real, imag} */,
  {32'h41c6e1f5, 32'hbfbbcd28} /* (23, 27, 24) {real, imag} */,
  {32'hbd225580, 32'h402bb5bf} /* (23, 27, 23) {real, imag} */,
  {32'hc1518ac2, 32'h3edc3ec0} /* (23, 27, 22) {real, imag} */,
  {32'hc1341078, 32'h4184a428} /* (23, 27, 21) {real, imag} */,
  {32'hc01814bd, 32'hbd3827e0} /* (23, 27, 20) {real, imag} */,
  {32'hc02c6413, 32'h40b97878} /* (23, 27, 19) {real, imag} */,
  {32'hbf0a9cc0, 32'h4023d4dd} /* (23, 27, 18) {real, imag} */,
  {32'hbf917420, 32'h40899dbe} /* (23, 27, 17) {real, imag} */,
  {32'h40346ed0, 32'hc11f71ca} /* (23, 27, 16) {real, imag} */,
  {32'hc0b4298b, 32'h3fc744bc} /* (23, 27, 15) {real, imag} */,
  {32'h3f45fcf8, 32'hc08d26e2} /* (23, 27, 14) {real, imag} */,
  {32'h40c3a10c, 32'hc180a834} /* (23, 27, 13) {real, imag} */,
  {32'h40052f14, 32'hc01a7d22} /* (23, 27, 12) {real, imag} */,
  {32'h409c1f36, 32'h4137d366} /* (23, 27, 11) {real, imag} */,
  {32'hc11e4626, 32'h403ba524} /* (23, 27, 10) {real, imag} */,
  {32'h4195c50e, 32'hc018f537} /* (23, 27, 9) {real, imag} */,
  {32'hc0178cf6, 32'hc0d7d9aa} /* (23, 27, 8) {real, imag} */,
  {32'h4003c90d, 32'h41849993} /* (23, 27, 7) {real, imag} */,
  {32'hc14b39b2, 32'h4059ee3c} /* (23, 27, 6) {real, imag} */,
  {32'hc218a6e6, 32'h411e20a0} /* (23, 27, 5) {real, imag} */,
  {32'h40fb3e3a, 32'h41cb11bb} /* (23, 27, 4) {real, imag} */,
  {32'h41d1db1b, 32'h41532b5d} /* (23, 27, 3) {real, imag} */,
  {32'hc27d2036, 32'hc145ac7f} /* (23, 27, 2) {real, imag} */,
  {32'h42d84026, 32'hc209b5bd} /* (23, 27, 1) {real, imag} */,
  {32'h42979ddc, 32'hc20a2077} /* (23, 27, 0) {real, imag} */,
  {32'h41678306, 32'hc141db32} /* (23, 26, 31) {real, imag} */,
  {32'hc1415c35, 32'h40281fbc} /* (23, 26, 30) {real, imag} */,
  {32'h412c603a, 32'h4115a49c} /* (23, 26, 29) {real, imag} */,
  {32'h419b5aee, 32'h41649fc4} /* (23, 26, 28) {real, imag} */,
  {32'hbbef5e00, 32'hc16bf90a} /* (23, 26, 27) {real, imag} */,
  {32'hc1c99020, 32'hbf002df0} /* (23, 26, 26) {real, imag} */,
  {32'hc10ddbfb, 32'hc15fafae} /* (23, 26, 25) {real, imag} */,
  {32'hc1820dad, 32'h40aebc9c} /* (23, 26, 24) {real, imag} */,
  {32'hbfcde19c, 32'hc0cd831d} /* (23, 26, 23) {real, imag} */,
  {32'hc0afed9e, 32'hc0ae63c2} /* (23, 26, 22) {real, imag} */,
  {32'hc13ebffc, 32'hc1559f47} /* (23, 26, 21) {real, imag} */,
  {32'h3fea1554, 32'h3fed0980} /* (23, 26, 20) {real, imag} */,
  {32'hc05ccd0a, 32'hc0515180} /* (23, 26, 19) {real, imag} */,
  {32'h3fdb7960, 32'hc10335c0} /* (23, 26, 18) {real, imag} */,
  {32'h40b17006, 32'hbfb00cce} /* (23, 26, 17) {real, imag} */,
  {32'h402053c4, 32'h4145b694} /* (23, 26, 16) {real, imag} */,
  {32'h408fde06, 32'h3fcb38dc} /* (23, 26, 15) {real, imag} */,
  {32'h41520c32, 32'h40a0bb34} /* (23, 26, 14) {real, imag} */,
  {32'hc13264af, 32'hc0a9ad21} /* (23, 26, 13) {real, imag} */,
  {32'h414671de, 32'h4090ceb2} /* (23, 26, 12) {real, imag} */,
  {32'hc17292ee, 32'h3e9ab3a0} /* (23, 26, 11) {real, imag} */,
  {32'hc1457b56, 32'h41b05815} /* (23, 26, 10) {real, imag} */,
  {32'h409e337f, 32'hc0e419b8} /* (23, 26, 9) {real, imag} */,
  {32'hbf9a8b74, 32'hc05f09be} /* (23, 26, 8) {real, imag} */,
  {32'h40e0ce3c, 32'h405513eb} /* (23, 26, 7) {real, imag} */,
  {32'hc1e68903, 32'hc00c0338} /* (23, 26, 6) {real, imag} */,
  {32'hc09f516d, 32'hc1b8e9c2} /* (23, 26, 5) {real, imag} */,
  {32'hbe2909c0, 32'hc1d65081} /* (23, 26, 4) {real, imag} */,
  {32'hc13c4c1c, 32'h41a384bc} /* (23, 26, 3) {real, imag} */,
  {32'hc0334f8c, 32'h4084adf7} /* (23, 26, 2) {real, imag} */,
  {32'h41343a3f, 32'h41c79094} /* (23, 26, 1) {real, imag} */,
  {32'h40a102da, 32'h40ae895c} /* (23, 26, 0) {real, imag} */,
  {32'hc13629ee, 32'h420501b4} /* (23, 25, 31) {real, imag} */,
  {32'h41cb8a6c, 32'h3f332fb0} /* (23, 25, 30) {real, imag} */,
  {32'hc141d150, 32'hc1aa09f7} /* (23, 25, 29) {real, imag} */,
  {32'h410ef746, 32'hbf8f6750} /* (23, 25, 28) {real, imag} */,
  {32'h4002a37c, 32'hc0927f6f} /* (23, 25, 27) {real, imag} */,
  {32'h4199dc3c, 32'hc0e8b651} /* (23, 25, 26) {real, imag} */,
  {32'h41493031, 32'h40a7d049} /* (23, 25, 25) {real, imag} */,
  {32'h41768fcc, 32'h3d9bca20} /* (23, 25, 24) {real, imag} */,
  {32'hc0d697fa, 32'h410e8c3e} /* (23, 25, 23) {real, imag} */,
  {32'hc0fa8098, 32'hc13e5339} /* (23, 25, 22) {real, imag} */,
  {32'h40acb3e1, 32'h41578a4d} /* (23, 25, 21) {real, imag} */,
  {32'hc1712f4b, 32'h4090fb74} /* (23, 25, 20) {real, imag} */,
  {32'h40f20ba2, 32'hbff4b1e0} /* (23, 25, 19) {real, imag} */,
  {32'hc0eac151, 32'h40151972} /* (23, 25, 18) {real, imag} */,
  {32'h4061d248, 32'h40117d8a} /* (23, 25, 17) {real, imag} */,
  {32'h40eefa2a, 32'h4174e8a6} /* (23, 25, 16) {real, imag} */,
  {32'h410ab6e3, 32'h417f4848} /* (23, 25, 15) {real, imag} */,
  {32'hc0ccd845, 32'hc030765c} /* (23, 25, 14) {real, imag} */,
  {32'h3fbe6590, 32'h3fe422bc} /* (23, 25, 13) {real, imag} */,
  {32'h41284ace, 32'h414451a2} /* (23, 25, 12) {real, imag} */,
  {32'hc002eabe, 32'hbfaed48a} /* (23, 25, 11) {real, imag} */,
  {32'h41011315, 32'hc04a9ef2} /* (23, 25, 10) {real, imag} */,
  {32'h4115f174, 32'hc070079c} /* (23, 25, 9) {real, imag} */,
  {32'h416f2485, 32'hc134965f} /* (23, 25, 8) {real, imag} */,
  {32'hc13d1f38, 32'hbffc6c08} /* (23, 25, 7) {real, imag} */,
  {32'hc0a6fd25, 32'hc1cdb741} /* (23, 25, 6) {real, imag} */,
  {32'hc1b08a3a, 32'hc059bd1e} /* (23, 25, 5) {real, imag} */,
  {32'h418a148e, 32'h3fef9068} /* (23, 25, 4) {real, imag} */,
  {32'h41301304, 32'hc15be9bf} /* (23, 25, 3) {real, imag} */,
  {32'hc0ed11b6, 32'hc133f151} /* (23, 25, 2) {real, imag} */,
  {32'hc211e3b0, 32'h41149aa7} /* (23, 25, 1) {real, imag} */,
  {32'h409e47b3, 32'h41eedda0} /* (23, 25, 0) {real, imag} */,
  {32'h4003f8d6, 32'hc19e10c6} /* (23, 24, 31) {real, imag} */,
  {32'hc18ff9e0, 32'h40a7689c} /* (23, 24, 30) {real, imag} */,
  {32'h40eb53a0, 32'h4193cd37} /* (23, 24, 29) {real, imag} */,
  {32'h40b057c6, 32'hc091b212} /* (23, 24, 28) {real, imag} */,
  {32'hc0f0d0f6, 32'h420079c3} /* (23, 24, 27) {real, imag} */,
  {32'h3f175200, 32'hc183ea75} /* (23, 24, 26) {real, imag} */,
  {32'h420d0358, 32'h409775a0} /* (23, 24, 25) {real, imag} */,
  {32'hc175b386, 32'h412563c2} /* (23, 24, 24) {real, imag} */,
  {32'hbfda6674, 32'h412c4477} /* (23, 24, 23) {real, imag} */,
  {32'h41c740e4, 32'hc155221a} /* (23, 24, 22) {real, imag} */,
  {32'h410c3290, 32'h4128ac84} /* (23, 24, 21) {real, imag} */,
  {32'hc1414446, 32'hc0702e25} /* (23, 24, 20) {real, imag} */,
  {32'hc16d2f37, 32'hc1447da2} /* (23, 24, 19) {real, imag} */,
  {32'hbfc9f93c, 32'h410ae0e8} /* (23, 24, 18) {real, imag} */,
  {32'h40646d53, 32'hc086d88c} /* (23, 24, 17) {real, imag} */,
  {32'h4111cdc1, 32'h40e58322} /* (23, 24, 16) {real, imag} */,
  {32'h403065b1, 32'h40d16526} /* (23, 24, 15) {real, imag} */,
  {32'hc064c3f6, 32'hc03825d6} /* (23, 24, 14) {real, imag} */,
  {32'h410944f9, 32'hc096ae51} /* (23, 24, 13) {real, imag} */,
  {32'hc0d312e0, 32'h40973606} /* (23, 24, 12) {real, imag} */,
  {32'h41264767, 32'h40dfe905} /* (23, 24, 11) {real, imag} */,
  {32'h40c2664c, 32'h4153b718} /* (23, 24, 10) {real, imag} */,
  {32'hc08f55d2, 32'hc13d71e5} /* (23, 24, 9) {real, imag} */,
  {32'hc187091e, 32'hc040aa8c} /* (23, 24, 8) {real, imag} */,
  {32'h40f7a234, 32'h418a31ef} /* (23, 24, 7) {real, imag} */,
  {32'h40b9efba, 32'h40cb6392} /* (23, 24, 6) {real, imag} */,
  {32'hc142072e, 32'hc133d818} /* (23, 24, 5) {real, imag} */,
  {32'h40d534c3, 32'h416b2516} /* (23, 24, 4) {real, imag} */,
  {32'h4046c4c9, 32'hc0cd7145} /* (23, 24, 3) {real, imag} */,
  {32'hc1a8028d, 32'h409ca0f0} /* (23, 24, 2) {real, imag} */,
  {32'h424aaac8, 32'hc18862db} /* (23, 24, 1) {real, imag} */,
  {32'h40ff9ee4, 32'hc1a6abbc} /* (23, 24, 0) {real, imag} */,
  {32'hc1de8423, 32'h41a44a91} /* (23, 23, 31) {real, imag} */,
  {32'hc18c1a68, 32'h40021c94} /* (23, 23, 30) {real, imag} */,
  {32'hc05f7302, 32'hc03c2280} /* (23, 23, 29) {real, imag} */,
  {32'hbf5e0670, 32'hc10e6080} /* (23, 23, 28) {real, imag} */,
  {32'hc188db91, 32'hc0445ba8} /* (23, 23, 27) {real, imag} */,
  {32'h404f040f, 32'h40817a2d} /* (23, 23, 26) {real, imag} */,
  {32'h40bdd510, 32'hc11b9214} /* (23, 23, 25) {real, imag} */,
  {32'h41b163be, 32'hc18497e0} /* (23, 23, 24) {real, imag} */,
  {32'hc0cc66d6, 32'hc141e3a6} /* (23, 23, 23) {real, imag} */,
  {32'h41d0fd49, 32'h3fda12e8} /* (23, 23, 22) {real, imag} */,
  {32'hc0b9bf76, 32'h408da08b} /* (23, 23, 21) {real, imag} */,
  {32'h41744ef3, 32'hc16cb563} /* (23, 23, 20) {real, imag} */,
  {32'h40d3b34e, 32'h40ca94c4} /* (23, 23, 19) {real, imag} */,
  {32'h407436f0, 32'h4074dd01} /* (23, 23, 18) {real, imag} */,
  {32'h4116dabc, 32'h410f19d0} /* (23, 23, 17) {real, imag} */,
  {32'h410fe848, 32'h40cf384c} /* (23, 23, 16) {real, imag} */,
  {32'hc1158493, 32'h40951e47} /* (23, 23, 15) {real, imag} */,
  {32'hc0c1c57c, 32'hc124b509} /* (23, 23, 14) {real, imag} */,
  {32'h4104e7d6, 32'h414691ab} /* (23, 23, 13) {real, imag} */,
  {32'h41598078, 32'h411193e7} /* (23, 23, 12) {real, imag} */,
  {32'hc0e603e4, 32'hc1106264} /* (23, 23, 11) {real, imag} */,
  {32'hbfaa2e0a, 32'hbfc28fb4} /* (23, 23, 10) {real, imag} */,
  {32'h41749e88, 32'hc09ccc58} /* (23, 23, 9) {real, imag} */,
  {32'h4075787c, 32'hc1652dac} /* (23, 23, 8) {real, imag} */,
  {32'h3f4bdd30, 32'hc008146d} /* (23, 23, 7) {real, imag} */,
  {32'h415c1db0, 32'h3fd1f408} /* (23, 23, 6) {real, imag} */,
  {32'hbfa4d36a, 32'hc16abbab} /* (23, 23, 5) {real, imag} */,
  {32'h4090384c, 32'hc14e81ca} /* (23, 23, 4) {real, imag} */,
  {32'hc1b2f509, 32'h41c0a547} /* (23, 23, 3) {real, imag} */,
  {32'h419a071a, 32'hc01d9124} /* (23, 23, 2) {real, imag} */,
  {32'h41a10013, 32'h41cba5f4} /* (23, 23, 1) {real, imag} */,
  {32'h3fbe8112, 32'h40d3e839} /* (23, 23, 0) {real, imag} */,
  {32'hc19fc695, 32'h3f745190} /* (23, 22, 31) {real, imag} */,
  {32'h3f49d92c, 32'hbf62e834} /* (23, 22, 30) {real, imag} */,
  {32'h412e8545, 32'h40e83a47} /* (23, 22, 29) {real, imag} */,
  {32'h3dfc5d00, 32'h41366238} /* (23, 22, 28) {real, imag} */,
  {32'h3fc89800, 32'hbea4ac40} /* (23, 22, 27) {real, imag} */,
  {32'hc0247d03, 32'hc16fec30} /* (23, 22, 26) {real, imag} */,
  {32'h40c5d82a, 32'hc0ea8747} /* (23, 22, 25) {real, imag} */,
  {32'hc118212b, 32'h3eb63370} /* (23, 22, 24) {real, imag} */,
  {32'h41351d48, 32'h41d2cad0} /* (23, 22, 23) {real, imag} */,
  {32'h4197c04d, 32'hc13261e2} /* (23, 22, 22) {real, imag} */,
  {32'hc11551a2, 32'hc0909df8} /* (23, 22, 21) {real, imag} */,
  {32'h4186a381, 32'h40a98d43} /* (23, 22, 20) {real, imag} */,
  {32'h406b2684, 32'hc181aac9} /* (23, 22, 19) {real, imag} */,
  {32'hc0ca4faa, 32'h3f585c40} /* (23, 22, 18) {real, imag} */,
  {32'hc060f2a2, 32'h40da4a65} /* (23, 22, 17) {real, imag} */,
  {32'hc16ccbdc, 32'h40cd517e} /* (23, 22, 16) {real, imag} */,
  {32'hbe4c13d0, 32'hc0b605a7} /* (23, 22, 15) {real, imag} */,
  {32'hc09a2e02, 32'hc0fe8862} /* (23, 22, 14) {real, imag} */,
  {32'h419ff176, 32'h412f7e65} /* (23, 22, 13) {real, imag} */,
  {32'h4004956e, 32'hbfdc7180} /* (23, 22, 12) {real, imag} */,
  {32'hc002cf88, 32'hc0e375e2} /* (23, 22, 11) {real, imag} */,
  {32'hc18efa9a, 32'h408e1bf4} /* (23, 22, 10) {real, imag} */,
  {32'hbf865ba4, 32'h40092bce} /* (23, 22, 9) {real, imag} */,
  {32'h4196431c, 32'h40f56f04} /* (23, 22, 8) {real, imag} */,
  {32'hc0380269, 32'hc1363736} /* (23, 22, 7) {real, imag} */,
  {32'h40e7568a, 32'hc0c9614d} /* (23, 22, 6) {real, imag} */,
  {32'hc18ed951, 32'hc1119af3} /* (23, 22, 5) {real, imag} */,
  {32'hc131ce43, 32'h41c25cd3} /* (23, 22, 4) {real, imag} */,
  {32'hc1b74276, 32'h41aa6572} /* (23, 22, 3) {real, imag} */,
  {32'h404528ef, 32'hc1d80256} /* (23, 22, 2) {real, imag} */,
  {32'hbd5a6a00, 32'h417a9897} /* (23, 22, 1) {real, imag} */,
  {32'h417f8c26, 32'h408da9b5} /* (23, 22, 0) {real, imag} */,
  {32'h411bcc05, 32'hc0b6a45c} /* (23, 21, 31) {real, imag} */,
  {32'hc0a13562, 32'h41064a30} /* (23, 21, 30) {real, imag} */,
  {32'hc021b0fc, 32'h4109bf44} /* (23, 21, 29) {real, imag} */,
  {32'hbf783680, 32'h4150c79f} /* (23, 21, 28) {real, imag} */,
  {32'hc1749d32, 32'h410df234} /* (23, 21, 27) {real, imag} */,
  {32'hc10801de, 32'h40bf5433} /* (23, 21, 26) {real, imag} */,
  {32'h40a73f40, 32'hc1424341} /* (23, 21, 25) {real, imag} */,
  {32'hc17fd908, 32'hc0a3317f} /* (23, 21, 24) {real, imag} */,
  {32'hc0a7df44, 32'h40b88676} /* (23, 21, 23) {real, imag} */,
  {32'hc12814f7, 32'h3e1ba020} /* (23, 21, 22) {real, imag} */,
  {32'h41a629bc, 32'hc10f51e8} /* (23, 21, 21) {real, imag} */,
  {32'h411d9f72, 32'h408c48a0} /* (23, 21, 20) {real, imag} */,
  {32'h417686ea, 32'hc0985315} /* (23, 21, 19) {real, imag} */,
  {32'hc1a46324, 32'h41b071cf} /* (23, 21, 18) {real, imag} */,
  {32'hc09d5ed1, 32'hc15d00a4} /* (23, 21, 17) {real, imag} */,
  {32'hc06dcba7, 32'h403a8d5e} /* (23, 21, 16) {real, imag} */,
  {32'hbf94be2c, 32'hbfa7a26f} /* (23, 21, 15) {real, imag} */,
  {32'hc185a0c4, 32'hc198019c} /* (23, 21, 14) {real, imag} */,
  {32'hc152d5b3, 32'hc121684a} /* (23, 21, 13) {real, imag} */,
  {32'hc0770446, 32'h40d00d26} /* (23, 21, 12) {real, imag} */,
  {32'hc116f9c2, 32'hc05746dc} /* (23, 21, 11) {real, imag} */,
  {32'h41128706, 32'h40821792} /* (23, 21, 10) {real, imag} */,
  {32'h4181ebcc, 32'h414e4f21} /* (23, 21, 9) {real, imag} */,
  {32'hc137d229, 32'h3f556248} /* (23, 21, 8) {real, imag} */,
  {32'hc0a9b6fb, 32'h3fde8bc0} /* (23, 21, 7) {real, imag} */,
  {32'hbfc52294, 32'h41b46e8d} /* (23, 21, 6) {real, imag} */,
  {32'hc15ec663, 32'h408475e2} /* (23, 21, 5) {real, imag} */,
  {32'h40508d85, 32'h4112469a} /* (23, 21, 4) {real, imag} */,
  {32'hc0d1b5aa, 32'hc1381fb4} /* (23, 21, 3) {real, imag} */,
  {32'hc087d698, 32'h41367c3a} /* (23, 21, 2) {real, imag} */,
  {32'h41954da5, 32'hc1bc4463} /* (23, 21, 1) {real, imag} */,
  {32'h40503828, 32'hc123d91e} /* (23, 21, 0) {real, imag} */,
  {32'hc0ed7d63, 32'hc0e15068} /* (23, 20, 31) {real, imag} */,
  {32'hc0912fae, 32'hc022d708} /* (23, 20, 30) {real, imag} */,
  {32'hc06abfcc, 32'h4112214f} /* (23, 20, 29) {real, imag} */,
  {32'h40f0ad78, 32'hbf570f3c} /* (23, 20, 28) {real, imag} */,
  {32'hc18bd314, 32'hc03435c0} /* (23, 20, 27) {real, imag} */,
  {32'hc0df2638, 32'hbfd44f78} /* (23, 20, 26) {real, imag} */,
  {32'h410c3f7c, 32'h40604710} /* (23, 20, 25) {real, imag} */,
  {32'h415e61be, 32'h419f1f38} /* (23, 20, 24) {real, imag} */,
  {32'hc1464232, 32'hc0082819} /* (23, 20, 23) {real, imag} */,
  {32'h40d2286a, 32'h4086b5f2} /* (23, 20, 22) {real, imag} */,
  {32'hbe4299d8, 32'hc19a112d} /* (23, 20, 21) {real, imag} */,
  {32'hc04cac5a, 32'hc130dbf5} /* (23, 20, 20) {real, imag} */,
  {32'hc10b13a8, 32'hc1093162} /* (23, 20, 19) {real, imag} */,
  {32'h3f06de9c, 32'hc11d5994} /* (23, 20, 18) {real, imag} */,
  {32'hc105fefd, 32'hc0e0b11c} /* (23, 20, 17) {real, imag} */,
  {32'h40365234, 32'h40eed2a4} /* (23, 20, 16) {real, imag} */,
  {32'hbfa319ae, 32'h40cbf318} /* (23, 20, 15) {real, imag} */,
  {32'hbf250280, 32'h4113ba91} /* (23, 20, 14) {real, imag} */,
  {32'h40cb35d0, 32'hc115cff6} /* (23, 20, 13) {real, imag} */,
  {32'hc16d116e, 32'hc13be564} /* (23, 20, 12) {real, imag} */,
  {32'hc19edfd8, 32'hc13581f4} /* (23, 20, 11) {real, imag} */,
  {32'hc12e0e46, 32'h413c00e9} /* (23, 20, 10) {real, imag} */,
  {32'h40d1b3c3, 32'hc0b2b777} /* (23, 20, 9) {real, imag} */,
  {32'hc18c1934, 32'h41304854} /* (23, 20, 8) {real, imag} */,
  {32'hbf77ee30, 32'hc087bc00} /* (23, 20, 7) {real, imag} */,
  {32'h41520aa8, 32'h3f230a9c} /* (23, 20, 6) {real, imag} */,
  {32'h3fd02188, 32'h41eadbe4} /* (23, 20, 5) {real, imag} */,
  {32'hc05888d1, 32'hc1113f30} /* (23, 20, 4) {real, imag} */,
  {32'h40efaa7a, 32'hc04229b1} /* (23, 20, 3) {real, imag} */,
  {32'hc00db6be, 32'h40466e59} /* (23, 20, 2) {real, imag} */,
  {32'hc18ed755, 32'h41039ec7} /* (23, 20, 1) {real, imag} */,
  {32'h3fc0d6f8, 32'h41a40fbd} /* (23, 20, 0) {real, imag} */,
  {32'h411b5912, 32'hc1266dfc} /* (23, 19, 31) {real, imag} */,
  {32'h40f05f88, 32'hc1b22541} /* (23, 19, 30) {real, imag} */,
  {32'hc0c53d6a, 32'hc0ca8099} /* (23, 19, 29) {real, imag} */,
  {32'h3f3ee2be, 32'hc10de438} /* (23, 19, 28) {real, imag} */,
  {32'h402fe6c2, 32'h3f5767cc} /* (23, 19, 27) {real, imag} */,
  {32'h3f32712e, 32'h40bdc21c} /* (23, 19, 26) {real, imag} */,
  {32'hc1747bac, 32'hc0f32a11} /* (23, 19, 25) {real, imag} */,
  {32'h3eb933d0, 32'h3dbb0000} /* (23, 19, 24) {real, imag} */,
  {32'hc0c0e140, 32'h4147743c} /* (23, 19, 23) {real, imag} */,
  {32'h40fc0caf, 32'hc1227a52} /* (23, 19, 22) {real, imag} */,
  {32'hc0f74a92, 32'hbfdd8e6a} /* (23, 19, 21) {real, imag} */,
  {32'h415c92d4, 32'hbf1fb838} /* (23, 19, 20) {real, imag} */,
  {32'hc02eab08, 32'h40e8d470} /* (23, 19, 19) {real, imag} */,
  {32'hbfb72488, 32'h4106d63b} /* (23, 19, 18) {real, imag} */,
  {32'hbfa90e36, 32'hc0ad8f02} /* (23, 19, 17) {real, imag} */,
  {32'h40bb5e0d, 32'hc0a65a76} /* (23, 19, 16) {real, imag} */,
  {32'hc01611eb, 32'hc02e3254} /* (23, 19, 15) {real, imag} */,
  {32'hc117e093, 32'hc0a941d2} /* (23, 19, 14) {real, imag} */,
  {32'hc0f9cc84, 32'hbef7ba78} /* (23, 19, 13) {real, imag} */,
  {32'h414e3db2, 32'hc11f7e3a} /* (23, 19, 12) {real, imag} */,
  {32'hc16262cf, 32'h4187098a} /* (23, 19, 11) {real, imag} */,
  {32'h400b25b8, 32'h40ca0a27} /* (23, 19, 10) {real, imag} */,
  {32'h418e5b4e, 32'hc0fd20e2} /* (23, 19, 9) {real, imag} */,
  {32'h3f969b5d, 32'hc00453f1} /* (23, 19, 8) {real, imag} */,
  {32'h40a24622, 32'hc1352820} /* (23, 19, 7) {real, imag} */,
  {32'h4142abae, 32'h417fef97} /* (23, 19, 6) {real, imag} */,
  {32'h41972d9b, 32'hc1080e04} /* (23, 19, 5) {real, imag} */,
  {32'h412ea246, 32'h3f6833f4} /* (23, 19, 4) {real, imag} */,
  {32'h40b95e8d, 32'h40b5e2c3} /* (23, 19, 3) {real, imag} */,
  {32'hc1ce7c2c, 32'hbfd16718} /* (23, 19, 2) {real, imag} */,
  {32'h40ea26fc, 32'hc13d4e17} /* (23, 19, 1) {real, imag} */,
  {32'hc0d37e0a, 32'h41670947} /* (23, 19, 0) {real, imag} */,
  {32'hc08b98d2, 32'hc120d4e4} /* (23, 18, 31) {real, imag} */,
  {32'hbf630540, 32'h4128b452} /* (23, 18, 30) {real, imag} */,
  {32'hbe7b7ff0, 32'h3ef27740} /* (23, 18, 29) {real, imag} */,
  {32'h40579092, 32'hc01cfe96} /* (23, 18, 28) {real, imag} */,
  {32'hc08510b3, 32'h414f0666} /* (23, 18, 27) {real, imag} */,
  {32'h413379a0, 32'h406b35fe} /* (23, 18, 26) {real, imag} */,
  {32'h40cb054c, 32'hc1127deb} /* (23, 18, 25) {real, imag} */,
  {32'hc09c417e, 32'h4103bfaa} /* (23, 18, 24) {real, imag} */,
  {32'hc01deeff, 32'hc02b4268} /* (23, 18, 23) {real, imag} */,
  {32'h412488a7, 32'h41216c4a} /* (23, 18, 22) {real, imag} */,
  {32'h411351dc, 32'hc089c932} /* (23, 18, 21) {real, imag} */,
  {32'hbfcb00c2, 32'hbe1001d8} /* (23, 18, 20) {real, imag} */,
  {32'h41319ea8, 32'h4157ce84} /* (23, 18, 19) {real, imag} */,
  {32'hc1324eb7, 32'hc0a3b68e} /* (23, 18, 18) {real, imag} */,
  {32'hc1143a89, 32'h4130bf8e} /* (23, 18, 17) {real, imag} */,
  {32'hc0b22127, 32'h40b0743b} /* (23, 18, 16) {real, imag} */,
  {32'h40ed2533, 32'hbf95cce8} /* (23, 18, 15) {real, imag} */,
  {32'h41245ecd, 32'h40765cb0} /* (23, 18, 14) {real, imag} */,
  {32'hc1120387, 32'h40f2f14b} /* (23, 18, 13) {real, imag} */,
  {32'h4108e2c9, 32'hc11304ad} /* (23, 18, 12) {real, imag} */,
  {32'hc178b687, 32'hc0992e73} /* (23, 18, 11) {real, imag} */,
  {32'hc0b6d886, 32'hc1a1a630} /* (23, 18, 10) {real, imag} */,
  {32'h41186e84, 32'hc104b105} /* (23, 18, 9) {real, imag} */,
  {32'h4038c3dc, 32'h3ff60cfa} /* (23, 18, 8) {real, imag} */,
  {32'h4101a9e6, 32'hc006ff0e} /* (23, 18, 7) {real, imag} */,
  {32'hc17be4ec, 32'hc061bb52} /* (23, 18, 6) {real, imag} */,
  {32'h3f3090a0, 32'hbe97b1c0} /* (23, 18, 5) {real, imag} */,
  {32'h40132bd4, 32'h40ba927f} /* (23, 18, 4) {real, imag} */,
  {32'h3f757172, 32'h3f8a25b4} /* (23, 18, 3) {real, imag} */,
  {32'h40b4f5e6, 32'hc08eb254} /* (23, 18, 2) {real, imag} */,
  {32'h40bad86f, 32'hc1822e1e} /* (23, 18, 1) {real, imag} */,
  {32'hc0cd8886, 32'hc08b148e} /* (23, 18, 0) {real, imag} */,
  {32'h40eab760, 32'h40da3be8} /* (23, 17, 31) {real, imag} */,
  {32'h411efce7, 32'hc0e92ebc} /* (23, 17, 30) {real, imag} */,
  {32'hc0f2e244, 32'hc0cc8a80} /* (23, 17, 29) {real, imag} */,
  {32'h3fb4be6c, 32'hc0dd1c41} /* (23, 17, 28) {real, imag} */,
  {32'h400c6cb3, 32'hc1487ca6} /* (23, 17, 27) {real, imag} */,
  {32'h41b947fd, 32'h3fd7bc60} /* (23, 17, 26) {real, imag} */,
  {32'h3f3cbeb0, 32'hc032224c} /* (23, 17, 25) {real, imag} */,
  {32'hc0095e00, 32'hc0ebd61a} /* (23, 17, 24) {real, imag} */,
  {32'h4094cfb4, 32'h4143ee50} /* (23, 17, 23) {real, imag} */,
  {32'hc0f5f204, 32'hc0967312} /* (23, 17, 22) {real, imag} */,
  {32'hc114d7e4, 32'h3fffff34} /* (23, 17, 21) {real, imag} */,
  {32'hc113adf6, 32'h410b053e} /* (23, 17, 20) {real, imag} */,
  {32'hc15bc0d9, 32'hbf8dee46} /* (23, 17, 19) {real, imag} */,
  {32'h40692bb7, 32'h402e3c02} /* (23, 17, 18) {real, imag} */,
  {32'h40c5c55f, 32'h4017ffad} /* (23, 17, 17) {real, imag} */,
  {32'h3fa65b1a, 32'hc0447d06} /* (23, 17, 16) {real, imag} */,
  {32'hc04299e3, 32'h3fa4a818} /* (23, 17, 15) {real, imag} */,
  {32'h41549fc6, 32'h40c6df48} /* (23, 17, 14) {real, imag} */,
  {32'hc1114fbd, 32'hc051cbe9} /* (23, 17, 13) {real, imag} */,
  {32'h4104eb9b, 32'hc0fd426b} /* (23, 17, 12) {real, imag} */,
  {32'h4091b278, 32'h40b16cbd} /* (23, 17, 11) {real, imag} */,
  {32'h41385939, 32'hbffd8700} /* (23, 17, 10) {real, imag} */,
  {32'hc0df5f71, 32'h418e477a} /* (23, 17, 9) {real, imag} */,
  {32'hc1275328, 32'h40bab348} /* (23, 17, 8) {real, imag} */,
  {32'h413b9648, 32'hc084a71e} /* (23, 17, 7) {real, imag} */,
  {32'hbf8d911c, 32'h40064c8e} /* (23, 17, 6) {real, imag} */,
  {32'h402d8f47, 32'hc103e321} /* (23, 17, 5) {real, imag} */,
  {32'hc0f6ad3a, 32'hbf6dacda} /* (23, 17, 4) {real, imag} */,
  {32'hc12f631d, 32'hc0a1e4dc} /* (23, 17, 3) {real, imag} */,
  {32'h4159de60, 32'hc13c52d5} /* (23, 17, 2) {real, imag} */,
  {32'hbfb34d9c, 32'h414d2207} /* (23, 17, 1) {real, imag} */,
  {32'hc198aa52, 32'h410d3607} /* (23, 17, 0) {real, imag} */,
  {32'h4092e74a, 32'h413f1b57} /* (23, 16, 31) {real, imag} */,
  {32'hc00ea486, 32'hc125a2ab} /* (23, 16, 30) {real, imag} */,
  {32'h40b565a6, 32'h3ff079c7} /* (23, 16, 29) {real, imag} */,
  {32'h4082fe6e, 32'h401b0f1e} /* (23, 16, 28) {real, imag} */,
  {32'hc089acdb, 32'hc0a718b0} /* (23, 16, 27) {real, imag} */,
  {32'h3f8e4a22, 32'hc10e3582} /* (23, 16, 26) {real, imag} */,
  {32'hc13da1bb, 32'h40d075bd} /* (23, 16, 25) {real, imag} */,
  {32'h3f09fa46, 32'h41555777} /* (23, 16, 24) {real, imag} */,
  {32'hc0ebe3ea, 32'h409c8bf6} /* (23, 16, 23) {real, imag} */,
  {32'hbe5b23c0, 32'hc07c8240} /* (23, 16, 22) {real, imag} */,
  {32'hc1306a22, 32'h410fd13c} /* (23, 16, 21) {real, imag} */,
  {32'hc07f98e8, 32'hc138a13c} /* (23, 16, 20) {real, imag} */,
  {32'h414548ce, 32'h41853cce} /* (23, 16, 19) {real, imag} */,
  {32'h410f0366, 32'h400dc819} /* (23, 16, 18) {real, imag} */,
  {32'hbf9aa0a3, 32'hc0a511e0} /* (23, 16, 17) {real, imag} */,
  {32'h41860335, 32'h00000000} /* (23, 16, 16) {real, imag} */,
  {32'hbf9aa0a3, 32'h40a511e0} /* (23, 16, 15) {real, imag} */,
  {32'h410f0366, 32'hc00dc819} /* (23, 16, 14) {real, imag} */,
  {32'h414548ce, 32'hc1853cce} /* (23, 16, 13) {real, imag} */,
  {32'hc07f98e8, 32'h4138a13c} /* (23, 16, 12) {real, imag} */,
  {32'hc1306a22, 32'hc10fd13c} /* (23, 16, 11) {real, imag} */,
  {32'hbe5b23c0, 32'h407c8240} /* (23, 16, 10) {real, imag} */,
  {32'hc0ebe3ea, 32'hc09c8bf6} /* (23, 16, 9) {real, imag} */,
  {32'h3f09fa46, 32'hc1555777} /* (23, 16, 8) {real, imag} */,
  {32'hc13da1bb, 32'hc0d075bd} /* (23, 16, 7) {real, imag} */,
  {32'h3f8e4a22, 32'h410e3582} /* (23, 16, 6) {real, imag} */,
  {32'hc089acdb, 32'h40a718b0} /* (23, 16, 5) {real, imag} */,
  {32'h4082fe6e, 32'hc01b0f1e} /* (23, 16, 4) {real, imag} */,
  {32'h40b565a6, 32'hbff079c7} /* (23, 16, 3) {real, imag} */,
  {32'hc00ea486, 32'h4125a2ab} /* (23, 16, 2) {real, imag} */,
  {32'h4092e74a, 32'hc13f1b57} /* (23, 16, 1) {real, imag} */,
  {32'h410a6e47, 32'h00000000} /* (23, 16, 0) {real, imag} */,
  {32'hbfb34d9c, 32'hc14d2207} /* (23, 15, 31) {real, imag} */,
  {32'h4159de60, 32'h413c52d5} /* (23, 15, 30) {real, imag} */,
  {32'hc12f631d, 32'h40a1e4dc} /* (23, 15, 29) {real, imag} */,
  {32'hc0f6ad3a, 32'h3f6dacda} /* (23, 15, 28) {real, imag} */,
  {32'h402d8f47, 32'h4103e321} /* (23, 15, 27) {real, imag} */,
  {32'hbf8d911c, 32'hc0064c8e} /* (23, 15, 26) {real, imag} */,
  {32'h413b9648, 32'h4084a71e} /* (23, 15, 25) {real, imag} */,
  {32'hc1275328, 32'hc0bab348} /* (23, 15, 24) {real, imag} */,
  {32'hc0df5f71, 32'hc18e477a} /* (23, 15, 23) {real, imag} */,
  {32'h41385939, 32'h3ffd8700} /* (23, 15, 22) {real, imag} */,
  {32'h4091b278, 32'hc0b16cbd} /* (23, 15, 21) {real, imag} */,
  {32'h4104eb9b, 32'h40fd426b} /* (23, 15, 20) {real, imag} */,
  {32'hc1114fbd, 32'h4051cbe9} /* (23, 15, 19) {real, imag} */,
  {32'h41549fc6, 32'hc0c6df48} /* (23, 15, 18) {real, imag} */,
  {32'hc04299e3, 32'hbfa4a818} /* (23, 15, 17) {real, imag} */,
  {32'h3fa65b1a, 32'h40447d06} /* (23, 15, 16) {real, imag} */,
  {32'h40c5c55f, 32'hc017ffad} /* (23, 15, 15) {real, imag} */,
  {32'h40692bb7, 32'hc02e3c02} /* (23, 15, 14) {real, imag} */,
  {32'hc15bc0d9, 32'h3f8dee46} /* (23, 15, 13) {real, imag} */,
  {32'hc113adf6, 32'hc10b053e} /* (23, 15, 12) {real, imag} */,
  {32'hc114d7e4, 32'hbfffff34} /* (23, 15, 11) {real, imag} */,
  {32'hc0f5f204, 32'h40967312} /* (23, 15, 10) {real, imag} */,
  {32'h4094cfb4, 32'hc143ee50} /* (23, 15, 9) {real, imag} */,
  {32'hc0095e00, 32'h40ebd61a} /* (23, 15, 8) {real, imag} */,
  {32'h3f3cbeb0, 32'h4032224c} /* (23, 15, 7) {real, imag} */,
  {32'h41b947fd, 32'hbfd7bc60} /* (23, 15, 6) {real, imag} */,
  {32'h400c6cb3, 32'h41487ca6} /* (23, 15, 5) {real, imag} */,
  {32'h3fb4be6c, 32'h40dd1c41} /* (23, 15, 4) {real, imag} */,
  {32'hc0f2e244, 32'h40cc8a80} /* (23, 15, 3) {real, imag} */,
  {32'h411efce7, 32'h40e92ebc} /* (23, 15, 2) {real, imag} */,
  {32'h40eab760, 32'hc0da3be8} /* (23, 15, 1) {real, imag} */,
  {32'hc198aa52, 32'hc10d3607} /* (23, 15, 0) {real, imag} */,
  {32'h40bad86f, 32'h41822e1e} /* (23, 14, 31) {real, imag} */,
  {32'h40b4f5e6, 32'h408eb254} /* (23, 14, 30) {real, imag} */,
  {32'h3f757172, 32'hbf8a25b4} /* (23, 14, 29) {real, imag} */,
  {32'h40132bd4, 32'hc0ba927f} /* (23, 14, 28) {real, imag} */,
  {32'h3f3090a0, 32'h3e97b1c0} /* (23, 14, 27) {real, imag} */,
  {32'hc17be4ec, 32'h4061bb52} /* (23, 14, 26) {real, imag} */,
  {32'h4101a9e6, 32'h4006ff0e} /* (23, 14, 25) {real, imag} */,
  {32'h4038c3dc, 32'hbff60cfa} /* (23, 14, 24) {real, imag} */,
  {32'h41186e84, 32'h4104b105} /* (23, 14, 23) {real, imag} */,
  {32'hc0b6d886, 32'h41a1a630} /* (23, 14, 22) {real, imag} */,
  {32'hc178b687, 32'h40992e73} /* (23, 14, 21) {real, imag} */,
  {32'h4108e2c9, 32'h411304ad} /* (23, 14, 20) {real, imag} */,
  {32'hc1120387, 32'hc0f2f14b} /* (23, 14, 19) {real, imag} */,
  {32'h41245ecd, 32'hc0765cb0} /* (23, 14, 18) {real, imag} */,
  {32'h40ed2533, 32'h3f95cce8} /* (23, 14, 17) {real, imag} */,
  {32'hc0b22127, 32'hc0b0743b} /* (23, 14, 16) {real, imag} */,
  {32'hc1143a89, 32'hc130bf8e} /* (23, 14, 15) {real, imag} */,
  {32'hc1324eb7, 32'h40a3b68e} /* (23, 14, 14) {real, imag} */,
  {32'h41319ea8, 32'hc157ce84} /* (23, 14, 13) {real, imag} */,
  {32'hbfcb00c2, 32'h3e1001d8} /* (23, 14, 12) {real, imag} */,
  {32'h411351dc, 32'h4089c932} /* (23, 14, 11) {real, imag} */,
  {32'h412488a7, 32'hc1216c4a} /* (23, 14, 10) {real, imag} */,
  {32'hc01deeff, 32'h402b4268} /* (23, 14, 9) {real, imag} */,
  {32'hc09c417e, 32'hc103bfaa} /* (23, 14, 8) {real, imag} */,
  {32'h40cb054c, 32'h41127deb} /* (23, 14, 7) {real, imag} */,
  {32'h413379a0, 32'hc06b35fe} /* (23, 14, 6) {real, imag} */,
  {32'hc08510b3, 32'hc14f0666} /* (23, 14, 5) {real, imag} */,
  {32'h40579092, 32'h401cfe96} /* (23, 14, 4) {real, imag} */,
  {32'hbe7b7ff0, 32'hbef27740} /* (23, 14, 3) {real, imag} */,
  {32'hbf630540, 32'hc128b452} /* (23, 14, 2) {real, imag} */,
  {32'hc08b98d2, 32'h4120d4e4} /* (23, 14, 1) {real, imag} */,
  {32'hc0cd8886, 32'h408b148e} /* (23, 14, 0) {real, imag} */,
  {32'h40ea26fc, 32'h413d4e17} /* (23, 13, 31) {real, imag} */,
  {32'hc1ce7c2c, 32'h3fd16718} /* (23, 13, 30) {real, imag} */,
  {32'h40b95e8d, 32'hc0b5e2c3} /* (23, 13, 29) {real, imag} */,
  {32'h412ea246, 32'hbf6833f4} /* (23, 13, 28) {real, imag} */,
  {32'h41972d9b, 32'h41080e04} /* (23, 13, 27) {real, imag} */,
  {32'h4142abae, 32'hc17fef97} /* (23, 13, 26) {real, imag} */,
  {32'h40a24622, 32'h41352820} /* (23, 13, 25) {real, imag} */,
  {32'h3f969b5d, 32'h400453f1} /* (23, 13, 24) {real, imag} */,
  {32'h418e5b4e, 32'h40fd20e2} /* (23, 13, 23) {real, imag} */,
  {32'h400b25b8, 32'hc0ca0a27} /* (23, 13, 22) {real, imag} */,
  {32'hc16262cf, 32'hc187098a} /* (23, 13, 21) {real, imag} */,
  {32'h414e3db2, 32'h411f7e3a} /* (23, 13, 20) {real, imag} */,
  {32'hc0f9cc84, 32'h3ef7ba78} /* (23, 13, 19) {real, imag} */,
  {32'hc117e093, 32'h40a941d2} /* (23, 13, 18) {real, imag} */,
  {32'hc01611eb, 32'h402e3254} /* (23, 13, 17) {real, imag} */,
  {32'h40bb5e0d, 32'h40a65a76} /* (23, 13, 16) {real, imag} */,
  {32'hbfa90e36, 32'h40ad8f02} /* (23, 13, 15) {real, imag} */,
  {32'hbfb72488, 32'hc106d63b} /* (23, 13, 14) {real, imag} */,
  {32'hc02eab08, 32'hc0e8d470} /* (23, 13, 13) {real, imag} */,
  {32'h415c92d4, 32'h3f1fb838} /* (23, 13, 12) {real, imag} */,
  {32'hc0f74a92, 32'h3fdd8e6a} /* (23, 13, 11) {real, imag} */,
  {32'h40fc0caf, 32'h41227a52} /* (23, 13, 10) {real, imag} */,
  {32'hc0c0e140, 32'hc147743c} /* (23, 13, 9) {real, imag} */,
  {32'h3eb933d0, 32'hbdbb0000} /* (23, 13, 8) {real, imag} */,
  {32'hc1747bac, 32'h40f32a11} /* (23, 13, 7) {real, imag} */,
  {32'h3f32712e, 32'hc0bdc21c} /* (23, 13, 6) {real, imag} */,
  {32'h402fe6c2, 32'hbf5767cc} /* (23, 13, 5) {real, imag} */,
  {32'h3f3ee2be, 32'h410de438} /* (23, 13, 4) {real, imag} */,
  {32'hc0c53d6a, 32'h40ca8099} /* (23, 13, 3) {real, imag} */,
  {32'h40f05f88, 32'h41b22541} /* (23, 13, 2) {real, imag} */,
  {32'h411b5912, 32'h41266dfc} /* (23, 13, 1) {real, imag} */,
  {32'hc0d37e0a, 32'hc1670947} /* (23, 13, 0) {real, imag} */,
  {32'hc18ed755, 32'hc1039ec7} /* (23, 12, 31) {real, imag} */,
  {32'hc00db6be, 32'hc0466e59} /* (23, 12, 30) {real, imag} */,
  {32'h40efaa7a, 32'h404229b1} /* (23, 12, 29) {real, imag} */,
  {32'hc05888d1, 32'h41113f30} /* (23, 12, 28) {real, imag} */,
  {32'h3fd02188, 32'hc1eadbe4} /* (23, 12, 27) {real, imag} */,
  {32'h41520aa8, 32'hbf230a9c} /* (23, 12, 26) {real, imag} */,
  {32'hbf77ee30, 32'h4087bc00} /* (23, 12, 25) {real, imag} */,
  {32'hc18c1934, 32'hc1304854} /* (23, 12, 24) {real, imag} */,
  {32'h40d1b3c3, 32'h40b2b777} /* (23, 12, 23) {real, imag} */,
  {32'hc12e0e46, 32'hc13c00e9} /* (23, 12, 22) {real, imag} */,
  {32'hc19edfd8, 32'h413581f4} /* (23, 12, 21) {real, imag} */,
  {32'hc16d116e, 32'h413be564} /* (23, 12, 20) {real, imag} */,
  {32'h40cb35d0, 32'h4115cff6} /* (23, 12, 19) {real, imag} */,
  {32'hbf250280, 32'hc113ba91} /* (23, 12, 18) {real, imag} */,
  {32'hbfa319ae, 32'hc0cbf318} /* (23, 12, 17) {real, imag} */,
  {32'h40365234, 32'hc0eed2a4} /* (23, 12, 16) {real, imag} */,
  {32'hc105fefd, 32'h40e0b11c} /* (23, 12, 15) {real, imag} */,
  {32'h3f06de9c, 32'h411d5994} /* (23, 12, 14) {real, imag} */,
  {32'hc10b13a8, 32'h41093162} /* (23, 12, 13) {real, imag} */,
  {32'hc04cac5a, 32'h4130dbf5} /* (23, 12, 12) {real, imag} */,
  {32'hbe4299d8, 32'h419a112d} /* (23, 12, 11) {real, imag} */,
  {32'h40d2286a, 32'hc086b5f2} /* (23, 12, 10) {real, imag} */,
  {32'hc1464232, 32'h40082819} /* (23, 12, 9) {real, imag} */,
  {32'h415e61be, 32'hc19f1f38} /* (23, 12, 8) {real, imag} */,
  {32'h410c3f7c, 32'hc0604710} /* (23, 12, 7) {real, imag} */,
  {32'hc0df2638, 32'h3fd44f78} /* (23, 12, 6) {real, imag} */,
  {32'hc18bd314, 32'h403435c0} /* (23, 12, 5) {real, imag} */,
  {32'h40f0ad78, 32'h3f570f3c} /* (23, 12, 4) {real, imag} */,
  {32'hc06abfcc, 32'hc112214f} /* (23, 12, 3) {real, imag} */,
  {32'hc0912fae, 32'h4022d708} /* (23, 12, 2) {real, imag} */,
  {32'hc0ed7d63, 32'h40e15068} /* (23, 12, 1) {real, imag} */,
  {32'h3fc0d6f8, 32'hc1a40fbd} /* (23, 12, 0) {real, imag} */,
  {32'h41954da5, 32'h41bc4463} /* (23, 11, 31) {real, imag} */,
  {32'hc087d698, 32'hc1367c3a} /* (23, 11, 30) {real, imag} */,
  {32'hc0d1b5aa, 32'h41381fb4} /* (23, 11, 29) {real, imag} */,
  {32'h40508d85, 32'hc112469a} /* (23, 11, 28) {real, imag} */,
  {32'hc15ec663, 32'hc08475e2} /* (23, 11, 27) {real, imag} */,
  {32'hbfc52294, 32'hc1b46e8d} /* (23, 11, 26) {real, imag} */,
  {32'hc0a9b6fb, 32'hbfde8bc0} /* (23, 11, 25) {real, imag} */,
  {32'hc137d229, 32'hbf556248} /* (23, 11, 24) {real, imag} */,
  {32'h4181ebcc, 32'hc14e4f21} /* (23, 11, 23) {real, imag} */,
  {32'h41128706, 32'hc0821792} /* (23, 11, 22) {real, imag} */,
  {32'hc116f9c2, 32'h405746dc} /* (23, 11, 21) {real, imag} */,
  {32'hc0770446, 32'hc0d00d26} /* (23, 11, 20) {real, imag} */,
  {32'hc152d5b3, 32'h4121684a} /* (23, 11, 19) {real, imag} */,
  {32'hc185a0c4, 32'h4198019c} /* (23, 11, 18) {real, imag} */,
  {32'hbf94be2c, 32'h3fa7a26f} /* (23, 11, 17) {real, imag} */,
  {32'hc06dcba7, 32'hc03a8d5e} /* (23, 11, 16) {real, imag} */,
  {32'hc09d5ed1, 32'h415d00a4} /* (23, 11, 15) {real, imag} */,
  {32'hc1a46324, 32'hc1b071cf} /* (23, 11, 14) {real, imag} */,
  {32'h417686ea, 32'h40985315} /* (23, 11, 13) {real, imag} */,
  {32'h411d9f72, 32'hc08c48a0} /* (23, 11, 12) {real, imag} */,
  {32'h41a629bc, 32'h410f51e8} /* (23, 11, 11) {real, imag} */,
  {32'hc12814f7, 32'hbe1ba020} /* (23, 11, 10) {real, imag} */,
  {32'hc0a7df44, 32'hc0b88676} /* (23, 11, 9) {real, imag} */,
  {32'hc17fd908, 32'h40a3317f} /* (23, 11, 8) {real, imag} */,
  {32'h40a73f40, 32'h41424341} /* (23, 11, 7) {real, imag} */,
  {32'hc10801de, 32'hc0bf5433} /* (23, 11, 6) {real, imag} */,
  {32'hc1749d32, 32'hc10df234} /* (23, 11, 5) {real, imag} */,
  {32'hbf783680, 32'hc150c79f} /* (23, 11, 4) {real, imag} */,
  {32'hc021b0fc, 32'hc109bf44} /* (23, 11, 3) {real, imag} */,
  {32'hc0a13562, 32'hc1064a30} /* (23, 11, 2) {real, imag} */,
  {32'h411bcc05, 32'h40b6a45c} /* (23, 11, 1) {real, imag} */,
  {32'h40503828, 32'h4123d91e} /* (23, 11, 0) {real, imag} */,
  {32'hbd5a6a00, 32'hc17a9897} /* (23, 10, 31) {real, imag} */,
  {32'h404528ef, 32'h41d80256} /* (23, 10, 30) {real, imag} */,
  {32'hc1b74276, 32'hc1aa6572} /* (23, 10, 29) {real, imag} */,
  {32'hc131ce43, 32'hc1c25cd3} /* (23, 10, 28) {real, imag} */,
  {32'hc18ed951, 32'h41119af3} /* (23, 10, 27) {real, imag} */,
  {32'h40e7568a, 32'h40c9614d} /* (23, 10, 26) {real, imag} */,
  {32'hc0380269, 32'h41363736} /* (23, 10, 25) {real, imag} */,
  {32'h4196431c, 32'hc0f56f04} /* (23, 10, 24) {real, imag} */,
  {32'hbf865ba4, 32'hc0092bce} /* (23, 10, 23) {real, imag} */,
  {32'hc18efa9a, 32'hc08e1bf4} /* (23, 10, 22) {real, imag} */,
  {32'hc002cf88, 32'h40e375e2} /* (23, 10, 21) {real, imag} */,
  {32'h4004956e, 32'h3fdc7180} /* (23, 10, 20) {real, imag} */,
  {32'h419ff176, 32'hc12f7e65} /* (23, 10, 19) {real, imag} */,
  {32'hc09a2e02, 32'h40fe8862} /* (23, 10, 18) {real, imag} */,
  {32'hbe4c13d0, 32'h40b605a7} /* (23, 10, 17) {real, imag} */,
  {32'hc16ccbdc, 32'hc0cd517e} /* (23, 10, 16) {real, imag} */,
  {32'hc060f2a2, 32'hc0da4a65} /* (23, 10, 15) {real, imag} */,
  {32'hc0ca4faa, 32'hbf585c40} /* (23, 10, 14) {real, imag} */,
  {32'h406b2684, 32'h4181aac9} /* (23, 10, 13) {real, imag} */,
  {32'h4186a381, 32'hc0a98d43} /* (23, 10, 12) {real, imag} */,
  {32'hc11551a2, 32'h40909df8} /* (23, 10, 11) {real, imag} */,
  {32'h4197c04d, 32'h413261e2} /* (23, 10, 10) {real, imag} */,
  {32'h41351d48, 32'hc1d2cad0} /* (23, 10, 9) {real, imag} */,
  {32'hc118212b, 32'hbeb63370} /* (23, 10, 8) {real, imag} */,
  {32'h40c5d82a, 32'h40ea8747} /* (23, 10, 7) {real, imag} */,
  {32'hc0247d03, 32'h416fec30} /* (23, 10, 6) {real, imag} */,
  {32'h3fc89800, 32'h3ea4ac40} /* (23, 10, 5) {real, imag} */,
  {32'h3dfc5d00, 32'hc1366238} /* (23, 10, 4) {real, imag} */,
  {32'h412e8545, 32'hc0e83a47} /* (23, 10, 3) {real, imag} */,
  {32'h3f49d92c, 32'h3f62e834} /* (23, 10, 2) {real, imag} */,
  {32'hc19fc695, 32'hbf745190} /* (23, 10, 1) {real, imag} */,
  {32'h417f8c26, 32'hc08da9b5} /* (23, 10, 0) {real, imag} */,
  {32'h41a10013, 32'hc1cba5f4} /* (23, 9, 31) {real, imag} */,
  {32'h419a071a, 32'h401d9124} /* (23, 9, 30) {real, imag} */,
  {32'hc1b2f509, 32'hc1c0a547} /* (23, 9, 29) {real, imag} */,
  {32'h4090384c, 32'h414e81ca} /* (23, 9, 28) {real, imag} */,
  {32'hbfa4d36a, 32'h416abbab} /* (23, 9, 27) {real, imag} */,
  {32'h415c1db0, 32'hbfd1f408} /* (23, 9, 26) {real, imag} */,
  {32'h3f4bdd30, 32'h4008146d} /* (23, 9, 25) {real, imag} */,
  {32'h4075787c, 32'h41652dac} /* (23, 9, 24) {real, imag} */,
  {32'h41749e88, 32'h409ccc58} /* (23, 9, 23) {real, imag} */,
  {32'hbfaa2e0a, 32'h3fc28fb4} /* (23, 9, 22) {real, imag} */,
  {32'hc0e603e4, 32'h41106264} /* (23, 9, 21) {real, imag} */,
  {32'h41598078, 32'hc11193e7} /* (23, 9, 20) {real, imag} */,
  {32'h4104e7d6, 32'hc14691ab} /* (23, 9, 19) {real, imag} */,
  {32'hc0c1c57c, 32'h4124b509} /* (23, 9, 18) {real, imag} */,
  {32'hc1158493, 32'hc0951e47} /* (23, 9, 17) {real, imag} */,
  {32'h410fe848, 32'hc0cf384c} /* (23, 9, 16) {real, imag} */,
  {32'h4116dabc, 32'hc10f19d0} /* (23, 9, 15) {real, imag} */,
  {32'h407436f0, 32'hc074dd01} /* (23, 9, 14) {real, imag} */,
  {32'h40d3b34e, 32'hc0ca94c4} /* (23, 9, 13) {real, imag} */,
  {32'h41744ef3, 32'h416cb563} /* (23, 9, 12) {real, imag} */,
  {32'hc0b9bf76, 32'hc08da08b} /* (23, 9, 11) {real, imag} */,
  {32'h41d0fd49, 32'hbfda12e8} /* (23, 9, 10) {real, imag} */,
  {32'hc0cc66d6, 32'h4141e3a6} /* (23, 9, 9) {real, imag} */,
  {32'h41b163be, 32'h418497e0} /* (23, 9, 8) {real, imag} */,
  {32'h40bdd510, 32'h411b9214} /* (23, 9, 7) {real, imag} */,
  {32'h404f040f, 32'hc0817a2d} /* (23, 9, 6) {real, imag} */,
  {32'hc188db91, 32'h40445ba8} /* (23, 9, 5) {real, imag} */,
  {32'hbf5e0670, 32'h410e6080} /* (23, 9, 4) {real, imag} */,
  {32'hc05f7302, 32'h403c2280} /* (23, 9, 3) {real, imag} */,
  {32'hc18c1a68, 32'hc0021c94} /* (23, 9, 2) {real, imag} */,
  {32'hc1de8423, 32'hc1a44a91} /* (23, 9, 1) {real, imag} */,
  {32'h3fbe8112, 32'hc0d3e839} /* (23, 9, 0) {real, imag} */,
  {32'h424aaac8, 32'h418862db} /* (23, 8, 31) {real, imag} */,
  {32'hc1a8028d, 32'hc09ca0f0} /* (23, 8, 30) {real, imag} */,
  {32'h4046c4c9, 32'h40cd7145} /* (23, 8, 29) {real, imag} */,
  {32'h40d534c3, 32'hc16b2516} /* (23, 8, 28) {real, imag} */,
  {32'hc142072e, 32'h4133d818} /* (23, 8, 27) {real, imag} */,
  {32'h40b9efba, 32'hc0cb6392} /* (23, 8, 26) {real, imag} */,
  {32'h40f7a234, 32'hc18a31ef} /* (23, 8, 25) {real, imag} */,
  {32'hc187091e, 32'h4040aa8c} /* (23, 8, 24) {real, imag} */,
  {32'hc08f55d2, 32'h413d71e5} /* (23, 8, 23) {real, imag} */,
  {32'h40c2664c, 32'hc153b718} /* (23, 8, 22) {real, imag} */,
  {32'h41264767, 32'hc0dfe905} /* (23, 8, 21) {real, imag} */,
  {32'hc0d312e0, 32'hc0973606} /* (23, 8, 20) {real, imag} */,
  {32'h410944f9, 32'h4096ae51} /* (23, 8, 19) {real, imag} */,
  {32'hc064c3f6, 32'h403825d6} /* (23, 8, 18) {real, imag} */,
  {32'h403065b1, 32'hc0d16526} /* (23, 8, 17) {real, imag} */,
  {32'h4111cdc1, 32'hc0e58322} /* (23, 8, 16) {real, imag} */,
  {32'h40646d53, 32'h4086d88c} /* (23, 8, 15) {real, imag} */,
  {32'hbfc9f93c, 32'hc10ae0e8} /* (23, 8, 14) {real, imag} */,
  {32'hc16d2f37, 32'h41447da2} /* (23, 8, 13) {real, imag} */,
  {32'hc1414446, 32'h40702e25} /* (23, 8, 12) {real, imag} */,
  {32'h410c3290, 32'hc128ac84} /* (23, 8, 11) {real, imag} */,
  {32'h41c740e4, 32'h4155221a} /* (23, 8, 10) {real, imag} */,
  {32'hbfda6674, 32'hc12c4477} /* (23, 8, 9) {real, imag} */,
  {32'hc175b386, 32'hc12563c2} /* (23, 8, 8) {real, imag} */,
  {32'h420d0358, 32'hc09775a0} /* (23, 8, 7) {real, imag} */,
  {32'h3f175200, 32'h4183ea75} /* (23, 8, 6) {real, imag} */,
  {32'hc0f0d0f6, 32'hc20079c3} /* (23, 8, 5) {real, imag} */,
  {32'h40b057c6, 32'h4091b212} /* (23, 8, 4) {real, imag} */,
  {32'h40eb53a0, 32'hc193cd37} /* (23, 8, 3) {real, imag} */,
  {32'hc18ff9e0, 32'hc0a7689c} /* (23, 8, 2) {real, imag} */,
  {32'h4003f8d6, 32'h419e10c6} /* (23, 8, 1) {real, imag} */,
  {32'h40ff9ee4, 32'h41a6abbc} /* (23, 8, 0) {real, imag} */,
  {32'hc211e3b0, 32'hc1149aa7} /* (23, 7, 31) {real, imag} */,
  {32'hc0ed11b6, 32'h4133f151} /* (23, 7, 30) {real, imag} */,
  {32'h41301304, 32'h415be9bf} /* (23, 7, 29) {real, imag} */,
  {32'h418a148e, 32'hbfef9068} /* (23, 7, 28) {real, imag} */,
  {32'hc1b08a3a, 32'h4059bd1e} /* (23, 7, 27) {real, imag} */,
  {32'hc0a6fd25, 32'h41cdb741} /* (23, 7, 26) {real, imag} */,
  {32'hc13d1f38, 32'h3ffc6c08} /* (23, 7, 25) {real, imag} */,
  {32'h416f2485, 32'h4134965f} /* (23, 7, 24) {real, imag} */,
  {32'h4115f174, 32'h4070079c} /* (23, 7, 23) {real, imag} */,
  {32'h41011315, 32'h404a9ef2} /* (23, 7, 22) {real, imag} */,
  {32'hc002eabe, 32'h3faed48a} /* (23, 7, 21) {real, imag} */,
  {32'h41284ace, 32'hc14451a2} /* (23, 7, 20) {real, imag} */,
  {32'h3fbe6590, 32'hbfe422bc} /* (23, 7, 19) {real, imag} */,
  {32'hc0ccd845, 32'h4030765c} /* (23, 7, 18) {real, imag} */,
  {32'h410ab6e3, 32'hc17f4848} /* (23, 7, 17) {real, imag} */,
  {32'h40eefa2a, 32'hc174e8a6} /* (23, 7, 16) {real, imag} */,
  {32'h4061d248, 32'hc0117d8a} /* (23, 7, 15) {real, imag} */,
  {32'hc0eac151, 32'hc0151972} /* (23, 7, 14) {real, imag} */,
  {32'h40f20ba2, 32'h3ff4b1e0} /* (23, 7, 13) {real, imag} */,
  {32'hc1712f4b, 32'hc090fb74} /* (23, 7, 12) {real, imag} */,
  {32'h40acb3e1, 32'hc1578a4d} /* (23, 7, 11) {real, imag} */,
  {32'hc0fa8098, 32'h413e5339} /* (23, 7, 10) {real, imag} */,
  {32'hc0d697fa, 32'hc10e8c3e} /* (23, 7, 9) {real, imag} */,
  {32'h41768fcc, 32'hbd9bca20} /* (23, 7, 8) {real, imag} */,
  {32'h41493031, 32'hc0a7d049} /* (23, 7, 7) {real, imag} */,
  {32'h4199dc3c, 32'h40e8b651} /* (23, 7, 6) {real, imag} */,
  {32'h4002a37c, 32'h40927f6f} /* (23, 7, 5) {real, imag} */,
  {32'h410ef746, 32'h3f8f6750} /* (23, 7, 4) {real, imag} */,
  {32'hc141d150, 32'h41aa09f7} /* (23, 7, 3) {real, imag} */,
  {32'h41cb8a6c, 32'hbf332fb0} /* (23, 7, 2) {real, imag} */,
  {32'hc13629ee, 32'hc20501b4} /* (23, 7, 1) {real, imag} */,
  {32'h409e47b3, 32'hc1eedda0} /* (23, 7, 0) {real, imag} */,
  {32'h41343a3f, 32'hc1c79094} /* (23, 6, 31) {real, imag} */,
  {32'hc0334f8c, 32'hc084adf7} /* (23, 6, 30) {real, imag} */,
  {32'hc13c4c1c, 32'hc1a384bc} /* (23, 6, 29) {real, imag} */,
  {32'hbe2909c0, 32'h41d65081} /* (23, 6, 28) {real, imag} */,
  {32'hc09f516d, 32'h41b8e9c2} /* (23, 6, 27) {real, imag} */,
  {32'hc1e68903, 32'h400c0338} /* (23, 6, 26) {real, imag} */,
  {32'h40e0ce3c, 32'hc05513eb} /* (23, 6, 25) {real, imag} */,
  {32'hbf9a8b74, 32'h405f09be} /* (23, 6, 24) {real, imag} */,
  {32'h409e337f, 32'h40e419b8} /* (23, 6, 23) {real, imag} */,
  {32'hc1457b56, 32'hc1b05815} /* (23, 6, 22) {real, imag} */,
  {32'hc17292ee, 32'hbe9ab3a0} /* (23, 6, 21) {real, imag} */,
  {32'h414671de, 32'hc090ceb2} /* (23, 6, 20) {real, imag} */,
  {32'hc13264af, 32'h40a9ad21} /* (23, 6, 19) {real, imag} */,
  {32'h41520c32, 32'hc0a0bb34} /* (23, 6, 18) {real, imag} */,
  {32'h408fde06, 32'hbfcb38dc} /* (23, 6, 17) {real, imag} */,
  {32'h402053c4, 32'hc145b694} /* (23, 6, 16) {real, imag} */,
  {32'h40b17006, 32'h3fb00cce} /* (23, 6, 15) {real, imag} */,
  {32'h3fdb7960, 32'h410335c0} /* (23, 6, 14) {real, imag} */,
  {32'hc05ccd0a, 32'h40515180} /* (23, 6, 13) {real, imag} */,
  {32'h3fea1554, 32'hbfed0980} /* (23, 6, 12) {real, imag} */,
  {32'hc13ebffc, 32'h41559f47} /* (23, 6, 11) {real, imag} */,
  {32'hc0afed9e, 32'h40ae63c2} /* (23, 6, 10) {real, imag} */,
  {32'hbfcde19c, 32'h40cd831d} /* (23, 6, 9) {real, imag} */,
  {32'hc1820dad, 32'hc0aebc9c} /* (23, 6, 8) {real, imag} */,
  {32'hc10ddbfb, 32'h415fafae} /* (23, 6, 7) {real, imag} */,
  {32'hc1c99020, 32'h3f002df0} /* (23, 6, 6) {real, imag} */,
  {32'hbbef5e00, 32'h416bf90a} /* (23, 6, 5) {real, imag} */,
  {32'h419b5aee, 32'hc1649fc4} /* (23, 6, 4) {real, imag} */,
  {32'h412c603a, 32'hc115a49c} /* (23, 6, 3) {real, imag} */,
  {32'hc1415c35, 32'hc0281fbc} /* (23, 6, 2) {real, imag} */,
  {32'h41678306, 32'h4141db32} /* (23, 6, 1) {real, imag} */,
  {32'h40a102da, 32'hc0ae895c} /* (23, 6, 0) {real, imag} */,
  {32'h42d84026, 32'h4209b5bd} /* (23, 5, 31) {real, imag} */,
  {32'hc27d2036, 32'h4145ac7f} /* (23, 5, 30) {real, imag} */,
  {32'h41d1db1b, 32'hc1532b5d} /* (23, 5, 29) {real, imag} */,
  {32'h40fb3e3a, 32'hc1cb11bb} /* (23, 5, 28) {real, imag} */,
  {32'hc218a6e6, 32'hc11e20a0} /* (23, 5, 27) {real, imag} */,
  {32'hc14b39b2, 32'hc059ee3c} /* (23, 5, 26) {real, imag} */,
  {32'h4003c90d, 32'hc1849993} /* (23, 5, 25) {real, imag} */,
  {32'hc0178cf6, 32'h40d7d9aa} /* (23, 5, 24) {real, imag} */,
  {32'h4195c50e, 32'h4018f537} /* (23, 5, 23) {real, imag} */,
  {32'hc11e4626, 32'hc03ba524} /* (23, 5, 22) {real, imag} */,
  {32'h409c1f36, 32'hc137d366} /* (23, 5, 21) {real, imag} */,
  {32'h40052f14, 32'h401a7d22} /* (23, 5, 20) {real, imag} */,
  {32'h40c3a10c, 32'h4180a834} /* (23, 5, 19) {real, imag} */,
  {32'h3f45fcf8, 32'h408d26e2} /* (23, 5, 18) {real, imag} */,
  {32'hc0b4298b, 32'hbfc744bc} /* (23, 5, 17) {real, imag} */,
  {32'h40346ed0, 32'h411f71ca} /* (23, 5, 16) {real, imag} */,
  {32'hbf917420, 32'hc0899dbe} /* (23, 5, 15) {real, imag} */,
  {32'hbf0a9cc0, 32'hc023d4dd} /* (23, 5, 14) {real, imag} */,
  {32'hc02c6413, 32'hc0b97878} /* (23, 5, 13) {real, imag} */,
  {32'hc01814bd, 32'h3d3827e0} /* (23, 5, 12) {real, imag} */,
  {32'hc1341078, 32'hc184a428} /* (23, 5, 11) {real, imag} */,
  {32'hc1518ac2, 32'hbedc3ec0} /* (23, 5, 10) {real, imag} */,
  {32'hbd225580, 32'hc02bb5bf} /* (23, 5, 9) {real, imag} */,
  {32'h41c6e1f5, 32'h3fbbcd28} /* (23, 5, 8) {real, imag} */,
  {32'h3e1a4540, 32'hbfb70114} /* (23, 5, 7) {real, imag} */,
  {32'h3eeb3bc0, 32'h417f234c} /* (23, 5, 6) {real, imag} */,
  {32'h3f1a0680, 32'hc1e1f99c} /* (23, 5, 5) {real, imag} */,
  {32'h40f41b86, 32'h423d769c} /* (23, 5, 4) {real, imag} */,
  {32'h409f5de4, 32'hc191ecb0} /* (23, 5, 3) {real, imag} */,
  {32'hc17ae3ee, 32'hc20f6100} /* (23, 5, 2) {real, imag} */,
  {32'h428039a0, 32'h42a4d11e} /* (23, 5, 1) {real, imag} */,
  {32'h42979ddc, 32'h420a2077} /* (23, 5, 0) {real, imag} */,
  {32'hc24c40d1, 32'hc2c23c90} /* (23, 4, 31) {real, imag} */,
  {32'h42be3f20, 32'h42b6ddde} /* (23, 4, 30) {real, imag} */,
  {32'h40f356ad, 32'hc0457254} /* (23, 4, 29) {real, imag} */,
  {32'hc2433705, 32'hc1777f69} /* (23, 4, 28) {real, imag} */,
  {32'h41d12176, 32'hc1d4c085} /* (23, 4, 27) {real, imag} */,
  {32'hc0942418, 32'hc0ae4926} /* (23, 4, 26) {real, imag} */,
  {32'hc14e9410, 32'hc00da686} /* (23, 4, 25) {real, imag} */,
  {32'h424a805e, 32'h408fce1c} /* (23, 4, 24) {real, imag} */,
  {32'hc039c4ba, 32'hbe500048} /* (23, 4, 23) {real, imag} */,
  {32'hc171ffd4, 32'h41027f1a} /* (23, 4, 22) {real, imag} */,
  {32'h3ec42a58, 32'hc10d2907} /* (23, 4, 21) {real, imag} */,
  {32'h410448f0, 32'h4155fba0} /* (23, 4, 20) {real, imag} */,
  {32'h41615fd6, 32'hc0cb687f} /* (23, 4, 19) {real, imag} */,
  {32'h3fd6d6cc, 32'h4115c101} /* (23, 4, 18) {real, imag} */,
  {32'h3f257258, 32'hc134ff53} /* (23, 4, 17) {real, imag} */,
  {32'hc017fd9a, 32'h40539c0b} /* (23, 4, 16) {real, imag} */,
  {32'h412fde39, 32'hc0adc509} /* (23, 4, 15) {real, imag} */,
  {32'h3e9399c8, 32'h415b53d6} /* (23, 4, 14) {real, imag} */,
  {32'hc033f2ec, 32'h40f2c11e} /* (23, 4, 13) {real, imag} */,
  {32'hc06f15c8, 32'h3f94386c} /* (23, 4, 12) {real, imag} */,
  {32'hc1621ae0, 32'h414690a3} /* (23, 4, 11) {real, imag} */,
  {32'h40fdbe28, 32'h410a49f0} /* (23, 4, 10) {real, imag} */,
  {32'hc0ef21ae, 32'hc12f7851} /* (23, 4, 9) {real, imag} */,
  {32'h408b4bbe, 32'hc14c0111} /* (23, 4, 8) {real, imag} */,
  {32'hc1c39506, 32'hc1049418} /* (23, 4, 7) {real, imag} */,
  {32'hc19cb234, 32'h40a4a876} /* (23, 4, 6) {real, imag} */,
  {32'h410a241c, 32'h40270af4} /* (23, 4, 5) {real, imag} */,
  {32'h4206d6d6, 32'hc2265bf0} /* (23, 4, 4) {real, imag} */,
  {32'h41702ed0, 32'hc1c49130} /* (23, 4, 3) {real, imag} */,
  {32'h42ec2057, 32'h42618a3b} /* (23, 4, 2) {real, imag} */,
  {32'hc304c3d7, 32'hc26f1274} /* (23, 4, 1) {real, imag} */,
  {32'hc29b529e, 32'h41a18e94} /* (23, 4, 0) {real, imag} */,
  {32'h4307fc76, 32'hc2aade2e} /* (23, 3, 31) {real, imag} */,
  {32'hc284e30c, 32'h42cca452} /* (23, 3, 30) {real, imag} */,
  {32'hc16b201a, 32'h4122248a} /* (23, 3, 29) {real, imag} */,
  {32'hc21632bb, 32'hc1d38c60} /* (23, 3, 28) {real, imag} */,
  {32'h423e318e, 32'h4044c28c} /* (23, 3, 27) {real, imag} */,
  {32'hc1210dfb, 32'h40b854ed} /* (23, 3, 26) {real, imag} */,
  {32'hbed1c5c0, 32'hc1f302c2} /* (23, 3, 25) {real, imag} */,
  {32'hc0f842c4, 32'h41518260} /* (23, 3, 24) {real, imag} */,
  {32'hc13a70ab, 32'hc169f307} /* (23, 3, 23) {real, imag} */,
  {32'hc044a30c, 32'hc00b2673} /* (23, 3, 22) {real, imag} */,
  {32'h3ff34252, 32'hc0dd369b} /* (23, 3, 21) {real, imag} */,
  {32'hc10803fc, 32'hc15798a4} /* (23, 3, 20) {real, imag} */,
  {32'hc0f5e146, 32'h412f8656} /* (23, 3, 19) {real, imag} */,
  {32'h40e61327, 32'h40c2aa06} /* (23, 3, 18) {real, imag} */,
  {32'hc11b4e51, 32'h407626b0} /* (23, 3, 17) {real, imag} */,
  {32'h4189be82, 32'h3f8e9e6c} /* (23, 3, 16) {real, imag} */,
  {32'h4091f61f, 32'hc05af65c} /* (23, 3, 15) {real, imag} */,
  {32'h3f6ab118, 32'h4121dce6} /* (23, 3, 14) {real, imag} */,
  {32'h403bc1ae, 32'h4009c567} /* (23, 3, 13) {real, imag} */,
  {32'hc1860867, 32'hc17bb03a} /* (23, 3, 12) {real, imag} */,
  {32'h411452f5, 32'hc0dfc04f} /* (23, 3, 11) {real, imag} */,
  {32'hc0b28a51, 32'h40efe7f5} /* (23, 3, 10) {real, imag} */,
  {32'h40047a64, 32'h3e970c38} /* (23, 3, 9) {real, imag} */,
  {32'hc1060738, 32'h4161a9de} /* (23, 3, 8) {real, imag} */,
  {32'hc135a23a, 32'hc1afadc0} /* (23, 3, 7) {real, imag} */,
  {32'hc1475569, 32'h41aba4e3} /* (23, 3, 6) {real, imag} */,
  {32'hc17f5bf6, 32'hc198e7ab} /* (23, 3, 5) {real, imag} */,
  {32'h4219a45a, 32'hc2171346} /* (23, 3, 4) {real, imag} */,
  {32'hc1098167, 32'hc0f2d87c} /* (23, 3, 3) {real, imag} */,
  {32'hc18fba7a, 32'h4314b7e2} /* (23, 3, 2) {real, imag} */,
  {32'hc2fa0378, 32'hc28b5b6e} /* (23, 3, 1) {real, imag} */,
  {32'h42b289dc, 32'h410fab8d} /* (23, 3, 0) {real, imag} */,
  {32'h448d8d54, 32'h428929ed} /* (23, 2, 31) {real, imag} */,
  {32'hc4004dd6, 32'h4318de2e} /* (23, 2, 30) {real, imag} */,
  {32'h4205622a, 32'hc1fe6136} /* (23, 2, 29) {real, imag} */,
  {32'h4210b104, 32'hc2a6d48d} /* (23, 2, 28) {real, imag} */,
  {32'hc26f603e, 32'h4170b745} /* (23, 2, 27) {real, imag} */,
  {32'hc14dc896, 32'h41a648f5} /* (23, 2, 26) {real, imag} */,
  {32'h409d8022, 32'h40c9aef5} /* (23, 2, 25) {real, imag} */,
  {32'hc08e63de, 32'h41875939} /* (23, 2, 24) {real, imag} */,
  {32'hc112a177, 32'h40ea2e14} /* (23, 2, 23) {real, imag} */,
  {32'h404a5c8e, 32'h410e57a6} /* (23, 2, 22) {real, imag} */,
  {32'hc0219e03, 32'hbf1d9d76} /* (23, 2, 21) {real, imag} */,
  {32'h40b49ca0, 32'h41035139} /* (23, 2, 20) {real, imag} */,
  {32'h40e81410, 32'h410996f8} /* (23, 2, 19) {real, imag} */,
  {32'h3f77215d, 32'h3f4684e0} /* (23, 2, 18) {real, imag} */,
  {32'hc116f083, 32'hc14a5172} /* (23, 2, 17) {real, imag} */,
  {32'hc10054e7, 32'h414cd86c} /* (23, 2, 16) {real, imag} */,
  {32'h414d39ba, 32'h41040d6c} /* (23, 2, 15) {real, imag} */,
  {32'hc0ddafee, 32'hbffc2230} /* (23, 2, 14) {real, imag} */,
  {32'hc08d3392, 32'hbf436538} /* (23, 2, 13) {real, imag} */,
  {32'hc0901495, 32'h4083563e} /* (23, 2, 12) {real, imag} */,
  {32'hc128cdde, 32'hc169f938} /* (23, 2, 11) {real, imag} */,
  {32'h407705b6, 32'h413f5da4} /* (23, 2, 10) {real, imag} */,
  {32'h4134e1ee, 32'h4149d1cb} /* (23, 2, 9) {real, imag} */,
  {32'hc1c7eb87, 32'h41c0f53e} /* (23, 2, 8) {real, imag} */,
  {32'h4192a0e2, 32'h4118f4de} /* (23, 2, 7) {real, imag} */,
  {32'hbfdb9b90, 32'h4094fb42} /* (23, 2, 6) {real, imag} */,
  {32'hc29969ca, 32'hc2895e65} /* (23, 2, 5) {real, imag} */,
  {32'h42bae243, 32'h426f8566} /* (23, 2, 4) {real, imag} */,
  {32'h40b051ae, 32'hc204bbfa} /* (23, 2, 3) {real, imag} */,
  {32'hc3b782d9, 32'h426039dd} /* (23, 2, 2) {real, imag} */,
  {32'h4423b111, 32'hc28030bb} /* (23, 2, 1) {real, imag} */,
  {32'h44136f1d, 32'h42debdb6} /* (23, 2, 0) {real, imag} */,
  {32'hc4bef642, 32'h43c64375} /* (23, 1, 31) {real, imag} */,
  {32'h43b97e08, 32'h42c7a4af} /* (23, 1, 30) {real, imag} */,
  {32'h423ed4c7, 32'hc2117ce6} /* (23, 1, 29) {real, imag} */,
  {32'hc2f497c3, 32'hc1bb464a} /* (23, 1, 28) {real, imag} */,
  {32'h43035292, 32'hc10a4b87} /* (23, 1, 27) {real, imag} */,
  {32'h41800e6c, 32'h408ba27f} /* (23, 1, 26) {real, imag} */,
  {32'hc188bbaa, 32'h41b2af03} /* (23, 1, 25) {real, imag} */,
  {32'h4164f898, 32'hc198423e} /* (23, 1, 24) {real, imag} */,
  {32'h410b3e58, 32'hc182ef78} /* (23, 1, 23) {real, imag} */,
  {32'hc135a73e, 32'hbe746030} /* (23, 1, 22) {real, imag} */,
  {32'h4154f591, 32'hc0e26385} /* (23, 1, 21) {real, imag} */,
  {32'hc03680a9, 32'h3fa71c0e} /* (23, 1, 20) {real, imag} */,
  {32'h3f431cb4, 32'h40a416b5} /* (23, 1, 19) {real, imag} */,
  {32'hc115d8c3, 32'hc101f154} /* (23, 1, 18) {real, imag} */,
  {32'h40261db8, 32'hc14b530e} /* (23, 1, 17) {real, imag} */,
  {32'hbf4096e4, 32'h3fb7c518} /* (23, 1, 16) {real, imag} */,
  {32'h40957fdf, 32'hc045ed62} /* (23, 1, 15) {real, imag} */,
  {32'hbdfaf530, 32'h40f11340} /* (23, 1, 14) {real, imag} */,
  {32'h3fc12f58, 32'hc11cd642} /* (23, 1, 13) {real, imag} */,
  {32'h401276c0, 32'hc00b597a} /* (23, 1, 12) {real, imag} */,
  {32'hc0957f2a, 32'h41c9ef1c} /* (23, 1, 11) {real, imag} */,
  {32'h410a7593, 32'hc025abe0} /* (23, 1, 10) {real, imag} */,
  {32'h41a2d8b8, 32'h40d60520} /* (23, 1, 9) {real, imag} */,
  {32'h4188e354, 32'h41847db0} /* (23, 1, 8) {real, imag} */,
  {32'hc19b6a79, 32'hc1713484} /* (23, 1, 7) {real, imag} */,
  {32'h41fa9161, 32'hc19f313e} /* (23, 1, 6) {real, imag} */,
  {32'h4289667e, 32'h423c3ea8} /* (23, 1, 5) {real, imag} */,
  {32'hc2779290, 32'hc24e75d0} /* (23, 1, 4) {real, imag} */,
  {32'h426795ba, 32'h41917c12} /* (23, 1, 3) {real, imag} */,
  {32'h4403b620, 32'h43f4792e} /* (23, 1, 2) {real, imag} */,
  {32'hc5068bfc, 32'hc497fdc2} /* (23, 1, 1) {real, imag} */,
  {32'hc4f7c643, 32'hc3749fae} /* (23, 1, 0) {real, imag} */,
  {32'hc4b17406, 32'h448d2b08} /* (23, 0, 31) {real, imag} */,
  {32'h43396d4a, 32'hc35bc84f} /* (23, 0, 30) {real, imag} */,
  {32'h416f21d6, 32'h4139f254} /* (23, 0, 29) {real, imag} */,
  {32'h424d64b2, 32'hc29f7024} /* (23, 0, 28) {real, imag} */,
  {32'h4268e6b6, 32'hc088d3c1} /* (23, 0, 27) {real, imag} */,
  {32'h410d7894, 32'h40e6c979} /* (23, 0, 26) {real, imag} */,
  {32'h41ddd128, 32'h418128b3} /* (23, 0, 25) {real, imag} */,
  {32'hc00af342, 32'h409b05bc} /* (23, 0, 24) {real, imag} */,
  {32'h4123112e, 32'h412db5c9} /* (23, 0, 23) {real, imag} */,
  {32'hc187c69d, 32'hc01a0468} /* (23, 0, 22) {real, imag} */,
  {32'h41845376, 32'h3d45ec80} /* (23, 0, 21) {real, imag} */,
  {32'hc13dec88, 32'h40caa794} /* (23, 0, 20) {real, imag} */,
  {32'hc1936f7e, 32'hbffe52d0} /* (23, 0, 19) {real, imag} */,
  {32'h3fbda822, 32'hc06dac72} /* (23, 0, 18) {real, imag} */,
  {32'h3f91129c, 32'h3f9982a4} /* (23, 0, 17) {real, imag} */,
  {32'hc090722e, 32'h00000000} /* (23, 0, 16) {real, imag} */,
  {32'h3f91129c, 32'hbf9982a4} /* (23, 0, 15) {real, imag} */,
  {32'h3fbda822, 32'h406dac72} /* (23, 0, 14) {real, imag} */,
  {32'hc1936f7e, 32'h3ffe52d0} /* (23, 0, 13) {real, imag} */,
  {32'hc13dec88, 32'hc0caa794} /* (23, 0, 12) {real, imag} */,
  {32'h41845376, 32'hbd45ec80} /* (23, 0, 11) {real, imag} */,
  {32'hc187c69d, 32'h401a0468} /* (23, 0, 10) {real, imag} */,
  {32'h4123112e, 32'hc12db5c9} /* (23, 0, 9) {real, imag} */,
  {32'hc00af342, 32'hc09b05bc} /* (23, 0, 8) {real, imag} */,
  {32'h41ddd128, 32'hc18128b3} /* (23, 0, 7) {real, imag} */,
  {32'h410d7894, 32'hc0e6c979} /* (23, 0, 6) {real, imag} */,
  {32'h4268e6b6, 32'h4088d3c1} /* (23, 0, 5) {real, imag} */,
  {32'h424d64b2, 32'h429f7024} /* (23, 0, 4) {real, imag} */,
  {32'h416f21d6, 32'hc139f254} /* (23, 0, 3) {real, imag} */,
  {32'h43396d4a, 32'h435bc84f} /* (23, 0, 2) {real, imag} */,
  {32'hc4b17406, 32'hc48d2b08} /* (23, 0, 1) {real, imag} */,
  {32'hc50b5d50, 32'h00000000} /* (23, 0, 0) {real, imag} */,
  {32'hc5188d2b, 32'h44a3f327} /* (22, 31, 31) {real, imag} */,
  {32'h44100e9d, 32'hc40e30d7} /* (22, 31, 30) {real, imag} */,
  {32'h42856b01, 32'hc1c10cc4} /* (22, 31, 29) {real, imag} */,
  {32'hc25493e2, 32'h428f9744} /* (22, 31, 28) {real, imag} */,
  {32'h42887c97, 32'hc26006c1} /* (22, 31, 27) {real, imag} */,
  {32'hc081a2c4, 32'h40c959ba} /* (22, 31, 26) {real, imag} */,
  {32'hc14586a9, 32'h422dcd14} /* (22, 31, 25) {real, imag} */,
  {32'h4099a629, 32'hc23cd0a4} /* (22, 31, 24) {real, imag} */,
  {32'h40cc8ed1, 32'h4145d99d} /* (22, 31, 23) {real, imag} */,
  {32'hc139412a, 32'hc14f3ee7} /* (22, 31, 22) {real, imag} */,
  {32'h4183ab84, 32'hc0ccfb0d} /* (22, 31, 21) {real, imag} */,
  {32'h4118f52a, 32'hc090004c} /* (22, 31, 20) {real, imag} */,
  {32'hc16ed590, 32'h40c06d60} /* (22, 31, 19) {real, imag} */,
  {32'h3ed43330, 32'hc1628776} /* (22, 31, 18) {real, imag} */,
  {32'hc090964e, 32'hc123f154} /* (22, 31, 17) {real, imag} */,
  {32'h40ad62ce, 32'h4098e40c} /* (22, 31, 16) {real, imag} */,
  {32'hc08e4226, 32'hc072ac55} /* (22, 31, 15) {real, imag} */,
  {32'h409ab3ec, 32'hc109683a} /* (22, 31, 14) {real, imag} */,
  {32'h40208910, 32'h40d1ebb4} /* (22, 31, 13) {real, imag} */,
  {32'h40cdcde5, 32'h40da1ffa} /* (22, 31, 12) {real, imag} */,
  {32'h40fe650b, 32'hc0f91436} /* (22, 31, 11) {real, imag} */,
  {32'h412eb0bd, 32'h410304c3} /* (22, 31, 10) {real, imag} */,
  {32'h4171c55c, 32'h41cfefc6} /* (22, 31, 9) {real, imag} */,
  {32'h4179f2c4, 32'h415d731e} /* (22, 31, 8) {real, imag} */,
  {32'hc18ec39c, 32'h414895c4} /* (22, 31, 7) {real, imag} */,
  {32'h41d6bc25, 32'h40542674} /* (22, 31, 6) {real, imag} */,
  {32'h430f695e, 32'h411fe67f} /* (22, 31, 5) {real, imag} */,
  {32'hc30cdf8f, 32'h4282e392} /* (22, 31, 4) {real, imag} */,
  {32'h41dc9d48, 32'h42892b77} /* (22, 31, 3) {real, imag} */,
  {32'h43e49f0c, 32'hc2aa096e} /* (22, 31, 2) {real, imag} */,
  {32'hc4d5cc2b, 32'hc3e59299} /* (22, 31, 1) {real, imag} */,
  {32'hc506879a, 32'h43971b6c} /* (22, 31, 0) {real, imag} */,
  {32'h44339153, 32'h42a62180} /* (22, 30, 31) {real, imag} */,
  {32'hc3cd8aca, 32'hc2b61d12} /* (22, 30, 30) {real, imag} */,
  {32'h40a6fc6c, 32'h4236204b} /* (22, 30, 29) {real, imag} */,
  {32'h42c03adf, 32'hc28b6ee7} /* (22, 30, 28) {real, imag} */,
  {32'hc2a34c60, 32'h42903032} /* (22, 30, 27) {real, imag} */,
  {32'hc0e2859a, 32'hc15ce178} /* (22, 30, 26) {real, imag} */,
  {32'h3f5f1538, 32'h4049f334} /* (22, 30, 25) {real, imag} */,
  {32'hc1ab67ca, 32'h41905571} /* (22, 30, 24) {real, imag} */,
  {32'h4089fac1, 32'h3fc8fcfc} /* (22, 30, 23) {real, imag} */,
  {32'h4159f63e, 32'hc1b283f3} /* (22, 30, 22) {real, imag} */,
  {32'hc092b6b3, 32'h41a96855} /* (22, 30, 21) {real, imag} */,
  {32'hc15b1b2a, 32'h4187bac5} /* (22, 30, 20) {real, imag} */,
  {32'h413d8a8e, 32'hc0ba691a} /* (22, 30, 19) {real, imag} */,
  {32'h415c3672, 32'hc01cd974} /* (22, 30, 18) {real, imag} */,
  {32'hbf9b4978, 32'hc032ef32} /* (22, 30, 17) {real, imag} */,
  {32'h3fa16b7e, 32'h3e81b444} /* (22, 30, 16) {real, imag} */,
  {32'h39b68000, 32'h40dd188a} /* (22, 30, 15) {real, imag} */,
  {32'hc052c0c6, 32'hc15f3a92} /* (22, 30, 14) {real, imag} */,
  {32'hc1926ad2, 32'hc1630a28} /* (22, 30, 13) {real, imag} */,
  {32'h412646c0, 32'hc1278714} /* (22, 30, 12) {real, imag} */,
  {32'h3ff429b4, 32'hc1106ed8} /* (22, 30, 11) {real, imag} */,
  {32'hc05e7c60, 32'hc12cb5f8} /* (22, 30, 10) {real, imag} */,
  {32'hc1086ef7, 32'h41058c64} /* (22, 30, 9) {real, imag} */,
  {32'hc12bd461, 32'hc10ba84c} /* (22, 30, 8) {real, imag} */,
  {32'h41e23c04, 32'h41620bc2} /* (22, 30, 7) {real, imag} */,
  {32'hc21428ad, 32'h40b43f0c} /* (22, 30, 6) {real, imag} */,
  {32'hc25e244b, 32'hc1e9443b} /* (22, 30, 5) {real, imag} */,
  {32'h420fa701, 32'h42c43e52} /* (22, 30, 4) {real, imag} */,
  {32'hc085e878, 32'h41b1d48c} /* (22, 30, 3) {real, imag} */,
  {32'hc40ac138, 32'hc3504f88} /* (22, 30, 2) {real, imag} */,
  {32'h449cedcb, 32'hc2199956} /* (22, 30, 1) {real, imag} */,
  {32'h441f47b8, 32'hc309dc98} /* (22, 30, 0) {real, imag} */,
  {32'hc304234c, 32'h42abcd6e} /* (22, 29, 31) {real, imag} */,
  {32'hc18e3b76, 32'hc30959f0} /* (22, 29, 30) {real, imag} */,
  {32'h40309af0, 32'h41a6b081} /* (22, 29, 29) {real, imag} */,
  {32'h41dc5fce, 32'h427481d2} /* (22, 29, 28) {real, imag} */,
  {32'hc1bd52a3, 32'h40e1d01e} /* (22, 29, 27) {real, imag} */,
  {32'h41716600, 32'hc0416bda} /* (22, 29, 26) {real, imag} */,
  {32'h40ef066d, 32'h4100565c} /* (22, 29, 25) {real, imag} */,
  {32'hc158a89a, 32'hc17847e9} /* (22, 29, 24) {real, imag} */,
  {32'hc12c692c, 32'h418d3c98} /* (22, 29, 23) {real, imag} */,
  {32'hc118ca58, 32'hc1ab1016} /* (22, 29, 22) {real, imag} */,
  {32'hc10190a6, 32'hbfe0d310} /* (22, 29, 21) {real, imag} */,
  {32'h41a0bde2, 32'h40958254} /* (22, 29, 20) {real, imag} */,
  {32'h40560d7b, 32'hc123a702} /* (22, 29, 19) {real, imag} */,
  {32'hc1288d5a, 32'hbfd6ae3c} /* (22, 29, 18) {real, imag} */,
  {32'hc12d7de3, 32'h3ff95bc0} /* (22, 29, 17) {real, imag} */,
  {32'h40a52e0e, 32'h40bc638a} /* (22, 29, 16) {real, imag} */,
  {32'hc0b893e3, 32'hc0924c06} /* (22, 29, 15) {real, imag} */,
  {32'h41484e6e, 32'hc02a3cf0} /* (22, 29, 14) {real, imag} */,
  {32'h411e469c, 32'hc117baa7} /* (22, 29, 13) {real, imag} */,
  {32'h412cb868, 32'h4124bee4} /* (22, 29, 12) {real, imag} */,
  {32'hbe7d4e98, 32'hc0df7e68} /* (22, 29, 11) {real, imag} */,
  {32'hc140f862, 32'h4139b9e8} /* (22, 29, 10) {real, imag} */,
  {32'hc0714d3c, 32'h4177f472} /* (22, 29, 9) {real, imag} */,
  {32'h41c94744, 32'hc0c34ee3} /* (22, 29, 8) {real, imag} */,
  {32'h41131b8f, 32'h4199069b} /* (22, 29, 7) {real, imag} */,
  {32'h4093ddb4, 32'h408605e2} /* (22, 29, 6) {real, imag} */,
  {32'h41a99642, 32'hc0f385f4} /* (22, 29, 5) {real, imag} */,
  {32'hc26afca8, 32'h41fa9d50} /* (22, 29, 4) {real, imag} */,
  {32'hc0216f84, 32'h408ddfa6} /* (22, 29, 3) {real, imag} */,
  {32'hc2be7f5b, 32'hc2db40fa} /* (22, 29, 2) {real, imag} */,
  {32'h43128d49, 32'h428e305d} /* (22, 29, 1) {real, imag} */,
  {32'h42850126, 32'h3f045a60} /* (22, 29, 0) {real, imag} */,
  {32'hc2e8461e, 32'h4214eb4a} /* (22, 28, 31) {real, imag} */,
  {32'h42d9f190, 32'hc284598b} /* (22, 28, 30) {real, imag} */,
  {32'h41273f7a, 32'h4107b3df} /* (22, 28, 29) {real, imag} */,
  {32'h418fd021, 32'h421d48d5} /* (22, 28, 28) {real, imag} */,
  {32'h402f07ec, 32'hc00149b0} /* (22, 28, 27) {real, imag} */,
  {32'hc171bdc2, 32'h4030a72c} /* (22, 28, 26) {real, imag} */,
  {32'hc09adeb2, 32'h3ed728f0} /* (22, 28, 25) {real, imag} */,
  {32'h418529ee, 32'h40ac7a72} /* (22, 28, 24) {real, imag} */,
  {32'h40ecd5c7, 32'h40c956e1} /* (22, 28, 23) {real, imag} */,
  {32'hbf512900, 32'hc17dd395} /* (22, 28, 22) {real, imag} */,
  {32'h41388ff7, 32'hc1730493} /* (22, 28, 21) {real, imag} */,
  {32'hc0c62c98, 32'h419dd60a} /* (22, 28, 20) {real, imag} */,
  {32'hc0fd0c50, 32'hc0cb30e0} /* (22, 28, 19) {real, imag} */,
  {32'h414e3398, 32'hc0642fb5} /* (22, 28, 18) {real, imag} */,
  {32'hc08239bd, 32'hc02717d0} /* (22, 28, 17) {real, imag} */,
  {32'hc070b3f8, 32'hc0199a83} /* (22, 28, 16) {real, imag} */,
  {32'hbda12eb8, 32'h3f1a0f30} /* (22, 28, 15) {real, imag} */,
  {32'h417568e6, 32'h40f9c769} /* (22, 28, 14) {real, imag} */,
  {32'hbf240991, 32'hc05c9c43} /* (22, 28, 13) {real, imag} */,
  {32'h3f79ade8, 32'h405f8728} /* (22, 28, 12) {real, imag} */,
  {32'hc1299460, 32'hc1326464} /* (22, 28, 11) {real, imag} */,
  {32'hc0856abc, 32'hc0b277ee} /* (22, 28, 10) {real, imag} */,
  {32'hc119c65e, 32'h416ad1b3} /* (22, 28, 9) {real, imag} */,
  {32'h41942800, 32'hc154c1ee} /* (22, 28, 8) {real, imag} */,
  {32'h411272a0, 32'h40a4770b} /* (22, 28, 7) {real, imag} */,
  {32'h409b4b7e, 32'h41230b76} /* (22, 28, 6) {real, imag} */,
  {32'h414c0331, 32'h413e7112} /* (22, 28, 5) {real, imag} */,
  {32'hc1a7e602, 32'h40c31b48} /* (22, 28, 4) {real, imag} */,
  {32'hc1d6fa5a, 32'hc0cf89b1} /* (22, 28, 3) {real, imag} */,
  {32'h42acce27, 32'hc2a58a7e} /* (22, 28, 2) {real, imag} */,
  {32'hc20ac486, 32'h42caa144} /* (22, 28, 1) {real, imag} */,
  {32'hc2a687b2, 32'hc1d23d72} /* (22, 28, 0) {real, imag} */,
  {32'h42c3ee42, 32'hc2bcd575} /* (22, 27, 31) {real, imag} */,
  {32'h40d77095, 32'h422206a0} /* (22, 27, 30) {real, imag} */,
  {32'hc027484b, 32'h40a225be} /* (22, 27, 29) {real, imag} */,
  {32'hc1260f44, 32'hc23f19b2} /* (22, 27, 28) {real, imag} */,
  {32'hc118e420, 32'h41ba9662} /* (22, 27, 27) {real, imag} */,
  {32'h4143ae9a, 32'hc009e92a} /* (22, 27, 26) {real, imag} */,
  {32'h411ca0d2, 32'h3f95b224} /* (22, 27, 25) {real, imag} */,
  {32'hbfb48140, 32'h3e547800} /* (22, 27, 24) {real, imag} */,
  {32'h40c5c1b3, 32'h3eaeb738} /* (22, 27, 23) {real, imag} */,
  {32'hc0a91a7e, 32'h4134a42a} /* (22, 27, 22) {real, imag} */,
  {32'hc0ada160, 32'h41816d7c} /* (22, 27, 21) {real, imag} */,
  {32'hc156c29c, 32'h40d8ed0f} /* (22, 27, 20) {real, imag} */,
  {32'h414e23aa, 32'h40ab34ff} /* (22, 27, 19) {real, imag} */,
  {32'h4131207a, 32'h40c04c78} /* (22, 27, 18) {real, imag} */,
  {32'hc01ba87c, 32'hc0c240c8} /* (22, 27, 17) {real, imag} */,
  {32'hc16a741c, 32'h41143956} /* (22, 27, 16) {real, imag} */,
  {32'h3fcbfbe1, 32'h402ad196} /* (22, 27, 15) {real, imag} */,
  {32'h41405570, 32'hbe810700} /* (22, 27, 14) {real, imag} */,
  {32'h40b45590, 32'h40a77a51} /* (22, 27, 13) {real, imag} */,
  {32'h41063ef1, 32'h41812952} /* (22, 27, 12) {real, imag} */,
  {32'hc021cc62, 32'hbff71508} /* (22, 27, 11) {real, imag} */,
  {32'hc1aaa39b, 32'hc0ebd3de} /* (22, 27, 10) {real, imag} */,
  {32'h41094d30, 32'h418040d8} /* (22, 27, 9) {real, imag} */,
  {32'hc149f456, 32'hbfdbddd0} /* (22, 27, 8) {real, imag} */,
  {32'hc0b9983c, 32'h40cead34} /* (22, 27, 7) {real, imag} */,
  {32'hbfd3cf8a, 32'hc1b48a86} /* (22, 27, 6) {real, imag} */,
  {32'hc2181e7b, 32'h404a6d3a} /* (22, 27, 5) {real, imag} */,
  {32'hc177b875, 32'h4070f3e8} /* (22, 27, 4) {real, imag} */,
  {32'hc0121dbf, 32'h40b32cc4} /* (22, 27, 3) {real, imag} */,
  {32'hc27955d3, 32'h4170a908} /* (22, 27, 2) {real, imag} */,
  {32'h42c21804, 32'hc1cd22ba} /* (22, 27, 1) {real, imag} */,
  {32'h428e3266, 32'hc221a283} /* (22, 27, 0) {real, imag} */,
  {32'h4146bbf4, 32'hc0d9f576} /* (22, 26, 31) {real, imag} */,
  {32'hc19c8e86, 32'hc038636c} /* (22, 26, 30) {real, imag} */,
  {32'h41be9294, 32'h420208b2} /* (22, 26, 29) {real, imag} */,
  {32'h41045c35, 32'hbfadbb34} /* (22, 26, 28) {real, imag} */,
  {32'hc1c8a185, 32'hc0fbd728} /* (22, 26, 27) {real, imag} */,
  {32'hc0a85a07, 32'h41823415} /* (22, 26, 26) {real, imag} */,
  {32'hc1703075, 32'h40f35a2e} /* (22, 26, 25) {real, imag} */,
  {32'h40b48b03, 32'h411f0ce4} /* (22, 26, 24) {real, imag} */,
  {32'h408b95f7, 32'h402cae22} /* (22, 26, 23) {real, imag} */,
  {32'hc19c00b5, 32'hbf43dbf0} /* (22, 26, 22) {real, imag} */,
  {32'hc1237747, 32'hc0ca14f6} /* (22, 26, 21) {real, imag} */,
  {32'h410f0d5f, 32'hc16b3741} /* (22, 26, 20) {real, imag} */,
  {32'h4108d128, 32'hc016f279} /* (22, 26, 19) {real, imag} */,
  {32'hc0f934d4, 32'hc121719e} /* (22, 26, 18) {real, imag} */,
  {32'hc0bd2b0a, 32'hc0e2332f} /* (22, 26, 17) {real, imag} */,
  {32'hc09e9fb3, 32'hc02735e0} /* (22, 26, 16) {real, imag} */,
  {32'h3fb89124, 32'h40f0202a} /* (22, 26, 15) {real, imag} */,
  {32'hc02a1d7a, 32'hc09ca880} /* (22, 26, 14) {real, imag} */,
  {32'hc00ff1e4, 32'hc146abe1} /* (22, 26, 13) {real, imag} */,
  {32'hc0831127, 32'h40f61efd} /* (22, 26, 12) {real, imag} */,
  {32'hbf0a1560, 32'h40cfb4f0} /* (22, 26, 11) {real, imag} */,
  {32'hc09d2bd2, 32'hc180d7e6} /* (22, 26, 10) {real, imag} */,
  {32'hc15ec086, 32'hc0427e68} /* (22, 26, 9) {real, imag} */,
  {32'h41027f05, 32'h4163b4f2} /* (22, 26, 8) {real, imag} */,
  {32'hc10cae06, 32'h3ed58d18} /* (22, 26, 7) {real, imag} */,
  {32'hc1955776, 32'hc1045686} /* (22, 26, 6) {real, imag} */,
  {32'hc055aec8, 32'h40bd3122} /* (22, 26, 5) {real, imag} */,
  {32'hc00926ec, 32'h41ac5217} /* (22, 26, 4) {real, imag} */,
  {32'h40d784e1, 32'hc15bcf7c} /* (22, 26, 3) {real, imag} */,
  {32'hc0daba98, 32'h40de9f77} /* (22, 26, 2) {real, imag} */,
  {32'h411730e6, 32'hc0f0ccd4} /* (22, 26, 1) {real, imag} */,
  {32'h3f5057f0, 32'hc12e6960} /* (22, 26, 0) {real, imag} */,
  {32'hc07e6088, 32'h419a0693} /* (22, 25, 31) {real, imag} */,
  {32'hc118243d, 32'h41123a1f} /* (22, 25, 30) {real, imag} */,
  {32'h413a04ed, 32'hc217fc00} /* (22, 25, 29) {real, imag} */,
  {32'h3f547e88, 32'h41556654} /* (22, 25, 28) {real, imag} */,
  {32'h409be992, 32'hc10778ad} /* (22, 25, 27) {real, imag} */,
  {32'h410207e4, 32'hc0adbc15} /* (22, 25, 26) {real, imag} */,
  {32'hc0a3cd84, 32'h41fb595c} /* (22, 25, 25) {real, imag} */,
  {32'h40c69615, 32'h415a709b} /* (22, 25, 24) {real, imag} */,
  {32'hc058415e, 32'h3fa84cfc} /* (22, 25, 23) {real, imag} */,
  {32'hc1241624, 32'hc1244048} /* (22, 25, 22) {real, imag} */,
  {32'hc1c12ec4, 32'hbf79bcb8} /* (22, 25, 21) {real, imag} */,
  {32'hc08dfb04, 32'hc0e2de5c} /* (22, 25, 20) {real, imag} */,
  {32'h403f3eb6, 32'hc039a450} /* (22, 25, 19) {real, imag} */,
  {32'hc0d31a67, 32'hbe02df40} /* (22, 25, 18) {real, imag} */,
  {32'h3fbda130, 32'hc10cc1ed} /* (22, 25, 17) {real, imag} */,
  {32'h4089a110, 32'hc0afb7e3} /* (22, 25, 16) {real, imag} */,
  {32'h410df84d, 32'h40e53efa} /* (22, 25, 15) {real, imag} */,
  {32'h410a371e, 32'h3fda6f24} /* (22, 25, 14) {real, imag} */,
  {32'hc17f67d8, 32'hc0ea6ede} /* (22, 25, 13) {real, imag} */,
  {32'h3f9dd128, 32'h418737ad} /* (22, 25, 12) {real, imag} */,
  {32'h41525f6f, 32'h3fb22162} /* (22, 25, 11) {real, imag} */,
  {32'hc0f33b7f, 32'h404a8c68} /* (22, 25, 10) {real, imag} */,
  {32'h416cc39c, 32'hc11bb4c1} /* (22, 25, 9) {real, imag} */,
  {32'hc1fede80, 32'hc058fada} /* (22, 25, 8) {real, imag} */,
  {32'h40b51048, 32'hbed960d0} /* (22, 25, 7) {real, imag} */,
  {32'hc1323ec0, 32'hc148946c} /* (22, 25, 6) {real, imag} */,
  {32'hc00dff9c, 32'hc0511860} /* (22, 25, 5) {real, imag} */,
  {32'h4198ee7e, 32'hc144ac83} /* (22, 25, 4) {real, imag} */,
  {32'h41accc00, 32'hc0ec65aa} /* (22, 25, 3) {real, imag} */,
  {32'h41138f8e, 32'hc04cb8a4} /* (22, 25, 2) {real, imag} */,
  {32'hc1ab9732, 32'h41994f12} /* (22, 25, 1) {real, imag} */,
  {32'hc09c0135, 32'h41886aca} /* (22, 25, 0) {real, imag} */,
  {32'h3fb09408, 32'hc100b8d0} /* (22, 24, 31) {real, imag} */,
  {32'hc08acbbc, 32'hc0325fbc} /* (22, 24, 30) {real, imag} */,
  {32'h3f975e78, 32'h4141ca30} /* (22, 24, 29) {real, imag} */,
  {32'h416855cc, 32'hc1974d68} /* (22, 24, 28) {real, imag} */,
  {32'hc1c3f168, 32'h4114d480} /* (22, 24, 27) {real, imag} */,
  {32'h400450a6, 32'hc0445bfa} /* (22, 24, 26) {real, imag} */,
  {32'h4188fee8, 32'h41158c42} /* (22, 24, 25) {real, imag} */,
  {32'hc15614ca, 32'h414e72d1} /* (22, 24, 24) {real, imag} */,
  {32'hbf601f88, 32'hc11013b2} /* (22, 24, 23) {real, imag} */,
  {32'hbf859606, 32'hc18c7c12} /* (22, 24, 22) {real, imag} */,
  {32'h41a82a69, 32'h40c89583} /* (22, 24, 21) {real, imag} */,
  {32'hc139c91a, 32'hbf44632c} /* (22, 24, 20) {real, imag} */,
  {32'hc1499845, 32'h41123204} /* (22, 24, 19) {real, imag} */,
  {32'h40bc1594, 32'h4185fac3} /* (22, 24, 18) {real, imag} */,
  {32'hbff4420c, 32'hbfa8dc81} /* (22, 24, 17) {real, imag} */,
  {32'hc15a6224, 32'hc002520a} /* (22, 24, 16) {real, imag} */,
  {32'hbe30d948, 32'h40351b24} /* (22, 24, 15) {real, imag} */,
  {32'hc075c764, 32'h40ddb011} /* (22, 24, 14) {real, imag} */,
  {32'hc1276f60, 32'h40e5f2ac} /* (22, 24, 13) {real, imag} */,
  {32'hc0b17df2, 32'hc0572944} /* (22, 24, 12) {real, imag} */,
  {32'hc0ef5480, 32'hc1344aa6} /* (22, 24, 11) {real, imag} */,
  {32'hc151c784, 32'h41188649} /* (22, 24, 10) {real, imag} */,
  {32'h41559cda, 32'hbf9fd8fa} /* (22, 24, 9) {real, imag} */,
  {32'hc0e48a0e, 32'h41159480} /* (22, 24, 8) {real, imag} */,
  {32'h41188029, 32'hc1a3d7ea} /* (22, 24, 7) {real, imag} */,
  {32'h3f458ecc, 32'h408f167a} /* (22, 24, 6) {real, imag} */,
  {32'hc1f767f4, 32'h40fd2656} /* (22, 24, 5) {real, imag} */,
  {32'h40c234ba, 32'h4116adec} /* (22, 24, 4) {real, imag} */,
  {32'hbe58e480, 32'hc12a1da8} /* (22, 24, 3) {real, imag} */,
  {32'hc1a65f70, 32'h4062ef98} /* (22, 24, 2) {real, imag} */,
  {32'h4221e523, 32'hc1accf87} /* (22, 24, 1) {real, imag} */,
  {32'h41c836bc, 32'h3f4e39f0} /* (22, 24, 0) {real, imag} */,
  {32'hc13668f0, 32'h41b41f1c} /* (22, 23, 31) {real, imag} */,
  {32'h40dea2d2, 32'hc0f26056} /* (22, 23, 30) {real, imag} */,
  {32'h40dbe485, 32'hc1ba0f44} /* (22, 23, 29) {real, imag} */,
  {32'h416ceb87, 32'h402d917e} /* (22, 23, 28) {real, imag} */,
  {32'hbf963938, 32'h3ec57f20} /* (22, 23, 27) {real, imag} */,
  {32'hc1dbf7b6, 32'h40f9aab9} /* (22, 23, 26) {real, imag} */,
  {32'h41788d0a, 32'hbf807fa8} /* (22, 23, 25) {real, imag} */,
  {32'h418d77de, 32'hc19e6f9a} /* (22, 23, 24) {real, imag} */,
  {32'h4194c7b8, 32'h4191d592} /* (22, 23, 23) {real, imag} */,
  {32'hc03e2834, 32'hc0da4ff6} /* (22, 23, 22) {real, imag} */,
  {32'h406d52fa, 32'hbf69c8f8} /* (22, 23, 21) {real, imag} */,
  {32'h41046a88, 32'h4183578a} /* (22, 23, 20) {real, imag} */,
  {32'hc168021e, 32'hbfd3443c} /* (22, 23, 19) {real, imag} */,
  {32'h3f036740, 32'h4114e742} /* (22, 23, 18) {real, imag} */,
  {32'h4196e4d8, 32'hbf7e2078} /* (22, 23, 17) {real, imag} */,
  {32'hc074b04e, 32'hbf9cc73a} /* (22, 23, 16) {real, imag} */,
  {32'hc099be2f, 32'hc134fd80} /* (22, 23, 15) {real, imag} */,
  {32'hc04e4362, 32'hc0d67db9} /* (22, 23, 14) {real, imag} */,
  {32'h40217952, 32'h414b4666} /* (22, 23, 13) {real, imag} */,
  {32'h40a544ea, 32'hc076113c} /* (22, 23, 12) {real, imag} */,
  {32'hc1050f30, 32'hc0ab1c36} /* (22, 23, 11) {real, imag} */,
  {32'h410717e4, 32'hc192538c} /* (22, 23, 10) {real, imag} */,
  {32'hc08c2066, 32'h403f9dd8} /* (22, 23, 9) {real, imag} */,
  {32'h4103cfa6, 32'h4074f100} /* (22, 23, 8) {real, imag} */,
  {32'hc147a8e8, 32'h4182cae7} /* (22, 23, 7) {real, imag} */,
  {32'hc13526f1, 32'hc10a7080} /* (22, 23, 6) {real, imag} */,
  {32'h415d8f46, 32'hbf54d198} /* (22, 23, 5) {real, imag} */,
  {32'h3f44a8c0, 32'hc1e9db56} /* (22, 23, 4) {real, imag} */,
  {32'h3d7a0bc0, 32'h40da0497} /* (22, 23, 3) {real, imag} */,
  {32'h413617ae, 32'hc1a6955a} /* (22, 23, 2) {real, imag} */,
  {32'h4160f5a0, 32'h40f71154} /* (22, 23, 1) {real, imag} */,
  {32'h3cc4c380, 32'hc18778a3} /* (22, 23, 0) {real, imag} */,
  {32'hc175f9f3, 32'h41a6a64c} /* (22, 22, 31) {real, imag} */,
  {32'h404d29c4, 32'hc1a0ae24} /* (22, 22, 30) {real, imag} */,
  {32'h4139e037, 32'h4151bce4} /* (22, 22, 29) {real, imag} */,
  {32'h3fee6e53, 32'h40db33ef} /* (22, 22, 28) {real, imag} */,
  {32'hc133cdb6, 32'hc166d7e3} /* (22, 22, 27) {real, imag} */,
  {32'h3eb146a0, 32'hc1863872} /* (22, 22, 26) {real, imag} */,
  {32'hc0a3abc2, 32'h40d7ceb0} /* (22, 22, 25) {real, imag} */,
  {32'hc0bae46b, 32'hc097de57} /* (22, 22, 24) {real, imag} */,
  {32'hc084a6f4, 32'hc102639c} /* (22, 22, 23) {real, imag} */,
  {32'hc19b12a4, 32'hbffc0af0} /* (22, 22, 22) {real, imag} */,
  {32'hc112c0aa, 32'h40c3c5e1} /* (22, 22, 21) {real, imag} */,
  {32'hc0e52cec, 32'h4130e0db} /* (22, 22, 20) {real, imag} */,
  {32'h4139aa2b, 32'hc199c92d} /* (22, 22, 19) {real, imag} */,
  {32'hbfc03668, 32'hbd6cd400} /* (22, 22, 18) {real, imag} */,
  {32'h3f179c48, 32'h40a8a8a4} /* (22, 22, 17) {real, imag} */,
  {32'hc018b262, 32'h4013c91f} /* (22, 22, 16) {real, imag} */,
  {32'hc1047320, 32'h3ff136c2} /* (22, 22, 15) {real, imag} */,
  {32'h4002ef9a, 32'hc103d3db} /* (22, 22, 14) {real, imag} */,
  {32'hc0bd6bb0, 32'hbe626800} /* (22, 22, 13) {real, imag} */,
  {32'h41c09cb0, 32'hc01956f0} /* (22, 22, 12) {real, imag} */,
  {32'hc11ffd89, 32'h40b2bc9e} /* (22, 22, 11) {real, imag} */,
  {32'h40814a0c, 32'h413c4d40} /* (22, 22, 10) {real, imag} */,
  {32'hbfd300a0, 32'hbfac69a0} /* (22, 22, 9) {real, imag} */,
  {32'h41285826, 32'h3d907600} /* (22, 22, 8) {real, imag} */,
  {32'hc0c36150, 32'h4077c867} /* (22, 22, 7) {real, imag} */,
  {32'hc060b63e, 32'h4059f8fc} /* (22, 22, 6) {real, imag} */,
  {32'h3ff08c98, 32'h41831928} /* (22, 22, 5) {real, imag} */,
  {32'hc1244114, 32'h41332a8a} /* (22, 22, 4) {real, imag} */,
  {32'hc0328002, 32'h41acd678} /* (22, 22, 3) {real, imag} */,
  {32'hc1068551, 32'hc0c3a112} /* (22, 22, 2) {real, imag} */,
  {32'h401e6ff8, 32'h417a19cb} /* (22, 22, 1) {real, imag} */,
  {32'hbf984f34, 32'h4155420c} /* (22, 22, 0) {real, imag} */,
  {32'hbf9a2989, 32'hc1e24284} /* (22, 21, 31) {real, imag} */,
  {32'h3fdc9170, 32'h4065075c} /* (22, 21, 30) {real, imag} */,
  {32'hc0207cf0, 32'h40b0bf5f} /* (22, 21, 29) {real, imag} */,
  {32'h41046f58, 32'hc1990675} /* (22, 21, 28) {real, imag} */,
  {32'hc15951da, 32'hc17686e0} /* (22, 21, 27) {real, imag} */,
  {32'hc1d55511, 32'hc0b7e8a2} /* (22, 21, 26) {real, imag} */,
  {32'hc062cce0, 32'h409dc849} /* (22, 21, 25) {real, imag} */,
  {32'hc0336229, 32'h411e395e} /* (22, 21, 24) {real, imag} */,
  {32'hc089ca3e, 32'hc205e66c} /* (22, 21, 23) {real, imag} */,
  {32'hbff56f12, 32'hc0a8c722} /* (22, 21, 22) {real, imag} */,
  {32'hc1878182, 32'h40898eb0} /* (22, 21, 21) {real, imag} */,
  {32'h412db0d6, 32'hc1b0bc9a} /* (22, 21, 20) {real, imag} */,
  {32'hc0f2b125, 32'hc15bb445} /* (22, 21, 19) {real, imag} */,
  {32'h40c881dd, 32'hc0c1d402} /* (22, 21, 18) {real, imag} */,
  {32'hbfd6a005, 32'h3edbad90} /* (22, 21, 17) {real, imag} */,
  {32'hbec119d0, 32'hc0dca602} /* (22, 21, 16) {real, imag} */,
  {32'h411f54d3, 32'h4033f33e} /* (22, 21, 15) {real, imag} */,
  {32'hc11df448, 32'hc14f0619} /* (22, 21, 14) {real, imag} */,
  {32'h403cd7b1, 32'h3f0a09f8} /* (22, 21, 13) {real, imag} */,
  {32'h40d8c2f0, 32'hbf5f94f8} /* (22, 21, 12) {real, imag} */,
  {32'hc0b78b1d, 32'h40886bf8} /* (22, 21, 11) {real, imag} */,
  {32'hc1aeded1, 32'h402a374c} /* (22, 21, 10) {real, imag} */,
  {32'hc15c7b3b, 32'hc18aaa5a} /* (22, 21, 9) {real, imag} */,
  {32'h41045016, 32'hbfa3fe18} /* (22, 21, 8) {real, imag} */,
  {32'hc0b5202e, 32'hc194c302} /* (22, 21, 7) {real, imag} */,
  {32'h3ef69840, 32'hc1247110} /* (22, 21, 6) {real, imag} */,
  {32'hbf48fa24, 32'h419ed968} /* (22, 21, 5) {real, imag} */,
  {32'hc0d9efb1, 32'h408aa936} /* (22, 21, 4) {real, imag} */,
  {32'h408ed08e, 32'h3fee7294} /* (22, 21, 3) {real, imag} */,
  {32'hc0c746e0, 32'h41c4c023} /* (22, 21, 2) {real, imag} */,
  {32'h41003910, 32'hc110caa4} /* (22, 21, 1) {real, imag} */,
  {32'h40da7052, 32'hc13e6be2} /* (22, 21, 0) {real, imag} */,
  {32'hbf3f298e, 32'hc0231ea6} /* (22, 20, 31) {real, imag} */,
  {32'h40baa854, 32'h4098a69a} /* (22, 20, 30) {real, imag} */,
  {32'hbd52b340, 32'h4100f2cc} /* (22, 20, 29) {real, imag} */,
  {32'h40146c24, 32'h408905b5} /* (22, 20, 28) {real, imag} */,
  {32'h40db55b6, 32'hc1c7d110} /* (22, 20, 27) {real, imag} */,
  {32'h4090c3e9, 32'h400b20bb} /* (22, 20, 26) {real, imag} */,
  {32'hc0ca6606, 32'hc11005a0} /* (22, 20, 25) {real, imag} */,
  {32'hc0e120ba, 32'hc12137f2} /* (22, 20, 24) {real, imag} */,
  {32'h413bdccc, 32'h3eb5eb60} /* (22, 20, 23) {real, imag} */,
  {32'h411349cc, 32'hbfa69958} /* (22, 20, 22) {real, imag} */,
  {32'h405847ee, 32'hc0f963ff} /* (22, 20, 21) {real, imag} */,
  {32'h41659c80, 32'h41270fd3} /* (22, 20, 20) {real, imag} */,
  {32'hbf9a288c, 32'hc1323004} /* (22, 20, 19) {real, imag} */,
  {32'h40c89104, 32'h418a4ec4} /* (22, 20, 18) {real, imag} */,
  {32'hc004ee7e, 32'hc07d8a6d} /* (22, 20, 17) {real, imag} */,
  {32'hc08b9f53, 32'hbe6770a0} /* (22, 20, 16) {real, imag} */,
  {32'hbf01b850, 32'hc02c93da} /* (22, 20, 15) {real, imag} */,
  {32'hc1841030, 32'h3f5bb260} /* (22, 20, 14) {real, imag} */,
  {32'h40bf90a8, 32'h418066df} /* (22, 20, 13) {real, imag} */,
  {32'hc1132aa9, 32'hc111ab0d} /* (22, 20, 12) {real, imag} */,
  {32'h3fbaa90e, 32'h403ef578} /* (22, 20, 11) {real, imag} */,
  {32'h41ad47d4, 32'hc10d8bab} /* (22, 20, 10) {real, imag} */,
  {32'h41264c5f, 32'hc0274ef4} /* (22, 20, 9) {real, imag} */,
  {32'hc13b331b, 32'hbfbac208} /* (22, 20, 8) {real, imag} */,
  {32'h4126b59c, 32'hbf052550} /* (22, 20, 7) {real, imag} */,
  {32'hbf92a0ab, 32'hc0a87980} /* (22, 20, 6) {real, imag} */,
  {32'h3ff4ae70, 32'hc09f767e} /* (22, 20, 5) {real, imag} */,
  {32'hc08ab043, 32'h4106a182} /* (22, 20, 4) {real, imag} */,
  {32'h410d3a37, 32'hc08e0852} /* (22, 20, 3) {real, imag} */,
  {32'h4112e6c2, 32'hc1248bdd} /* (22, 20, 2) {real, imag} */,
  {32'hc1914350, 32'h40ca5c70} /* (22, 20, 1) {real, imag} */,
  {32'hbff8ad4c, 32'h40c70210} /* (22, 20, 0) {real, imag} */,
  {32'hc0b14100, 32'h410f3d34} /* (22, 19, 31) {real, imag} */,
  {32'h4131538c, 32'h4144299c} /* (22, 19, 30) {real, imag} */,
  {32'h41731b75, 32'h402e944b} /* (22, 19, 29) {real, imag} */,
  {32'hbe95eb20, 32'hc15858fd} /* (22, 19, 28) {real, imag} */,
  {32'hc19d1002, 32'h418f1c1a} /* (22, 19, 27) {real, imag} */,
  {32'h40fc1072, 32'hc01cc652} /* (22, 19, 26) {real, imag} */,
  {32'hc0187574, 32'h405fab3e} /* (22, 19, 25) {real, imag} */,
  {32'hc1314535, 32'hc08bf5d7} /* (22, 19, 24) {real, imag} */,
  {32'h40ef804a, 32'hc155309f} /* (22, 19, 23) {real, imag} */,
  {32'h4024dc1e, 32'hc0107e38} /* (22, 19, 22) {real, imag} */,
  {32'hc188bc3a, 32'hc049dec6} /* (22, 19, 21) {real, imag} */,
  {32'hc109523c, 32'h3fce48a8} /* (22, 19, 20) {real, imag} */,
  {32'hc114d4be, 32'h40c2a0b3} /* (22, 19, 19) {real, imag} */,
  {32'hc160ce38, 32'hc1000e17} /* (22, 19, 18) {real, imag} */,
  {32'hbf62bf8c, 32'hc13e36c6} /* (22, 19, 17) {real, imag} */,
  {32'h3fe8508d, 32'h41097fa4} /* (22, 19, 16) {real, imag} */,
  {32'hc09520c0, 32'hc02ff77c} /* (22, 19, 15) {real, imag} */,
  {32'h40175ead, 32'h413473ad} /* (22, 19, 14) {real, imag} */,
  {32'hc04d6036, 32'h4126c6cc} /* (22, 19, 13) {real, imag} */,
  {32'hc079fca0, 32'hbf86846a} /* (22, 19, 12) {real, imag} */,
  {32'h416b47ea, 32'hc0471e26} /* (22, 19, 11) {real, imag} */,
  {32'hc0891f76, 32'hc151736a} /* (22, 19, 10) {real, imag} */,
  {32'h4148e99e, 32'h417a423e} /* (22, 19, 9) {real, imag} */,
  {32'h4107601c, 32'hbef63180} /* (22, 19, 8) {real, imag} */,
  {32'hbed9d370, 32'hc1836c9f} /* (22, 19, 7) {real, imag} */,
  {32'hc0b31ccc, 32'hc1319a3f} /* (22, 19, 6) {real, imag} */,
  {32'h412d9cec, 32'h4148f865} /* (22, 19, 5) {real, imag} */,
  {32'hc157fe86, 32'hc0ee942a} /* (22, 19, 4) {real, imag} */,
  {32'hc182b3ad, 32'h40ad6a6c} /* (22, 19, 3) {real, imag} */,
  {32'hc1308ebf, 32'h410850e4} /* (22, 19, 2) {real, imag} */,
  {32'h4159f7e2, 32'h411ecddb} /* (22, 19, 1) {real, imag} */,
  {32'hc0814c90, 32'hc113c642} /* (22, 19, 0) {real, imag} */,
  {32'hc163b868, 32'hc1944b45} /* (22, 18, 31) {real, imag} */,
  {32'hc11d4bed, 32'hc08aa5ef} /* (22, 18, 30) {real, imag} */,
  {32'h41054de0, 32'h40a23bc4} /* (22, 18, 29) {real, imag} */,
  {32'hbf4bf5bc, 32'hc0dfd2fe} /* (22, 18, 28) {real, imag} */,
  {32'h40761a04, 32'h41199bf6} /* (22, 18, 27) {real, imag} */,
  {32'hc0cdd18e, 32'h416cdec0} /* (22, 18, 26) {real, imag} */,
  {32'hc150af6e, 32'h40aad8f6} /* (22, 18, 25) {real, imag} */,
  {32'h4143ccd7, 32'h3f323337} /* (22, 18, 24) {real, imag} */,
  {32'h3f113e6c, 32'hc0d8c696} /* (22, 18, 23) {real, imag} */,
  {32'hc1435194, 32'h4066e04c} /* (22, 18, 22) {real, imag} */,
  {32'hc07042ec, 32'hbfbc0da8} /* (22, 18, 21) {real, imag} */,
  {32'hc10c66ec, 32'h41a41999} /* (22, 18, 20) {real, imag} */,
  {32'hc1307f3c, 32'hc14777f2} /* (22, 18, 19) {real, imag} */,
  {32'h40aa3b1b, 32'hc123939a} /* (22, 18, 18) {real, imag} */,
  {32'h41034ab7, 32'hc1353bd4} /* (22, 18, 17) {real, imag} */,
  {32'h4052a88a, 32'hc073e58a} /* (22, 18, 16) {real, imag} */,
  {32'hc046e2b8, 32'h409c3470} /* (22, 18, 15) {real, imag} */,
  {32'hbf8f83c4, 32'hbef03258} /* (22, 18, 14) {real, imag} */,
  {32'hc1114e7d, 32'h40443ffa} /* (22, 18, 13) {real, imag} */,
  {32'h4055e85a, 32'hc156bdcd} /* (22, 18, 12) {real, imag} */,
  {32'hbf510c30, 32'hc05a6584} /* (22, 18, 11) {real, imag} */,
  {32'h41619a92, 32'h411c7aa4} /* (22, 18, 10) {real, imag} */,
  {32'hc0eaf2e9, 32'h4092c309} /* (22, 18, 9) {real, imag} */,
  {32'hc16f6275, 32'hbf7507b4} /* (22, 18, 8) {real, imag} */,
  {32'h4157cdca, 32'h41bf3b3a} /* (22, 18, 7) {real, imag} */,
  {32'h41182fe2, 32'h414071b4} /* (22, 18, 6) {real, imag} */,
  {32'h3ffaea97, 32'h413aca4a} /* (22, 18, 5) {real, imag} */,
  {32'h402348eb, 32'hc0b079c0} /* (22, 18, 4) {real, imag} */,
  {32'h4020255c, 32'h40ef72f5} /* (22, 18, 3) {real, imag} */,
  {32'hc1258f32, 32'h41832756} /* (22, 18, 2) {real, imag} */,
  {32'h3f9ff0c4, 32'hc093cfda} /* (22, 18, 1) {real, imag} */,
  {32'hc13d81dd, 32'hc183976a} /* (22, 18, 0) {real, imag} */,
  {32'hc125d50e, 32'h41365aa2} /* (22, 17, 31) {real, imag} */,
  {32'h40f9d3c4, 32'h40757818} /* (22, 17, 30) {real, imag} */,
  {32'hbee78170, 32'hbfc73a22} /* (22, 17, 29) {real, imag} */,
  {32'hbfbb6932, 32'h4121daeb} /* (22, 17, 28) {real, imag} */,
  {32'hc0b7cda5, 32'h41610e3c} /* (22, 17, 27) {real, imag} */,
  {32'hbfbf0512, 32'hc09e947e} /* (22, 17, 26) {real, imag} */,
  {32'h40852eb8, 32'hc0cb68c7} /* (22, 17, 25) {real, imag} */,
  {32'h41425e20, 32'h4039bcb2} /* (22, 17, 24) {real, imag} */,
  {32'hc0d7633f, 32'hbfa14494} /* (22, 17, 23) {real, imag} */,
  {32'hc1cb4da4, 32'hc1310cfd} /* (22, 17, 22) {real, imag} */,
  {32'hc0d1cd00, 32'h3ffa89d8} /* (22, 17, 21) {real, imag} */,
  {32'h419e4bf4, 32'hbffd180b} /* (22, 17, 20) {real, imag} */,
  {32'h40af5f65, 32'hc0c535e4} /* (22, 17, 19) {real, imag} */,
  {32'h409e5804, 32'hc15cb78e} /* (22, 17, 18) {real, imag} */,
  {32'h408ced19, 32'h3f3eae18} /* (22, 17, 17) {real, imag} */,
  {32'h3f965807, 32'h407f78ce} /* (22, 17, 16) {real, imag} */,
  {32'h40119180, 32'h3f38dc98} /* (22, 17, 15) {real, imag} */,
  {32'h402b4fc7, 32'h407959e8} /* (22, 17, 14) {real, imag} */,
  {32'h3f6f723c, 32'hc1a77284} /* (22, 17, 13) {real, imag} */,
  {32'hc17454c0, 32'h4102299e} /* (22, 17, 12) {real, imag} */,
  {32'h415572b2, 32'hc03f4ede} /* (22, 17, 11) {real, imag} */,
  {32'hc0d66142, 32'h40524d18} /* (22, 17, 10) {real, imag} */,
  {32'h411dfe92, 32'h3ebf0700} /* (22, 17, 9) {real, imag} */,
  {32'h4127402d, 32'hc0249580} /* (22, 17, 8) {real, imag} */,
  {32'h40ee22dd, 32'h4180adbe} /* (22, 17, 7) {real, imag} */,
  {32'hc0983b81, 32'h3d1f4d80} /* (22, 17, 6) {real, imag} */,
  {32'hc0f1bd51, 32'hbfb40f08} /* (22, 17, 5) {real, imag} */,
  {32'hc06ce1e4, 32'hbefe66d0} /* (22, 17, 4) {real, imag} */,
  {32'hc107bf94, 32'hc0380996} /* (22, 17, 3) {real, imag} */,
  {32'hc0cd3e52, 32'hc177e92c} /* (22, 17, 2) {real, imag} */,
  {32'h40aae46a, 32'hbe90d380} /* (22, 17, 1) {real, imag} */,
  {32'hc073f2b1, 32'hbefa2a88} /* (22, 17, 0) {real, imag} */,
  {32'h40c5dad2, 32'hc074aee8} /* (22, 16, 31) {real, imag} */,
  {32'h40a9db77, 32'h40d08986} /* (22, 16, 30) {real, imag} */,
  {32'hc043fad8, 32'h4114e719} /* (22, 16, 29) {real, imag} */,
  {32'hc053a227, 32'h402ce7da} /* (22, 16, 28) {real, imag} */,
  {32'h3d7556c0, 32'hbea4b968} /* (22, 16, 27) {real, imag} */,
  {32'h408d85a8, 32'h3f02b89a} /* (22, 16, 26) {real, imag} */,
  {32'hc0820115, 32'hbffb7207} /* (22, 16, 25) {real, imag} */,
  {32'h3fe2e398, 32'hc0e306ad} /* (22, 16, 24) {real, imag} */,
  {32'hc09dceaa, 32'h402b25c6} /* (22, 16, 23) {real, imag} */,
  {32'hc1493698, 32'h401755ac} /* (22, 16, 22) {real, imag} */,
  {32'h40c54cd6, 32'hc0ea132a} /* (22, 16, 21) {real, imag} */,
  {32'hc0cdb665, 32'h410704b5} /* (22, 16, 20) {real, imag} */,
  {32'h4055ba7b, 32'h40a3d5f0} /* (22, 16, 19) {real, imag} */,
  {32'h4153d9d6, 32'h411ab7be} /* (22, 16, 18) {real, imag} */,
  {32'hbf383838, 32'h3f5e4ca4} /* (22, 16, 17) {real, imag} */,
  {32'hc0d81f1d, 32'h00000000} /* (22, 16, 16) {real, imag} */,
  {32'hbf383838, 32'hbf5e4ca4} /* (22, 16, 15) {real, imag} */,
  {32'h4153d9d6, 32'hc11ab7be} /* (22, 16, 14) {real, imag} */,
  {32'h4055ba7b, 32'hc0a3d5f0} /* (22, 16, 13) {real, imag} */,
  {32'hc0cdb665, 32'hc10704b5} /* (22, 16, 12) {real, imag} */,
  {32'h40c54cd6, 32'h40ea132a} /* (22, 16, 11) {real, imag} */,
  {32'hc1493698, 32'hc01755ac} /* (22, 16, 10) {real, imag} */,
  {32'hc09dceaa, 32'hc02b25c6} /* (22, 16, 9) {real, imag} */,
  {32'h3fe2e398, 32'h40e306ad} /* (22, 16, 8) {real, imag} */,
  {32'hc0820115, 32'h3ffb7207} /* (22, 16, 7) {real, imag} */,
  {32'h408d85a8, 32'hbf02b89a} /* (22, 16, 6) {real, imag} */,
  {32'h3d7556c0, 32'h3ea4b968} /* (22, 16, 5) {real, imag} */,
  {32'hc053a227, 32'hc02ce7da} /* (22, 16, 4) {real, imag} */,
  {32'hc043fad8, 32'hc114e719} /* (22, 16, 3) {real, imag} */,
  {32'h40a9db77, 32'hc0d08986} /* (22, 16, 2) {real, imag} */,
  {32'h40c5dad2, 32'h4074aee8} /* (22, 16, 1) {real, imag} */,
  {32'h4177ec54, 32'h00000000} /* (22, 16, 0) {real, imag} */,
  {32'h40aae46a, 32'h3e90d380} /* (22, 15, 31) {real, imag} */,
  {32'hc0cd3e52, 32'h4177e92c} /* (22, 15, 30) {real, imag} */,
  {32'hc107bf94, 32'h40380996} /* (22, 15, 29) {real, imag} */,
  {32'hc06ce1e4, 32'h3efe66d0} /* (22, 15, 28) {real, imag} */,
  {32'hc0f1bd51, 32'h3fb40f08} /* (22, 15, 27) {real, imag} */,
  {32'hc0983b81, 32'hbd1f4d80} /* (22, 15, 26) {real, imag} */,
  {32'h40ee22dd, 32'hc180adbe} /* (22, 15, 25) {real, imag} */,
  {32'h4127402d, 32'h40249580} /* (22, 15, 24) {real, imag} */,
  {32'h411dfe92, 32'hbebf0700} /* (22, 15, 23) {real, imag} */,
  {32'hc0d66142, 32'hc0524d18} /* (22, 15, 22) {real, imag} */,
  {32'h415572b2, 32'h403f4ede} /* (22, 15, 21) {real, imag} */,
  {32'hc17454c0, 32'hc102299e} /* (22, 15, 20) {real, imag} */,
  {32'h3f6f723c, 32'h41a77284} /* (22, 15, 19) {real, imag} */,
  {32'h402b4fc7, 32'hc07959e8} /* (22, 15, 18) {real, imag} */,
  {32'h40119180, 32'hbf38dc98} /* (22, 15, 17) {real, imag} */,
  {32'h3f965807, 32'hc07f78ce} /* (22, 15, 16) {real, imag} */,
  {32'h408ced19, 32'hbf3eae18} /* (22, 15, 15) {real, imag} */,
  {32'h409e5804, 32'h415cb78e} /* (22, 15, 14) {real, imag} */,
  {32'h40af5f65, 32'h40c535e4} /* (22, 15, 13) {real, imag} */,
  {32'h419e4bf4, 32'h3ffd180b} /* (22, 15, 12) {real, imag} */,
  {32'hc0d1cd00, 32'hbffa89d8} /* (22, 15, 11) {real, imag} */,
  {32'hc1cb4da4, 32'h41310cfd} /* (22, 15, 10) {real, imag} */,
  {32'hc0d7633f, 32'h3fa14494} /* (22, 15, 9) {real, imag} */,
  {32'h41425e20, 32'hc039bcb2} /* (22, 15, 8) {real, imag} */,
  {32'h40852eb8, 32'h40cb68c7} /* (22, 15, 7) {real, imag} */,
  {32'hbfbf0512, 32'h409e947e} /* (22, 15, 6) {real, imag} */,
  {32'hc0b7cda5, 32'hc1610e3c} /* (22, 15, 5) {real, imag} */,
  {32'hbfbb6932, 32'hc121daeb} /* (22, 15, 4) {real, imag} */,
  {32'hbee78170, 32'h3fc73a22} /* (22, 15, 3) {real, imag} */,
  {32'h40f9d3c4, 32'hc0757818} /* (22, 15, 2) {real, imag} */,
  {32'hc125d50e, 32'hc1365aa2} /* (22, 15, 1) {real, imag} */,
  {32'hc073f2b1, 32'h3efa2a88} /* (22, 15, 0) {real, imag} */,
  {32'h3f9ff0c4, 32'h4093cfda} /* (22, 14, 31) {real, imag} */,
  {32'hc1258f32, 32'hc1832756} /* (22, 14, 30) {real, imag} */,
  {32'h4020255c, 32'hc0ef72f5} /* (22, 14, 29) {real, imag} */,
  {32'h402348eb, 32'h40b079c0} /* (22, 14, 28) {real, imag} */,
  {32'h3ffaea97, 32'hc13aca4a} /* (22, 14, 27) {real, imag} */,
  {32'h41182fe2, 32'hc14071b4} /* (22, 14, 26) {real, imag} */,
  {32'h4157cdca, 32'hc1bf3b3a} /* (22, 14, 25) {real, imag} */,
  {32'hc16f6275, 32'h3f7507b4} /* (22, 14, 24) {real, imag} */,
  {32'hc0eaf2e9, 32'hc092c309} /* (22, 14, 23) {real, imag} */,
  {32'h41619a92, 32'hc11c7aa4} /* (22, 14, 22) {real, imag} */,
  {32'hbf510c30, 32'h405a6584} /* (22, 14, 21) {real, imag} */,
  {32'h4055e85a, 32'h4156bdcd} /* (22, 14, 20) {real, imag} */,
  {32'hc1114e7d, 32'hc0443ffa} /* (22, 14, 19) {real, imag} */,
  {32'hbf8f83c4, 32'h3ef03258} /* (22, 14, 18) {real, imag} */,
  {32'hc046e2b8, 32'hc09c3470} /* (22, 14, 17) {real, imag} */,
  {32'h4052a88a, 32'h4073e58a} /* (22, 14, 16) {real, imag} */,
  {32'h41034ab7, 32'h41353bd4} /* (22, 14, 15) {real, imag} */,
  {32'h40aa3b1b, 32'h4123939a} /* (22, 14, 14) {real, imag} */,
  {32'hc1307f3c, 32'h414777f2} /* (22, 14, 13) {real, imag} */,
  {32'hc10c66ec, 32'hc1a41999} /* (22, 14, 12) {real, imag} */,
  {32'hc07042ec, 32'h3fbc0da8} /* (22, 14, 11) {real, imag} */,
  {32'hc1435194, 32'hc066e04c} /* (22, 14, 10) {real, imag} */,
  {32'h3f113e6c, 32'h40d8c696} /* (22, 14, 9) {real, imag} */,
  {32'h4143ccd7, 32'hbf323337} /* (22, 14, 8) {real, imag} */,
  {32'hc150af6e, 32'hc0aad8f6} /* (22, 14, 7) {real, imag} */,
  {32'hc0cdd18e, 32'hc16cdec0} /* (22, 14, 6) {real, imag} */,
  {32'h40761a04, 32'hc1199bf6} /* (22, 14, 5) {real, imag} */,
  {32'hbf4bf5bc, 32'h40dfd2fe} /* (22, 14, 4) {real, imag} */,
  {32'h41054de0, 32'hc0a23bc4} /* (22, 14, 3) {real, imag} */,
  {32'hc11d4bed, 32'h408aa5ef} /* (22, 14, 2) {real, imag} */,
  {32'hc163b868, 32'h41944b45} /* (22, 14, 1) {real, imag} */,
  {32'hc13d81dd, 32'h4183976a} /* (22, 14, 0) {real, imag} */,
  {32'h4159f7e2, 32'hc11ecddb} /* (22, 13, 31) {real, imag} */,
  {32'hc1308ebf, 32'hc10850e4} /* (22, 13, 30) {real, imag} */,
  {32'hc182b3ad, 32'hc0ad6a6c} /* (22, 13, 29) {real, imag} */,
  {32'hc157fe86, 32'h40ee942a} /* (22, 13, 28) {real, imag} */,
  {32'h412d9cec, 32'hc148f865} /* (22, 13, 27) {real, imag} */,
  {32'hc0b31ccc, 32'h41319a3f} /* (22, 13, 26) {real, imag} */,
  {32'hbed9d370, 32'h41836c9f} /* (22, 13, 25) {real, imag} */,
  {32'h4107601c, 32'h3ef63180} /* (22, 13, 24) {real, imag} */,
  {32'h4148e99e, 32'hc17a423e} /* (22, 13, 23) {real, imag} */,
  {32'hc0891f76, 32'h4151736a} /* (22, 13, 22) {real, imag} */,
  {32'h416b47ea, 32'h40471e26} /* (22, 13, 21) {real, imag} */,
  {32'hc079fca0, 32'h3f86846a} /* (22, 13, 20) {real, imag} */,
  {32'hc04d6036, 32'hc126c6cc} /* (22, 13, 19) {real, imag} */,
  {32'h40175ead, 32'hc13473ad} /* (22, 13, 18) {real, imag} */,
  {32'hc09520c0, 32'h402ff77c} /* (22, 13, 17) {real, imag} */,
  {32'h3fe8508d, 32'hc1097fa4} /* (22, 13, 16) {real, imag} */,
  {32'hbf62bf8c, 32'h413e36c6} /* (22, 13, 15) {real, imag} */,
  {32'hc160ce38, 32'h41000e17} /* (22, 13, 14) {real, imag} */,
  {32'hc114d4be, 32'hc0c2a0b3} /* (22, 13, 13) {real, imag} */,
  {32'hc109523c, 32'hbfce48a8} /* (22, 13, 12) {real, imag} */,
  {32'hc188bc3a, 32'h4049dec6} /* (22, 13, 11) {real, imag} */,
  {32'h4024dc1e, 32'h40107e38} /* (22, 13, 10) {real, imag} */,
  {32'h40ef804a, 32'h4155309f} /* (22, 13, 9) {real, imag} */,
  {32'hc1314535, 32'h408bf5d7} /* (22, 13, 8) {real, imag} */,
  {32'hc0187574, 32'hc05fab3e} /* (22, 13, 7) {real, imag} */,
  {32'h40fc1072, 32'h401cc652} /* (22, 13, 6) {real, imag} */,
  {32'hc19d1002, 32'hc18f1c1a} /* (22, 13, 5) {real, imag} */,
  {32'hbe95eb20, 32'h415858fd} /* (22, 13, 4) {real, imag} */,
  {32'h41731b75, 32'hc02e944b} /* (22, 13, 3) {real, imag} */,
  {32'h4131538c, 32'hc144299c} /* (22, 13, 2) {real, imag} */,
  {32'hc0b14100, 32'hc10f3d34} /* (22, 13, 1) {real, imag} */,
  {32'hc0814c90, 32'h4113c642} /* (22, 13, 0) {real, imag} */,
  {32'hc1914350, 32'hc0ca5c70} /* (22, 12, 31) {real, imag} */,
  {32'h4112e6c2, 32'h41248bdd} /* (22, 12, 30) {real, imag} */,
  {32'h410d3a37, 32'h408e0852} /* (22, 12, 29) {real, imag} */,
  {32'hc08ab043, 32'hc106a182} /* (22, 12, 28) {real, imag} */,
  {32'h3ff4ae70, 32'h409f767e} /* (22, 12, 27) {real, imag} */,
  {32'hbf92a0ab, 32'h40a87980} /* (22, 12, 26) {real, imag} */,
  {32'h4126b59c, 32'h3f052550} /* (22, 12, 25) {real, imag} */,
  {32'hc13b331b, 32'h3fbac208} /* (22, 12, 24) {real, imag} */,
  {32'h41264c5f, 32'h40274ef4} /* (22, 12, 23) {real, imag} */,
  {32'h41ad47d4, 32'h410d8bab} /* (22, 12, 22) {real, imag} */,
  {32'h3fbaa90e, 32'hc03ef578} /* (22, 12, 21) {real, imag} */,
  {32'hc1132aa9, 32'h4111ab0d} /* (22, 12, 20) {real, imag} */,
  {32'h40bf90a8, 32'hc18066df} /* (22, 12, 19) {real, imag} */,
  {32'hc1841030, 32'hbf5bb260} /* (22, 12, 18) {real, imag} */,
  {32'hbf01b850, 32'h402c93da} /* (22, 12, 17) {real, imag} */,
  {32'hc08b9f53, 32'h3e6770a0} /* (22, 12, 16) {real, imag} */,
  {32'hc004ee7e, 32'h407d8a6d} /* (22, 12, 15) {real, imag} */,
  {32'h40c89104, 32'hc18a4ec4} /* (22, 12, 14) {real, imag} */,
  {32'hbf9a288c, 32'h41323004} /* (22, 12, 13) {real, imag} */,
  {32'h41659c80, 32'hc1270fd3} /* (22, 12, 12) {real, imag} */,
  {32'h405847ee, 32'h40f963ff} /* (22, 12, 11) {real, imag} */,
  {32'h411349cc, 32'h3fa69958} /* (22, 12, 10) {real, imag} */,
  {32'h413bdccc, 32'hbeb5eb60} /* (22, 12, 9) {real, imag} */,
  {32'hc0e120ba, 32'h412137f2} /* (22, 12, 8) {real, imag} */,
  {32'hc0ca6606, 32'h411005a0} /* (22, 12, 7) {real, imag} */,
  {32'h4090c3e9, 32'hc00b20bb} /* (22, 12, 6) {real, imag} */,
  {32'h40db55b6, 32'h41c7d110} /* (22, 12, 5) {real, imag} */,
  {32'h40146c24, 32'hc08905b5} /* (22, 12, 4) {real, imag} */,
  {32'hbd52b340, 32'hc100f2cc} /* (22, 12, 3) {real, imag} */,
  {32'h40baa854, 32'hc098a69a} /* (22, 12, 2) {real, imag} */,
  {32'hbf3f298e, 32'h40231ea6} /* (22, 12, 1) {real, imag} */,
  {32'hbff8ad4c, 32'hc0c70210} /* (22, 12, 0) {real, imag} */,
  {32'h41003910, 32'h4110caa4} /* (22, 11, 31) {real, imag} */,
  {32'hc0c746e0, 32'hc1c4c023} /* (22, 11, 30) {real, imag} */,
  {32'h408ed08e, 32'hbfee7294} /* (22, 11, 29) {real, imag} */,
  {32'hc0d9efb1, 32'hc08aa936} /* (22, 11, 28) {real, imag} */,
  {32'hbf48fa24, 32'hc19ed968} /* (22, 11, 27) {real, imag} */,
  {32'h3ef69840, 32'h41247110} /* (22, 11, 26) {real, imag} */,
  {32'hc0b5202e, 32'h4194c302} /* (22, 11, 25) {real, imag} */,
  {32'h41045016, 32'h3fa3fe18} /* (22, 11, 24) {real, imag} */,
  {32'hc15c7b3b, 32'h418aaa5a} /* (22, 11, 23) {real, imag} */,
  {32'hc1aeded1, 32'hc02a374c} /* (22, 11, 22) {real, imag} */,
  {32'hc0b78b1d, 32'hc0886bf8} /* (22, 11, 21) {real, imag} */,
  {32'h40d8c2f0, 32'h3f5f94f8} /* (22, 11, 20) {real, imag} */,
  {32'h403cd7b1, 32'hbf0a09f8} /* (22, 11, 19) {real, imag} */,
  {32'hc11df448, 32'h414f0619} /* (22, 11, 18) {real, imag} */,
  {32'h411f54d3, 32'hc033f33e} /* (22, 11, 17) {real, imag} */,
  {32'hbec119d0, 32'h40dca602} /* (22, 11, 16) {real, imag} */,
  {32'hbfd6a005, 32'hbedbad90} /* (22, 11, 15) {real, imag} */,
  {32'h40c881dd, 32'h40c1d402} /* (22, 11, 14) {real, imag} */,
  {32'hc0f2b125, 32'h415bb445} /* (22, 11, 13) {real, imag} */,
  {32'h412db0d6, 32'h41b0bc9a} /* (22, 11, 12) {real, imag} */,
  {32'hc1878182, 32'hc0898eb0} /* (22, 11, 11) {real, imag} */,
  {32'hbff56f12, 32'h40a8c722} /* (22, 11, 10) {real, imag} */,
  {32'hc089ca3e, 32'h4205e66c} /* (22, 11, 9) {real, imag} */,
  {32'hc0336229, 32'hc11e395e} /* (22, 11, 8) {real, imag} */,
  {32'hc062cce0, 32'hc09dc849} /* (22, 11, 7) {real, imag} */,
  {32'hc1d55511, 32'h40b7e8a2} /* (22, 11, 6) {real, imag} */,
  {32'hc15951da, 32'h417686e0} /* (22, 11, 5) {real, imag} */,
  {32'h41046f58, 32'h41990675} /* (22, 11, 4) {real, imag} */,
  {32'hc0207cf0, 32'hc0b0bf5f} /* (22, 11, 3) {real, imag} */,
  {32'h3fdc9170, 32'hc065075c} /* (22, 11, 2) {real, imag} */,
  {32'hbf9a2989, 32'h41e24284} /* (22, 11, 1) {real, imag} */,
  {32'h40da7052, 32'h413e6be2} /* (22, 11, 0) {real, imag} */,
  {32'h401e6ff8, 32'hc17a19cb} /* (22, 10, 31) {real, imag} */,
  {32'hc1068551, 32'h40c3a112} /* (22, 10, 30) {real, imag} */,
  {32'hc0328002, 32'hc1acd678} /* (22, 10, 29) {real, imag} */,
  {32'hc1244114, 32'hc1332a8a} /* (22, 10, 28) {real, imag} */,
  {32'h3ff08c98, 32'hc1831928} /* (22, 10, 27) {real, imag} */,
  {32'hc060b63e, 32'hc059f8fc} /* (22, 10, 26) {real, imag} */,
  {32'hc0c36150, 32'hc077c867} /* (22, 10, 25) {real, imag} */,
  {32'h41285826, 32'hbd907600} /* (22, 10, 24) {real, imag} */,
  {32'hbfd300a0, 32'h3fac69a0} /* (22, 10, 23) {real, imag} */,
  {32'h40814a0c, 32'hc13c4d40} /* (22, 10, 22) {real, imag} */,
  {32'hc11ffd89, 32'hc0b2bc9e} /* (22, 10, 21) {real, imag} */,
  {32'h41c09cb0, 32'h401956f0} /* (22, 10, 20) {real, imag} */,
  {32'hc0bd6bb0, 32'h3e626800} /* (22, 10, 19) {real, imag} */,
  {32'h4002ef9a, 32'h4103d3db} /* (22, 10, 18) {real, imag} */,
  {32'hc1047320, 32'hbff136c2} /* (22, 10, 17) {real, imag} */,
  {32'hc018b262, 32'hc013c91f} /* (22, 10, 16) {real, imag} */,
  {32'h3f179c48, 32'hc0a8a8a4} /* (22, 10, 15) {real, imag} */,
  {32'hbfc03668, 32'h3d6cd400} /* (22, 10, 14) {real, imag} */,
  {32'h4139aa2b, 32'h4199c92d} /* (22, 10, 13) {real, imag} */,
  {32'hc0e52cec, 32'hc130e0db} /* (22, 10, 12) {real, imag} */,
  {32'hc112c0aa, 32'hc0c3c5e1} /* (22, 10, 11) {real, imag} */,
  {32'hc19b12a4, 32'h3ffc0af0} /* (22, 10, 10) {real, imag} */,
  {32'hc084a6f4, 32'h4102639c} /* (22, 10, 9) {real, imag} */,
  {32'hc0bae46b, 32'h4097de57} /* (22, 10, 8) {real, imag} */,
  {32'hc0a3abc2, 32'hc0d7ceb0} /* (22, 10, 7) {real, imag} */,
  {32'h3eb146a0, 32'h41863872} /* (22, 10, 6) {real, imag} */,
  {32'hc133cdb6, 32'h4166d7e3} /* (22, 10, 5) {real, imag} */,
  {32'h3fee6e53, 32'hc0db33ef} /* (22, 10, 4) {real, imag} */,
  {32'h4139e037, 32'hc151bce4} /* (22, 10, 3) {real, imag} */,
  {32'h404d29c4, 32'h41a0ae24} /* (22, 10, 2) {real, imag} */,
  {32'hc175f9f3, 32'hc1a6a64c} /* (22, 10, 1) {real, imag} */,
  {32'hbf984f34, 32'hc155420c} /* (22, 10, 0) {real, imag} */,
  {32'h4160f5a0, 32'hc0f71154} /* (22, 9, 31) {real, imag} */,
  {32'h413617ae, 32'h41a6955a} /* (22, 9, 30) {real, imag} */,
  {32'h3d7a0bc0, 32'hc0da0497} /* (22, 9, 29) {real, imag} */,
  {32'h3f44a8c0, 32'h41e9db56} /* (22, 9, 28) {real, imag} */,
  {32'h415d8f46, 32'h3f54d198} /* (22, 9, 27) {real, imag} */,
  {32'hc13526f1, 32'h410a7080} /* (22, 9, 26) {real, imag} */,
  {32'hc147a8e8, 32'hc182cae7} /* (22, 9, 25) {real, imag} */,
  {32'h4103cfa6, 32'hc074f100} /* (22, 9, 24) {real, imag} */,
  {32'hc08c2066, 32'hc03f9dd8} /* (22, 9, 23) {real, imag} */,
  {32'h410717e4, 32'h4192538c} /* (22, 9, 22) {real, imag} */,
  {32'hc1050f30, 32'h40ab1c36} /* (22, 9, 21) {real, imag} */,
  {32'h40a544ea, 32'h4076113c} /* (22, 9, 20) {real, imag} */,
  {32'h40217952, 32'hc14b4666} /* (22, 9, 19) {real, imag} */,
  {32'hc04e4362, 32'h40d67db9} /* (22, 9, 18) {real, imag} */,
  {32'hc099be2f, 32'h4134fd80} /* (22, 9, 17) {real, imag} */,
  {32'hc074b04e, 32'h3f9cc73a} /* (22, 9, 16) {real, imag} */,
  {32'h4196e4d8, 32'h3f7e2078} /* (22, 9, 15) {real, imag} */,
  {32'h3f036740, 32'hc114e742} /* (22, 9, 14) {real, imag} */,
  {32'hc168021e, 32'h3fd3443c} /* (22, 9, 13) {real, imag} */,
  {32'h41046a88, 32'hc183578a} /* (22, 9, 12) {real, imag} */,
  {32'h406d52fa, 32'h3f69c8f8} /* (22, 9, 11) {real, imag} */,
  {32'hc03e2834, 32'h40da4ff6} /* (22, 9, 10) {real, imag} */,
  {32'h4194c7b8, 32'hc191d592} /* (22, 9, 9) {real, imag} */,
  {32'h418d77de, 32'h419e6f9a} /* (22, 9, 8) {real, imag} */,
  {32'h41788d0a, 32'h3f807fa8} /* (22, 9, 7) {real, imag} */,
  {32'hc1dbf7b6, 32'hc0f9aab9} /* (22, 9, 6) {real, imag} */,
  {32'hbf963938, 32'hbec57f20} /* (22, 9, 5) {real, imag} */,
  {32'h416ceb87, 32'hc02d917e} /* (22, 9, 4) {real, imag} */,
  {32'h40dbe485, 32'h41ba0f44} /* (22, 9, 3) {real, imag} */,
  {32'h40dea2d2, 32'h40f26056} /* (22, 9, 2) {real, imag} */,
  {32'hc13668f0, 32'hc1b41f1c} /* (22, 9, 1) {real, imag} */,
  {32'h3cc4c380, 32'h418778a3} /* (22, 9, 0) {real, imag} */,
  {32'h4221e523, 32'h41accf87} /* (22, 8, 31) {real, imag} */,
  {32'hc1a65f70, 32'hc062ef98} /* (22, 8, 30) {real, imag} */,
  {32'hbe58e480, 32'h412a1da8} /* (22, 8, 29) {real, imag} */,
  {32'h40c234ba, 32'hc116adec} /* (22, 8, 28) {real, imag} */,
  {32'hc1f767f4, 32'hc0fd2656} /* (22, 8, 27) {real, imag} */,
  {32'h3f458ecc, 32'hc08f167a} /* (22, 8, 26) {real, imag} */,
  {32'h41188029, 32'h41a3d7ea} /* (22, 8, 25) {real, imag} */,
  {32'hc0e48a0e, 32'hc1159480} /* (22, 8, 24) {real, imag} */,
  {32'h41559cda, 32'h3f9fd8fa} /* (22, 8, 23) {real, imag} */,
  {32'hc151c784, 32'hc1188649} /* (22, 8, 22) {real, imag} */,
  {32'hc0ef5480, 32'h41344aa6} /* (22, 8, 21) {real, imag} */,
  {32'hc0b17df2, 32'h40572944} /* (22, 8, 20) {real, imag} */,
  {32'hc1276f60, 32'hc0e5f2ac} /* (22, 8, 19) {real, imag} */,
  {32'hc075c764, 32'hc0ddb011} /* (22, 8, 18) {real, imag} */,
  {32'hbe30d948, 32'hc0351b24} /* (22, 8, 17) {real, imag} */,
  {32'hc15a6224, 32'h4002520a} /* (22, 8, 16) {real, imag} */,
  {32'hbff4420c, 32'h3fa8dc81} /* (22, 8, 15) {real, imag} */,
  {32'h40bc1594, 32'hc185fac3} /* (22, 8, 14) {real, imag} */,
  {32'hc1499845, 32'hc1123204} /* (22, 8, 13) {real, imag} */,
  {32'hc139c91a, 32'h3f44632c} /* (22, 8, 12) {real, imag} */,
  {32'h41a82a69, 32'hc0c89583} /* (22, 8, 11) {real, imag} */,
  {32'hbf859606, 32'h418c7c12} /* (22, 8, 10) {real, imag} */,
  {32'hbf601f88, 32'h411013b2} /* (22, 8, 9) {real, imag} */,
  {32'hc15614ca, 32'hc14e72d1} /* (22, 8, 8) {real, imag} */,
  {32'h4188fee8, 32'hc1158c42} /* (22, 8, 7) {real, imag} */,
  {32'h400450a6, 32'h40445bfa} /* (22, 8, 6) {real, imag} */,
  {32'hc1c3f168, 32'hc114d480} /* (22, 8, 5) {real, imag} */,
  {32'h416855cc, 32'h41974d68} /* (22, 8, 4) {real, imag} */,
  {32'h3f975e78, 32'hc141ca30} /* (22, 8, 3) {real, imag} */,
  {32'hc08acbbc, 32'h40325fbc} /* (22, 8, 2) {real, imag} */,
  {32'h3fb09408, 32'h4100b8d0} /* (22, 8, 1) {real, imag} */,
  {32'h41c836bc, 32'hbf4e39f0} /* (22, 8, 0) {real, imag} */,
  {32'hc1ab9732, 32'hc1994f12} /* (22, 7, 31) {real, imag} */,
  {32'h41138f8e, 32'h404cb8a4} /* (22, 7, 30) {real, imag} */,
  {32'h41accc00, 32'h40ec65aa} /* (22, 7, 29) {real, imag} */,
  {32'h4198ee7e, 32'h4144ac83} /* (22, 7, 28) {real, imag} */,
  {32'hc00dff9c, 32'h40511860} /* (22, 7, 27) {real, imag} */,
  {32'hc1323ec0, 32'h4148946c} /* (22, 7, 26) {real, imag} */,
  {32'h40b51048, 32'h3ed960d0} /* (22, 7, 25) {real, imag} */,
  {32'hc1fede80, 32'h4058fada} /* (22, 7, 24) {real, imag} */,
  {32'h416cc39c, 32'h411bb4c1} /* (22, 7, 23) {real, imag} */,
  {32'hc0f33b7f, 32'hc04a8c68} /* (22, 7, 22) {real, imag} */,
  {32'h41525f6f, 32'hbfb22162} /* (22, 7, 21) {real, imag} */,
  {32'h3f9dd128, 32'hc18737ad} /* (22, 7, 20) {real, imag} */,
  {32'hc17f67d8, 32'h40ea6ede} /* (22, 7, 19) {real, imag} */,
  {32'h410a371e, 32'hbfda6f24} /* (22, 7, 18) {real, imag} */,
  {32'h410df84d, 32'hc0e53efa} /* (22, 7, 17) {real, imag} */,
  {32'h4089a110, 32'h40afb7e3} /* (22, 7, 16) {real, imag} */,
  {32'h3fbda130, 32'h410cc1ed} /* (22, 7, 15) {real, imag} */,
  {32'hc0d31a67, 32'h3e02df40} /* (22, 7, 14) {real, imag} */,
  {32'h403f3eb6, 32'h4039a450} /* (22, 7, 13) {real, imag} */,
  {32'hc08dfb04, 32'h40e2de5c} /* (22, 7, 12) {real, imag} */,
  {32'hc1c12ec4, 32'h3f79bcb8} /* (22, 7, 11) {real, imag} */,
  {32'hc1241624, 32'h41244048} /* (22, 7, 10) {real, imag} */,
  {32'hc058415e, 32'hbfa84cfc} /* (22, 7, 9) {real, imag} */,
  {32'h40c69615, 32'hc15a709b} /* (22, 7, 8) {real, imag} */,
  {32'hc0a3cd84, 32'hc1fb595c} /* (22, 7, 7) {real, imag} */,
  {32'h410207e4, 32'h40adbc15} /* (22, 7, 6) {real, imag} */,
  {32'h409be992, 32'h410778ad} /* (22, 7, 5) {real, imag} */,
  {32'h3f547e88, 32'hc1556654} /* (22, 7, 4) {real, imag} */,
  {32'h413a04ed, 32'h4217fc00} /* (22, 7, 3) {real, imag} */,
  {32'hc118243d, 32'hc1123a1f} /* (22, 7, 2) {real, imag} */,
  {32'hc07e6088, 32'hc19a0693} /* (22, 7, 1) {real, imag} */,
  {32'hc09c0135, 32'hc1886aca} /* (22, 7, 0) {real, imag} */,
  {32'h411730e6, 32'h40f0ccd4} /* (22, 6, 31) {real, imag} */,
  {32'hc0daba98, 32'hc0de9f77} /* (22, 6, 30) {real, imag} */,
  {32'h40d784e1, 32'h415bcf7c} /* (22, 6, 29) {real, imag} */,
  {32'hc00926ec, 32'hc1ac5217} /* (22, 6, 28) {real, imag} */,
  {32'hc055aec8, 32'hc0bd3122} /* (22, 6, 27) {real, imag} */,
  {32'hc1955776, 32'h41045686} /* (22, 6, 26) {real, imag} */,
  {32'hc10cae06, 32'hbed58d18} /* (22, 6, 25) {real, imag} */,
  {32'h41027f05, 32'hc163b4f2} /* (22, 6, 24) {real, imag} */,
  {32'hc15ec086, 32'h40427e68} /* (22, 6, 23) {real, imag} */,
  {32'hc09d2bd2, 32'h4180d7e6} /* (22, 6, 22) {real, imag} */,
  {32'hbf0a1560, 32'hc0cfb4f0} /* (22, 6, 21) {real, imag} */,
  {32'hc0831127, 32'hc0f61efd} /* (22, 6, 20) {real, imag} */,
  {32'hc00ff1e4, 32'h4146abe1} /* (22, 6, 19) {real, imag} */,
  {32'hc02a1d7a, 32'h409ca880} /* (22, 6, 18) {real, imag} */,
  {32'h3fb89124, 32'hc0f0202a} /* (22, 6, 17) {real, imag} */,
  {32'hc09e9fb3, 32'h402735e0} /* (22, 6, 16) {real, imag} */,
  {32'hc0bd2b0a, 32'h40e2332f} /* (22, 6, 15) {real, imag} */,
  {32'hc0f934d4, 32'h4121719e} /* (22, 6, 14) {real, imag} */,
  {32'h4108d128, 32'h4016f279} /* (22, 6, 13) {real, imag} */,
  {32'h410f0d5f, 32'h416b3741} /* (22, 6, 12) {real, imag} */,
  {32'hc1237747, 32'h40ca14f6} /* (22, 6, 11) {real, imag} */,
  {32'hc19c00b5, 32'h3f43dbf0} /* (22, 6, 10) {real, imag} */,
  {32'h408b95f7, 32'hc02cae22} /* (22, 6, 9) {real, imag} */,
  {32'h40b48b03, 32'hc11f0ce4} /* (22, 6, 8) {real, imag} */,
  {32'hc1703075, 32'hc0f35a2e} /* (22, 6, 7) {real, imag} */,
  {32'hc0a85a07, 32'hc1823415} /* (22, 6, 6) {real, imag} */,
  {32'hc1c8a185, 32'h40fbd728} /* (22, 6, 5) {real, imag} */,
  {32'h41045c35, 32'h3fadbb34} /* (22, 6, 4) {real, imag} */,
  {32'h41be9294, 32'hc20208b2} /* (22, 6, 3) {real, imag} */,
  {32'hc19c8e86, 32'h4038636c} /* (22, 6, 2) {real, imag} */,
  {32'h4146bbf4, 32'h40d9f576} /* (22, 6, 1) {real, imag} */,
  {32'h3f5057f0, 32'h412e6960} /* (22, 6, 0) {real, imag} */,
  {32'h42c21804, 32'h41cd22ba} /* (22, 5, 31) {real, imag} */,
  {32'hc27955d3, 32'hc170a908} /* (22, 5, 30) {real, imag} */,
  {32'hc0121dbf, 32'hc0b32cc4} /* (22, 5, 29) {real, imag} */,
  {32'hc177b875, 32'hc070f3e8} /* (22, 5, 28) {real, imag} */,
  {32'hc2181e7b, 32'hc04a6d3a} /* (22, 5, 27) {real, imag} */,
  {32'hbfd3cf8a, 32'h41b48a86} /* (22, 5, 26) {real, imag} */,
  {32'hc0b9983c, 32'hc0cead34} /* (22, 5, 25) {real, imag} */,
  {32'hc149f456, 32'h3fdbddd0} /* (22, 5, 24) {real, imag} */,
  {32'h41094d30, 32'hc18040d8} /* (22, 5, 23) {real, imag} */,
  {32'hc1aaa39b, 32'h40ebd3de} /* (22, 5, 22) {real, imag} */,
  {32'hc021cc62, 32'h3ff71508} /* (22, 5, 21) {real, imag} */,
  {32'h41063ef1, 32'hc1812952} /* (22, 5, 20) {real, imag} */,
  {32'h40b45590, 32'hc0a77a51} /* (22, 5, 19) {real, imag} */,
  {32'h41405570, 32'h3e810700} /* (22, 5, 18) {real, imag} */,
  {32'h3fcbfbe1, 32'hc02ad196} /* (22, 5, 17) {real, imag} */,
  {32'hc16a741c, 32'hc1143956} /* (22, 5, 16) {real, imag} */,
  {32'hc01ba87c, 32'h40c240c8} /* (22, 5, 15) {real, imag} */,
  {32'h4131207a, 32'hc0c04c78} /* (22, 5, 14) {real, imag} */,
  {32'h414e23aa, 32'hc0ab34ff} /* (22, 5, 13) {real, imag} */,
  {32'hc156c29c, 32'hc0d8ed0f} /* (22, 5, 12) {real, imag} */,
  {32'hc0ada160, 32'hc1816d7c} /* (22, 5, 11) {real, imag} */,
  {32'hc0a91a7e, 32'hc134a42a} /* (22, 5, 10) {real, imag} */,
  {32'h40c5c1b3, 32'hbeaeb738} /* (22, 5, 9) {real, imag} */,
  {32'hbfb48140, 32'hbe547800} /* (22, 5, 8) {real, imag} */,
  {32'h411ca0d2, 32'hbf95b224} /* (22, 5, 7) {real, imag} */,
  {32'h4143ae9a, 32'h4009e92a} /* (22, 5, 6) {real, imag} */,
  {32'hc118e420, 32'hc1ba9662} /* (22, 5, 5) {real, imag} */,
  {32'hc1260f44, 32'h423f19b2} /* (22, 5, 4) {real, imag} */,
  {32'hc027484b, 32'hc0a225be} /* (22, 5, 3) {real, imag} */,
  {32'h40d77095, 32'hc22206a0} /* (22, 5, 2) {real, imag} */,
  {32'h42c3ee42, 32'h42bcd575} /* (22, 5, 1) {real, imag} */,
  {32'h428e3266, 32'h4221a283} /* (22, 5, 0) {real, imag} */,
  {32'hc20ac486, 32'hc2caa144} /* (22, 4, 31) {real, imag} */,
  {32'h42acce27, 32'h42a58a7e} /* (22, 4, 30) {real, imag} */,
  {32'hc1d6fa5a, 32'h40cf89b1} /* (22, 4, 29) {real, imag} */,
  {32'hc1a7e602, 32'hc0c31b48} /* (22, 4, 28) {real, imag} */,
  {32'h414c0331, 32'hc13e7112} /* (22, 4, 27) {real, imag} */,
  {32'h409b4b7e, 32'hc1230b76} /* (22, 4, 26) {real, imag} */,
  {32'h411272a0, 32'hc0a4770b} /* (22, 4, 25) {real, imag} */,
  {32'h41942800, 32'h4154c1ee} /* (22, 4, 24) {real, imag} */,
  {32'hc119c65e, 32'hc16ad1b3} /* (22, 4, 23) {real, imag} */,
  {32'hc0856abc, 32'h40b277ee} /* (22, 4, 22) {real, imag} */,
  {32'hc1299460, 32'h41326464} /* (22, 4, 21) {real, imag} */,
  {32'h3f79ade8, 32'hc05f8728} /* (22, 4, 20) {real, imag} */,
  {32'hbf240991, 32'h405c9c43} /* (22, 4, 19) {real, imag} */,
  {32'h417568e6, 32'hc0f9c769} /* (22, 4, 18) {real, imag} */,
  {32'hbda12eb8, 32'hbf1a0f30} /* (22, 4, 17) {real, imag} */,
  {32'hc070b3f8, 32'h40199a83} /* (22, 4, 16) {real, imag} */,
  {32'hc08239bd, 32'h402717d0} /* (22, 4, 15) {real, imag} */,
  {32'h414e3398, 32'h40642fb5} /* (22, 4, 14) {real, imag} */,
  {32'hc0fd0c50, 32'h40cb30e0} /* (22, 4, 13) {real, imag} */,
  {32'hc0c62c98, 32'hc19dd60a} /* (22, 4, 12) {real, imag} */,
  {32'h41388ff7, 32'h41730493} /* (22, 4, 11) {real, imag} */,
  {32'hbf512900, 32'h417dd395} /* (22, 4, 10) {real, imag} */,
  {32'h40ecd5c7, 32'hc0c956e1} /* (22, 4, 9) {real, imag} */,
  {32'h418529ee, 32'hc0ac7a72} /* (22, 4, 8) {real, imag} */,
  {32'hc09adeb2, 32'hbed728f0} /* (22, 4, 7) {real, imag} */,
  {32'hc171bdc2, 32'hc030a72c} /* (22, 4, 6) {real, imag} */,
  {32'h402f07ec, 32'h400149b0} /* (22, 4, 5) {real, imag} */,
  {32'h418fd021, 32'hc21d48d5} /* (22, 4, 4) {real, imag} */,
  {32'h41273f7a, 32'hc107b3df} /* (22, 4, 3) {real, imag} */,
  {32'h42d9f190, 32'h4284598b} /* (22, 4, 2) {real, imag} */,
  {32'hc2e8461e, 32'hc214eb4a} /* (22, 4, 1) {real, imag} */,
  {32'hc2a687b2, 32'h41d23d72} /* (22, 4, 0) {real, imag} */,
  {32'h43128d49, 32'hc28e305d} /* (22, 3, 31) {real, imag} */,
  {32'hc2be7f5b, 32'h42db40fa} /* (22, 3, 30) {real, imag} */,
  {32'hc0216f84, 32'hc08ddfa6} /* (22, 3, 29) {real, imag} */,
  {32'hc26afca8, 32'hc1fa9d50} /* (22, 3, 28) {real, imag} */,
  {32'h41a99642, 32'h40f385f4} /* (22, 3, 27) {real, imag} */,
  {32'h4093ddb4, 32'hc08605e2} /* (22, 3, 26) {real, imag} */,
  {32'h41131b8f, 32'hc199069b} /* (22, 3, 25) {real, imag} */,
  {32'h41c94744, 32'h40c34ee3} /* (22, 3, 24) {real, imag} */,
  {32'hc0714d3c, 32'hc177f472} /* (22, 3, 23) {real, imag} */,
  {32'hc140f862, 32'hc139b9e8} /* (22, 3, 22) {real, imag} */,
  {32'hbe7d4e98, 32'h40df7e68} /* (22, 3, 21) {real, imag} */,
  {32'h412cb868, 32'hc124bee4} /* (22, 3, 20) {real, imag} */,
  {32'h411e469c, 32'h4117baa7} /* (22, 3, 19) {real, imag} */,
  {32'h41484e6e, 32'h402a3cf0} /* (22, 3, 18) {real, imag} */,
  {32'hc0b893e3, 32'h40924c06} /* (22, 3, 17) {real, imag} */,
  {32'h40a52e0e, 32'hc0bc638a} /* (22, 3, 16) {real, imag} */,
  {32'hc12d7de3, 32'hbff95bc0} /* (22, 3, 15) {real, imag} */,
  {32'hc1288d5a, 32'h3fd6ae3c} /* (22, 3, 14) {real, imag} */,
  {32'h40560d7b, 32'h4123a702} /* (22, 3, 13) {real, imag} */,
  {32'h41a0bde2, 32'hc0958254} /* (22, 3, 12) {real, imag} */,
  {32'hc10190a6, 32'h3fe0d310} /* (22, 3, 11) {real, imag} */,
  {32'hc118ca58, 32'h41ab1016} /* (22, 3, 10) {real, imag} */,
  {32'hc12c692c, 32'hc18d3c98} /* (22, 3, 9) {real, imag} */,
  {32'hc158a89a, 32'h417847e9} /* (22, 3, 8) {real, imag} */,
  {32'h40ef066d, 32'hc100565c} /* (22, 3, 7) {real, imag} */,
  {32'h41716600, 32'h40416bda} /* (22, 3, 6) {real, imag} */,
  {32'hc1bd52a3, 32'hc0e1d01e} /* (22, 3, 5) {real, imag} */,
  {32'h41dc5fce, 32'hc27481d2} /* (22, 3, 4) {real, imag} */,
  {32'h40309af0, 32'hc1a6b081} /* (22, 3, 3) {real, imag} */,
  {32'hc18e3b76, 32'h430959f0} /* (22, 3, 2) {real, imag} */,
  {32'hc304234c, 32'hc2abcd6e} /* (22, 3, 1) {real, imag} */,
  {32'h42850126, 32'hbf045a60} /* (22, 3, 0) {real, imag} */,
  {32'h449cedcb, 32'h42199956} /* (22, 2, 31) {real, imag} */,
  {32'hc40ac138, 32'h43504f88} /* (22, 2, 30) {real, imag} */,
  {32'hc085e878, 32'hc1b1d48c} /* (22, 2, 29) {real, imag} */,
  {32'h420fa701, 32'hc2c43e52} /* (22, 2, 28) {real, imag} */,
  {32'hc25e244b, 32'h41e9443b} /* (22, 2, 27) {real, imag} */,
  {32'hc21428ad, 32'hc0b43f0c} /* (22, 2, 26) {real, imag} */,
  {32'h41e23c04, 32'hc1620bc2} /* (22, 2, 25) {real, imag} */,
  {32'hc12bd461, 32'h410ba84c} /* (22, 2, 24) {real, imag} */,
  {32'hc1086ef7, 32'hc1058c64} /* (22, 2, 23) {real, imag} */,
  {32'hc05e7c60, 32'h412cb5f8} /* (22, 2, 22) {real, imag} */,
  {32'h3ff429b4, 32'h41106ed8} /* (22, 2, 21) {real, imag} */,
  {32'h412646c0, 32'h41278714} /* (22, 2, 20) {real, imag} */,
  {32'hc1926ad2, 32'h41630a28} /* (22, 2, 19) {real, imag} */,
  {32'hc052c0c6, 32'h415f3a92} /* (22, 2, 18) {real, imag} */,
  {32'h39b68000, 32'hc0dd188a} /* (22, 2, 17) {real, imag} */,
  {32'h3fa16b7e, 32'hbe81b444} /* (22, 2, 16) {real, imag} */,
  {32'hbf9b4978, 32'h4032ef32} /* (22, 2, 15) {real, imag} */,
  {32'h415c3672, 32'h401cd974} /* (22, 2, 14) {real, imag} */,
  {32'h413d8a8e, 32'h40ba691a} /* (22, 2, 13) {real, imag} */,
  {32'hc15b1b2a, 32'hc187bac5} /* (22, 2, 12) {real, imag} */,
  {32'hc092b6b3, 32'hc1a96855} /* (22, 2, 11) {real, imag} */,
  {32'h4159f63e, 32'h41b283f3} /* (22, 2, 10) {real, imag} */,
  {32'h4089fac1, 32'hbfc8fcfc} /* (22, 2, 9) {real, imag} */,
  {32'hc1ab67ca, 32'hc1905571} /* (22, 2, 8) {real, imag} */,
  {32'h3f5f1538, 32'hc049f334} /* (22, 2, 7) {real, imag} */,
  {32'hc0e2859a, 32'h415ce178} /* (22, 2, 6) {real, imag} */,
  {32'hc2a34c60, 32'hc2903032} /* (22, 2, 5) {real, imag} */,
  {32'h42c03adf, 32'h428b6ee7} /* (22, 2, 4) {real, imag} */,
  {32'h40a6fc6c, 32'hc236204b} /* (22, 2, 3) {real, imag} */,
  {32'hc3cd8aca, 32'h42b61d12} /* (22, 2, 2) {real, imag} */,
  {32'h44339153, 32'hc2a62180} /* (22, 2, 1) {real, imag} */,
  {32'h441f47b8, 32'h4309dc98} /* (22, 2, 0) {real, imag} */,
  {32'hc4d5cc2b, 32'h43e59299} /* (22, 1, 31) {real, imag} */,
  {32'h43e49f0c, 32'h42aa096e} /* (22, 1, 30) {real, imag} */,
  {32'h41dc9d48, 32'hc2892b77} /* (22, 1, 29) {real, imag} */,
  {32'hc30cdf8f, 32'hc282e392} /* (22, 1, 28) {real, imag} */,
  {32'h430f695e, 32'hc11fe67f} /* (22, 1, 27) {real, imag} */,
  {32'h41d6bc25, 32'hc0542674} /* (22, 1, 26) {real, imag} */,
  {32'hc18ec39c, 32'hc14895c4} /* (22, 1, 25) {real, imag} */,
  {32'h4179f2c4, 32'hc15d731e} /* (22, 1, 24) {real, imag} */,
  {32'h4171c55c, 32'hc1cfefc6} /* (22, 1, 23) {real, imag} */,
  {32'h412eb0bd, 32'hc10304c3} /* (22, 1, 22) {real, imag} */,
  {32'h40fe650b, 32'h40f91436} /* (22, 1, 21) {real, imag} */,
  {32'h40cdcde5, 32'hc0da1ffa} /* (22, 1, 20) {real, imag} */,
  {32'h40208910, 32'hc0d1ebb4} /* (22, 1, 19) {real, imag} */,
  {32'h409ab3ec, 32'h4109683a} /* (22, 1, 18) {real, imag} */,
  {32'hc08e4226, 32'h4072ac55} /* (22, 1, 17) {real, imag} */,
  {32'h40ad62ce, 32'hc098e40c} /* (22, 1, 16) {real, imag} */,
  {32'hc090964e, 32'h4123f154} /* (22, 1, 15) {real, imag} */,
  {32'h3ed43330, 32'h41628776} /* (22, 1, 14) {real, imag} */,
  {32'hc16ed590, 32'hc0c06d60} /* (22, 1, 13) {real, imag} */,
  {32'h4118f52a, 32'h4090004c} /* (22, 1, 12) {real, imag} */,
  {32'h4183ab84, 32'h40ccfb0d} /* (22, 1, 11) {real, imag} */,
  {32'hc139412a, 32'h414f3ee7} /* (22, 1, 10) {real, imag} */,
  {32'h40cc8ed1, 32'hc145d99d} /* (22, 1, 9) {real, imag} */,
  {32'h4099a629, 32'h423cd0a4} /* (22, 1, 8) {real, imag} */,
  {32'hc14586a9, 32'hc22dcd14} /* (22, 1, 7) {real, imag} */,
  {32'hc081a2c4, 32'hc0c959ba} /* (22, 1, 6) {real, imag} */,
  {32'h42887c97, 32'h426006c1} /* (22, 1, 5) {real, imag} */,
  {32'hc25493e2, 32'hc28f9744} /* (22, 1, 4) {real, imag} */,
  {32'h42856b01, 32'h41c10cc4} /* (22, 1, 3) {real, imag} */,
  {32'h44100e9d, 32'h440e30d7} /* (22, 1, 2) {real, imag} */,
  {32'hc5188d2b, 32'hc4a3f327} /* (22, 1, 1) {real, imag} */,
  {32'hc506879a, 32'hc3971b6c} /* (22, 1, 0) {real, imag} */,
  {32'hc4c03ee8, 32'h44995acc} /* (22, 0, 31) {real, imag} */,
  {32'h43332310, 32'hc38b3bc4} /* (22, 0, 30) {real, imag} */,
  {32'h3e3b6500, 32'hc1352c96} /* (22, 0, 29) {real, imag} */,
  {32'h42049fdf, 32'hc2890194} /* (22, 0, 28) {real, imag} */,
  {32'h429772d6, 32'h3ffd81d8} /* (22, 0, 27) {real, imag} */,
  {32'hc146c26a, 32'hc16d4910} /* (22, 0, 26) {real, imag} */,
  {32'h41b2a2ce, 32'hbf825010} /* (22, 0, 25) {real, imag} */,
  {32'h401d9b94, 32'hc208ff76} /* (22, 0, 24) {real, imag} */,
  {32'h4160a356, 32'hc0a04a88} /* (22, 0, 23) {real, imag} */,
  {32'h41173167, 32'h410021ce} /* (22, 0, 22) {real, imag} */,
  {32'h40c919b8, 32'hc183c30f} /* (22, 0, 21) {real, imag} */,
  {32'hc0e850fd, 32'h407ce99f} /* (22, 0, 20) {real, imag} */,
  {32'h3ffbcaf1, 32'hc0eeb7ee} /* (22, 0, 19) {real, imag} */,
  {32'hc15193f8, 32'hc027ad29} /* (22, 0, 18) {real, imag} */,
  {32'h4005fbec, 32'h41093e9a} /* (22, 0, 17) {real, imag} */,
  {32'h40329ff8, 32'h00000000} /* (22, 0, 16) {real, imag} */,
  {32'h4005fbec, 32'hc1093e9a} /* (22, 0, 15) {real, imag} */,
  {32'hc15193f8, 32'h4027ad29} /* (22, 0, 14) {real, imag} */,
  {32'h3ffbcaf1, 32'h40eeb7ee} /* (22, 0, 13) {real, imag} */,
  {32'hc0e850fd, 32'hc07ce99f} /* (22, 0, 12) {real, imag} */,
  {32'h40c919b8, 32'h4183c30f} /* (22, 0, 11) {real, imag} */,
  {32'h41173167, 32'hc10021ce} /* (22, 0, 10) {real, imag} */,
  {32'h4160a356, 32'h40a04a88} /* (22, 0, 9) {real, imag} */,
  {32'h401d9b94, 32'h4208ff76} /* (22, 0, 8) {real, imag} */,
  {32'h41b2a2ce, 32'h3f825010} /* (22, 0, 7) {real, imag} */,
  {32'hc146c26a, 32'h416d4910} /* (22, 0, 6) {real, imag} */,
  {32'h429772d6, 32'hbffd81d8} /* (22, 0, 5) {real, imag} */,
  {32'h42049fdf, 32'h42890194} /* (22, 0, 4) {real, imag} */,
  {32'h3e3b6500, 32'h41352c96} /* (22, 0, 3) {real, imag} */,
  {32'h43332310, 32'h438b3bc4} /* (22, 0, 2) {real, imag} */,
  {32'hc4c03ee8, 32'hc4995acc} /* (22, 0, 1) {real, imag} */,
  {32'hc51598fc, 32'h00000000} /* (22, 0, 0) {real, imag} */,
  {32'hc51ee7a3, 32'h44aa4da7} /* (21, 31, 31) {real, imag} */,
  {32'h440f4c17, 32'hc4104db4} /* (21, 31, 30) {real, imag} */,
  {32'h426163fa, 32'hc1a846d6} /* (21, 31, 29) {real, imag} */,
  {32'hc1c67fe8, 32'h429162c8} /* (21, 31, 28) {real, imag} */,
  {32'h42854e6c, 32'hc280f509} /* (21, 31, 27) {real, imag} */,
  {32'hc115ca7d, 32'h40d7d8f4} /* (21, 31, 26) {real, imag} */,
  {32'h4061fdc8, 32'h41ce4f79} /* (21, 31, 25) {real, imag} */,
  {32'h40d77b58, 32'hc234bb8a} /* (21, 31, 24) {real, imag} */,
  {32'h4218a2bd, 32'hc11d4159} /* (21, 31, 23) {real, imag} */,
  {32'hc1727c7c, 32'h4067abec} /* (21, 31, 22) {real, imag} */,
  {32'h40c3dd87, 32'hc1d59e6a} /* (21, 31, 21) {real, imag} */,
  {32'h404d9fd2, 32'hc1a121f0} /* (21, 31, 20) {real, imag} */,
  {32'hbf87e6e0, 32'h417b8434} /* (21, 31, 19) {real, imag} */,
  {32'hc110b2e6, 32'hc11142ca} /* (21, 31, 18) {real, imag} */,
  {32'hc087d492, 32'h40e822ca} /* (21, 31, 17) {real, imag} */,
  {32'hbf58c234, 32'h40cda5c6} /* (21, 31, 16) {real, imag} */,
  {32'h41863785, 32'hbf85abc0} /* (21, 31, 15) {real, imag} */,
  {32'h408bc460, 32'hc0a21341} /* (21, 31, 14) {real, imag} */,
  {32'hbfb4d968, 32'h412ac105} /* (21, 31, 13) {real, imag} */,
  {32'h413ec4fc, 32'hc03892db} /* (21, 31, 12) {real, imag} */,
  {32'h41f002f3, 32'hc0d28a8b} /* (21, 31, 11) {real, imag} */,
  {32'h41ffed07, 32'h4054a3f8} /* (21, 31, 10) {real, imag} */,
  {32'h41a87ea4, 32'h4176d706} /* (21, 31, 9) {real, imag} */,
  {32'h404a2924, 32'h41880721} /* (21, 31, 8) {real, imag} */,
  {32'h40bc3e07, 32'h41966f83} /* (21, 31, 7) {real, imag} */,
  {32'h41134a2f, 32'h41e0eaff} /* (21, 31, 6) {real, imag} */,
  {32'h43076ed6, 32'h416832f8} /* (21, 31, 5) {real, imag} */,
  {32'hc2dc6d9a, 32'h42c9a8ce} /* (21, 31, 4) {real, imag} */,
  {32'h407047d0, 32'h426920f2} /* (21, 31, 3) {real, imag} */,
  {32'h43f436ba, 32'hc1ab5ccb} /* (21, 31, 2) {real, imag} */,
  {32'hc4e15558, 32'hc3f3fda5} /* (21, 31, 1) {real, imag} */,
  {32'hc50a002c, 32'h43a856a6} /* (21, 31, 0) {real, imag} */,
  {32'h4443ca46, 32'h42d46b7e} /* (21, 30, 31) {real, imag} */,
  {32'hc3c92148, 32'hc2bbd477} /* (21, 30, 30) {real, imag} */,
  {32'h405090d0, 32'h41d58fc4} /* (21, 30, 29) {real, imag} */,
  {32'h42c42db8, 32'hc1a83ce5} /* (21, 30, 28) {real, imag} */,
  {32'hc2adfe11, 32'h4269ac94} /* (21, 30, 27) {real, imag} */,
  {32'h407b8667, 32'hc132b07d} /* (21, 30, 26) {real, imag} */,
  {32'h3fe8248e, 32'h41386ddf} /* (21, 30, 25) {real, imag} */,
  {32'hc1729192, 32'h41f64f98} /* (21, 30, 24) {real, imag} */,
  {32'h41683a34, 32'h40a6cceb} /* (21, 30, 23) {real, imag} */,
  {32'h41376366, 32'h407cbe30} /* (21, 30, 22) {real, imag} */,
  {32'h3f1ecd74, 32'h41919470} /* (21, 30, 21) {real, imag} */,
  {32'h4105be9e, 32'hc018c694} /* (21, 30, 20) {real, imag} */,
  {32'hc09167ec, 32'hc120187a} /* (21, 30, 19) {real, imag} */,
  {32'h40e2beec, 32'h41c15f93} /* (21, 30, 18) {real, imag} */,
  {32'hc053f85c, 32'hc0b4ccda} /* (21, 30, 17) {real, imag} */,
  {32'hc100017b, 32'hbfb73352} /* (21, 30, 16) {real, imag} */,
  {32'h3f8e6650, 32'h4141acdc} /* (21, 30, 15) {real, imag} */,
  {32'hc19d12a0, 32'hc0c620c8} /* (21, 30, 14) {real, imag} */,
  {32'hc017e177, 32'h40861f04} /* (21, 30, 13) {real, imag} */,
  {32'h4113a82e, 32'h40949d28} /* (21, 30, 12) {real, imag} */,
  {32'h3fbad3fc, 32'hc09abe48} /* (21, 30, 11) {real, imag} */,
  {32'hc160899b, 32'h3e80c098} /* (21, 30, 10) {real, imag} */,
  {32'hc16d993a, 32'hc0233836} /* (21, 30, 9) {real, imag} */,
  {32'hc1f90397, 32'hc23aeb5f} /* (21, 30, 8) {real, imag} */,
  {32'h41c0fc76, 32'h419a725e} /* (21, 30, 7) {real, imag} */,
  {32'hbfbdb5d8, 32'hc1674c88} /* (21, 30, 6) {real, imag} */,
  {32'hc2276feb, 32'hc1eac712} /* (21, 30, 5) {real, imag} */,
  {32'h40a32870, 32'h427e464c} /* (21, 30, 4) {real, imag} */,
  {32'hbf250508, 32'hc0ed6e25} /* (21, 30, 3) {real, imag} */,
  {32'hc4143477, 32'hc36680f3} /* (21, 30, 2) {real, imag} */,
  {32'h44a46bad, 32'hc1875c0a} /* (21, 30, 1) {real, imag} */,
  {32'h4424705c, 32'hc3073b9c} /* (21, 30, 0) {real, imag} */,
  {32'hc308adde, 32'h42b7548c} /* (21, 29, 31) {real, imag} */,
  {32'hc1052833, 32'hc2e586ac} /* (21, 29, 30) {real, imag} */,
  {32'h424ac748, 32'hc11a2c5a} /* (21, 29, 29) {real, imag} */,
  {32'h42312b07, 32'h42324670} /* (21, 29, 28) {real, imag} */,
  {32'hc10b83c6, 32'h40639be2} /* (21, 29, 27) {real, imag} */,
  {32'hbfa49684, 32'h401a418a} /* (21, 29, 26) {real, imag} */,
  {32'h419dc7dc, 32'h41352d3f} /* (21, 29, 25) {real, imag} */,
  {32'hc183c27e, 32'hc1592208} /* (21, 29, 24) {real, imag} */,
  {32'hc1da58ce, 32'hbfec76c4} /* (21, 29, 23) {real, imag} */,
  {32'h40d1a864, 32'hc13d6069} /* (21, 29, 22) {real, imag} */,
  {32'hc06e3a9a, 32'hc0bf8c20} /* (21, 29, 21) {real, imag} */,
  {32'hbfb73850, 32'hc12b0e13} /* (21, 29, 20) {real, imag} */,
  {32'h404fdacc, 32'h3f23a002} /* (21, 29, 19) {real, imag} */,
  {32'hbefc3aa0, 32'hc1473263} /* (21, 29, 18) {real, imag} */,
  {32'h411a784b, 32'hbf065550} /* (21, 29, 17) {real, imag} */,
  {32'h418005d1, 32'hc02f0124} /* (21, 29, 16) {real, imag} */,
  {32'h3f76f1b8, 32'hbfa8d270} /* (21, 29, 15) {real, imag} */,
  {32'hc0e1615e, 32'h41473e02} /* (21, 29, 14) {real, imag} */,
  {32'h417cfb7d, 32'h411d4fff} /* (21, 29, 13) {real, imag} */,
  {32'h418a5966, 32'hc195f017} /* (21, 29, 12) {real, imag} */,
  {32'h4131061a, 32'hc1a00dd0} /* (21, 29, 11) {real, imag} */,
  {32'hc0efc6db, 32'h41cb9a10} /* (21, 29, 10) {real, imag} */,
  {32'hbf952e9c, 32'h41ad83df} /* (21, 29, 9) {real, imag} */,
  {32'h41b6d850, 32'hc0dd6283} /* (21, 29, 8) {real, imag} */,
  {32'hc1d3e032, 32'h409bda4a} /* (21, 29, 7) {real, imag} */,
  {32'h410e44fc, 32'h41da7e81} /* (21, 29, 6) {real, imag} */,
  {32'h417fad59, 32'h40720d54} /* (21, 29, 5) {real, imag} */,
  {32'hc2447536, 32'h421809de} /* (21, 29, 4) {real, imag} */,
  {32'hc11a8dcb, 32'hc07924b9} /* (21, 29, 3) {real, imag} */,
  {32'hc2cf5563, 32'hc2c5f0e9} /* (21, 29, 2) {real, imag} */,
  {32'h4313f214, 32'h42a111e1} /* (21, 29, 1) {real, imag} */,
  {32'h4240fea0, 32'hc13207d2} /* (21, 29, 0) {real, imag} */,
  {32'hc30e25c0, 32'h426c4de8} /* (21, 28, 31) {real, imag} */,
  {32'h42f36fd0, 32'hc270705c} /* (21, 28, 30) {real, imag} */,
  {32'hc06aabe0, 32'h4218af4a} /* (21, 28, 29) {real, imag} */,
  {32'h41cf7a63, 32'h420587ad} /* (21, 28, 28) {real, imag} */,
  {32'h41bcfe58, 32'hc110531e} /* (21, 28, 27) {real, imag} */,
  {32'hbf8863c8, 32'hbf982d08} /* (21, 28, 26) {real, imag} */,
  {32'hc190d2e4, 32'hc09e8fe7} /* (21, 28, 25) {real, imag} */,
  {32'h41b19a4d, 32'hc13b8a99} /* (21, 28, 24) {real, imag} */,
  {32'h403a87e8, 32'hbfe14bb4} /* (21, 28, 23) {real, imag} */,
  {32'h409cdff2, 32'h408616f5} /* (21, 28, 22) {real, imag} */,
  {32'h4198bac7, 32'hc0879407} /* (21, 28, 21) {real, imag} */,
  {32'hc0e39be7, 32'hbfb75a0f} /* (21, 28, 20) {real, imag} */,
  {32'hc10e3c3a, 32'h41b15bb6} /* (21, 28, 19) {real, imag} */,
  {32'h3e2af9e0, 32'h4101ceea} /* (21, 28, 18) {real, imag} */,
  {32'h404a15a4, 32'h3e453428} /* (21, 28, 17) {real, imag} */,
  {32'hc0b700a2, 32'hbfddcf24} /* (21, 28, 16) {real, imag} */,
  {32'h3fb1349c, 32'hc0529ae4} /* (21, 28, 15) {real, imag} */,
  {32'h418a62ac, 32'hc1602be6} /* (21, 28, 14) {real, imag} */,
  {32'hc0c1e5b0, 32'hc19a8f9a} /* (21, 28, 13) {real, imag} */,
  {32'h418a8a6d, 32'hc18f7464} /* (21, 28, 12) {real, imag} */,
  {32'hc18c8005, 32'h41055968} /* (21, 28, 11) {real, imag} */,
  {32'hc1157701, 32'hc01548d7} /* (21, 28, 10) {real, imag} */,
  {32'hc1150669, 32'h40863eb5} /* (21, 28, 9) {real, imag} */,
  {32'h414f046c, 32'hc0f53f05} /* (21, 28, 8) {real, imag} */,
  {32'h4116f032, 32'hc19d6c32} /* (21, 28, 7) {real, imag} */,
  {32'h41204934, 32'h41a774f2} /* (21, 28, 6) {real, imag} */,
  {32'h405ffa2e, 32'h41c7ef34} /* (21, 28, 5) {real, imag} */,
  {32'hc1926db6, 32'hc1b739ac} /* (21, 28, 4) {real, imag} */,
  {32'h40b570c2, 32'hbe945e20} /* (21, 28, 3) {real, imag} */,
  {32'h42c1bff3, 32'hc26864da} /* (21, 28, 2) {real, imag} */,
  {32'hc1f6f992, 32'h42d9fc9f} /* (21, 28, 1) {real, imag} */,
  {32'hc283df29, 32'hc2280a95} /* (21, 28, 0) {real, imag} */,
  {32'h4281da38, 32'hc28106c8} /* (21, 27, 31) {real, imag} */,
  {32'hc17f4f69, 32'h423ca04f} /* (21, 27, 30) {real, imag} */,
  {32'h41123773, 32'hc114306c} /* (21, 27, 29) {real, imag} */,
  {32'hc163baf0, 32'hc194d418} /* (21, 27, 28) {real, imag} */,
  {32'hc1939dd8, 32'h4181563d} /* (21, 27, 27) {real, imag} */,
  {32'h40f9787c, 32'h41236fe8} /* (21, 27, 26) {real, imag} */,
  {32'h42074d8c, 32'hc14d9639} /* (21, 27, 25) {real, imag} */,
  {32'hc0cda84b, 32'h40412ed0} /* (21, 27, 24) {real, imag} */,
  {32'h40fe9a15, 32'h417a41a2} /* (21, 27, 23) {real, imag} */,
  {32'h41067b40, 32'hc0c7d274} /* (21, 27, 22) {real, imag} */,
  {32'hc10f9e70, 32'h4192d404} /* (21, 27, 21) {real, imag} */,
  {32'hc0aa43d0, 32'h41040ba6} /* (21, 27, 20) {real, imag} */,
  {32'h40a62d48, 32'h3f2a5670} /* (21, 27, 19) {real, imag} */,
  {32'hc1133b91, 32'h40213344} /* (21, 27, 18) {real, imag} */,
  {32'hc0cee78c, 32'hbdb69a00} /* (21, 27, 17) {real, imag} */,
  {32'hc0ac0092, 32'hc04b97be} /* (21, 27, 16) {real, imag} */,
  {32'h40ab4179, 32'h411c60db} /* (21, 27, 15) {real, imag} */,
  {32'hbfc49b52, 32'hc060551e} /* (21, 27, 14) {real, imag} */,
  {32'hc00e23e8, 32'hbfedb4dc} /* (21, 27, 13) {real, imag} */,
  {32'h4125506a, 32'hc102bb36} /* (21, 27, 12) {real, imag} */,
  {32'hbed0e568, 32'h40d7b5ce} /* (21, 27, 11) {real, imag} */,
  {32'hc0bd7857, 32'h3d404700} /* (21, 27, 10) {real, imag} */,
  {32'h3ff5a488, 32'hc0d32f05} /* (21, 27, 9) {real, imag} */,
  {32'hc0aa8644, 32'hc0a47504} /* (21, 27, 8) {real, imag} */,
  {32'h410d6142, 32'hbfa8dfde} /* (21, 27, 7) {real, imag} */,
  {32'hc1d9b72e, 32'hc037449e} /* (21, 27, 6) {real, imag} */,
  {32'hc1f38dee, 32'h4047c98c} /* (21, 27, 5) {real, imag} */,
  {32'h4195423c, 32'h40e2c888} /* (21, 27, 4) {real, imag} */,
  {32'h3fe74b80, 32'hc14f53e4} /* (21, 27, 3) {real, imag} */,
  {32'hc203cf70, 32'h4153c5f0} /* (21, 27, 2) {real, imag} */,
  {32'h42bd67e2, 32'hc1618323} /* (21, 27, 1) {real, imag} */,
  {32'h42162774, 32'hc295cd98} /* (21, 27, 0) {real, imag} */,
  {32'hc050f7c8, 32'hc12c6f77} /* (21, 26, 31) {real, imag} */,
  {32'h408e3884, 32'hc1b83a26} /* (21, 26, 30) {real, imag} */,
  {32'h419b20b3, 32'h41a50a81} /* (21, 26, 29) {real, imag} */,
  {32'hc08c1600, 32'hc01647d1} /* (21, 26, 28) {real, imag} */,
  {32'hc1b87360, 32'hc0bee95d} /* (21, 26, 27) {real, imag} */,
  {32'hc150a914, 32'h4190b2ee} /* (21, 26, 26) {real, imag} */,
  {32'hc0f65d1e, 32'h4015ea8a} /* (21, 26, 25) {real, imag} */,
  {32'hc0852d8a, 32'h41af788c} /* (21, 26, 24) {real, imag} */,
  {32'h3f464030, 32'hc162f9c7} /* (21, 26, 23) {real, imag} */,
  {32'h3e56bf00, 32'hc198492c} /* (21, 26, 22) {real, imag} */,
  {32'hc191e8c2, 32'h418066cb} /* (21, 26, 21) {real, imag} */,
  {32'hc11b616e, 32'hc085f412} /* (21, 26, 20) {real, imag} */,
  {32'hbfad5b67, 32'h4173bb01} /* (21, 26, 19) {real, imag} */,
  {32'h40c125ea, 32'hc098adb0} /* (21, 26, 18) {real, imag} */,
  {32'h3d740f60, 32'hbff96d5e} /* (21, 26, 17) {real, imag} */,
  {32'hc0c23fd4, 32'h40d62aad} /* (21, 26, 16) {real, imag} */,
  {32'h418630e9, 32'hc0ee77d2} /* (21, 26, 15) {real, imag} */,
  {32'hc083c696, 32'hc17db580} /* (21, 26, 14) {real, imag} */,
  {32'hc10adb2e, 32'h412a702b} /* (21, 26, 13) {real, imag} */,
  {32'hc16c2d95, 32'h3eb54f10} /* (21, 26, 12) {real, imag} */,
  {32'hc0e038eb, 32'h3fe60c80} /* (21, 26, 11) {real, imag} */,
  {32'h401c7640, 32'h41369056} /* (21, 26, 10) {real, imag} */,
  {32'hc10dd212, 32'hc177ff78} /* (21, 26, 9) {real, imag} */,
  {32'hc10009c6, 32'hc0e6a97b} /* (21, 26, 8) {real, imag} */,
  {32'hc09f4018, 32'h4121a559} /* (21, 26, 7) {real, imag} */,
  {32'h414a7d0e, 32'h4182638a} /* (21, 26, 6) {real, imag} */,
  {32'hc0fe644c, 32'h41baaf9d} /* (21, 26, 5) {real, imag} */,
  {32'h41ade48c, 32'h41a0a7f5} /* (21, 26, 4) {real, imag} */,
  {32'h40fe0aa5, 32'hc084667a} /* (21, 26, 3) {real, imag} */,
  {32'h3f85c200, 32'h40870388} /* (21, 26, 2) {real, imag} */,
  {32'hc10be10a, 32'hc2029357} /* (21, 26, 1) {real, imag} */,
  {32'hc0d33a47, 32'hc095f1e1} /* (21, 26, 0) {real, imag} */,
  {32'h40d05b28, 32'h40605b6f} /* (21, 25, 31) {real, imag} */,
  {32'h411c4d14, 32'hc0def07c} /* (21, 25, 30) {real, imag} */,
  {32'h41d6105b, 32'hc1626cce} /* (21, 25, 29) {real, imag} */,
  {32'h3ece6d40, 32'h4135830d} /* (21, 25, 28) {real, imag} */,
  {32'h41d5ed6c, 32'h4105035a} /* (21, 25, 27) {real, imag} */,
  {32'hc0e30ddf, 32'hc195c674} /* (21, 25, 26) {real, imag} */,
  {32'hc1b968ae, 32'h3f755d90} /* (21, 25, 25) {real, imag} */,
  {32'hc0f139bd, 32'hbebeeef8} /* (21, 25, 24) {real, imag} */,
  {32'hc094d9b7, 32'hc047f028} /* (21, 25, 23) {real, imag} */,
  {32'hc0cd5d66, 32'h40d10976} /* (21, 25, 22) {real, imag} */,
  {32'hc1af4b36, 32'hc162ea48} /* (21, 25, 21) {real, imag} */,
  {32'hc0843ab3, 32'h40cbe7ea} /* (21, 25, 20) {real, imag} */,
  {32'hc012808e, 32'hc0cae15b} /* (21, 25, 19) {real, imag} */,
  {32'hc16d2434, 32'hc040cdb8} /* (21, 25, 18) {real, imag} */,
  {32'h3e89fca4, 32'hc03591fe} /* (21, 25, 17) {real, imag} */,
  {32'hc0639f69, 32'h4150b56d} /* (21, 25, 16) {real, imag} */,
  {32'hc11b595c, 32'hc093efb4} /* (21, 25, 15) {real, imag} */,
  {32'h3ff04e38, 32'h40b30e13} /* (21, 25, 14) {real, imag} */,
  {32'h403b437c, 32'hc13cbfeb} /* (21, 25, 13) {real, imag} */,
  {32'hc0977cb0, 32'h3ebdbeac} /* (21, 25, 12) {real, imag} */,
  {32'h3f443f28, 32'h419437f4} /* (21, 25, 11) {real, imag} */,
  {32'hc19df8cb, 32'hc0aa2584} /* (21, 25, 10) {real, imag} */,
  {32'hc0974642, 32'h40c1b15f} /* (21, 25, 9) {real, imag} */,
  {32'hc09a5dd2, 32'hc1812ca6} /* (21, 25, 8) {real, imag} */,
  {32'hc12e164c, 32'hc160b147} /* (21, 25, 7) {real, imag} */,
  {32'hc11b75ba, 32'hc1b209f8} /* (21, 25, 6) {real, imag} */,
  {32'hc1375d73, 32'hc0a01ec5} /* (21, 25, 5) {real, imag} */,
  {32'h419e85c6, 32'hc080a594} /* (21, 25, 4) {real, imag} */,
  {32'h4059f536, 32'h40888e9b} /* (21, 25, 3) {real, imag} */,
  {32'h418d938f, 32'h41c7321b} /* (21, 25, 2) {real, imag} */,
  {32'h3ed23780, 32'h4167c94c} /* (21, 25, 1) {real, imag} */,
  {32'hc1c6c9e7, 32'h41ec1c8e} /* (21, 25, 0) {real, imag} */,
  {32'h41986e44, 32'hc149bbf2} /* (21, 24, 31) {real, imag} */,
  {32'hc19bbb3f, 32'h40e784d0} /* (21, 24, 30) {real, imag} */,
  {32'h41720080, 32'h40e0fefd} /* (21, 24, 29) {real, imag} */,
  {32'h418738b9, 32'h407bc962} /* (21, 24, 28) {real, imag} */,
  {32'hc2087754, 32'h406ac1d4} /* (21, 24, 27) {real, imag} */,
  {32'h4035b7cc, 32'hbf2bac00} /* (21, 24, 26) {real, imag} */,
  {32'hc01552f4, 32'h40caac96} /* (21, 24, 25) {real, imag} */,
  {32'hbf4a14e0, 32'hc00cafc2} /* (21, 24, 24) {real, imag} */,
  {32'hbff1f840, 32'h400c10d8} /* (21, 24, 23) {real, imag} */,
  {32'hc18db8f6, 32'hc1c2438e} /* (21, 24, 22) {real, imag} */,
  {32'hbe299a40, 32'h41c9d051} /* (21, 24, 21) {real, imag} */,
  {32'h40c4c29a, 32'h4134c39a} /* (21, 24, 20) {real, imag} */,
  {32'h3f10f380, 32'h40f81da0} /* (21, 24, 19) {real, imag} */,
  {32'hc0ebb5b3, 32'hc0051572} /* (21, 24, 18) {real, imag} */,
  {32'hc0dd22dc, 32'hc0ac4711} /* (21, 24, 17) {real, imag} */,
  {32'h3f87269c, 32'h408a9782} /* (21, 24, 16) {real, imag} */,
  {32'h4004d4cc, 32'hbf177110} /* (21, 24, 15) {real, imag} */,
  {32'hc050c5dc, 32'hc12a805a} /* (21, 24, 14) {real, imag} */,
  {32'h4062e398, 32'h41541651} /* (21, 24, 13) {real, imag} */,
  {32'h40a3eb8b, 32'hbfbfc9b4} /* (21, 24, 12) {real, imag} */,
  {32'hc0709a8e, 32'hc1c95788} /* (21, 24, 11) {real, imag} */,
  {32'hbe078d80, 32'h403ab0d8} /* (21, 24, 10) {real, imag} */,
  {32'h411c3a13, 32'hc11e78b7} /* (21, 24, 9) {real, imag} */,
  {32'hc0998693, 32'h41828a0c} /* (21, 24, 8) {real, imag} */,
  {32'h40f742b3, 32'h407803d0} /* (21, 24, 7) {real, imag} */,
  {32'h41f3339a, 32'h3e641a00} /* (21, 24, 6) {real, imag} */,
  {32'hc1d4a9fe, 32'h4191bb49} /* (21, 24, 5) {real, imag} */,
  {32'h4075ec40, 32'hc113132b} /* (21, 24, 4) {real, imag} */,
  {32'h410451b2, 32'hbf7c6b18} /* (21, 24, 3) {real, imag} */,
  {32'hc1bb04cd, 32'h4151d501} /* (21, 24, 2) {real, imag} */,
  {32'h42156bc1, 32'hc2052325} /* (21, 24, 1) {real, imag} */,
  {32'h411e3e58, 32'h40c24b1c} /* (21, 24, 0) {real, imag} */,
  {32'hc1ac64f8, 32'h403de9dc} /* (21, 23, 31) {real, imag} */,
  {32'hbf882fbc, 32'hc132c967} /* (21, 23, 30) {real, imag} */,
  {32'h41528adf, 32'h4131aa87} /* (21, 23, 29) {real, imag} */,
  {32'hc1736f04, 32'hc01dd7ef} /* (21, 23, 28) {real, imag} */,
  {32'h41bdea61, 32'hc0a89747} /* (21, 23, 27) {real, imag} */,
  {32'hc1496e07, 32'h41d16a40} /* (21, 23, 26) {real, imag} */,
  {32'h40c15b7c, 32'h41a23ddc} /* (21, 23, 25) {real, imag} */,
  {32'hc17b1608, 32'hc0cae552} /* (21, 23, 24) {real, imag} */,
  {32'h41b4f97a, 32'h40d51398} /* (21, 23, 23) {real, imag} */,
  {32'h411e3e20, 32'h40d701c7} /* (21, 23, 22) {real, imag} */,
  {32'h3ea11430, 32'hc163c516} /* (21, 23, 21) {real, imag} */,
  {32'hc1a5acbf, 32'hc0541d60} /* (21, 23, 20) {real, imag} */,
  {32'hc0ac8392, 32'hc0e0bb37} /* (21, 23, 19) {real, imag} */,
  {32'h3e9be448, 32'hc13ab478} /* (21, 23, 18) {real, imag} */,
  {32'h4087eb8a, 32'h40402015} /* (21, 23, 17) {real, imag} */,
  {32'hbdf5cd40, 32'hc091f94f} /* (21, 23, 16) {real, imag} */,
  {32'hc08b4b3c, 32'h419cc79e} /* (21, 23, 15) {real, imag} */,
  {32'h4125d6c7, 32'hc068cd36} /* (21, 23, 14) {real, imag} */,
  {32'hc00c7c80, 32'h40245668} /* (21, 23, 13) {real, imag} */,
  {32'h400e5c44, 32'hc09bce5e} /* (21, 23, 12) {real, imag} */,
  {32'hc10307d3, 32'hc03a3544} /* (21, 23, 11) {real, imag} */,
  {32'hc0b3ce7f, 32'h4187346a} /* (21, 23, 10) {real, imag} */,
  {32'hbf1f4ce4, 32'h3e0e1080} /* (21, 23, 9) {real, imag} */,
  {32'hc08f7c11, 32'hc1852dbd} /* (21, 23, 8) {real, imag} */,
  {32'hc0cae2a4, 32'hc09009c5} /* (21, 23, 7) {real, imag} */,
  {32'hc0784c4c, 32'hbfb77e14} /* (21, 23, 6) {real, imag} */,
  {32'h404e0378, 32'h40d6bc65} /* (21, 23, 5) {real, imag} */,
  {32'hbfd625e8, 32'h419cf116} /* (21, 23, 4) {real, imag} */,
  {32'hc126acbc, 32'h41748036} /* (21, 23, 3) {real, imag} */,
  {32'hc076b3be, 32'hc11d2e84} /* (21, 23, 2) {real, imag} */,
  {32'h4171b561, 32'hc17e8fca} /* (21, 23, 1) {real, imag} */,
  {32'h4186b3e3, 32'hc1228e66} /* (21, 23, 0) {real, imag} */,
  {32'hc1f0e694, 32'h41693db2} /* (21, 22, 31) {real, imag} */,
  {32'h40d91e1a, 32'h3fb69548} /* (21, 22, 30) {real, imag} */,
  {32'h3ffb40cc, 32'h3f16cf28} /* (21, 22, 29) {real, imag} */,
  {32'h40541328, 32'hc145d2b8} /* (21, 22, 28) {real, imag} */,
  {32'hc173fd64, 32'h41680ed3} /* (21, 22, 27) {real, imag} */,
  {32'h415c72fa, 32'h41836d7c} /* (21, 22, 26) {real, imag} */,
  {32'hc0ffe706, 32'hc06e3219} /* (21, 22, 25) {real, imag} */,
  {32'hc0f42492, 32'h410457b8} /* (21, 22, 24) {real, imag} */,
  {32'hbfb3ded0, 32'h3fbab364} /* (21, 22, 23) {real, imag} */,
  {32'h4152a866, 32'hc16fb632} /* (21, 22, 22) {real, imag} */,
  {32'hc061d9e0, 32'hc00c6cec} /* (21, 22, 21) {real, imag} */,
  {32'hc038167c, 32'hc18d67e8} /* (21, 22, 20) {real, imag} */,
  {32'hc0685b45, 32'h3fc28370} /* (21, 22, 19) {real, imag} */,
  {32'hbfe102ce, 32'h40c69c80} /* (21, 22, 18) {real, imag} */,
  {32'h40c8acb2, 32'h3ecbd1d0} /* (21, 22, 17) {real, imag} */,
  {32'h41890f35, 32'h40d3e9ba} /* (21, 22, 16) {real, imag} */,
  {32'hc111b11a, 32'hc14b3cc0} /* (21, 22, 15) {real, imag} */,
  {32'h3cf81c40, 32'h40f1a102} /* (21, 22, 14) {real, imag} */,
  {32'hc0dcbcd7, 32'h4084ae55} /* (21, 22, 13) {real, imag} */,
  {32'hbf14d074, 32'h416fb11a} /* (21, 22, 12) {real, imag} */,
  {32'h41a24b53, 32'h40fabfb4} /* (21, 22, 11) {real, imag} */,
  {32'h3e5d9fb0, 32'h410d12f5} /* (21, 22, 10) {real, imag} */,
  {32'hc1539aa6, 32'h40c63d94} /* (21, 22, 9) {real, imag} */,
  {32'h412fb52a, 32'hc0a6163e} /* (21, 22, 8) {real, imag} */,
  {32'hc18b2b00, 32'h406ad684} /* (21, 22, 7) {real, imag} */,
  {32'h41203376, 32'hc13e7db1} /* (21, 22, 6) {real, imag} */,
  {32'h41106aeb, 32'hc0a4f73b} /* (21, 22, 5) {real, imag} */,
  {32'hc1229643, 32'hc05db6ef} /* (21, 22, 4) {real, imag} */,
  {32'h403c7839, 32'h3fade910} /* (21, 22, 3) {real, imag} */,
  {32'h4151c0ef, 32'hc1a89d7b} /* (21, 22, 2) {real, imag} */,
  {32'h413d8b1c, 32'h41f60b3e} /* (21, 22, 1) {real, imag} */,
  {32'hc1dad4c8, 32'h40cac227} /* (21, 22, 0) {real, imag} */,
  {32'h3ffa5853, 32'hc199bf30} /* (21, 21, 31) {real, imag} */,
  {32'h40f8aa08, 32'h41254854} /* (21, 21, 30) {real, imag} */,
  {32'h41331ef5, 32'h41838600} /* (21, 21, 29) {real, imag} */,
  {32'hc115f8b0, 32'hc08c445e} /* (21, 21, 28) {real, imag} */,
  {32'h41535014, 32'h3fd4a4b0} /* (21, 21, 27) {real, imag} */,
  {32'h4145a0c2, 32'hc0e652a7} /* (21, 21, 26) {real, imag} */,
  {32'h4111a605, 32'h3fcbac38} /* (21, 21, 25) {real, imag} */,
  {32'h416dbfbf, 32'h3ddc8180} /* (21, 21, 24) {real, imag} */,
  {32'h414baa62, 32'h411a7108} /* (21, 21, 23) {real, imag} */,
  {32'h408a3b45, 32'h3fd722d8} /* (21, 21, 22) {real, imag} */,
  {32'hc1864264, 32'h3f299afc} /* (21, 21, 21) {real, imag} */,
  {32'hc144da70, 32'hc12bc2bd} /* (21, 21, 20) {real, imag} */,
  {32'hc0197313, 32'hc06049f6} /* (21, 21, 19) {real, imag} */,
  {32'h3df89b40, 32'hc096a9c6} /* (21, 21, 18) {real, imag} */,
  {32'h40083876, 32'h4104a76e} /* (21, 21, 17) {real, imag} */,
  {32'hc15caec6, 32'hc11c11e5} /* (21, 21, 16) {real, imag} */,
  {32'hc083a6ec, 32'h40af1030} /* (21, 21, 15) {real, imag} */,
  {32'h41684bbe, 32'h41913ff1} /* (21, 21, 14) {real, imag} */,
  {32'h4134ea39, 32'hc0ef7f97} /* (21, 21, 13) {real, imag} */,
  {32'h40b21faa, 32'hbece1ec0} /* (21, 21, 12) {real, imag} */,
  {32'hc0fccd98, 32'hc11b2a41} /* (21, 21, 11) {real, imag} */,
  {32'h41579ee8, 32'h40f8d3b0} /* (21, 21, 10) {real, imag} */,
  {32'h3f879a6c, 32'h3fc24928} /* (21, 21, 9) {real, imag} */,
  {32'h4125f604, 32'h4066f3b2} /* (21, 21, 8) {real, imag} */,
  {32'hc0fa8bf8, 32'hc0600e0c} /* (21, 21, 7) {real, imag} */,
  {32'hc17904e3, 32'h40cd8ff0} /* (21, 21, 6) {real, imag} */,
  {32'hc02072f2, 32'hc130e5fe} /* (21, 21, 5) {real, imag} */,
  {32'hc1a73d46, 32'hc08f4f5f} /* (21, 21, 4) {real, imag} */,
  {32'h4011d856, 32'hc080797b} /* (21, 21, 3) {real, imag} */,
  {32'hc1cade5b, 32'hc01c217d} /* (21, 21, 2) {real, imag} */,
  {32'h41201852, 32'hc069af7e} /* (21, 21, 1) {real, imag} */,
  {32'h413ecdfb, 32'hc1a917ed} /* (21, 21, 0) {real, imag} */,
  {32'h4050d53d, 32'h40a28556} /* (21, 20, 31) {real, imag} */,
  {32'h405416f6, 32'h40c470b4} /* (21, 20, 30) {real, imag} */,
  {32'hc0d5dadd, 32'hc0a2dad7} /* (21, 20, 29) {real, imag} */,
  {32'h41088516, 32'h4044c705} /* (21, 20, 28) {real, imag} */,
  {32'h4103ad56, 32'h401a7554} /* (21, 20, 27) {real, imag} */,
  {32'h410e0ffa, 32'hc03b274c} /* (21, 20, 26) {real, imag} */,
  {32'hc1a023c8, 32'hc0372dbc} /* (21, 20, 25) {real, imag} */,
  {32'hc143acc6, 32'hc13351a6} /* (21, 20, 24) {real, imag} */,
  {32'h40da209b, 32'h40efd856} /* (21, 20, 23) {real, imag} */,
  {32'hc02fe40e, 32'hc0eb3ab6} /* (21, 20, 22) {real, imag} */,
  {32'hc18bdb46, 32'hc01bb139} /* (21, 20, 21) {real, imag} */,
  {32'h41754a2c, 32'hc170b9b0} /* (21, 20, 20) {real, imag} */,
  {32'h40dbc5a7, 32'hc03b9e45} /* (21, 20, 19) {real, imag} */,
  {32'h40b9a501, 32'hbf9eb0f8} /* (21, 20, 18) {real, imag} */,
  {32'h40da2d46, 32'h413b5ea0} /* (21, 20, 17) {real, imag} */,
  {32'hc0d1ea52, 32'hc0cf51a4} /* (21, 20, 16) {real, imag} */,
  {32'h41622385, 32'hc12e5653} /* (21, 20, 15) {real, imag} */,
  {32'h4101ce7e, 32'h41628062} /* (21, 20, 14) {real, imag} */,
  {32'h401a5cd7, 32'h400409fe} /* (21, 20, 13) {real, imag} */,
  {32'h40d54c5c, 32'h4192df42} /* (21, 20, 12) {real, imag} */,
  {32'h41efbce0, 32'hc0a2bd34} /* (21, 20, 11) {real, imag} */,
  {32'h404d7a84, 32'hbecc0a0c} /* (21, 20, 10) {real, imag} */,
  {32'h4176d3e8, 32'h4037c210} /* (21, 20, 9) {real, imag} */,
  {32'h40281c7c, 32'hc12dca3f} /* (21, 20, 8) {real, imag} */,
  {32'h411e026b, 32'h3e4cf3e0} /* (21, 20, 7) {real, imag} */,
  {32'hc1b8cb9c, 32'hc0bc2390} /* (21, 20, 6) {real, imag} */,
  {32'h3f819ee2, 32'h4141e1db} /* (21, 20, 5) {real, imag} */,
  {32'hc0a73185, 32'hc0d0b578} /* (21, 20, 4) {real, imag} */,
  {32'h3f3f81d4, 32'h412a7a2a} /* (21, 20, 3) {real, imag} */,
  {32'hc16ef9f8, 32'h4078f5c0} /* (21, 20, 2) {real, imag} */,
  {32'hc08aa9d4, 32'hbf7815f8} /* (21, 20, 1) {real, imag} */,
  {32'h41c9bc09, 32'hc129d1c4} /* (21, 20, 0) {real, imag} */,
  {32'hc1b92bb0, 32'h41164d96} /* (21, 19, 31) {real, imag} */,
  {32'hc14e4ac1, 32'h3e4ef6c0} /* (21, 19, 30) {real, imag} */,
  {32'hc1132e18, 32'h3fd078b6} /* (21, 19, 29) {real, imag} */,
  {32'h413de89d, 32'h410b7ac3} /* (21, 19, 28) {real, imag} */,
  {32'h4123eeb4, 32'h4190c37e} /* (21, 19, 27) {real, imag} */,
  {32'hc132b89e, 32'hc1bfb61a} /* (21, 19, 26) {real, imag} */,
  {32'hbc7e5c00, 32'h40bf9283} /* (21, 19, 25) {real, imag} */,
  {32'h418fc9c8, 32'hc144021e} /* (21, 19, 24) {real, imag} */,
  {32'hc04f3b62, 32'h4041f490} /* (21, 19, 23) {real, imag} */,
  {32'hc158e6e0, 32'hc0d54c50} /* (21, 19, 22) {real, imag} */,
  {32'h4121ccf5, 32'h41a6c184} /* (21, 19, 21) {real, imag} */,
  {32'hc10cef3e, 32'hc1456134} /* (21, 19, 20) {real, imag} */,
  {32'h4130e958, 32'h3fdfa6d0} /* (21, 19, 19) {real, imag} */,
  {32'h419cff7f, 32'hc0c2c5f0} /* (21, 19, 18) {real, imag} */,
  {32'h3f2a46b6, 32'h3fdbb3c0} /* (21, 19, 17) {real, imag} */,
  {32'hc13792a9, 32'h403834fc} /* (21, 19, 16) {real, imag} */,
  {32'hc0a24e52, 32'h40dcc876} /* (21, 19, 15) {real, imag} */,
  {32'h410453f5, 32'hc107564b} /* (21, 19, 14) {real, imag} */,
  {32'hc12b57ff, 32'hc0e5f7ca} /* (21, 19, 13) {real, imag} */,
  {32'h40777974, 32'hc0311f74} /* (21, 19, 12) {real, imag} */,
  {32'h3fed0438, 32'hc0a9e829} /* (21, 19, 11) {real, imag} */,
  {32'h41343332, 32'hbf2834a8} /* (21, 19, 10) {real, imag} */,
  {32'h40c62d96, 32'h40a4c1a2} /* (21, 19, 9) {real, imag} */,
  {32'h40e00d04, 32'h417de83a} /* (21, 19, 8) {real, imag} */,
  {32'hc0a72ef9, 32'hc17cd96e} /* (21, 19, 7) {real, imag} */,
  {32'hc1a99d4e, 32'h409f4bd1} /* (21, 19, 6) {real, imag} */,
  {32'hc0568c1b, 32'h408c65f3} /* (21, 19, 5) {real, imag} */,
  {32'hc0925ba1, 32'h40c47b43} /* (21, 19, 4) {real, imag} */,
  {32'h41205238, 32'hc18398e4} /* (21, 19, 3) {real, imag} */,
  {32'hc19653eb, 32'h404ccd78} /* (21, 19, 2) {real, imag} */,
  {32'h410e1954, 32'hc057b80c} /* (21, 19, 1) {real, imag} */,
  {32'hc105b42f, 32'h3ffff12c} /* (21, 19, 0) {real, imag} */,
  {32'hc0e3447a, 32'hbe18d2c0} /* (21, 18, 31) {real, imag} */,
  {32'hc0b8d353, 32'hc00094ff} /* (21, 18, 30) {real, imag} */,
  {32'h4060e670, 32'h3fb59948} /* (21, 18, 29) {real, imag} */,
  {32'h40381b2c, 32'hc02d413c} /* (21, 18, 28) {real, imag} */,
  {32'hc0ea76c5, 32'h40d7e048} /* (21, 18, 27) {real, imag} */,
  {32'hc0fb3f8d, 32'h3ec1cd4c} /* (21, 18, 26) {real, imag} */,
  {32'hc16c80f0, 32'hc0d6b64c} /* (21, 18, 25) {real, imag} */,
  {32'h413dd722, 32'h3e30f320} /* (21, 18, 24) {real, imag} */,
  {32'hc10debd2, 32'hc18ec8ed} /* (21, 18, 23) {real, imag} */,
  {32'h404ed554, 32'hc151d598} /* (21, 18, 22) {real, imag} */,
  {32'h411e0c5a, 32'hc05c9eb8} /* (21, 18, 21) {real, imag} */,
  {32'h41b0c67d, 32'h415087e4} /* (21, 18, 20) {real, imag} */,
  {32'h403f3104, 32'hc0d41ce2} /* (21, 18, 19) {real, imag} */,
  {32'hc0491cd0, 32'h40e6abbb} /* (21, 18, 18) {real, imag} */,
  {32'h4071874a, 32'h417703d2} /* (21, 18, 17) {real, imag} */,
  {32'hbf8dd91c, 32'h409b7f06} /* (21, 18, 16) {real, imag} */,
  {32'hc183cd7d, 32'h3f9548a8} /* (21, 18, 15) {real, imag} */,
  {32'h4106f027, 32'hc0575cda} /* (21, 18, 14) {real, imag} */,
  {32'hc031b4a2, 32'hc14fdd0b} /* (21, 18, 13) {real, imag} */,
  {32'hc12e6808, 32'h407dc60b} /* (21, 18, 12) {real, imag} */,
  {32'hc15b3e08, 32'hc0dd6808} /* (21, 18, 11) {real, imag} */,
  {32'hc167251c, 32'hc010e9d8} /* (21, 18, 10) {real, imag} */,
  {32'hc017d881, 32'h40c96d20} /* (21, 18, 9) {real, imag} */,
  {32'hc15f24ac, 32'h40fcdbc3} /* (21, 18, 8) {real, imag} */,
  {32'h3ea46134, 32'hc160f968} /* (21, 18, 7) {real, imag} */,
  {32'hbf7b7c78, 32'hc15517f9} /* (21, 18, 6) {real, imag} */,
  {32'hc036d4b6, 32'h40114870} /* (21, 18, 5) {real, imag} */,
  {32'h41426593, 32'h3f71c950} /* (21, 18, 4) {real, imag} */,
  {32'h411e0726, 32'h4091b13e} /* (21, 18, 3) {real, imag} */,
  {32'hc10add00, 32'h40149a74} /* (21, 18, 2) {real, imag} */,
  {32'h40f2a63a, 32'hc1879689} /* (21, 18, 1) {real, imag} */,
  {32'hc0e848e2, 32'hc1797276} /* (21, 18, 0) {real, imag} */,
  {32'h40a66ace, 32'hc0ee319a} /* (21, 17, 31) {real, imag} */,
  {32'h41029f17, 32'hc10edd29} /* (21, 17, 30) {real, imag} */,
  {32'h3f6eedf8, 32'h409cd37a} /* (21, 17, 29) {real, imag} */,
  {32'hc152df54, 32'hc0aa5e72} /* (21, 17, 28) {real, imag} */,
  {32'hc13ef61c, 32'h40c52c81} /* (21, 17, 27) {real, imag} */,
  {32'hbf10627c, 32'h3fc12628} /* (21, 17, 26) {real, imag} */,
  {32'hbf92ed96, 32'h3f854af0} /* (21, 17, 25) {real, imag} */,
  {32'hc109b7d9, 32'h4073c8f9} /* (21, 17, 24) {real, imag} */,
  {32'hc0b0f7ce, 32'hc09caaa6} /* (21, 17, 23) {real, imag} */,
  {32'h4180b474, 32'h4098440f} /* (21, 17, 22) {real, imag} */,
  {32'h409745dd, 32'hc17db58e} /* (21, 17, 21) {real, imag} */,
  {32'h41031d19, 32'h408bd5c3} /* (21, 17, 20) {real, imag} */,
  {32'hc00a344a, 32'h40bb83fa} /* (21, 17, 19) {real, imag} */,
  {32'hc06fac64, 32'h40e65399} /* (21, 17, 18) {real, imag} */,
  {32'h40180bc4, 32'hc14b03f1} /* (21, 17, 17) {real, imag} */,
  {32'hc10fdc35, 32'h411bf7d1} /* (21, 17, 16) {real, imag} */,
  {32'h40f9a65b, 32'hc168c672} /* (21, 17, 15) {real, imag} */,
  {32'h3febcdf8, 32'hc07f792c} /* (21, 17, 14) {real, imag} */,
  {32'hbfaca420, 32'h40bd52ca} /* (21, 17, 13) {real, imag} */,
  {32'h40167124, 32'h40234208} /* (21, 17, 12) {real, imag} */,
  {32'hc18968f4, 32'hc1485712} /* (21, 17, 11) {real, imag} */,
  {32'hc153e3bc, 32'h40e794e5} /* (21, 17, 10) {real, imag} */,
  {32'h410e07b5, 32'h3ebf8bb0} /* (21, 17, 9) {real, imag} */,
  {32'hc11c109c, 32'h40825cec} /* (21, 17, 8) {real, imag} */,
  {32'hbf9c5f84, 32'h40ae5b57} /* (21, 17, 7) {real, imag} */,
  {32'hc0a8ffbd, 32'hc04037ad} /* (21, 17, 6) {real, imag} */,
  {32'hc0789d30, 32'h40b23947} /* (21, 17, 5) {real, imag} */,
  {32'h40796fe4, 32'hbd7c8a40} /* (21, 17, 4) {real, imag} */,
  {32'h4094546c, 32'hc0621393} /* (21, 17, 3) {real, imag} */,
  {32'hc05d4069, 32'h4052980f} /* (21, 17, 2) {real, imag} */,
  {32'h4114ec56, 32'h403f8abc} /* (21, 17, 1) {real, imag} */,
  {32'h40de4622, 32'h40e8eed8} /* (21, 17, 0) {real, imag} */,
  {32'h405cb700, 32'h3fa53ea5} /* (21, 16, 31) {real, imag} */,
  {32'h40426d33, 32'hc0cfed72} /* (21, 16, 30) {real, imag} */,
  {32'hbfb037fd, 32'hc0b099b7} /* (21, 16, 29) {real, imag} */,
  {32'hc154b3ee, 32'hc0883c57} /* (21, 16, 28) {real, imag} */,
  {32'hbf49ad3c, 32'hc12f6c18} /* (21, 16, 27) {real, imag} */,
  {32'hc0e6b13d, 32'hc00f2c91} /* (21, 16, 26) {real, imag} */,
  {32'hbf26ee7a, 32'hc0804ccc} /* (21, 16, 25) {real, imag} */,
  {32'h402c2e4c, 32'h3e0f2390} /* (21, 16, 24) {real, imag} */,
  {32'hbf103a08, 32'h40c7bc36} /* (21, 16, 23) {real, imag} */,
  {32'h40fbdecb, 32'hbeea0fae} /* (21, 16, 22) {real, imag} */,
  {32'hc00cfb3c, 32'hc064e78c} /* (21, 16, 21) {real, imag} */,
  {32'h407fbb09, 32'hc1042226} /* (21, 16, 20) {real, imag} */,
  {32'hc0dda24e, 32'hc0fcaad3} /* (21, 16, 19) {real, imag} */,
  {32'h4034d51c, 32'hc045ca76} /* (21, 16, 18) {real, imag} */,
  {32'h3f9d5bb5, 32'hbf6eead0} /* (21, 16, 17) {real, imag} */,
  {32'hc0587578, 32'h00000000} /* (21, 16, 16) {real, imag} */,
  {32'h3f9d5bb5, 32'h3f6eead0} /* (21, 16, 15) {real, imag} */,
  {32'h4034d51c, 32'h4045ca76} /* (21, 16, 14) {real, imag} */,
  {32'hc0dda24e, 32'h40fcaad3} /* (21, 16, 13) {real, imag} */,
  {32'h407fbb09, 32'h41042226} /* (21, 16, 12) {real, imag} */,
  {32'hc00cfb3c, 32'h4064e78c} /* (21, 16, 11) {real, imag} */,
  {32'h40fbdecb, 32'h3eea0fae} /* (21, 16, 10) {real, imag} */,
  {32'hbf103a08, 32'hc0c7bc36} /* (21, 16, 9) {real, imag} */,
  {32'h402c2e4c, 32'hbe0f2390} /* (21, 16, 8) {real, imag} */,
  {32'hbf26ee7a, 32'h40804ccc} /* (21, 16, 7) {real, imag} */,
  {32'hc0e6b13d, 32'h400f2c91} /* (21, 16, 6) {real, imag} */,
  {32'hbf49ad3c, 32'h412f6c18} /* (21, 16, 5) {real, imag} */,
  {32'hc154b3ee, 32'h40883c57} /* (21, 16, 4) {real, imag} */,
  {32'hbfb037fd, 32'h40b099b7} /* (21, 16, 3) {real, imag} */,
  {32'h40426d33, 32'h40cfed72} /* (21, 16, 2) {real, imag} */,
  {32'h405cb700, 32'hbfa53ea5} /* (21, 16, 1) {real, imag} */,
  {32'h410d583c, 32'h00000000} /* (21, 16, 0) {real, imag} */,
  {32'h4114ec56, 32'hc03f8abc} /* (21, 15, 31) {real, imag} */,
  {32'hc05d4069, 32'hc052980f} /* (21, 15, 30) {real, imag} */,
  {32'h4094546c, 32'h40621393} /* (21, 15, 29) {real, imag} */,
  {32'h40796fe4, 32'h3d7c8a40} /* (21, 15, 28) {real, imag} */,
  {32'hc0789d30, 32'hc0b23947} /* (21, 15, 27) {real, imag} */,
  {32'hc0a8ffbd, 32'h404037ad} /* (21, 15, 26) {real, imag} */,
  {32'hbf9c5f84, 32'hc0ae5b57} /* (21, 15, 25) {real, imag} */,
  {32'hc11c109c, 32'hc0825cec} /* (21, 15, 24) {real, imag} */,
  {32'h410e07b5, 32'hbebf8bb0} /* (21, 15, 23) {real, imag} */,
  {32'hc153e3bc, 32'hc0e794e5} /* (21, 15, 22) {real, imag} */,
  {32'hc18968f4, 32'h41485712} /* (21, 15, 21) {real, imag} */,
  {32'h40167124, 32'hc0234208} /* (21, 15, 20) {real, imag} */,
  {32'hbfaca420, 32'hc0bd52ca} /* (21, 15, 19) {real, imag} */,
  {32'h3febcdf8, 32'h407f792c} /* (21, 15, 18) {real, imag} */,
  {32'h40f9a65b, 32'h4168c672} /* (21, 15, 17) {real, imag} */,
  {32'hc10fdc35, 32'hc11bf7d1} /* (21, 15, 16) {real, imag} */,
  {32'h40180bc4, 32'h414b03f1} /* (21, 15, 15) {real, imag} */,
  {32'hc06fac64, 32'hc0e65399} /* (21, 15, 14) {real, imag} */,
  {32'hc00a344a, 32'hc0bb83fa} /* (21, 15, 13) {real, imag} */,
  {32'h41031d19, 32'hc08bd5c3} /* (21, 15, 12) {real, imag} */,
  {32'h409745dd, 32'h417db58e} /* (21, 15, 11) {real, imag} */,
  {32'h4180b474, 32'hc098440f} /* (21, 15, 10) {real, imag} */,
  {32'hc0b0f7ce, 32'h409caaa6} /* (21, 15, 9) {real, imag} */,
  {32'hc109b7d9, 32'hc073c8f9} /* (21, 15, 8) {real, imag} */,
  {32'hbf92ed96, 32'hbf854af0} /* (21, 15, 7) {real, imag} */,
  {32'hbf10627c, 32'hbfc12628} /* (21, 15, 6) {real, imag} */,
  {32'hc13ef61c, 32'hc0c52c81} /* (21, 15, 5) {real, imag} */,
  {32'hc152df54, 32'h40aa5e72} /* (21, 15, 4) {real, imag} */,
  {32'h3f6eedf8, 32'hc09cd37a} /* (21, 15, 3) {real, imag} */,
  {32'h41029f17, 32'h410edd29} /* (21, 15, 2) {real, imag} */,
  {32'h40a66ace, 32'h40ee319a} /* (21, 15, 1) {real, imag} */,
  {32'h40de4622, 32'hc0e8eed8} /* (21, 15, 0) {real, imag} */,
  {32'h40f2a63a, 32'h41879689} /* (21, 14, 31) {real, imag} */,
  {32'hc10add00, 32'hc0149a74} /* (21, 14, 30) {real, imag} */,
  {32'h411e0726, 32'hc091b13e} /* (21, 14, 29) {real, imag} */,
  {32'h41426593, 32'hbf71c950} /* (21, 14, 28) {real, imag} */,
  {32'hc036d4b6, 32'hc0114870} /* (21, 14, 27) {real, imag} */,
  {32'hbf7b7c78, 32'h415517f9} /* (21, 14, 26) {real, imag} */,
  {32'h3ea46134, 32'h4160f968} /* (21, 14, 25) {real, imag} */,
  {32'hc15f24ac, 32'hc0fcdbc3} /* (21, 14, 24) {real, imag} */,
  {32'hc017d881, 32'hc0c96d20} /* (21, 14, 23) {real, imag} */,
  {32'hc167251c, 32'h4010e9d8} /* (21, 14, 22) {real, imag} */,
  {32'hc15b3e08, 32'h40dd6808} /* (21, 14, 21) {real, imag} */,
  {32'hc12e6808, 32'hc07dc60b} /* (21, 14, 20) {real, imag} */,
  {32'hc031b4a2, 32'h414fdd0b} /* (21, 14, 19) {real, imag} */,
  {32'h4106f027, 32'h40575cda} /* (21, 14, 18) {real, imag} */,
  {32'hc183cd7d, 32'hbf9548a8} /* (21, 14, 17) {real, imag} */,
  {32'hbf8dd91c, 32'hc09b7f06} /* (21, 14, 16) {real, imag} */,
  {32'h4071874a, 32'hc17703d2} /* (21, 14, 15) {real, imag} */,
  {32'hc0491cd0, 32'hc0e6abbb} /* (21, 14, 14) {real, imag} */,
  {32'h403f3104, 32'h40d41ce2} /* (21, 14, 13) {real, imag} */,
  {32'h41b0c67d, 32'hc15087e4} /* (21, 14, 12) {real, imag} */,
  {32'h411e0c5a, 32'h405c9eb8} /* (21, 14, 11) {real, imag} */,
  {32'h404ed554, 32'h4151d598} /* (21, 14, 10) {real, imag} */,
  {32'hc10debd2, 32'h418ec8ed} /* (21, 14, 9) {real, imag} */,
  {32'h413dd722, 32'hbe30f320} /* (21, 14, 8) {real, imag} */,
  {32'hc16c80f0, 32'h40d6b64c} /* (21, 14, 7) {real, imag} */,
  {32'hc0fb3f8d, 32'hbec1cd4c} /* (21, 14, 6) {real, imag} */,
  {32'hc0ea76c5, 32'hc0d7e048} /* (21, 14, 5) {real, imag} */,
  {32'h40381b2c, 32'h402d413c} /* (21, 14, 4) {real, imag} */,
  {32'h4060e670, 32'hbfb59948} /* (21, 14, 3) {real, imag} */,
  {32'hc0b8d353, 32'h400094ff} /* (21, 14, 2) {real, imag} */,
  {32'hc0e3447a, 32'h3e18d2c0} /* (21, 14, 1) {real, imag} */,
  {32'hc0e848e2, 32'h41797276} /* (21, 14, 0) {real, imag} */,
  {32'h410e1954, 32'h4057b80c} /* (21, 13, 31) {real, imag} */,
  {32'hc19653eb, 32'hc04ccd78} /* (21, 13, 30) {real, imag} */,
  {32'h41205238, 32'h418398e4} /* (21, 13, 29) {real, imag} */,
  {32'hc0925ba1, 32'hc0c47b43} /* (21, 13, 28) {real, imag} */,
  {32'hc0568c1b, 32'hc08c65f3} /* (21, 13, 27) {real, imag} */,
  {32'hc1a99d4e, 32'hc09f4bd1} /* (21, 13, 26) {real, imag} */,
  {32'hc0a72ef9, 32'h417cd96e} /* (21, 13, 25) {real, imag} */,
  {32'h40e00d04, 32'hc17de83a} /* (21, 13, 24) {real, imag} */,
  {32'h40c62d96, 32'hc0a4c1a2} /* (21, 13, 23) {real, imag} */,
  {32'h41343332, 32'h3f2834a8} /* (21, 13, 22) {real, imag} */,
  {32'h3fed0438, 32'h40a9e829} /* (21, 13, 21) {real, imag} */,
  {32'h40777974, 32'h40311f74} /* (21, 13, 20) {real, imag} */,
  {32'hc12b57ff, 32'h40e5f7ca} /* (21, 13, 19) {real, imag} */,
  {32'h410453f5, 32'h4107564b} /* (21, 13, 18) {real, imag} */,
  {32'hc0a24e52, 32'hc0dcc876} /* (21, 13, 17) {real, imag} */,
  {32'hc13792a9, 32'hc03834fc} /* (21, 13, 16) {real, imag} */,
  {32'h3f2a46b6, 32'hbfdbb3c0} /* (21, 13, 15) {real, imag} */,
  {32'h419cff7f, 32'h40c2c5f0} /* (21, 13, 14) {real, imag} */,
  {32'h4130e958, 32'hbfdfa6d0} /* (21, 13, 13) {real, imag} */,
  {32'hc10cef3e, 32'h41456134} /* (21, 13, 12) {real, imag} */,
  {32'h4121ccf5, 32'hc1a6c184} /* (21, 13, 11) {real, imag} */,
  {32'hc158e6e0, 32'h40d54c50} /* (21, 13, 10) {real, imag} */,
  {32'hc04f3b62, 32'hc041f490} /* (21, 13, 9) {real, imag} */,
  {32'h418fc9c8, 32'h4144021e} /* (21, 13, 8) {real, imag} */,
  {32'hbc7e5c00, 32'hc0bf9283} /* (21, 13, 7) {real, imag} */,
  {32'hc132b89e, 32'h41bfb61a} /* (21, 13, 6) {real, imag} */,
  {32'h4123eeb4, 32'hc190c37e} /* (21, 13, 5) {real, imag} */,
  {32'h413de89d, 32'hc10b7ac3} /* (21, 13, 4) {real, imag} */,
  {32'hc1132e18, 32'hbfd078b6} /* (21, 13, 3) {real, imag} */,
  {32'hc14e4ac1, 32'hbe4ef6c0} /* (21, 13, 2) {real, imag} */,
  {32'hc1b92bb0, 32'hc1164d96} /* (21, 13, 1) {real, imag} */,
  {32'hc105b42f, 32'hbffff12c} /* (21, 13, 0) {real, imag} */,
  {32'hc08aa9d4, 32'h3f7815f8} /* (21, 12, 31) {real, imag} */,
  {32'hc16ef9f8, 32'hc078f5c0} /* (21, 12, 30) {real, imag} */,
  {32'h3f3f81d4, 32'hc12a7a2a} /* (21, 12, 29) {real, imag} */,
  {32'hc0a73185, 32'h40d0b578} /* (21, 12, 28) {real, imag} */,
  {32'h3f819ee2, 32'hc141e1db} /* (21, 12, 27) {real, imag} */,
  {32'hc1b8cb9c, 32'h40bc2390} /* (21, 12, 26) {real, imag} */,
  {32'h411e026b, 32'hbe4cf3e0} /* (21, 12, 25) {real, imag} */,
  {32'h40281c7c, 32'h412dca3f} /* (21, 12, 24) {real, imag} */,
  {32'h4176d3e8, 32'hc037c210} /* (21, 12, 23) {real, imag} */,
  {32'h404d7a84, 32'h3ecc0a0c} /* (21, 12, 22) {real, imag} */,
  {32'h41efbce0, 32'h40a2bd34} /* (21, 12, 21) {real, imag} */,
  {32'h40d54c5c, 32'hc192df42} /* (21, 12, 20) {real, imag} */,
  {32'h401a5cd7, 32'hc00409fe} /* (21, 12, 19) {real, imag} */,
  {32'h4101ce7e, 32'hc1628062} /* (21, 12, 18) {real, imag} */,
  {32'h41622385, 32'h412e5653} /* (21, 12, 17) {real, imag} */,
  {32'hc0d1ea52, 32'h40cf51a4} /* (21, 12, 16) {real, imag} */,
  {32'h40da2d46, 32'hc13b5ea0} /* (21, 12, 15) {real, imag} */,
  {32'h40b9a501, 32'h3f9eb0f8} /* (21, 12, 14) {real, imag} */,
  {32'h40dbc5a7, 32'h403b9e45} /* (21, 12, 13) {real, imag} */,
  {32'h41754a2c, 32'h4170b9b0} /* (21, 12, 12) {real, imag} */,
  {32'hc18bdb46, 32'h401bb139} /* (21, 12, 11) {real, imag} */,
  {32'hc02fe40e, 32'h40eb3ab6} /* (21, 12, 10) {real, imag} */,
  {32'h40da209b, 32'hc0efd856} /* (21, 12, 9) {real, imag} */,
  {32'hc143acc6, 32'h413351a6} /* (21, 12, 8) {real, imag} */,
  {32'hc1a023c8, 32'h40372dbc} /* (21, 12, 7) {real, imag} */,
  {32'h410e0ffa, 32'h403b274c} /* (21, 12, 6) {real, imag} */,
  {32'h4103ad56, 32'hc01a7554} /* (21, 12, 5) {real, imag} */,
  {32'h41088516, 32'hc044c705} /* (21, 12, 4) {real, imag} */,
  {32'hc0d5dadd, 32'h40a2dad7} /* (21, 12, 3) {real, imag} */,
  {32'h405416f6, 32'hc0c470b4} /* (21, 12, 2) {real, imag} */,
  {32'h4050d53d, 32'hc0a28556} /* (21, 12, 1) {real, imag} */,
  {32'h41c9bc09, 32'h4129d1c4} /* (21, 12, 0) {real, imag} */,
  {32'h41201852, 32'h4069af7e} /* (21, 11, 31) {real, imag} */,
  {32'hc1cade5b, 32'h401c217d} /* (21, 11, 30) {real, imag} */,
  {32'h4011d856, 32'h4080797b} /* (21, 11, 29) {real, imag} */,
  {32'hc1a73d46, 32'h408f4f5f} /* (21, 11, 28) {real, imag} */,
  {32'hc02072f2, 32'h4130e5fe} /* (21, 11, 27) {real, imag} */,
  {32'hc17904e3, 32'hc0cd8ff0} /* (21, 11, 26) {real, imag} */,
  {32'hc0fa8bf8, 32'h40600e0c} /* (21, 11, 25) {real, imag} */,
  {32'h4125f604, 32'hc066f3b2} /* (21, 11, 24) {real, imag} */,
  {32'h3f879a6c, 32'hbfc24928} /* (21, 11, 23) {real, imag} */,
  {32'h41579ee8, 32'hc0f8d3b0} /* (21, 11, 22) {real, imag} */,
  {32'hc0fccd98, 32'h411b2a41} /* (21, 11, 21) {real, imag} */,
  {32'h40b21faa, 32'h3ece1ec0} /* (21, 11, 20) {real, imag} */,
  {32'h4134ea39, 32'h40ef7f97} /* (21, 11, 19) {real, imag} */,
  {32'h41684bbe, 32'hc1913ff1} /* (21, 11, 18) {real, imag} */,
  {32'hc083a6ec, 32'hc0af1030} /* (21, 11, 17) {real, imag} */,
  {32'hc15caec6, 32'h411c11e5} /* (21, 11, 16) {real, imag} */,
  {32'h40083876, 32'hc104a76e} /* (21, 11, 15) {real, imag} */,
  {32'h3df89b40, 32'h4096a9c6} /* (21, 11, 14) {real, imag} */,
  {32'hc0197313, 32'h406049f6} /* (21, 11, 13) {real, imag} */,
  {32'hc144da70, 32'h412bc2bd} /* (21, 11, 12) {real, imag} */,
  {32'hc1864264, 32'hbf299afc} /* (21, 11, 11) {real, imag} */,
  {32'h408a3b45, 32'hbfd722d8} /* (21, 11, 10) {real, imag} */,
  {32'h414baa62, 32'hc11a7108} /* (21, 11, 9) {real, imag} */,
  {32'h416dbfbf, 32'hbddc8180} /* (21, 11, 8) {real, imag} */,
  {32'h4111a605, 32'hbfcbac38} /* (21, 11, 7) {real, imag} */,
  {32'h4145a0c2, 32'h40e652a7} /* (21, 11, 6) {real, imag} */,
  {32'h41535014, 32'hbfd4a4b0} /* (21, 11, 5) {real, imag} */,
  {32'hc115f8b0, 32'h408c445e} /* (21, 11, 4) {real, imag} */,
  {32'h41331ef5, 32'hc1838600} /* (21, 11, 3) {real, imag} */,
  {32'h40f8aa08, 32'hc1254854} /* (21, 11, 2) {real, imag} */,
  {32'h3ffa5853, 32'h4199bf30} /* (21, 11, 1) {real, imag} */,
  {32'h413ecdfb, 32'h41a917ed} /* (21, 11, 0) {real, imag} */,
  {32'h413d8b1c, 32'hc1f60b3e} /* (21, 10, 31) {real, imag} */,
  {32'h4151c0ef, 32'h41a89d7b} /* (21, 10, 30) {real, imag} */,
  {32'h403c7839, 32'hbfade910} /* (21, 10, 29) {real, imag} */,
  {32'hc1229643, 32'h405db6ef} /* (21, 10, 28) {real, imag} */,
  {32'h41106aeb, 32'h40a4f73b} /* (21, 10, 27) {real, imag} */,
  {32'h41203376, 32'h413e7db1} /* (21, 10, 26) {real, imag} */,
  {32'hc18b2b00, 32'hc06ad684} /* (21, 10, 25) {real, imag} */,
  {32'h412fb52a, 32'h40a6163e} /* (21, 10, 24) {real, imag} */,
  {32'hc1539aa6, 32'hc0c63d94} /* (21, 10, 23) {real, imag} */,
  {32'h3e5d9fb0, 32'hc10d12f5} /* (21, 10, 22) {real, imag} */,
  {32'h41a24b53, 32'hc0fabfb4} /* (21, 10, 21) {real, imag} */,
  {32'hbf14d074, 32'hc16fb11a} /* (21, 10, 20) {real, imag} */,
  {32'hc0dcbcd7, 32'hc084ae55} /* (21, 10, 19) {real, imag} */,
  {32'h3cf81c40, 32'hc0f1a102} /* (21, 10, 18) {real, imag} */,
  {32'hc111b11a, 32'h414b3cc0} /* (21, 10, 17) {real, imag} */,
  {32'h41890f35, 32'hc0d3e9ba} /* (21, 10, 16) {real, imag} */,
  {32'h40c8acb2, 32'hbecbd1d0} /* (21, 10, 15) {real, imag} */,
  {32'hbfe102ce, 32'hc0c69c80} /* (21, 10, 14) {real, imag} */,
  {32'hc0685b45, 32'hbfc28370} /* (21, 10, 13) {real, imag} */,
  {32'hc038167c, 32'h418d67e8} /* (21, 10, 12) {real, imag} */,
  {32'hc061d9e0, 32'h400c6cec} /* (21, 10, 11) {real, imag} */,
  {32'h4152a866, 32'h416fb632} /* (21, 10, 10) {real, imag} */,
  {32'hbfb3ded0, 32'hbfbab364} /* (21, 10, 9) {real, imag} */,
  {32'hc0f42492, 32'hc10457b8} /* (21, 10, 8) {real, imag} */,
  {32'hc0ffe706, 32'h406e3219} /* (21, 10, 7) {real, imag} */,
  {32'h415c72fa, 32'hc1836d7c} /* (21, 10, 6) {real, imag} */,
  {32'hc173fd64, 32'hc1680ed3} /* (21, 10, 5) {real, imag} */,
  {32'h40541328, 32'h4145d2b8} /* (21, 10, 4) {real, imag} */,
  {32'h3ffb40cc, 32'hbf16cf28} /* (21, 10, 3) {real, imag} */,
  {32'h40d91e1a, 32'hbfb69548} /* (21, 10, 2) {real, imag} */,
  {32'hc1f0e694, 32'hc1693db2} /* (21, 10, 1) {real, imag} */,
  {32'hc1dad4c8, 32'hc0cac227} /* (21, 10, 0) {real, imag} */,
  {32'h4171b561, 32'h417e8fca} /* (21, 9, 31) {real, imag} */,
  {32'hc076b3be, 32'h411d2e84} /* (21, 9, 30) {real, imag} */,
  {32'hc126acbc, 32'hc1748036} /* (21, 9, 29) {real, imag} */,
  {32'hbfd625e8, 32'hc19cf116} /* (21, 9, 28) {real, imag} */,
  {32'h404e0378, 32'hc0d6bc65} /* (21, 9, 27) {real, imag} */,
  {32'hc0784c4c, 32'h3fb77e14} /* (21, 9, 26) {real, imag} */,
  {32'hc0cae2a4, 32'h409009c5} /* (21, 9, 25) {real, imag} */,
  {32'hc08f7c11, 32'h41852dbd} /* (21, 9, 24) {real, imag} */,
  {32'hbf1f4ce4, 32'hbe0e1080} /* (21, 9, 23) {real, imag} */,
  {32'hc0b3ce7f, 32'hc187346a} /* (21, 9, 22) {real, imag} */,
  {32'hc10307d3, 32'h403a3544} /* (21, 9, 21) {real, imag} */,
  {32'h400e5c44, 32'h409bce5e} /* (21, 9, 20) {real, imag} */,
  {32'hc00c7c80, 32'hc0245668} /* (21, 9, 19) {real, imag} */,
  {32'h4125d6c7, 32'h4068cd36} /* (21, 9, 18) {real, imag} */,
  {32'hc08b4b3c, 32'hc19cc79e} /* (21, 9, 17) {real, imag} */,
  {32'hbdf5cd40, 32'h4091f94f} /* (21, 9, 16) {real, imag} */,
  {32'h4087eb8a, 32'hc0402015} /* (21, 9, 15) {real, imag} */,
  {32'h3e9be448, 32'h413ab478} /* (21, 9, 14) {real, imag} */,
  {32'hc0ac8392, 32'h40e0bb37} /* (21, 9, 13) {real, imag} */,
  {32'hc1a5acbf, 32'h40541d60} /* (21, 9, 12) {real, imag} */,
  {32'h3ea11430, 32'h4163c516} /* (21, 9, 11) {real, imag} */,
  {32'h411e3e20, 32'hc0d701c7} /* (21, 9, 10) {real, imag} */,
  {32'h41b4f97a, 32'hc0d51398} /* (21, 9, 9) {real, imag} */,
  {32'hc17b1608, 32'h40cae552} /* (21, 9, 8) {real, imag} */,
  {32'h40c15b7c, 32'hc1a23ddc} /* (21, 9, 7) {real, imag} */,
  {32'hc1496e07, 32'hc1d16a40} /* (21, 9, 6) {real, imag} */,
  {32'h41bdea61, 32'h40a89747} /* (21, 9, 5) {real, imag} */,
  {32'hc1736f04, 32'h401dd7ef} /* (21, 9, 4) {real, imag} */,
  {32'h41528adf, 32'hc131aa87} /* (21, 9, 3) {real, imag} */,
  {32'hbf882fbc, 32'h4132c967} /* (21, 9, 2) {real, imag} */,
  {32'hc1ac64f8, 32'hc03de9dc} /* (21, 9, 1) {real, imag} */,
  {32'h4186b3e3, 32'h41228e66} /* (21, 9, 0) {real, imag} */,
  {32'h42156bc1, 32'h42052325} /* (21, 8, 31) {real, imag} */,
  {32'hc1bb04cd, 32'hc151d501} /* (21, 8, 30) {real, imag} */,
  {32'h410451b2, 32'h3f7c6b18} /* (21, 8, 29) {real, imag} */,
  {32'h4075ec40, 32'h4113132b} /* (21, 8, 28) {real, imag} */,
  {32'hc1d4a9fe, 32'hc191bb49} /* (21, 8, 27) {real, imag} */,
  {32'h41f3339a, 32'hbe641a00} /* (21, 8, 26) {real, imag} */,
  {32'h40f742b3, 32'hc07803d0} /* (21, 8, 25) {real, imag} */,
  {32'hc0998693, 32'hc1828a0c} /* (21, 8, 24) {real, imag} */,
  {32'h411c3a13, 32'h411e78b7} /* (21, 8, 23) {real, imag} */,
  {32'hbe078d80, 32'hc03ab0d8} /* (21, 8, 22) {real, imag} */,
  {32'hc0709a8e, 32'h41c95788} /* (21, 8, 21) {real, imag} */,
  {32'h40a3eb8b, 32'h3fbfc9b4} /* (21, 8, 20) {real, imag} */,
  {32'h4062e398, 32'hc1541651} /* (21, 8, 19) {real, imag} */,
  {32'hc050c5dc, 32'h412a805a} /* (21, 8, 18) {real, imag} */,
  {32'h4004d4cc, 32'h3f177110} /* (21, 8, 17) {real, imag} */,
  {32'h3f87269c, 32'hc08a9782} /* (21, 8, 16) {real, imag} */,
  {32'hc0dd22dc, 32'h40ac4711} /* (21, 8, 15) {real, imag} */,
  {32'hc0ebb5b3, 32'h40051572} /* (21, 8, 14) {real, imag} */,
  {32'h3f10f380, 32'hc0f81da0} /* (21, 8, 13) {real, imag} */,
  {32'h40c4c29a, 32'hc134c39a} /* (21, 8, 12) {real, imag} */,
  {32'hbe299a40, 32'hc1c9d051} /* (21, 8, 11) {real, imag} */,
  {32'hc18db8f6, 32'h41c2438e} /* (21, 8, 10) {real, imag} */,
  {32'hbff1f840, 32'hc00c10d8} /* (21, 8, 9) {real, imag} */,
  {32'hbf4a14e0, 32'h400cafc2} /* (21, 8, 8) {real, imag} */,
  {32'hc01552f4, 32'hc0caac96} /* (21, 8, 7) {real, imag} */,
  {32'h4035b7cc, 32'h3f2bac00} /* (21, 8, 6) {real, imag} */,
  {32'hc2087754, 32'hc06ac1d4} /* (21, 8, 5) {real, imag} */,
  {32'h418738b9, 32'hc07bc962} /* (21, 8, 4) {real, imag} */,
  {32'h41720080, 32'hc0e0fefd} /* (21, 8, 3) {real, imag} */,
  {32'hc19bbb3f, 32'hc0e784d0} /* (21, 8, 2) {real, imag} */,
  {32'h41986e44, 32'h4149bbf2} /* (21, 8, 1) {real, imag} */,
  {32'h411e3e58, 32'hc0c24b1c} /* (21, 8, 0) {real, imag} */,
  {32'h3ed23780, 32'hc167c94c} /* (21, 7, 31) {real, imag} */,
  {32'h418d938f, 32'hc1c7321b} /* (21, 7, 30) {real, imag} */,
  {32'h4059f536, 32'hc0888e9b} /* (21, 7, 29) {real, imag} */,
  {32'h419e85c6, 32'h4080a594} /* (21, 7, 28) {real, imag} */,
  {32'hc1375d73, 32'h40a01ec5} /* (21, 7, 27) {real, imag} */,
  {32'hc11b75ba, 32'h41b209f8} /* (21, 7, 26) {real, imag} */,
  {32'hc12e164c, 32'h4160b147} /* (21, 7, 25) {real, imag} */,
  {32'hc09a5dd2, 32'h41812ca6} /* (21, 7, 24) {real, imag} */,
  {32'hc0974642, 32'hc0c1b15f} /* (21, 7, 23) {real, imag} */,
  {32'hc19df8cb, 32'h40aa2584} /* (21, 7, 22) {real, imag} */,
  {32'h3f443f28, 32'hc19437f4} /* (21, 7, 21) {real, imag} */,
  {32'hc0977cb0, 32'hbebdbeac} /* (21, 7, 20) {real, imag} */,
  {32'h403b437c, 32'h413cbfeb} /* (21, 7, 19) {real, imag} */,
  {32'h3ff04e38, 32'hc0b30e13} /* (21, 7, 18) {real, imag} */,
  {32'hc11b595c, 32'h4093efb4} /* (21, 7, 17) {real, imag} */,
  {32'hc0639f69, 32'hc150b56d} /* (21, 7, 16) {real, imag} */,
  {32'h3e89fca4, 32'h403591fe} /* (21, 7, 15) {real, imag} */,
  {32'hc16d2434, 32'h4040cdb8} /* (21, 7, 14) {real, imag} */,
  {32'hc012808e, 32'h40cae15b} /* (21, 7, 13) {real, imag} */,
  {32'hc0843ab3, 32'hc0cbe7ea} /* (21, 7, 12) {real, imag} */,
  {32'hc1af4b36, 32'h4162ea48} /* (21, 7, 11) {real, imag} */,
  {32'hc0cd5d66, 32'hc0d10976} /* (21, 7, 10) {real, imag} */,
  {32'hc094d9b7, 32'h4047f028} /* (21, 7, 9) {real, imag} */,
  {32'hc0f139bd, 32'h3ebeeef8} /* (21, 7, 8) {real, imag} */,
  {32'hc1b968ae, 32'hbf755d90} /* (21, 7, 7) {real, imag} */,
  {32'hc0e30ddf, 32'h4195c674} /* (21, 7, 6) {real, imag} */,
  {32'h41d5ed6c, 32'hc105035a} /* (21, 7, 5) {real, imag} */,
  {32'h3ece6d40, 32'hc135830d} /* (21, 7, 4) {real, imag} */,
  {32'h41d6105b, 32'h41626cce} /* (21, 7, 3) {real, imag} */,
  {32'h411c4d14, 32'h40def07c} /* (21, 7, 2) {real, imag} */,
  {32'h40d05b28, 32'hc0605b6f} /* (21, 7, 1) {real, imag} */,
  {32'hc1c6c9e7, 32'hc1ec1c8e} /* (21, 7, 0) {real, imag} */,
  {32'hc10be10a, 32'h42029357} /* (21, 6, 31) {real, imag} */,
  {32'h3f85c200, 32'hc0870388} /* (21, 6, 30) {real, imag} */,
  {32'h40fe0aa5, 32'h4084667a} /* (21, 6, 29) {real, imag} */,
  {32'h41ade48c, 32'hc1a0a7f5} /* (21, 6, 28) {real, imag} */,
  {32'hc0fe644c, 32'hc1baaf9d} /* (21, 6, 27) {real, imag} */,
  {32'h414a7d0e, 32'hc182638a} /* (21, 6, 26) {real, imag} */,
  {32'hc09f4018, 32'hc121a559} /* (21, 6, 25) {real, imag} */,
  {32'hc10009c6, 32'h40e6a97b} /* (21, 6, 24) {real, imag} */,
  {32'hc10dd212, 32'h4177ff78} /* (21, 6, 23) {real, imag} */,
  {32'h401c7640, 32'hc1369056} /* (21, 6, 22) {real, imag} */,
  {32'hc0e038eb, 32'hbfe60c80} /* (21, 6, 21) {real, imag} */,
  {32'hc16c2d95, 32'hbeb54f10} /* (21, 6, 20) {real, imag} */,
  {32'hc10adb2e, 32'hc12a702b} /* (21, 6, 19) {real, imag} */,
  {32'hc083c696, 32'h417db580} /* (21, 6, 18) {real, imag} */,
  {32'h418630e9, 32'h40ee77d2} /* (21, 6, 17) {real, imag} */,
  {32'hc0c23fd4, 32'hc0d62aad} /* (21, 6, 16) {real, imag} */,
  {32'h3d740f60, 32'h3ff96d5e} /* (21, 6, 15) {real, imag} */,
  {32'h40c125ea, 32'h4098adb0} /* (21, 6, 14) {real, imag} */,
  {32'hbfad5b67, 32'hc173bb01} /* (21, 6, 13) {real, imag} */,
  {32'hc11b616e, 32'h4085f412} /* (21, 6, 12) {real, imag} */,
  {32'hc191e8c2, 32'hc18066cb} /* (21, 6, 11) {real, imag} */,
  {32'h3e56bf00, 32'h4198492c} /* (21, 6, 10) {real, imag} */,
  {32'h3f464030, 32'h4162f9c7} /* (21, 6, 9) {real, imag} */,
  {32'hc0852d8a, 32'hc1af788c} /* (21, 6, 8) {real, imag} */,
  {32'hc0f65d1e, 32'hc015ea8a} /* (21, 6, 7) {real, imag} */,
  {32'hc150a914, 32'hc190b2ee} /* (21, 6, 6) {real, imag} */,
  {32'hc1b87360, 32'h40bee95d} /* (21, 6, 5) {real, imag} */,
  {32'hc08c1600, 32'h401647d1} /* (21, 6, 4) {real, imag} */,
  {32'h419b20b3, 32'hc1a50a81} /* (21, 6, 3) {real, imag} */,
  {32'h408e3884, 32'h41b83a26} /* (21, 6, 2) {real, imag} */,
  {32'hc050f7c8, 32'h412c6f77} /* (21, 6, 1) {real, imag} */,
  {32'hc0d33a47, 32'h4095f1e1} /* (21, 6, 0) {real, imag} */,
  {32'h42bd67e2, 32'h41618323} /* (21, 5, 31) {real, imag} */,
  {32'hc203cf70, 32'hc153c5f0} /* (21, 5, 30) {real, imag} */,
  {32'h3fe74b80, 32'h414f53e4} /* (21, 5, 29) {real, imag} */,
  {32'h4195423c, 32'hc0e2c888} /* (21, 5, 28) {real, imag} */,
  {32'hc1f38dee, 32'hc047c98c} /* (21, 5, 27) {real, imag} */,
  {32'hc1d9b72e, 32'h4037449e} /* (21, 5, 26) {real, imag} */,
  {32'h410d6142, 32'h3fa8dfde} /* (21, 5, 25) {real, imag} */,
  {32'hc0aa8644, 32'h40a47504} /* (21, 5, 24) {real, imag} */,
  {32'h3ff5a488, 32'h40d32f05} /* (21, 5, 23) {real, imag} */,
  {32'hc0bd7857, 32'hbd404700} /* (21, 5, 22) {real, imag} */,
  {32'hbed0e568, 32'hc0d7b5ce} /* (21, 5, 21) {real, imag} */,
  {32'h4125506a, 32'h4102bb36} /* (21, 5, 20) {real, imag} */,
  {32'hc00e23e8, 32'h3fedb4dc} /* (21, 5, 19) {real, imag} */,
  {32'hbfc49b52, 32'h4060551e} /* (21, 5, 18) {real, imag} */,
  {32'h40ab4179, 32'hc11c60db} /* (21, 5, 17) {real, imag} */,
  {32'hc0ac0092, 32'h404b97be} /* (21, 5, 16) {real, imag} */,
  {32'hc0cee78c, 32'h3db69a00} /* (21, 5, 15) {real, imag} */,
  {32'hc1133b91, 32'hc0213344} /* (21, 5, 14) {real, imag} */,
  {32'h40a62d48, 32'hbf2a5670} /* (21, 5, 13) {real, imag} */,
  {32'hc0aa43d0, 32'hc1040ba6} /* (21, 5, 12) {real, imag} */,
  {32'hc10f9e70, 32'hc192d404} /* (21, 5, 11) {real, imag} */,
  {32'h41067b40, 32'h40c7d274} /* (21, 5, 10) {real, imag} */,
  {32'h40fe9a15, 32'hc17a41a2} /* (21, 5, 9) {real, imag} */,
  {32'hc0cda84b, 32'hc0412ed0} /* (21, 5, 8) {real, imag} */,
  {32'h42074d8c, 32'h414d9639} /* (21, 5, 7) {real, imag} */,
  {32'h40f9787c, 32'hc1236fe8} /* (21, 5, 6) {real, imag} */,
  {32'hc1939dd8, 32'hc181563d} /* (21, 5, 5) {real, imag} */,
  {32'hc163baf0, 32'h4194d418} /* (21, 5, 4) {real, imag} */,
  {32'h41123773, 32'h4114306c} /* (21, 5, 3) {real, imag} */,
  {32'hc17f4f69, 32'hc23ca04f} /* (21, 5, 2) {real, imag} */,
  {32'h4281da38, 32'h428106c8} /* (21, 5, 1) {real, imag} */,
  {32'h42162774, 32'h4295cd98} /* (21, 5, 0) {real, imag} */,
  {32'hc1f6f992, 32'hc2d9fc9f} /* (21, 4, 31) {real, imag} */,
  {32'h42c1bff3, 32'h426864da} /* (21, 4, 30) {real, imag} */,
  {32'h40b570c2, 32'h3e945e20} /* (21, 4, 29) {real, imag} */,
  {32'hc1926db6, 32'h41b739ac} /* (21, 4, 28) {real, imag} */,
  {32'h405ffa2e, 32'hc1c7ef34} /* (21, 4, 27) {real, imag} */,
  {32'h41204934, 32'hc1a774f2} /* (21, 4, 26) {real, imag} */,
  {32'h4116f032, 32'h419d6c32} /* (21, 4, 25) {real, imag} */,
  {32'h414f046c, 32'h40f53f05} /* (21, 4, 24) {real, imag} */,
  {32'hc1150669, 32'hc0863eb5} /* (21, 4, 23) {real, imag} */,
  {32'hc1157701, 32'h401548d7} /* (21, 4, 22) {real, imag} */,
  {32'hc18c8005, 32'hc1055968} /* (21, 4, 21) {real, imag} */,
  {32'h418a8a6d, 32'h418f7464} /* (21, 4, 20) {real, imag} */,
  {32'hc0c1e5b0, 32'h419a8f9a} /* (21, 4, 19) {real, imag} */,
  {32'h418a62ac, 32'h41602be6} /* (21, 4, 18) {real, imag} */,
  {32'h3fb1349c, 32'h40529ae4} /* (21, 4, 17) {real, imag} */,
  {32'hc0b700a2, 32'h3fddcf24} /* (21, 4, 16) {real, imag} */,
  {32'h404a15a4, 32'hbe453428} /* (21, 4, 15) {real, imag} */,
  {32'h3e2af9e0, 32'hc101ceea} /* (21, 4, 14) {real, imag} */,
  {32'hc10e3c3a, 32'hc1b15bb6} /* (21, 4, 13) {real, imag} */,
  {32'hc0e39be7, 32'h3fb75a0f} /* (21, 4, 12) {real, imag} */,
  {32'h4198bac7, 32'h40879407} /* (21, 4, 11) {real, imag} */,
  {32'h409cdff2, 32'hc08616f5} /* (21, 4, 10) {real, imag} */,
  {32'h403a87e8, 32'h3fe14bb4} /* (21, 4, 9) {real, imag} */,
  {32'h41b19a4d, 32'h413b8a99} /* (21, 4, 8) {real, imag} */,
  {32'hc190d2e4, 32'h409e8fe7} /* (21, 4, 7) {real, imag} */,
  {32'hbf8863c8, 32'h3f982d08} /* (21, 4, 6) {real, imag} */,
  {32'h41bcfe58, 32'h4110531e} /* (21, 4, 5) {real, imag} */,
  {32'h41cf7a63, 32'hc20587ad} /* (21, 4, 4) {real, imag} */,
  {32'hc06aabe0, 32'hc218af4a} /* (21, 4, 3) {real, imag} */,
  {32'h42f36fd0, 32'h4270705c} /* (21, 4, 2) {real, imag} */,
  {32'hc30e25c0, 32'hc26c4de8} /* (21, 4, 1) {real, imag} */,
  {32'hc283df29, 32'h42280a95} /* (21, 4, 0) {real, imag} */,
  {32'h4313f214, 32'hc2a111e1} /* (21, 3, 31) {real, imag} */,
  {32'hc2cf5563, 32'h42c5f0e9} /* (21, 3, 30) {real, imag} */,
  {32'hc11a8dcb, 32'h407924b9} /* (21, 3, 29) {real, imag} */,
  {32'hc2447536, 32'hc21809de} /* (21, 3, 28) {real, imag} */,
  {32'h417fad59, 32'hc0720d54} /* (21, 3, 27) {real, imag} */,
  {32'h410e44fc, 32'hc1da7e81} /* (21, 3, 26) {real, imag} */,
  {32'hc1d3e032, 32'hc09bda4a} /* (21, 3, 25) {real, imag} */,
  {32'h41b6d850, 32'h40dd6283} /* (21, 3, 24) {real, imag} */,
  {32'hbf952e9c, 32'hc1ad83df} /* (21, 3, 23) {real, imag} */,
  {32'hc0efc6db, 32'hc1cb9a10} /* (21, 3, 22) {real, imag} */,
  {32'h4131061a, 32'h41a00dd0} /* (21, 3, 21) {real, imag} */,
  {32'h418a5966, 32'h4195f017} /* (21, 3, 20) {real, imag} */,
  {32'h417cfb7d, 32'hc11d4fff} /* (21, 3, 19) {real, imag} */,
  {32'hc0e1615e, 32'hc1473e02} /* (21, 3, 18) {real, imag} */,
  {32'h3f76f1b8, 32'h3fa8d270} /* (21, 3, 17) {real, imag} */,
  {32'h418005d1, 32'h402f0124} /* (21, 3, 16) {real, imag} */,
  {32'h411a784b, 32'h3f065550} /* (21, 3, 15) {real, imag} */,
  {32'hbefc3aa0, 32'h41473263} /* (21, 3, 14) {real, imag} */,
  {32'h404fdacc, 32'hbf23a002} /* (21, 3, 13) {real, imag} */,
  {32'hbfb73850, 32'h412b0e13} /* (21, 3, 12) {real, imag} */,
  {32'hc06e3a9a, 32'h40bf8c20} /* (21, 3, 11) {real, imag} */,
  {32'h40d1a864, 32'h413d6069} /* (21, 3, 10) {real, imag} */,
  {32'hc1da58ce, 32'h3fec76c4} /* (21, 3, 9) {real, imag} */,
  {32'hc183c27e, 32'h41592208} /* (21, 3, 8) {real, imag} */,
  {32'h419dc7dc, 32'hc1352d3f} /* (21, 3, 7) {real, imag} */,
  {32'hbfa49684, 32'hc01a418a} /* (21, 3, 6) {real, imag} */,
  {32'hc10b83c6, 32'hc0639be2} /* (21, 3, 5) {real, imag} */,
  {32'h42312b07, 32'hc2324670} /* (21, 3, 4) {real, imag} */,
  {32'h424ac748, 32'h411a2c5a} /* (21, 3, 3) {real, imag} */,
  {32'hc1052833, 32'h42e586ac} /* (21, 3, 2) {real, imag} */,
  {32'hc308adde, 32'hc2b7548c} /* (21, 3, 1) {real, imag} */,
  {32'h4240fea0, 32'h413207d2} /* (21, 3, 0) {real, imag} */,
  {32'h44a46bad, 32'h41875c0a} /* (21, 2, 31) {real, imag} */,
  {32'hc4143477, 32'h436680f3} /* (21, 2, 30) {real, imag} */,
  {32'hbf250508, 32'h40ed6e25} /* (21, 2, 29) {real, imag} */,
  {32'h40a32870, 32'hc27e464c} /* (21, 2, 28) {real, imag} */,
  {32'hc2276feb, 32'h41eac712} /* (21, 2, 27) {real, imag} */,
  {32'hbfbdb5d8, 32'h41674c88} /* (21, 2, 26) {real, imag} */,
  {32'h41c0fc76, 32'hc19a725e} /* (21, 2, 25) {real, imag} */,
  {32'hc1f90397, 32'h423aeb5f} /* (21, 2, 24) {real, imag} */,
  {32'hc16d993a, 32'h40233836} /* (21, 2, 23) {real, imag} */,
  {32'hc160899b, 32'hbe80c098} /* (21, 2, 22) {real, imag} */,
  {32'h3fbad3fc, 32'h409abe48} /* (21, 2, 21) {real, imag} */,
  {32'h4113a82e, 32'hc0949d28} /* (21, 2, 20) {real, imag} */,
  {32'hc017e177, 32'hc0861f04} /* (21, 2, 19) {real, imag} */,
  {32'hc19d12a0, 32'h40c620c8} /* (21, 2, 18) {real, imag} */,
  {32'h3f8e6650, 32'hc141acdc} /* (21, 2, 17) {real, imag} */,
  {32'hc100017b, 32'h3fb73352} /* (21, 2, 16) {real, imag} */,
  {32'hc053f85c, 32'h40b4ccda} /* (21, 2, 15) {real, imag} */,
  {32'h40e2beec, 32'hc1c15f93} /* (21, 2, 14) {real, imag} */,
  {32'hc09167ec, 32'h4120187a} /* (21, 2, 13) {real, imag} */,
  {32'h4105be9e, 32'h4018c694} /* (21, 2, 12) {real, imag} */,
  {32'h3f1ecd74, 32'hc1919470} /* (21, 2, 11) {real, imag} */,
  {32'h41376366, 32'hc07cbe30} /* (21, 2, 10) {real, imag} */,
  {32'h41683a34, 32'hc0a6cceb} /* (21, 2, 9) {real, imag} */,
  {32'hc1729192, 32'hc1f64f98} /* (21, 2, 8) {real, imag} */,
  {32'h3fe8248e, 32'hc1386ddf} /* (21, 2, 7) {real, imag} */,
  {32'h407b8667, 32'h4132b07d} /* (21, 2, 6) {real, imag} */,
  {32'hc2adfe11, 32'hc269ac94} /* (21, 2, 5) {real, imag} */,
  {32'h42c42db8, 32'h41a83ce5} /* (21, 2, 4) {real, imag} */,
  {32'h405090d0, 32'hc1d58fc4} /* (21, 2, 3) {real, imag} */,
  {32'hc3c92148, 32'h42bbd477} /* (21, 2, 2) {real, imag} */,
  {32'h4443ca46, 32'hc2d46b7e} /* (21, 2, 1) {real, imag} */,
  {32'h4424705c, 32'h43073b9c} /* (21, 2, 0) {real, imag} */,
  {32'hc4e15558, 32'h43f3fda5} /* (21, 1, 31) {real, imag} */,
  {32'h43f436ba, 32'h41ab5ccb} /* (21, 1, 30) {real, imag} */,
  {32'h407047d0, 32'hc26920f2} /* (21, 1, 29) {real, imag} */,
  {32'hc2dc6d9a, 32'hc2c9a8ce} /* (21, 1, 28) {real, imag} */,
  {32'h43076ed6, 32'hc16832f8} /* (21, 1, 27) {real, imag} */,
  {32'h41134a2f, 32'hc1e0eaff} /* (21, 1, 26) {real, imag} */,
  {32'h40bc3e07, 32'hc1966f83} /* (21, 1, 25) {real, imag} */,
  {32'h404a2924, 32'hc1880721} /* (21, 1, 24) {real, imag} */,
  {32'h41a87ea4, 32'hc176d706} /* (21, 1, 23) {real, imag} */,
  {32'h41ffed07, 32'hc054a3f8} /* (21, 1, 22) {real, imag} */,
  {32'h41f002f3, 32'h40d28a8b} /* (21, 1, 21) {real, imag} */,
  {32'h413ec4fc, 32'h403892db} /* (21, 1, 20) {real, imag} */,
  {32'hbfb4d968, 32'hc12ac105} /* (21, 1, 19) {real, imag} */,
  {32'h408bc460, 32'h40a21341} /* (21, 1, 18) {real, imag} */,
  {32'h41863785, 32'h3f85abc0} /* (21, 1, 17) {real, imag} */,
  {32'hbf58c234, 32'hc0cda5c6} /* (21, 1, 16) {real, imag} */,
  {32'hc087d492, 32'hc0e822ca} /* (21, 1, 15) {real, imag} */,
  {32'hc110b2e6, 32'h411142ca} /* (21, 1, 14) {real, imag} */,
  {32'hbf87e6e0, 32'hc17b8434} /* (21, 1, 13) {real, imag} */,
  {32'h404d9fd2, 32'h41a121f0} /* (21, 1, 12) {real, imag} */,
  {32'h40c3dd87, 32'h41d59e6a} /* (21, 1, 11) {real, imag} */,
  {32'hc1727c7c, 32'hc067abec} /* (21, 1, 10) {real, imag} */,
  {32'h4218a2bd, 32'h411d4159} /* (21, 1, 9) {real, imag} */,
  {32'h40d77b58, 32'h4234bb8a} /* (21, 1, 8) {real, imag} */,
  {32'h4061fdc8, 32'hc1ce4f79} /* (21, 1, 7) {real, imag} */,
  {32'hc115ca7d, 32'hc0d7d8f4} /* (21, 1, 6) {real, imag} */,
  {32'h42854e6c, 32'h4280f509} /* (21, 1, 5) {real, imag} */,
  {32'hc1c67fe8, 32'hc29162c8} /* (21, 1, 4) {real, imag} */,
  {32'h426163fa, 32'h41a846d6} /* (21, 1, 3) {real, imag} */,
  {32'h440f4c17, 32'h44104db4} /* (21, 1, 2) {real, imag} */,
  {32'hc51ee7a3, 32'hc4aa4da7} /* (21, 1, 1) {real, imag} */,
  {32'hc50a002c, 32'hc3a856a6} /* (21, 1, 0) {real, imag} */,
  {32'hc4c4a908, 32'h449a1a0d} /* (21, 0, 31) {real, imag} */,
  {32'h4343e9a1, 32'hc3a10a2c} /* (21, 0, 30) {real, imag} */,
  {32'hc0b1fe24, 32'hc0738e28} /* (21, 0, 29) {real, imag} */,
  {32'hbe5d2e00, 32'hc2835dc0} /* (21, 0, 28) {real, imag} */,
  {32'h42a00ea0, 32'hc080cdd4} /* (21, 0, 27) {real, imag} */,
  {32'hc142f0fe, 32'hc14368f9} /* (21, 0, 26) {real, imag} */,
  {32'h416bdc93, 32'h41e8391c} /* (21, 0, 25) {real, imag} */,
  {32'h40d0c002, 32'hc1aa21d3} /* (21, 0, 24) {real, imag} */,
  {32'h40ccff6e, 32'h41d13dec} /* (21, 0, 23) {real, imag} */,
  {32'h4147efb0, 32'hc1365d92} /* (21, 0, 22) {real, imag} */,
  {32'hc169e5da, 32'hbfdf9992} /* (21, 0, 21) {real, imag} */,
  {32'hc0fe1e0f, 32'hc14edc24} /* (21, 0, 20) {real, imag} */,
  {32'h40b61723, 32'h3fd7c418} /* (21, 0, 19) {real, imag} */,
  {32'h40b62747, 32'hc0c656ad} /* (21, 0, 18) {real, imag} */,
  {32'hc13bfcb5, 32'h40205f4e} /* (21, 0, 17) {real, imag} */,
  {32'h41621bba, 32'h00000000} /* (21, 0, 16) {real, imag} */,
  {32'hc13bfcb5, 32'hc0205f4e} /* (21, 0, 15) {real, imag} */,
  {32'h40b62747, 32'h40c656ad} /* (21, 0, 14) {real, imag} */,
  {32'h40b61723, 32'hbfd7c418} /* (21, 0, 13) {real, imag} */,
  {32'hc0fe1e0f, 32'h414edc24} /* (21, 0, 12) {real, imag} */,
  {32'hc169e5da, 32'h3fdf9992} /* (21, 0, 11) {real, imag} */,
  {32'h4147efb0, 32'h41365d92} /* (21, 0, 10) {real, imag} */,
  {32'h40ccff6e, 32'hc1d13dec} /* (21, 0, 9) {real, imag} */,
  {32'h40d0c002, 32'h41aa21d3} /* (21, 0, 8) {real, imag} */,
  {32'h416bdc93, 32'hc1e8391c} /* (21, 0, 7) {real, imag} */,
  {32'hc142f0fe, 32'h414368f9} /* (21, 0, 6) {real, imag} */,
  {32'h42a00ea0, 32'h4080cdd4} /* (21, 0, 5) {real, imag} */,
  {32'hbe5d2e00, 32'h42835dc0} /* (21, 0, 4) {real, imag} */,
  {32'hc0b1fe24, 32'h40738e28} /* (21, 0, 3) {real, imag} */,
  {32'h4343e9a1, 32'h43a10a2c} /* (21, 0, 2) {real, imag} */,
  {32'hc4c4a908, 32'hc49a1a0d} /* (21, 0, 1) {real, imag} */,
  {32'hc514e715, 32'h00000000} /* (21, 0, 0) {real, imag} */,
  {32'hc51b5d9d, 32'h44a444ab} /* (20, 31, 31) {real, imag} */,
  {32'h440b9b13, 32'hc414fd1c} /* (20, 31, 30) {real, imag} */,
  {32'h426e8cc4, 32'hc1cb97e1} /* (20, 31, 29) {real, imag} */,
  {32'hc1c7bd5a, 32'h42a4b38c} /* (20, 31, 28) {real, imag} */,
  {32'h4270ad2f, 32'hc245485f} /* (20, 31, 27) {real, imag} */,
  {32'h3fc6d2f0, 32'hc0bbc3fa} /* (20, 31, 26) {real, imag} */,
  {32'hc21a6639, 32'h418c1a32} /* (20, 31, 25) {real, imag} */,
  {32'h418a1dde, 32'hc1e990b1} /* (20, 31, 24) {real, imag} */,
  {32'h404cb25f, 32'h3ee3c4f0} /* (20, 31, 23) {real, imag} */,
  {32'h41b470f4, 32'hc08a0fe3} /* (20, 31, 22) {real, imag} */,
  {32'hc08c7bdc, 32'hc1bdf1d7} /* (20, 31, 21) {real, imag} */,
  {32'hc10e1ace, 32'hc0d7b255} /* (20, 31, 20) {real, imag} */,
  {32'hc0884d52, 32'hc100f278} /* (20, 31, 19) {real, imag} */,
  {32'h3fc87e42, 32'hc158a142} /* (20, 31, 18) {real, imag} */,
  {32'h40fe1e08, 32'h408d20ab} /* (20, 31, 17) {real, imag} */,
  {32'hbec2fef8, 32'h40851dc0} /* (20, 31, 16) {real, imag} */,
  {32'hc0cdefa8, 32'h40b69388} /* (20, 31, 15) {real, imag} */,
  {32'h40a3aa64, 32'h417a716a} /* (20, 31, 14) {real, imag} */,
  {32'h3fd45798, 32'h3fadc170} /* (20, 31, 13) {real, imag} */,
  {32'hc0dddfab, 32'hc09de5f7} /* (20, 31, 12) {real, imag} */,
  {32'h412b1f1e, 32'hc08791f8} /* (20, 31, 11) {real, imag} */,
  {32'h40a23ff6, 32'h416f6e2e} /* (20, 31, 10) {real, imag} */,
  {32'h3e57de40, 32'h401a6e88} /* (20, 31, 9) {real, imag} */,
  {32'hc109d17b, 32'h41c2817c} /* (20, 31, 8) {real, imag} */,
  {32'hc1738d96, 32'hc18c1ed6} /* (20, 31, 7) {real, imag} */,
  {32'h41d5c249, 32'h41239f03} /* (20, 31, 6) {real, imag} */,
  {32'h4307550d, 32'hc1116d18} /* (20, 31, 5) {real, imag} */,
  {32'hc2934257, 32'h42b8bb86} /* (20, 31, 4) {real, imag} */,
  {32'hc1e0731e, 32'h41e59471} /* (20, 31, 3) {real, imag} */,
  {32'h43edbc2f, 32'hc19f65a7} /* (20, 31, 2) {real, imag} */,
  {32'hc4db3350, 32'hc3f56ab8} /* (20, 31, 1) {real, imag} */,
  {32'hc5057347, 32'h43a791d7} /* (20, 31, 0) {real, imag} */,
  {32'h44448726, 32'h42ee840f} /* (20, 30, 31) {real, imag} */,
  {32'hc3d0d7c1, 32'hc2ace058} /* (20, 30, 30) {real, imag} */,
  {32'h411c25e9, 32'h404395a6} /* (20, 30, 29) {real, imag} */,
  {32'h42ff0aeb, 32'hc0d426f8} /* (20, 30, 28) {real, imag} */,
  {32'hc2a03008, 32'h42b1db17} /* (20, 30, 27) {real, imag} */,
  {32'hc10ce8cd, 32'h415d3819} /* (20, 30, 26) {real, imag} */,
  {32'h411e8ae0, 32'hc0930a32} /* (20, 30, 25) {real, imag} */,
  {32'hc1d65898, 32'h421925f4} /* (20, 30, 24) {real, imag} */,
  {32'hbf8ac0e0, 32'hc12d17b2} /* (20, 30, 23) {real, imag} */,
  {32'h4157d422, 32'hc13ee3ac} /* (20, 30, 22) {real, imag} */,
  {32'h4126570a, 32'h412930d0} /* (20, 30, 21) {real, imag} */,
  {32'h3fd586a4, 32'hc02b00d8} /* (20, 30, 20) {real, imag} */,
  {32'hc104a2fa, 32'h40d52e63} /* (20, 30, 19) {real, imag} */,
  {32'hc16530b4, 32'h4008d8ac} /* (20, 30, 18) {real, imag} */,
  {32'h413014c1, 32'h40ed1a6a} /* (20, 30, 17) {real, imag} */,
  {32'hbf7aeb0e, 32'h40a2dc2a} /* (20, 30, 16) {real, imag} */,
  {32'hc0fb4408, 32'h414f9bee} /* (20, 30, 15) {real, imag} */,
  {32'hbef16b12, 32'h40bbe3d3} /* (20, 30, 14) {real, imag} */,
  {32'hc109cf30, 32'hbf4c6fc4} /* (20, 30, 13) {real, imag} */,
  {32'h40f9e3a8, 32'h40543d10} /* (20, 30, 12) {real, imag} */,
  {32'h3f491000, 32'hc168af79} /* (20, 30, 11) {real, imag} */,
  {32'hc18ec44e, 32'h4156af92} /* (20, 30, 10) {real, imag} */,
  {32'h3f9ca65c, 32'h40c8728b} /* (20, 30, 9) {real, imag} */,
  {32'hc1200584, 32'hc2243d57} /* (20, 30, 8) {real, imag} */,
  {32'h4181bcec, 32'h41af8576} /* (20, 30, 7) {real, imag} */,
  {32'h4194ceed, 32'hc1411471} /* (20, 30, 6) {real, imag} */,
  {32'hc26226ad, 32'hc0161cf0} /* (20, 30, 5) {real, imag} */,
  {32'h41aa320d, 32'h424b2e18} /* (20, 30, 4) {real, imag} */,
  {32'h42124ba8, 32'h416193bb} /* (20, 30, 3) {real, imag} */,
  {32'hc417a590, 32'hc357c390} /* (20, 30, 2) {real, imag} */,
  {32'h44a0d4b0, 32'hc0993e6e} /* (20, 30, 1) {real, imag} */,
  {32'h44275dce, 32'hc2ecb550} /* (20, 30, 0) {real, imag} */,
  {32'hc318e2c7, 32'h42a891b5} /* (20, 29, 31) {real, imag} */,
  {32'h41c8b5de, 32'hc309d2aa} /* (20, 29, 30) {real, imag} */,
  {32'h421f48b2, 32'hc188b819} /* (20, 29, 29) {real, imag} */,
  {32'h4218e171, 32'h41058c4c} /* (20, 29, 28) {real, imag} */,
  {32'hc1a14155, 32'h3f62f0e0} /* (20, 29, 27) {real, imag} */,
  {32'h3ebfbb60, 32'h411544ba} /* (20, 29, 26) {real, imag} */,
  {32'h419d71f9, 32'hbfdd5c38} /* (20, 29, 25) {real, imag} */,
  {32'hc101bb3a, 32'hc18aabef} /* (20, 29, 24) {real, imag} */,
  {32'hc17f68e8, 32'h40e5a600} /* (20, 29, 23) {real, imag} */,
  {32'h416c316a, 32'hc102bb29} /* (20, 29, 22) {real, imag} */,
  {32'hc03e104c, 32'hc08d39ee} /* (20, 29, 21) {real, imag} */,
  {32'h414e70ba, 32'hc044cb48} /* (20, 29, 20) {real, imag} */,
  {32'hc01e7d7e, 32'hc11596ec} /* (20, 29, 19) {real, imag} */,
  {32'h40c6d120, 32'h3f036050} /* (20, 29, 18) {real, imag} */,
  {32'hc10762ae, 32'hbef098e0} /* (20, 29, 17) {real, imag} */,
  {32'hbec7b3fa, 32'h402fec0c} /* (20, 29, 16) {real, imag} */,
  {32'hbf32d772, 32'h406fcf01} /* (20, 29, 15) {real, imag} */,
  {32'hc061520e, 32'hc036ab12} /* (20, 29, 14) {real, imag} */,
  {32'hc112c8d0, 32'hc0908d64} /* (20, 29, 13) {real, imag} */,
  {32'h40a34a6a, 32'hc077d575} /* (20, 29, 12) {real, imag} */,
  {32'hc0f01982, 32'hc0a2894e} /* (20, 29, 11) {real, imag} */,
  {32'hc03df5ce, 32'h40ac98f4} /* (20, 29, 10) {real, imag} */,
  {32'hbfeb2830, 32'h414616a7} /* (20, 29, 9) {real, imag} */,
  {32'hc0da3a72, 32'h40560d08} /* (20, 29, 8) {real, imag} */,
  {32'hc1c28a8f, 32'hc0bb0f46} /* (20, 29, 7) {real, imag} */,
  {32'hbf166be4, 32'h40709e5c} /* (20, 29, 6) {real, imag} */,
  {32'hc058f320, 32'h411bab82} /* (20, 29, 5) {real, imag} */,
  {32'hc1dd0ef2, 32'h4214668c} /* (20, 29, 4) {real, imag} */,
  {32'hc1a9dbc1, 32'h4087c5f6} /* (20, 29, 3) {real, imag} */,
  {32'hc286b455, 32'hc3049385} /* (20, 29, 2) {real, imag} */,
  {32'h42e8e9b9, 32'h42de163e} /* (20, 29, 1) {real, imag} */,
  {32'h412447d1, 32'hc174ecd2} /* (20, 29, 0) {real, imag} */,
  {32'hc3066ec0, 32'h42790c92} /* (20, 28, 31) {real, imag} */,
  {32'h430011c4, 32'hc2a10ec4} /* (20, 28, 30) {real, imag} */,
  {32'hc1d8ac38, 32'h422305c0} /* (20, 28, 29) {real, imag} */,
  {32'h400116ac, 32'h4189d6f4} /* (20, 28, 28) {real, imag} */,
  {32'h41bea895, 32'hc1e192d6} /* (20, 28, 27) {real, imag} */,
  {32'hc1857b17, 32'hc195999a} /* (20, 28, 26) {real, imag} */,
  {32'hc093965c, 32'h41e34184} /* (20, 28, 25) {real, imag} */,
  {32'h3ffb73e3, 32'hbe7df100} /* (20, 28, 24) {real, imag} */,
  {32'hbeffff20, 32'h412ed022} /* (20, 28, 23) {real, imag} */,
  {32'hc1038bb5, 32'h408a5a56} /* (20, 28, 22) {real, imag} */,
  {32'hc17686de, 32'hc0f8d113} /* (20, 28, 21) {real, imag} */,
  {32'hc117bc6a, 32'hc181bf96} /* (20, 28, 20) {real, imag} */,
  {32'h40e9202a, 32'h3e901850} /* (20, 28, 19) {real, imag} */,
  {32'hc080aefa, 32'hc1415543} /* (20, 28, 18) {real, imag} */,
  {32'hc061d383, 32'h411fb0e2} /* (20, 28, 17) {real, imag} */,
  {32'h40357c39, 32'hc0cb8f34} /* (20, 28, 16) {real, imag} */,
  {32'hc114ea90, 32'hc1422195} /* (20, 28, 15) {real, imag} */,
  {32'hc107f912, 32'hc0a17f4c} /* (20, 28, 14) {real, imag} */,
  {32'h4164f95c, 32'h41710963} /* (20, 28, 13) {real, imag} */,
  {32'hc09231e4, 32'hc0edc38c} /* (20, 28, 12) {real, imag} */,
  {32'h4145f0c8, 32'h41385300} /* (20, 28, 11) {real, imag} */,
  {32'h41172054, 32'h3fbe34d6} /* (20, 28, 10) {real, imag} */,
  {32'hc1071c90, 32'h40d9c3c8} /* (20, 28, 9) {real, imag} */,
  {32'h41ce0c7c, 32'h40b95d3c} /* (20, 28, 8) {real, imag} */,
  {32'h40df4006, 32'hc1740a7e} /* (20, 28, 7) {real, imag} */,
  {32'hc1d7da59, 32'h41e7de52} /* (20, 28, 6) {real, imag} */,
  {32'h41b765e3, 32'h41ce5344} /* (20, 28, 5) {real, imag} */,
  {32'hc1d5c348, 32'h3eea1da8} /* (20, 28, 4) {real, imag} */,
  {32'hc01be250, 32'hc093553a} /* (20, 28, 3) {real, imag} */,
  {32'h42815489, 32'hc28ed1b3} /* (20, 28, 2) {real, imag} */,
  {32'hc1fc09eb, 32'h4300e973} /* (20, 28, 1) {real, imag} */,
  {32'hc2868616, 32'h4095598b} /* (20, 28, 0) {real, imag} */,
  {32'h421a6ddc, 32'hc2b178a3} /* (20, 27, 31) {real, imag} */,
  {32'hc1e0b282, 32'h42499bde} /* (20, 27, 30) {real, imag} */,
  {32'h418625f8, 32'hc11b65bc} /* (20, 27, 29) {real, imag} */,
  {32'h41bd3304, 32'hc06b6e60} /* (20, 27, 28) {real, imag} */,
  {32'hc1255955, 32'h413c26ca} /* (20, 27, 27) {real, imag} */,
  {32'h41b4610c, 32'h4067c73b} /* (20, 27, 26) {real, imag} */,
  {32'h4010dc34, 32'hc1730297} /* (20, 27, 25) {real, imag} */,
  {32'h411aa1d9, 32'hc11c5f98} /* (20, 27, 24) {real, imag} */,
  {32'hc105d81a, 32'h418468f1} /* (20, 27, 23) {real, imag} */,
  {32'h4153f76e, 32'hc146893e} /* (20, 27, 22) {real, imag} */,
  {32'h4145ee58, 32'h41cfcdd4} /* (20, 27, 21) {real, imag} */,
  {32'hc08a4af9, 32'h418a0554} /* (20, 27, 20) {real, imag} */,
  {32'hc08c5f61, 32'h3fb36870} /* (20, 27, 19) {real, imag} */,
  {32'hc0990c06, 32'hc010121c} /* (20, 27, 18) {real, imag} */,
  {32'h4035c1a8, 32'hc01208f5} /* (20, 27, 17) {real, imag} */,
  {32'h4022dbc4, 32'hc0efe0ca} /* (20, 27, 16) {real, imag} */,
  {32'hc107e1d6, 32'hc052079c} /* (20, 27, 15) {real, imag} */,
  {32'hc09e455f, 32'hc0ad570c} /* (20, 27, 14) {real, imag} */,
  {32'hc11acfd9, 32'h414750d3} /* (20, 27, 13) {real, imag} */,
  {32'h40a519d0, 32'h3fb02335} /* (20, 27, 12) {real, imag} */,
  {32'h4081416a, 32'hc05805d9} /* (20, 27, 11) {real, imag} */,
  {32'hc203a9a4, 32'h3f9cbb0c} /* (20, 27, 10) {real, imag} */,
  {32'hc14aae46, 32'hc1079192} /* (20, 27, 9) {real, imag} */,
  {32'hc0f03c4d, 32'hc1cbfb54} /* (20, 27, 8) {real, imag} */,
  {32'hbfdba644, 32'hc139b508} /* (20, 27, 7) {real, imag} */,
  {32'hc0c5aa50, 32'h3f850c74} /* (20, 27, 6) {real, imag} */,
  {32'hc1a160f1, 32'h3fad75a8} /* (20, 27, 5) {real, imag} */,
  {32'hc03dee38, 32'hc0923b9c} /* (20, 27, 4) {real, imag} */,
  {32'h41c7ef15, 32'hc1d7e91f} /* (20, 27, 3) {real, imag} */,
  {32'hc2556600, 32'hc0bfd076} /* (20, 27, 2) {real, imag} */,
  {32'h42ba0310, 32'h40624920} /* (20, 27, 1) {real, imag} */,
  {32'h424aa5ed, 32'hc28a429f} /* (20, 27, 0) {real, imag} */,
  {32'hc1b6c592, 32'h3e610f00} /* (20, 26, 31) {real, imag} */,
  {32'h40e45a5f, 32'hc0e92969} /* (20, 26, 30) {real, imag} */,
  {32'h40910e23, 32'h41f4a99a} /* (20, 26, 29) {real, imag} */,
  {32'hc0ffce53, 32'hc17d8094} /* (20, 26, 28) {real, imag} */,
  {32'h40a565ee, 32'h40fb9868} /* (20, 26, 27) {real, imag} */,
  {32'h408559c4, 32'h41535b39} /* (20, 26, 26) {real, imag} */,
  {32'hc1d075bc, 32'hc17e7a82} /* (20, 26, 25) {real, imag} */,
  {32'hc033aaf6, 32'h3ff2ef68} /* (20, 26, 24) {real, imag} */,
  {32'hc102f89e, 32'hc16cf436} /* (20, 26, 23) {real, imag} */,
  {32'h3dff7b80, 32'hc0e3bbb7} /* (20, 26, 22) {real, imag} */,
  {32'h405634a1, 32'hbffde8e2} /* (20, 26, 21) {real, imag} */,
  {32'h4105b0c4, 32'h40a54d4b} /* (20, 26, 20) {real, imag} */,
  {32'h40cfc910, 32'h419489d4} /* (20, 26, 19) {real, imag} */,
  {32'hc135d137, 32'hc128f46a} /* (20, 26, 18) {real, imag} */,
  {32'h40ac34dc, 32'h4129451f} /* (20, 26, 17) {real, imag} */,
  {32'h3e8752e0, 32'h3f9f5c36} /* (20, 26, 16) {real, imag} */,
  {32'hc084114e, 32'h415e10e1} /* (20, 26, 15) {real, imag} */,
  {32'h4058208e, 32'hc0a98e76} /* (20, 26, 14) {real, imag} */,
  {32'hc10cc962, 32'h40fdca5c} /* (20, 26, 13) {real, imag} */,
  {32'h417412c6, 32'hc0bcb469} /* (20, 26, 12) {real, imag} */,
  {32'hc126caae, 32'h408cb0e0} /* (20, 26, 11) {real, imag} */,
  {32'hc09890a2, 32'h41bb9990} /* (20, 26, 10) {real, imag} */,
  {32'h413c6376, 32'hc191d0f9} /* (20, 26, 9) {real, imag} */,
  {32'hc195c302, 32'h4139b449} /* (20, 26, 8) {real, imag} */,
  {32'hc1583296, 32'h4128ae2c} /* (20, 26, 7) {real, imag} */,
  {32'h40ad2e0f, 32'h418fbd76} /* (20, 26, 6) {real, imag} */,
  {32'h3f580858, 32'h41153ec2} /* (20, 26, 5) {real, imag} */,
  {32'h414383ac, 32'hc121ed42} /* (20, 26, 4) {real, imag} */,
  {32'hc0dfb65a, 32'h3e081540} /* (20, 26, 3) {real, imag} */,
  {32'hc0162bd0, 32'h3f756dc8} /* (20, 26, 2) {real, imag} */,
  {32'hbff39f8c, 32'hc1191200} /* (20, 26, 1) {real, imag} */,
  {32'h4199724f, 32'h4065857e} /* (20, 26, 0) {real, imag} */,
  {32'h416d0924, 32'h419174d8} /* (20, 25, 31) {real, imag} */,
  {32'hc04a37b0, 32'hc0c4d278} /* (20, 25, 30) {real, imag} */,
  {32'h418dde7a, 32'hc0a23f08} /* (20, 25, 29) {real, imag} */,
  {32'h41ae3b3a, 32'hc1219f87} /* (20, 25, 28) {real, imag} */,
  {32'h3ffa5e7c, 32'hc16ab43b} /* (20, 25, 27) {real, imag} */,
  {32'h40c48faa, 32'h41948d34} /* (20, 25, 26) {real, imag} */,
  {32'hc1b7ba0b, 32'hc08fbeb4} /* (20, 25, 25) {real, imag} */,
  {32'hc11fde34, 32'hc0ebe86f} /* (20, 25, 24) {real, imag} */,
  {32'h41806bbd, 32'h40a6c641} /* (20, 25, 23) {real, imag} */,
  {32'h416bfdc6, 32'h411d07d0} /* (20, 25, 22) {real, imag} */,
  {32'hc14d1408, 32'hc10425f6} /* (20, 25, 21) {real, imag} */,
  {32'h41192869, 32'hc111330f} /* (20, 25, 20) {real, imag} */,
  {32'hc05e5b02, 32'h3fa6a740} /* (20, 25, 19) {real, imag} */,
  {32'hc124b591, 32'hc0a71608} /* (20, 25, 18) {real, imag} */,
  {32'hc07c8079, 32'hc125d4f3} /* (20, 25, 17) {real, imag} */,
  {32'h400ad124, 32'hc0a32f4a} /* (20, 25, 16) {real, imag} */,
  {32'h40aa63db, 32'hc0fd1d1a} /* (20, 25, 15) {real, imag} */,
  {32'h4091360c, 32'h4105fe47} /* (20, 25, 14) {real, imag} */,
  {32'hc0098602, 32'hc09bc936} /* (20, 25, 13) {real, imag} */,
  {32'hc1263f12, 32'hbf217af8} /* (20, 25, 12) {real, imag} */,
  {32'hc1611412, 32'hbe54ade0} /* (20, 25, 11) {real, imag} */,
  {32'h40b65848, 32'h4055844c} /* (20, 25, 10) {real, imag} */,
  {32'hbeba6850, 32'hc14da967} /* (20, 25, 9) {real, imag} */,
  {32'h418aa836, 32'hc115f140} /* (20, 25, 8) {real, imag} */,
  {32'h3f7fd1e0, 32'hc1c3b334} /* (20, 25, 7) {real, imag} */,
  {32'hbf8d60a7, 32'hc0499b02} /* (20, 25, 6) {real, imag} */,
  {32'hc12df262, 32'hc127e1a2} /* (20, 25, 5) {real, imag} */,
  {32'hc1530690, 32'h411aa057} /* (20, 25, 4) {real, imag} */,
  {32'h415274b2, 32'h4106fd42} /* (20, 25, 3) {real, imag} */,
  {32'hbf04b02c, 32'h3fab59c0} /* (20, 25, 2) {real, imag} */,
  {32'hc194538c, 32'h42047887} /* (20, 25, 1) {real, imag} */,
  {32'hc0eb5726, 32'h412c5a7c} /* (20, 25, 0) {real, imag} */,
  {32'h41b28eb0, 32'hc1bd2269} /* (20, 24, 31) {real, imag} */,
  {32'hc21bd865, 32'h41632e1e} /* (20, 24, 30) {real, imag} */,
  {32'hc1952b94, 32'hc0fefd92} /* (20, 24, 29) {real, imag} */,
  {32'h3fd9e370, 32'hc0a3b2f8} /* (20, 24, 28) {real, imag} */,
  {32'hc1ad4317, 32'h41a6517e} /* (20, 24, 27) {real, imag} */,
  {32'hbfdb9698, 32'hc0926f15} /* (20, 24, 26) {real, imag} */,
  {32'hc18fd401, 32'hc0c6e073} /* (20, 24, 25) {real, imag} */,
  {32'hc1a74173, 32'h3e890f20} /* (20, 24, 24) {real, imag} */,
  {32'hc1565319, 32'hc0c87fce} /* (20, 24, 23) {real, imag} */,
  {32'hc119c774, 32'hc1e02b54} /* (20, 24, 22) {real, imag} */,
  {32'h41037d76, 32'h3fcab458} /* (20, 24, 21) {real, imag} */,
  {32'hc03085c3, 32'h411250c0} /* (20, 24, 20) {real, imag} */,
  {32'h408b5016, 32'hc0ff4639} /* (20, 24, 19) {real, imag} */,
  {32'h3d9b65c0, 32'hc06aafba} /* (20, 24, 18) {real, imag} */,
  {32'hc112b41e, 32'hbf33b8e8} /* (20, 24, 17) {real, imag} */,
  {32'hc04a899b, 32'hc058e90e} /* (20, 24, 16) {real, imag} */,
  {32'hc0076cdd, 32'hbfbaf460} /* (20, 24, 15) {real, imag} */,
  {32'hc0510810, 32'hbe65fe24} /* (20, 24, 14) {real, imag} */,
  {32'h41708ddc, 32'hc046578a} /* (20, 24, 13) {real, imag} */,
  {32'hc1b66b68, 32'hc079e564} /* (20, 24, 12) {real, imag} */,
  {32'hc13c547c, 32'h4101a1d0} /* (20, 24, 11) {real, imag} */,
  {32'hc0150460, 32'hc1bd0c72} /* (20, 24, 10) {real, imag} */,
  {32'hbebf0c20, 32'h4157cc25} /* (20, 24, 9) {real, imag} */,
  {32'h40e8dfb5, 32'h4169b4fd} /* (20, 24, 8) {real, imag} */,
  {32'h401bd033, 32'h40f893ec} /* (20, 24, 7) {real, imag} */,
  {32'h40a41e9d, 32'h41434443} /* (20, 24, 6) {real, imag} */,
  {32'hc209ad76, 32'h4028b10b} /* (20, 24, 5) {real, imag} */,
  {32'h40baa97f, 32'hc0d51a45} /* (20, 24, 4) {real, imag} */,
  {32'h413db43e, 32'h415a03ea} /* (20, 24, 3) {real, imag} */,
  {32'hc0d2b89c, 32'h40c70603} /* (20, 24, 2) {real, imag} */,
  {32'h425576b6, 32'hc22a2995} /* (20, 24, 1) {real, imag} */,
  {32'h41996922, 32'h41093043} /* (20, 24, 0) {real, imag} */,
  {32'hc19e807e, 32'h41943045} /* (20, 23, 31) {real, imag} */,
  {32'hc1d9495c, 32'hc0f49d68} /* (20, 23, 30) {real, imag} */,
  {32'h412c8f42, 32'h4151eab5} /* (20, 23, 29) {real, imag} */,
  {32'hc057d4b7, 32'hc04998da} /* (20, 23, 28) {real, imag} */,
  {32'hc099fd8a, 32'hc085e56e} /* (20, 23, 27) {real, imag} */,
  {32'hbe8ec480, 32'hc123e896} /* (20, 23, 26) {real, imag} */,
  {32'h405f0ea6, 32'h402b067d} /* (20, 23, 25) {real, imag} */,
  {32'h412da96f, 32'hc144532d} /* (20, 23, 24) {real, imag} */,
  {32'h40c84159, 32'hc1babc62} /* (20, 23, 23) {real, imag} */,
  {32'hc0acc0fc, 32'h40ef74b1} /* (20, 23, 22) {real, imag} */,
  {32'h4180427d, 32'h409b8a6b} /* (20, 23, 21) {real, imag} */,
  {32'h4158f37f, 32'h40c27bc4} /* (20, 23, 20) {real, imag} */,
  {32'hc1122090, 32'h410dd33c} /* (20, 23, 19) {real, imag} */,
  {32'h3f1a3024, 32'h41961592} /* (20, 23, 18) {real, imag} */,
  {32'h4010260b, 32'hc0325d72} /* (20, 23, 17) {real, imag} */,
  {32'hc1577ccb, 32'h4052d33d} /* (20, 23, 16) {real, imag} */,
  {32'hbede0b84, 32'h40b8d622} /* (20, 23, 15) {real, imag} */,
  {32'hc154b4d6, 32'hc05db367} /* (20, 23, 14) {real, imag} */,
  {32'hc0d8d528, 32'hc10f312d} /* (20, 23, 13) {real, imag} */,
  {32'h4160ada0, 32'h412ec94c} /* (20, 23, 12) {real, imag} */,
  {32'hc08f57c5, 32'h4021eb32} /* (20, 23, 11) {real, imag} */,
  {32'hc1676224, 32'hc1ab7b67} /* (20, 23, 10) {real, imag} */,
  {32'hc027bc41, 32'h40195d68} /* (20, 23, 9) {real, imag} */,
  {32'h404b6008, 32'h3e978a40} /* (20, 23, 8) {real, imag} */,
  {32'h413878ec, 32'hc0c2edf5} /* (20, 23, 7) {real, imag} */,
  {32'hc143f1db, 32'hc1844168} /* (20, 23, 6) {real, imag} */,
  {32'hc0f68727, 32'hc0eb5e42} /* (20, 23, 5) {real, imag} */,
  {32'hc177257c, 32'h4041e740} /* (20, 23, 4) {real, imag} */,
  {32'h40d62968, 32'h40ed1324} /* (20, 23, 3) {real, imag} */,
  {32'hc0fed538, 32'h400b0454} /* (20, 23, 2) {real, imag} */,
  {32'h4172084f, 32'hc15d4f54} /* (20, 23, 1) {real, imag} */,
  {32'h418f1d57, 32'h40dfec7e} /* (20, 23, 0) {real, imag} */,
  {32'hc0779cbc, 32'hc117fe50} /* (20, 22, 31) {real, imag} */,
  {32'h3f614158, 32'hc0f97ec8} /* (20, 22, 30) {real, imag} */,
  {32'h4193f7bf, 32'hc1903d2e} /* (20, 22, 29) {real, imag} */,
  {32'hc01c89e8, 32'h41ceb1e9} /* (20, 22, 28) {real, imag} */,
  {32'hc1342ffc, 32'h40a6b3cb} /* (20, 22, 27) {real, imag} */,
  {32'hc0d481f9, 32'hbe81b310} /* (20, 22, 26) {real, imag} */,
  {32'h409aa905, 32'hbee29f20} /* (20, 22, 25) {real, imag} */,
  {32'h40bb37fe, 32'hc133f34c} /* (20, 22, 24) {real, imag} */,
  {32'hc1823fed, 32'hbf31f9d8} /* (20, 22, 23) {real, imag} */,
  {32'h40bd58e9, 32'hbfc77aa8} /* (20, 22, 22) {real, imag} */,
  {32'h419d25e4, 32'hc0a11c13} /* (20, 22, 21) {real, imag} */,
  {32'hc1ce18f8, 32'h3fc8fda4} /* (20, 22, 20) {real, imag} */,
  {32'hc03fa56e, 32'hc11b6206} /* (20, 22, 19) {real, imag} */,
  {32'h40997842, 32'hc158fe88} /* (20, 22, 18) {real, imag} */,
  {32'hbebd8420, 32'hc08ad5d5} /* (20, 22, 17) {real, imag} */,
  {32'h3fd564f0, 32'hc08ea540} /* (20, 22, 16) {real, imag} */,
  {32'hbf409cee, 32'h4127f827} /* (20, 22, 15) {real, imag} */,
  {32'hc0dcab4e, 32'hc0ea10af} /* (20, 22, 14) {real, imag} */,
  {32'h40964507, 32'hc0a7cb7c} /* (20, 22, 13) {real, imag} */,
  {32'h40906be9, 32'hc0a9207a} /* (20, 22, 12) {real, imag} */,
  {32'hbf361020, 32'hc1a73318} /* (20, 22, 11) {real, imag} */,
  {32'h4083457b, 32'h410925e2} /* (20, 22, 10) {real, imag} */,
  {32'hc08fce1e, 32'hc1acafbd} /* (20, 22, 9) {real, imag} */,
  {32'h41b23d2e, 32'h409741af} /* (20, 22, 8) {real, imag} */,
  {32'h40991872, 32'h403e4b28} /* (20, 22, 7) {real, imag} */,
  {32'hc16b6b10, 32'h412b28e6} /* (20, 22, 6) {real, imag} */,
  {32'h41393084, 32'h419b80df} /* (20, 22, 5) {real, imag} */,
  {32'hc11a9840, 32'h418a06da} /* (20, 22, 4) {real, imag} */,
  {32'hc196c596, 32'h3f1de3f4} /* (20, 22, 3) {real, imag} */,
  {32'hc12c9115, 32'hc1446e40} /* (20, 22, 2) {real, imag} */,
  {32'h4055ffce, 32'h3ef9ff20} /* (20, 22, 1) {real, imag} */,
  {32'h4101d95e, 32'h40f73817} /* (20, 22, 0) {real, imag} */,
  {32'h417fc744, 32'hc178a518} /* (20, 21, 31) {real, imag} */,
  {32'hc1837d69, 32'h4161abf5} /* (20, 21, 30) {real, imag} */,
  {32'hc0059f30, 32'h41673b40} /* (20, 21, 29) {real, imag} */,
  {32'hc149f244, 32'h401f8b90} /* (20, 21, 28) {real, imag} */,
  {32'hc12904f1, 32'h3ffffeb4} /* (20, 21, 27) {real, imag} */,
  {32'h409c2eb3, 32'h40d6ea06} /* (20, 21, 26) {real, imag} */,
  {32'h40820afa, 32'hc1a50bb4} /* (20, 21, 25) {real, imag} */,
  {32'hc1749eee, 32'h40b329c9} /* (20, 21, 24) {real, imag} */,
  {32'hc17a0ea9, 32'h419616c6} /* (20, 21, 23) {real, imag} */,
  {32'hc0eebb33, 32'h40541ac4} /* (20, 21, 22) {real, imag} */,
  {32'h40b694b9, 32'h40af870a} /* (20, 21, 21) {real, imag} */,
  {32'hc0644378, 32'h3f7e0750} /* (20, 21, 20) {real, imag} */,
  {32'hbde6ddb0, 32'hc0373a3c} /* (20, 21, 19) {real, imag} */,
  {32'hc0fd1eaa, 32'h41119cea} /* (20, 21, 18) {real, imag} */,
  {32'h41199130, 32'hbf9e4172} /* (20, 21, 17) {real, imag} */,
  {32'hc0720fc0, 32'hbf9c089a} /* (20, 21, 16) {real, imag} */,
  {32'hc1078307, 32'hc1a1241f} /* (20, 21, 15) {real, imag} */,
  {32'h414db8c8, 32'h3f0ee064} /* (20, 21, 14) {real, imag} */,
  {32'hbe256840, 32'h40e731a8} /* (20, 21, 13) {real, imag} */,
  {32'hc0933330, 32'h4068cdfa} /* (20, 21, 12) {real, imag} */,
  {32'h4002f1c0, 32'h413f757c} /* (20, 21, 11) {real, imag} */,
  {32'hc08e4b82, 32'h410d0ce1} /* (20, 21, 10) {real, imag} */,
  {32'h416a664f, 32'h415dc5cf} /* (20, 21, 9) {real, imag} */,
  {32'hc1217a93, 32'h403cc7a1} /* (20, 21, 8) {real, imag} */,
  {32'hc1b2b481, 32'h4035a5c0} /* (20, 21, 7) {real, imag} */,
  {32'hc1834b62, 32'h41625048} /* (20, 21, 6) {real, imag} */,
  {32'hbf37e13c, 32'hc01d215a} /* (20, 21, 5) {real, imag} */,
  {32'hc0d6eb4a, 32'h4196368c} /* (20, 21, 4) {real, imag} */,
  {32'hc0f3ffdc, 32'hbf943577} /* (20, 21, 3) {real, imag} */,
  {32'hbf6f5630, 32'hbee6d300} /* (20, 21, 2) {real, imag} */,
  {32'h418e061a, 32'hc1a63a66} /* (20, 21, 1) {real, imag} */,
  {32'h41673e20, 32'hc1416aeb} /* (20, 21, 0) {real, imag} */,
  {32'hc060d1f5, 32'hc0e199c4} /* (20, 20, 31) {real, imag} */,
  {32'h3f6bbc38, 32'hc1980fda} /* (20, 20, 30) {real, imag} */,
  {32'hc15aed6e, 32'h417bcee9} /* (20, 20, 29) {real, imag} */,
  {32'h3fe76ecb, 32'h41055e21} /* (20, 20, 28) {real, imag} */,
  {32'hc0d2581a, 32'h4090eca0} /* (20, 20, 27) {real, imag} */,
  {32'hc12425aa, 32'hc0922e48} /* (20, 20, 26) {real, imag} */,
  {32'h41cc3823, 32'h40d40565} /* (20, 20, 25) {real, imag} */,
  {32'h4112ea43, 32'hc1ad8baf} /* (20, 20, 24) {real, imag} */,
  {32'hc0dd6814, 32'hc118d146} /* (20, 20, 23) {real, imag} */,
  {32'hbfd9c428, 32'h41503b95} /* (20, 20, 22) {real, imag} */,
  {32'hc08fc422, 32'hbe55ab40} /* (20, 20, 21) {real, imag} */,
  {32'hc0a70450, 32'hc186fa40} /* (20, 20, 20) {real, imag} */,
  {32'h40df5084, 32'hc088f9f3} /* (20, 20, 19) {real, imag} */,
  {32'h40536183, 32'hbff25a7c} /* (20, 20, 18) {real, imag} */,
  {32'h40a996a4, 32'h40271970} /* (20, 20, 17) {real, imag} */,
  {32'hc05892e6, 32'h4127d392} /* (20, 20, 16) {real, imag} */,
  {32'h41364af0, 32'hc0603a0f} /* (20, 20, 15) {real, imag} */,
  {32'hbf1232d8, 32'h40415230} /* (20, 20, 14) {real, imag} */,
  {32'hbf60cc28, 32'hc12d475f} /* (20, 20, 13) {real, imag} */,
  {32'h4144a79c, 32'hc0f83d26} /* (20, 20, 12) {real, imag} */,
  {32'hc10dfcec, 32'h4050d9d5} /* (20, 20, 11) {real, imag} */,
  {32'hc12ec521, 32'h416f0b4c} /* (20, 20, 10) {real, imag} */,
  {32'h41287d1e, 32'hc15c99c8} /* (20, 20, 9) {real, imag} */,
  {32'h4131b9d6, 32'hc00d8ce5} /* (20, 20, 8) {real, imag} */,
  {32'h40ff4545, 32'hc1b1ac6d} /* (20, 20, 7) {real, imag} */,
  {32'h40ad4968, 32'hc11869a1} /* (20, 20, 6) {real, imag} */,
  {32'hc0d778ca, 32'hbf19d0d8} /* (20, 20, 5) {real, imag} */,
  {32'h41867514, 32'h403071f9} /* (20, 20, 4) {real, imag} */,
  {32'h407b1c18, 32'hc09d0008} /* (20, 20, 3) {real, imag} */,
  {32'hc1995553, 32'h40de776a} /* (20, 20, 2) {real, imag} */,
  {32'hc1113700, 32'hbffe883c} /* (20, 20, 1) {real, imag} */,
  {32'hbfffd774, 32'h40703531} /* (20, 20, 0) {real, imag} */,
  {32'hc104051e, 32'h3f1d0394} /* (20, 19, 31) {real, imag} */,
  {32'h41118f1f, 32'h4112943a} /* (20, 19, 30) {real, imag} */,
  {32'h3faae097, 32'hc11fc451} /* (20, 19, 29) {real, imag} */,
  {32'h408a9e38, 32'h4000fa7c} /* (20, 19, 28) {real, imag} */,
  {32'hc0e9cc58, 32'hc1560b12} /* (20, 19, 27) {real, imag} */,
  {32'h414f681e, 32'hbff7ceca} /* (20, 19, 26) {real, imag} */,
  {32'hc13905bb, 32'hc12872f5} /* (20, 19, 25) {real, imag} */,
  {32'h4128bb3c, 32'hc1008b09} /* (20, 19, 24) {real, imag} */,
  {32'h40d73663, 32'hc0a6e9d2} /* (20, 19, 23) {real, imag} */,
  {32'h40c7dbd1, 32'h40f312c6} /* (20, 19, 22) {real, imag} */,
  {32'hc1adbe52, 32'h4153e8b4} /* (20, 19, 21) {real, imag} */,
  {32'hc0e72b62, 32'h4125ff9d} /* (20, 19, 20) {real, imag} */,
  {32'hc0a6722d, 32'h3efc5280} /* (20, 19, 19) {real, imag} */,
  {32'h40fc8e6e, 32'h410cdacb} /* (20, 19, 18) {real, imag} */,
  {32'hc14f404a, 32'h410cef46} /* (20, 19, 17) {real, imag} */,
  {32'h412802fa, 32'h40fb73f8} /* (20, 19, 16) {real, imag} */,
  {32'h40d52468, 32'hbfefcfa9} /* (20, 19, 15) {real, imag} */,
  {32'hc0ed47b8, 32'h415ff0ac} /* (20, 19, 14) {real, imag} */,
  {32'h4096fd16, 32'h4072d863} /* (20, 19, 13) {real, imag} */,
  {32'hc1a4757d, 32'h41d13359} /* (20, 19, 12) {real, imag} */,
  {32'h40861072, 32'h41368904} /* (20, 19, 11) {real, imag} */,
  {32'hc135112e, 32'hc0692d3c} /* (20, 19, 10) {real, imag} */,
  {32'h4102b7da, 32'hc0b0d6cd} /* (20, 19, 9) {real, imag} */,
  {32'hc0db4e72, 32'hc1577998} /* (20, 19, 8) {real, imag} */,
  {32'h403fc495, 32'h4140f357} /* (20, 19, 7) {real, imag} */,
  {32'hc0a01a77, 32'hbf2f6ca2} /* (20, 19, 6) {real, imag} */,
  {32'h40a1eec7, 32'h41028af7} /* (20, 19, 5) {real, imag} */,
  {32'hc11d89e4, 32'h410052a6} /* (20, 19, 4) {real, imag} */,
  {32'h40ea6a76, 32'hc0829b20} /* (20, 19, 3) {real, imag} */,
  {32'hc08ce87f, 32'hc0b0bfaf} /* (20, 19, 2) {real, imag} */,
  {32'h3eb2c170, 32'h40df20b9} /* (20, 19, 1) {real, imag} */,
  {32'hc115487a, 32'h40faca54} /* (20, 19, 0) {real, imag} */,
  {32'hc16f8674, 32'hc1158c69} /* (20, 18, 31) {real, imag} */,
  {32'hbe172930, 32'h40b11de0} /* (20, 18, 30) {real, imag} */,
  {32'h40ec414d, 32'h3ed97940} /* (20, 18, 29) {real, imag} */,
  {32'hbf9aabc0, 32'h4174bf74} /* (20, 18, 28) {real, imag} */,
  {32'h41051322, 32'hc0ade898} /* (20, 18, 27) {real, imag} */,
  {32'hc10f1d4c, 32'h40d49906} /* (20, 18, 26) {real, imag} */,
  {32'h4101c1c3, 32'hc111b35f} /* (20, 18, 25) {real, imag} */,
  {32'h4125e9f1, 32'h3fa291c5} /* (20, 18, 24) {real, imag} */,
  {32'h3ffe3a64, 32'h41428b8c} /* (20, 18, 23) {real, imag} */,
  {32'h4184259a, 32'hc08f0c70} /* (20, 18, 22) {real, imag} */,
  {32'hc0198e22, 32'hc0d1ac39} /* (20, 18, 21) {real, imag} */,
  {32'h4024dfde, 32'hc13f9972} /* (20, 18, 20) {real, imag} */,
  {32'h404dc0ac, 32'hc0308fe2} /* (20, 18, 19) {real, imag} */,
  {32'h3f35f0ac, 32'h409cfb83} /* (20, 18, 18) {real, imag} */,
  {32'hbf056176, 32'hc0f8f2c6} /* (20, 18, 17) {real, imag} */,
  {32'h409fd6d5, 32'hc0ce4c56} /* (20, 18, 16) {real, imag} */,
  {32'h4128fe52, 32'h40a96904} /* (20, 18, 15) {real, imag} */,
  {32'h403ea7e0, 32'h4113e2b4} /* (20, 18, 14) {real, imag} */,
  {32'hc1903e28, 32'hc162024c} /* (20, 18, 13) {real, imag} */,
  {32'h41682fd3, 32'hc15c606e} /* (20, 18, 12) {real, imag} */,
  {32'h4087be00, 32'h404baf9a} /* (20, 18, 11) {real, imag} */,
  {32'hc122efe9, 32'h40716341} /* (20, 18, 10) {real, imag} */,
  {32'h4114f344, 32'hc0c206e0} /* (20, 18, 9) {real, imag} */,
  {32'hc10e90de, 32'h416bb45c} /* (20, 18, 8) {real, imag} */,
  {32'h40dc5094, 32'hbe524020} /* (20, 18, 7) {real, imag} */,
  {32'hbeff05d0, 32'h401374db} /* (20, 18, 6) {real, imag} */,
  {32'h3d623f00, 32'h401beff0} /* (20, 18, 5) {real, imag} */,
  {32'h414d78d5, 32'h409544ec} /* (20, 18, 4) {real, imag} */,
  {32'hbe11d4b4, 32'hbf99f54b} /* (20, 18, 3) {real, imag} */,
  {32'hc12ca460, 32'h3fa717a0} /* (20, 18, 2) {real, imag} */,
  {32'hbfa30144, 32'hc15afaef} /* (20, 18, 1) {real, imag} */,
  {32'hbdcec550, 32'hc1709d26} /* (20, 18, 0) {real, imag} */,
  {32'h40e40a98, 32'h4017ff4a} /* (20, 17, 31) {real, imag} */,
  {32'h414e845e, 32'h3ebe7f38} /* (20, 17, 30) {real, imag} */,
  {32'h400ee998, 32'h40e67586} /* (20, 17, 29) {real, imag} */,
  {32'h3fc8fd87, 32'hc0aa93e6} /* (20, 17, 28) {real, imag} */,
  {32'hbfd6296e, 32'hbec94e88} /* (20, 17, 27) {real, imag} */,
  {32'hc13e5cea, 32'h410ea8aa} /* (20, 17, 26) {real, imag} */,
  {32'hc0b386e2, 32'hbea441e0} /* (20, 17, 25) {real, imag} */,
  {32'h3f68d978, 32'hc1196046} /* (20, 17, 24) {real, imag} */,
  {32'hc064446e, 32'h3f78ea00} /* (20, 17, 23) {real, imag} */,
  {32'h40e2f4ee, 32'h3f0e7364} /* (20, 17, 22) {real, imag} */,
  {32'h40896802, 32'hc035da11} /* (20, 17, 21) {real, imag} */,
  {32'hc10846b9, 32'hc135d999} /* (20, 17, 20) {real, imag} */,
  {32'hbf41552c, 32'hc0a6d6a1} /* (20, 17, 19) {real, imag} */,
  {32'hbf536e50, 32'h40030168} /* (20, 17, 18) {real, imag} */,
  {32'hc0ec6d02, 32'h410511a4} /* (20, 17, 17) {real, imag} */,
  {32'hc00078b1, 32'h4104c500} /* (20, 17, 16) {real, imag} */,
  {32'hc147b25d, 32'hc08b29c1} /* (20, 17, 15) {real, imag} */,
  {32'hc151ea94, 32'h40ae1372} /* (20, 17, 14) {real, imag} */,
  {32'hc12f8a34, 32'h411253df} /* (20, 17, 13) {real, imag} */,
  {32'hc094c5a0, 32'hbf38d480} /* (20, 17, 12) {real, imag} */,
  {32'h411860da, 32'h4124e572} /* (20, 17, 11) {real, imag} */,
  {32'hc17fea06, 32'hc11f9b9f} /* (20, 17, 10) {real, imag} */,
  {32'hc104903e, 32'hc14417f3} /* (20, 17, 9) {real, imag} */,
  {32'hc124cfd0, 32'hc153f637} /* (20, 17, 8) {real, imag} */,
  {32'h3edd0950, 32'h40a66c38} /* (20, 17, 7) {real, imag} */,
  {32'hc0abfff4, 32'h4131c06c} /* (20, 17, 6) {real, imag} */,
  {32'hc03890be, 32'hbfda4717} /* (20, 17, 5) {real, imag} */,
  {32'hc110d1b0, 32'hc132e37f} /* (20, 17, 4) {real, imag} */,
  {32'hc1901476, 32'hc12c9f35} /* (20, 17, 3) {real, imag} */,
  {32'h4087cca0, 32'hbfe99f40} /* (20, 17, 2) {real, imag} */,
  {32'hc0653982, 32'h40dfd27f} /* (20, 17, 1) {real, imag} */,
  {32'h3fd790b8, 32'h4108c6cd} /* (20, 17, 0) {real, imag} */,
  {32'hc1493c4d, 32'h3f27cfda} /* (20, 16, 31) {real, imag} */,
  {32'h41003c0a, 32'hbe3dc870} /* (20, 16, 30) {real, imag} */,
  {32'h3de731a0, 32'hc0c1c9cf} /* (20, 16, 29) {real, imag} */,
  {32'hc0240029, 32'hc00fde18} /* (20, 16, 28) {real, imag} */,
  {32'h4011d80a, 32'hc057d4aa} /* (20, 16, 27) {real, imag} */,
  {32'h41021b04, 32'hc132cd78} /* (20, 16, 26) {real, imag} */,
  {32'hc10cb490, 32'h40a58422} /* (20, 16, 25) {real, imag} */,
  {32'hbfaa080c, 32'h3c69ab00} /* (20, 16, 24) {real, imag} */,
  {32'h3eec1548, 32'h407cfe5e} /* (20, 16, 23) {real, imag} */,
  {32'hc117ab87, 32'h408fb979} /* (20, 16, 22) {real, imag} */,
  {32'hc08afeea, 32'h41010373} /* (20, 16, 21) {real, imag} */,
  {32'h3f90979f, 32'hc1953760} /* (20, 16, 20) {real, imag} */,
  {32'h411b3d96, 32'h40c3294e} /* (20, 16, 19) {real, imag} */,
  {32'hc08ddc74, 32'h4108f533} /* (20, 16, 18) {real, imag} */,
  {32'h3ffff234, 32'hbff01c47} /* (20, 16, 17) {real, imag} */,
  {32'hc0766ca0, 32'h00000000} /* (20, 16, 16) {real, imag} */,
  {32'h3ffff234, 32'h3ff01c47} /* (20, 16, 15) {real, imag} */,
  {32'hc08ddc74, 32'hc108f533} /* (20, 16, 14) {real, imag} */,
  {32'h411b3d96, 32'hc0c3294e} /* (20, 16, 13) {real, imag} */,
  {32'h3f90979f, 32'h41953760} /* (20, 16, 12) {real, imag} */,
  {32'hc08afeea, 32'hc1010373} /* (20, 16, 11) {real, imag} */,
  {32'hc117ab87, 32'hc08fb979} /* (20, 16, 10) {real, imag} */,
  {32'h3eec1548, 32'hc07cfe5e} /* (20, 16, 9) {real, imag} */,
  {32'hbfaa080c, 32'hbc69ab00} /* (20, 16, 8) {real, imag} */,
  {32'hc10cb490, 32'hc0a58422} /* (20, 16, 7) {real, imag} */,
  {32'h41021b04, 32'h4132cd78} /* (20, 16, 6) {real, imag} */,
  {32'h4011d80a, 32'h4057d4aa} /* (20, 16, 5) {real, imag} */,
  {32'hc0240029, 32'h400fde18} /* (20, 16, 4) {real, imag} */,
  {32'h3de731a0, 32'h40c1c9cf} /* (20, 16, 3) {real, imag} */,
  {32'h41003c0a, 32'h3e3dc870} /* (20, 16, 2) {real, imag} */,
  {32'hc1493c4d, 32'hbf27cfda} /* (20, 16, 1) {real, imag} */,
  {32'h3fdad272, 32'h00000000} /* (20, 16, 0) {real, imag} */,
  {32'hc0653982, 32'hc0dfd27f} /* (20, 15, 31) {real, imag} */,
  {32'h4087cca0, 32'h3fe99f40} /* (20, 15, 30) {real, imag} */,
  {32'hc1901476, 32'h412c9f35} /* (20, 15, 29) {real, imag} */,
  {32'hc110d1b0, 32'h4132e37f} /* (20, 15, 28) {real, imag} */,
  {32'hc03890be, 32'h3fda4717} /* (20, 15, 27) {real, imag} */,
  {32'hc0abfff4, 32'hc131c06c} /* (20, 15, 26) {real, imag} */,
  {32'h3edd0950, 32'hc0a66c38} /* (20, 15, 25) {real, imag} */,
  {32'hc124cfd0, 32'h4153f637} /* (20, 15, 24) {real, imag} */,
  {32'hc104903e, 32'h414417f3} /* (20, 15, 23) {real, imag} */,
  {32'hc17fea06, 32'h411f9b9f} /* (20, 15, 22) {real, imag} */,
  {32'h411860da, 32'hc124e572} /* (20, 15, 21) {real, imag} */,
  {32'hc094c5a0, 32'h3f38d480} /* (20, 15, 20) {real, imag} */,
  {32'hc12f8a34, 32'hc11253df} /* (20, 15, 19) {real, imag} */,
  {32'hc151ea94, 32'hc0ae1372} /* (20, 15, 18) {real, imag} */,
  {32'hc147b25d, 32'h408b29c1} /* (20, 15, 17) {real, imag} */,
  {32'hc00078b1, 32'hc104c500} /* (20, 15, 16) {real, imag} */,
  {32'hc0ec6d02, 32'hc10511a4} /* (20, 15, 15) {real, imag} */,
  {32'hbf536e50, 32'hc0030168} /* (20, 15, 14) {real, imag} */,
  {32'hbf41552c, 32'h40a6d6a1} /* (20, 15, 13) {real, imag} */,
  {32'hc10846b9, 32'h4135d999} /* (20, 15, 12) {real, imag} */,
  {32'h40896802, 32'h4035da11} /* (20, 15, 11) {real, imag} */,
  {32'h40e2f4ee, 32'hbf0e7364} /* (20, 15, 10) {real, imag} */,
  {32'hc064446e, 32'hbf78ea00} /* (20, 15, 9) {real, imag} */,
  {32'h3f68d978, 32'h41196046} /* (20, 15, 8) {real, imag} */,
  {32'hc0b386e2, 32'h3ea441e0} /* (20, 15, 7) {real, imag} */,
  {32'hc13e5cea, 32'hc10ea8aa} /* (20, 15, 6) {real, imag} */,
  {32'hbfd6296e, 32'h3ec94e88} /* (20, 15, 5) {real, imag} */,
  {32'h3fc8fd87, 32'h40aa93e6} /* (20, 15, 4) {real, imag} */,
  {32'h400ee998, 32'hc0e67586} /* (20, 15, 3) {real, imag} */,
  {32'h414e845e, 32'hbebe7f38} /* (20, 15, 2) {real, imag} */,
  {32'h40e40a98, 32'hc017ff4a} /* (20, 15, 1) {real, imag} */,
  {32'h3fd790b8, 32'hc108c6cd} /* (20, 15, 0) {real, imag} */,
  {32'hbfa30144, 32'h415afaef} /* (20, 14, 31) {real, imag} */,
  {32'hc12ca460, 32'hbfa717a0} /* (20, 14, 30) {real, imag} */,
  {32'hbe11d4b4, 32'h3f99f54b} /* (20, 14, 29) {real, imag} */,
  {32'h414d78d5, 32'hc09544ec} /* (20, 14, 28) {real, imag} */,
  {32'h3d623f00, 32'hc01beff0} /* (20, 14, 27) {real, imag} */,
  {32'hbeff05d0, 32'hc01374db} /* (20, 14, 26) {real, imag} */,
  {32'h40dc5094, 32'h3e524020} /* (20, 14, 25) {real, imag} */,
  {32'hc10e90de, 32'hc16bb45c} /* (20, 14, 24) {real, imag} */,
  {32'h4114f344, 32'h40c206e0} /* (20, 14, 23) {real, imag} */,
  {32'hc122efe9, 32'hc0716341} /* (20, 14, 22) {real, imag} */,
  {32'h4087be00, 32'hc04baf9a} /* (20, 14, 21) {real, imag} */,
  {32'h41682fd3, 32'h415c606e} /* (20, 14, 20) {real, imag} */,
  {32'hc1903e28, 32'h4162024c} /* (20, 14, 19) {real, imag} */,
  {32'h403ea7e0, 32'hc113e2b4} /* (20, 14, 18) {real, imag} */,
  {32'h4128fe52, 32'hc0a96904} /* (20, 14, 17) {real, imag} */,
  {32'h409fd6d5, 32'h40ce4c56} /* (20, 14, 16) {real, imag} */,
  {32'hbf056176, 32'h40f8f2c6} /* (20, 14, 15) {real, imag} */,
  {32'h3f35f0ac, 32'hc09cfb83} /* (20, 14, 14) {real, imag} */,
  {32'h404dc0ac, 32'h40308fe2} /* (20, 14, 13) {real, imag} */,
  {32'h4024dfde, 32'h413f9972} /* (20, 14, 12) {real, imag} */,
  {32'hc0198e22, 32'h40d1ac39} /* (20, 14, 11) {real, imag} */,
  {32'h4184259a, 32'h408f0c70} /* (20, 14, 10) {real, imag} */,
  {32'h3ffe3a64, 32'hc1428b8c} /* (20, 14, 9) {real, imag} */,
  {32'h4125e9f1, 32'hbfa291c5} /* (20, 14, 8) {real, imag} */,
  {32'h4101c1c3, 32'h4111b35f} /* (20, 14, 7) {real, imag} */,
  {32'hc10f1d4c, 32'hc0d49906} /* (20, 14, 6) {real, imag} */,
  {32'h41051322, 32'h40ade898} /* (20, 14, 5) {real, imag} */,
  {32'hbf9aabc0, 32'hc174bf74} /* (20, 14, 4) {real, imag} */,
  {32'h40ec414d, 32'hbed97940} /* (20, 14, 3) {real, imag} */,
  {32'hbe172930, 32'hc0b11de0} /* (20, 14, 2) {real, imag} */,
  {32'hc16f8674, 32'h41158c69} /* (20, 14, 1) {real, imag} */,
  {32'hbdcec550, 32'h41709d26} /* (20, 14, 0) {real, imag} */,
  {32'h3eb2c170, 32'hc0df20b9} /* (20, 13, 31) {real, imag} */,
  {32'hc08ce87f, 32'h40b0bfaf} /* (20, 13, 30) {real, imag} */,
  {32'h40ea6a76, 32'h40829b20} /* (20, 13, 29) {real, imag} */,
  {32'hc11d89e4, 32'hc10052a6} /* (20, 13, 28) {real, imag} */,
  {32'h40a1eec7, 32'hc1028af7} /* (20, 13, 27) {real, imag} */,
  {32'hc0a01a77, 32'h3f2f6ca2} /* (20, 13, 26) {real, imag} */,
  {32'h403fc495, 32'hc140f357} /* (20, 13, 25) {real, imag} */,
  {32'hc0db4e72, 32'h41577998} /* (20, 13, 24) {real, imag} */,
  {32'h4102b7da, 32'h40b0d6cd} /* (20, 13, 23) {real, imag} */,
  {32'hc135112e, 32'h40692d3c} /* (20, 13, 22) {real, imag} */,
  {32'h40861072, 32'hc1368904} /* (20, 13, 21) {real, imag} */,
  {32'hc1a4757d, 32'hc1d13359} /* (20, 13, 20) {real, imag} */,
  {32'h4096fd16, 32'hc072d863} /* (20, 13, 19) {real, imag} */,
  {32'hc0ed47b8, 32'hc15ff0ac} /* (20, 13, 18) {real, imag} */,
  {32'h40d52468, 32'h3fefcfa9} /* (20, 13, 17) {real, imag} */,
  {32'h412802fa, 32'hc0fb73f8} /* (20, 13, 16) {real, imag} */,
  {32'hc14f404a, 32'hc10cef46} /* (20, 13, 15) {real, imag} */,
  {32'h40fc8e6e, 32'hc10cdacb} /* (20, 13, 14) {real, imag} */,
  {32'hc0a6722d, 32'hbefc5280} /* (20, 13, 13) {real, imag} */,
  {32'hc0e72b62, 32'hc125ff9d} /* (20, 13, 12) {real, imag} */,
  {32'hc1adbe52, 32'hc153e8b4} /* (20, 13, 11) {real, imag} */,
  {32'h40c7dbd1, 32'hc0f312c6} /* (20, 13, 10) {real, imag} */,
  {32'h40d73663, 32'h40a6e9d2} /* (20, 13, 9) {real, imag} */,
  {32'h4128bb3c, 32'h41008b09} /* (20, 13, 8) {real, imag} */,
  {32'hc13905bb, 32'h412872f5} /* (20, 13, 7) {real, imag} */,
  {32'h414f681e, 32'h3ff7ceca} /* (20, 13, 6) {real, imag} */,
  {32'hc0e9cc58, 32'h41560b12} /* (20, 13, 5) {real, imag} */,
  {32'h408a9e38, 32'hc000fa7c} /* (20, 13, 4) {real, imag} */,
  {32'h3faae097, 32'h411fc451} /* (20, 13, 3) {real, imag} */,
  {32'h41118f1f, 32'hc112943a} /* (20, 13, 2) {real, imag} */,
  {32'hc104051e, 32'hbf1d0394} /* (20, 13, 1) {real, imag} */,
  {32'hc115487a, 32'hc0faca54} /* (20, 13, 0) {real, imag} */,
  {32'hc1113700, 32'h3ffe883c} /* (20, 12, 31) {real, imag} */,
  {32'hc1995553, 32'hc0de776a} /* (20, 12, 30) {real, imag} */,
  {32'h407b1c18, 32'h409d0008} /* (20, 12, 29) {real, imag} */,
  {32'h41867514, 32'hc03071f9} /* (20, 12, 28) {real, imag} */,
  {32'hc0d778ca, 32'h3f19d0d8} /* (20, 12, 27) {real, imag} */,
  {32'h40ad4968, 32'h411869a1} /* (20, 12, 26) {real, imag} */,
  {32'h40ff4545, 32'h41b1ac6d} /* (20, 12, 25) {real, imag} */,
  {32'h4131b9d6, 32'h400d8ce5} /* (20, 12, 24) {real, imag} */,
  {32'h41287d1e, 32'h415c99c8} /* (20, 12, 23) {real, imag} */,
  {32'hc12ec521, 32'hc16f0b4c} /* (20, 12, 22) {real, imag} */,
  {32'hc10dfcec, 32'hc050d9d5} /* (20, 12, 21) {real, imag} */,
  {32'h4144a79c, 32'h40f83d26} /* (20, 12, 20) {real, imag} */,
  {32'hbf60cc28, 32'h412d475f} /* (20, 12, 19) {real, imag} */,
  {32'hbf1232d8, 32'hc0415230} /* (20, 12, 18) {real, imag} */,
  {32'h41364af0, 32'h40603a0f} /* (20, 12, 17) {real, imag} */,
  {32'hc05892e6, 32'hc127d392} /* (20, 12, 16) {real, imag} */,
  {32'h40a996a4, 32'hc0271970} /* (20, 12, 15) {real, imag} */,
  {32'h40536183, 32'h3ff25a7c} /* (20, 12, 14) {real, imag} */,
  {32'h40df5084, 32'h4088f9f3} /* (20, 12, 13) {real, imag} */,
  {32'hc0a70450, 32'h4186fa40} /* (20, 12, 12) {real, imag} */,
  {32'hc08fc422, 32'h3e55ab40} /* (20, 12, 11) {real, imag} */,
  {32'hbfd9c428, 32'hc1503b95} /* (20, 12, 10) {real, imag} */,
  {32'hc0dd6814, 32'h4118d146} /* (20, 12, 9) {real, imag} */,
  {32'h4112ea43, 32'h41ad8baf} /* (20, 12, 8) {real, imag} */,
  {32'h41cc3823, 32'hc0d40565} /* (20, 12, 7) {real, imag} */,
  {32'hc12425aa, 32'h40922e48} /* (20, 12, 6) {real, imag} */,
  {32'hc0d2581a, 32'hc090eca0} /* (20, 12, 5) {real, imag} */,
  {32'h3fe76ecb, 32'hc1055e21} /* (20, 12, 4) {real, imag} */,
  {32'hc15aed6e, 32'hc17bcee9} /* (20, 12, 3) {real, imag} */,
  {32'h3f6bbc38, 32'h41980fda} /* (20, 12, 2) {real, imag} */,
  {32'hc060d1f5, 32'h40e199c4} /* (20, 12, 1) {real, imag} */,
  {32'hbfffd774, 32'hc0703531} /* (20, 12, 0) {real, imag} */,
  {32'h418e061a, 32'h41a63a66} /* (20, 11, 31) {real, imag} */,
  {32'hbf6f5630, 32'h3ee6d300} /* (20, 11, 30) {real, imag} */,
  {32'hc0f3ffdc, 32'h3f943577} /* (20, 11, 29) {real, imag} */,
  {32'hc0d6eb4a, 32'hc196368c} /* (20, 11, 28) {real, imag} */,
  {32'hbf37e13c, 32'h401d215a} /* (20, 11, 27) {real, imag} */,
  {32'hc1834b62, 32'hc1625048} /* (20, 11, 26) {real, imag} */,
  {32'hc1b2b481, 32'hc035a5c0} /* (20, 11, 25) {real, imag} */,
  {32'hc1217a93, 32'hc03cc7a1} /* (20, 11, 24) {real, imag} */,
  {32'h416a664f, 32'hc15dc5cf} /* (20, 11, 23) {real, imag} */,
  {32'hc08e4b82, 32'hc10d0ce1} /* (20, 11, 22) {real, imag} */,
  {32'h4002f1c0, 32'hc13f757c} /* (20, 11, 21) {real, imag} */,
  {32'hc0933330, 32'hc068cdfa} /* (20, 11, 20) {real, imag} */,
  {32'hbe256840, 32'hc0e731a8} /* (20, 11, 19) {real, imag} */,
  {32'h414db8c8, 32'hbf0ee064} /* (20, 11, 18) {real, imag} */,
  {32'hc1078307, 32'h41a1241f} /* (20, 11, 17) {real, imag} */,
  {32'hc0720fc0, 32'h3f9c089a} /* (20, 11, 16) {real, imag} */,
  {32'h41199130, 32'h3f9e4172} /* (20, 11, 15) {real, imag} */,
  {32'hc0fd1eaa, 32'hc1119cea} /* (20, 11, 14) {real, imag} */,
  {32'hbde6ddb0, 32'h40373a3c} /* (20, 11, 13) {real, imag} */,
  {32'hc0644378, 32'hbf7e0750} /* (20, 11, 12) {real, imag} */,
  {32'h40b694b9, 32'hc0af870a} /* (20, 11, 11) {real, imag} */,
  {32'hc0eebb33, 32'hc0541ac4} /* (20, 11, 10) {real, imag} */,
  {32'hc17a0ea9, 32'hc19616c6} /* (20, 11, 9) {real, imag} */,
  {32'hc1749eee, 32'hc0b329c9} /* (20, 11, 8) {real, imag} */,
  {32'h40820afa, 32'h41a50bb4} /* (20, 11, 7) {real, imag} */,
  {32'h409c2eb3, 32'hc0d6ea06} /* (20, 11, 6) {real, imag} */,
  {32'hc12904f1, 32'hbffffeb4} /* (20, 11, 5) {real, imag} */,
  {32'hc149f244, 32'hc01f8b90} /* (20, 11, 4) {real, imag} */,
  {32'hc0059f30, 32'hc1673b40} /* (20, 11, 3) {real, imag} */,
  {32'hc1837d69, 32'hc161abf5} /* (20, 11, 2) {real, imag} */,
  {32'h417fc744, 32'h4178a518} /* (20, 11, 1) {real, imag} */,
  {32'h41673e20, 32'h41416aeb} /* (20, 11, 0) {real, imag} */,
  {32'h4055ffce, 32'hbef9ff20} /* (20, 10, 31) {real, imag} */,
  {32'hc12c9115, 32'h41446e40} /* (20, 10, 30) {real, imag} */,
  {32'hc196c596, 32'hbf1de3f4} /* (20, 10, 29) {real, imag} */,
  {32'hc11a9840, 32'hc18a06da} /* (20, 10, 28) {real, imag} */,
  {32'h41393084, 32'hc19b80df} /* (20, 10, 27) {real, imag} */,
  {32'hc16b6b10, 32'hc12b28e6} /* (20, 10, 26) {real, imag} */,
  {32'h40991872, 32'hc03e4b28} /* (20, 10, 25) {real, imag} */,
  {32'h41b23d2e, 32'hc09741af} /* (20, 10, 24) {real, imag} */,
  {32'hc08fce1e, 32'h41acafbd} /* (20, 10, 23) {real, imag} */,
  {32'h4083457b, 32'hc10925e2} /* (20, 10, 22) {real, imag} */,
  {32'hbf361020, 32'h41a73318} /* (20, 10, 21) {real, imag} */,
  {32'h40906be9, 32'h40a9207a} /* (20, 10, 20) {real, imag} */,
  {32'h40964507, 32'h40a7cb7c} /* (20, 10, 19) {real, imag} */,
  {32'hc0dcab4e, 32'h40ea10af} /* (20, 10, 18) {real, imag} */,
  {32'hbf409cee, 32'hc127f827} /* (20, 10, 17) {real, imag} */,
  {32'h3fd564f0, 32'h408ea540} /* (20, 10, 16) {real, imag} */,
  {32'hbebd8420, 32'h408ad5d5} /* (20, 10, 15) {real, imag} */,
  {32'h40997842, 32'h4158fe88} /* (20, 10, 14) {real, imag} */,
  {32'hc03fa56e, 32'h411b6206} /* (20, 10, 13) {real, imag} */,
  {32'hc1ce18f8, 32'hbfc8fda4} /* (20, 10, 12) {real, imag} */,
  {32'h419d25e4, 32'h40a11c13} /* (20, 10, 11) {real, imag} */,
  {32'h40bd58e9, 32'h3fc77aa8} /* (20, 10, 10) {real, imag} */,
  {32'hc1823fed, 32'h3f31f9d8} /* (20, 10, 9) {real, imag} */,
  {32'h40bb37fe, 32'h4133f34c} /* (20, 10, 8) {real, imag} */,
  {32'h409aa905, 32'h3ee29f20} /* (20, 10, 7) {real, imag} */,
  {32'hc0d481f9, 32'h3e81b310} /* (20, 10, 6) {real, imag} */,
  {32'hc1342ffc, 32'hc0a6b3cb} /* (20, 10, 5) {real, imag} */,
  {32'hc01c89e8, 32'hc1ceb1e9} /* (20, 10, 4) {real, imag} */,
  {32'h4193f7bf, 32'h41903d2e} /* (20, 10, 3) {real, imag} */,
  {32'h3f614158, 32'h40f97ec8} /* (20, 10, 2) {real, imag} */,
  {32'hc0779cbc, 32'h4117fe50} /* (20, 10, 1) {real, imag} */,
  {32'h4101d95e, 32'hc0f73817} /* (20, 10, 0) {real, imag} */,
  {32'h4172084f, 32'h415d4f54} /* (20, 9, 31) {real, imag} */,
  {32'hc0fed538, 32'hc00b0454} /* (20, 9, 30) {real, imag} */,
  {32'h40d62968, 32'hc0ed1324} /* (20, 9, 29) {real, imag} */,
  {32'hc177257c, 32'hc041e740} /* (20, 9, 28) {real, imag} */,
  {32'hc0f68727, 32'h40eb5e42} /* (20, 9, 27) {real, imag} */,
  {32'hc143f1db, 32'h41844168} /* (20, 9, 26) {real, imag} */,
  {32'h413878ec, 32'h40c2edf5} /* (20, 9, 25) {real, imag} */,
  {32'h404b6008, 32'hbe978a40} /* (20, 9, 24) {real, imag} */,
  {32'hc027bc41, 32'hc0195d68} /* (20, 9, 23) {real, imag} */,
  {32'hc1676224, 32'h41ab7b67} /* (20, 9, 22) {real, imag} */,
  {32'hc08f57c5, 32'hc021eb32} /* (20, 9, 21) {real, imag} */,
  {32'h4160ada0, 32'hc12ec94c} /* (20, 9, 20) {real, imag} */,
  {32'hc0d8d528, 32'h410f312d} /* (20, 9, 19) {real, imag} */,
  {32'hc154b4d6, 32'h405db367} /* (20, 9, 18) {real, imag} */,
  {32'hbede0b84, 32'hc0b8d622} /* (20, 9, 17) {real, imag} */,
  {32'hc1577ccb, 32'hc052d33d} /* (20, 9, 16) {real, imag} */,
  {32'h4010260b, 32'h40325d72} /* (20, 9, 15) {real, imag} */,
  {32'h3f1a3024, 32'hc1961592} /* (20, 9, 14) {real, imag} */,
  {32'hc1122090, 32'hc10dd33c} /* (20, 9, 13) {real, imag} */,
  {32'h4158f37f, 32'hc0c27bc4} /* (20, 9, 12) {real, imag} */,
  {32'h4180427d, 32'hc09b8a6b} /* (20, 9, 11) {real, imag} */,
  {32'hc0acc0fc, 32'hc0ef74b1} /* (20, 9, 10) {real, imag} */,
  {32'h40c84159, 32'h41babc62} /* (20, 9, 9) {real, imag} */,
  {32'h412da96f, 32'h4144532d} /* (20, 9, 8) {real, imag} */,
  {32'h405f0ea6, 32'hc02b067d} /* (20, 9, 7) {real, imag} */,
  {32'hbe8ec480, 32'h4123e896} /* (20, 9, 6) {real, imag} */,
  {32'hc099fd8a, 32'h4085e56e} /* (20, 9, 5) {real, imag} */,
  {32'hc057d4b7, 32'h404998da} /* (20, 9, 4) {real, imag} */,
  {32'h412c8f42, 32'hc151eab5} /* (20, 9, 3) {real, imag} */,
  {32'hc1d9495c, 32'h40f49d68} /* (20, 9, 2) {real, imag} */,
  {32'hc19e807e, 32'hc1943045} /* (20, 9, 1) {real, imag} */,
  {32'h418f1d57, 32'hc0dfec7e} /* (20, 9, 0) {real, imag} */,
  {32'h425576b6, 32'h422a2995} /* (20, 8, 31) {real, imag} */,
  {32'hc0d2b89c, 32'hc0c70603} /* (20, 8, 30) {real, imag} */,
  {32'h413db43e, 32'hc15a03ea} /* (20, 8, 29) {real, imag} */,
  {32'h40baa97f, 32'h40d51a45} /* (20, 8, 28) {real, imag} */,
  {32'hc209ad76, 32'hc028b10b} /* (20, 8, 27) {real, imag} */,
  {32'h40a41e9d, 32'hc1434443} /* (20, 8, 26) {real, imag} */,
  {32'h401bd033, 32'hc0f893ec} /* (20, 8, 25) {real, imag} */,
  {32'h40e8dfb5, 32'hc169b4fd} /* (20, 8, 24) {real, imag} */,
  {32'hbebf0c20, 32'hc157cc25} /* (20, 8, 23) {real, imag} */,
  {32'hc0150460, 32'h41bd0c72} /* (20, 8, 22) {real, imag} */,
  {32'hc13c547c, 32'hc101a1d0} /* (20, 8, 21) {real, imag} */,
  {32'hc1b66b68, 32'h4079e564} /* (20, 8, 20) {real, imag} */,
  {32'h41708ddc, 32'h4046578a} /* (20, 8, 19) {real, imag} */,
  {32'hc0510810, 32'h3e65fe24} /* (20, 8, 18) {real, imag} */,
  {32'hc0076cdd, 32'h3fbaf460} /* (20, 8, 17) {real, imag} */,
  {32'hc04a899b, 32'h4058e90e} /* (20, 8, 16) {real, imag} */,
  {32'hc112b41e, 32'h3f33b8e8} /* (20, 8, 15) {real, imag} */,
  {32'h3d9b65c0, 32'h406aafba} /* (20, 8, 14) {real, imag} */,
  {32'h408b5016, 32'h40ff4639} /* (20, 8, 13) {real, imag} */,
  {32'hc03085c3, 32'hc11250c0} /* (20, 8, 12) {real, imag} */,
  {32'h41037d76, 32'hbfcab458} /* (20, 8, 11) {real, imag} */,
  {32'hc119c774, 32'h41e02b54} /* (20, 8, 10) {real, imag} */,
  {32'hc1565319, 32'h40c87fce} /* (20, 8, 9) {real, imag} */,
  {32'hc1a74173, 32'hbe890f20} /* (20, 8, 8) {real, imag} */,
  {32'hc18fd401, 32'h40c6e073} /* (20, 8, 7) {real, imag} */,
  {32'hbfdb9698, 32'h40926f15} /* (20, 8, 6) {real, imag} */,
  {32'hc1ad4317, 32'hc1a6517e} /* (20, 8, 5) {real, imag} */,
  {32'h3fd9e370, 32'h40a3b2f8} /* (20, 8, 4) {real, imag} */,
  {32'hc1952b94, 32'h40fefd92} /* (20, 8, 3) {real, imag} */,
  {32'hc21bd865, 32'hc1632e1e} /* (20, 8, 2) {real, imag} */,
  {32'h41b28eb0, 32'h41bd2269} /* (20, 8, 1) {real, imag} */,
  {32'h41996922, 32'hc1093043} /* (20, 8, 0) {real, imag} */,
  {32'hc194538c, 32'hc2047887} /* (20, 7, 31) {real, imag} */,
  {32'hbf04b02c, 32'hbfab59c0} /* (20, 7, 30) {real, imag} */,
  {32'h415274b2, 32'hc106fd42} /* (20, 7, 29) {real, imag} */,
  {32'hc1530690, 32'hc11aa057} /* (20, 7, 28) {real, imag} */,
  {32'hc12df262, 32'h4127e1a2} /* (20, 7, 27) {real, imag} */,
  {32'hbf8d60a7, 32'h40499b02} /* (20, 7, 26) {real, imag} */,
  {32'h3f7fd1e0, 32'h41c3b334} /* (20, 7, 25) {real, imag} */,
  {32'h418aa836, 32'h4115f140} /* (20, 7, 24) {real, imag} */,
  {32'hbeba6850, 32'h414da967} /* (20, 7, 23) {real, imag} */,
  {32'h40b65848, 32'hc055844c} /* (20, 7, 22) {real, imag} */,
  {32'hc1611412, 32'h3e54ade0} /* (20, 7, 21) {real, imag} */,
  {32'hc1263f12, 32'h3f217af8} /* (20, 7, 20) {real, imag} */,
  {32'hc0098602, 32'h409bc936} /* (20, 7, 19) {real, imag} */,
  {32'h4091360c, 32'hc105fe47} /* (20, 7, 18) {real, imag} */,
  {32'h40aa63db, 32'h40fd1d1a} /* (20, 7, 17) {real, imag} */,
  {32'h400ad124, 32'h40a32f4a} /* (20, 7, 16) {real, imag} */,
  {32'hc07c8079, 32'h4125d4f3} /* (20, 7, 15) {real, imag} */,
  {32'hc124b591, 32'h40a71608} /* (20, 7, 14) {real, imag} */,
  {32'hc05e5b02, 32'hbfa6a740} /* (20, 7, 13) {real, imag} */,
  {32'h41192869, 32'h4111330f} /* (20, 7, 12) {real, imag} */,
  {32'hc14d1408, 32'h410425f6} /* (20, 7, 11) {real, imag} */,
  {32'h416bfdc6, 32'hc11d07d0} /* (20, 7, 10) {real, imag} */,
  {32'h41806bbd, 32'hc0a6c641} /* (20, 7, 9) {real, imag} */,
  {32'hc11fde34, 32'h40ebe86f} /* (20, 7, 8) {real, imag} */,
  {32'hc1b7ba0b, 32'h408fbeb4} /* (20, 7, 7) {real, imag} */,
  {32'h40c48faa, 32'hc1948d34} /* (20, 7, 6) {real, imag} */,
  {32'h3ffa5e7c, 32'h416ab43b} /* (20, 7, 5) {real, imag} */,
  {32'h41ae3b3a, 32'h41219f87} /* (20, 7, 4) {real, imag} */,
  {32'h418dde7a, 32'h40a23f08} /* (20, 7, 3) {real, imag} */,
  {32'hc04a37b0, 32'h40c4d278} /* (20, 7, 2) {real, imag} */,
  {32'h416d0924, 32'hc19174d8} /* (20, 7, 1) {real, imag} */,
  {32'hc0eb5726, 32'hc12c5a7c} /* (20, 7, 0) {real, imag} */,
  {32'hbff39f8c, 32'h41191200} /* (20, 6, 31) {real, imag} */,
  {32'hc0162bd0, 32'hbf756dc8} /* (20, 6, 30) {real, imag} */,
  {32'hc0dfb65a, 32'hbe081540} /* (20, 6, 29) {real, imag} */,
  {32'h414383ac, 32'h4121ed42} /* (20, 6, 28) {real, imag} */,
  {32'h3f580858, 32'hc1153ec2} /* (20, 6, 27) {real, imag} */,
  {32'h40ad2e0f, 32'hc18fbd76} /* (20, 6, 26) {real, imag} */,
  {32'hc1583296, 32'hc128ae2c} /* (20, 6, 25) {real, imag} */,
  {32'hc195c302, 32'hc139b449} /* (20, 6, 24) {real, imag} */,
  {32'h413c6376, 32'h4191d0f9} /* (20, 6, 23) {real, imag} */,
  {32'hc09890a2, 32'hc1bb9990} /* (20, 6, 22) {real, imag} */,
  {32'hc126caae, 32'hc08cb0e0} /* (20, 6, 21) {real, imag} */,
  {32'h417412c6, 32'h40bcb469} /* (20, 6, 20) {real, imag} */,
  {32'hc10cc962, 32'hc0fdca5c} /* (20, 6, 19) {real, imag} */,
  {32'h4058208e, 32'h40a98e76} /* (20, 6, 18) {real, imag} */,
  {32'hc084114e, 32'hc15e10e1} /* (20, 6, 17) {real, imag} */,
  {32'h3e8752e0, 32'hbf9f5c36} /* (20, 6, 16) {real, imag} */,
  {32'h40ac34dc, 32'hc129451f} /* (20, 6, 15) {real, imag} */,
  {32'hc135d137, 32'h4128f46a} /* (20, 6, 14) {real, imag} */,
  {32'h40cfc910, 32'hc19489d4} /* (20, 6, 13) {real, imag} */,
  {32'h4105b0c4, 32'hc0a54d4b} /* (20, 6, 12) {real, imag} */,
  {32'h405634a1, 32'h3ffde8e2} /* (20, 6, 11) {real, imag} */,
  {32'h3dff7b80, 32'h40e3bbb7} /* (20, 6, 10) {real, imag} */,
  {32'hc102f89e, 32'h416cf436} /* (20, 6, 9) {real, imag} */,
  {32'hc033aaf6, 32'hbff2ef68} /* (20, 6, 8) {real, imag} */,
  {32'hc1d075bc, 32'h417e7a82} /* (20, 6, 7) {real, imag} */,
  {32'h408559c4, 32'hc1535b39} /* (20, 6, 6) {real, imag} */,
  {32'h40a565ee, 32'hc0fb9868} /* (20, 6, 5) {real, imag} */,
  {32'hc0ffce53, 32'h417d8094} /* (20, 6, 4) {real, imag} */,
  {32'h40910e23, 32'hc1f4a99a} /* (20, 6, 3) {real, imag} */,
  {32'h40e45a5f, 32'h40e92969} /* (20, 6, 2) {real, imag} */,
  {32'hc1b6c592, 32'hbe610f00} /* (20, 6, 1) {real, imag} */,
  {32'h4199724f, 32'hc065857e} /* (20, 6, 0) {real, imag} */,
  {32'h42ba0310, 32'hc0624920} /* (20, 5, 31) {real, imag} */,
  {32'hc2556600, 32'h40bfd076} /* (20, 5, 30) {real, imag} */,
  {32'h41c7ef15, 32'h41d7e91f} /* (20, 5, 29) {real, imag} */,
  {32'hc03dee38, 32'h40923b9c} /* (20, 5, 28) {real, imag} */,
  {32'hc1a160f1, 32'hbfad75a8} /* (20, 5, 27) {real, imag} */,
  {32'hc0c5aa50, 32'hbf850c74} /* (20, 5, 26) {real, imag} */,
  {32'hbfdba644, 32'h4139b508} /* (20, 5, 25) {real, imag} */,
  {32'hc0f03c4d, 32'h41cbfb54} /* (20, 5, 24) {real, imag} */,
  {32'hc14aae46, 32'h41079192} /* (20, 5, 23) {real, imag} */,
  {32'hc203a9a4, 32'hbf9cbb0c} /* (20, 5, 22) {real, imag} */,
  {32'h4081416a, 32'h405805d9} /* (20, 5, 21) {real, imag} */,
  {32'h40a519d0, 32'hbfb02335} /* (20, 5, 20) {real, imag} */,
  {32'hc11acfd9, 32'hc14750d3} /* (20, 5, 19) {real, imag} */,
  {32'hc09e455f, 32'h40ad570c} /* (20, 5, 18) {real, imag} */,
  {32'hc107e1d6, 32'h4052079c} /* (20, 5, 17) {real, imag} */,
  {32'h4022dbc4, 32'h40efe0ca} /* (20, 5, 16) {real, imag} */,
  {32'h4035c1a8, 32'h401208f5} /* (20, 5, 15) {real, imag} */,
  {32'hc0990c06, 32'h4010121c} /* (20, 5, 14) {real, imag} */,
  {32'hc08c5f61, 32'hbfb36870} /* (20, 5, 13) {real, imag} */,
  {32'hc08a4af9, 32'hc18a0554} /* (20, 5, 12) {real, imag} */,
  {32'h4145ee58, 32'hc1cfcdd4} /* (20, 5, 11) {real, imag} */,
  {32'h4153f76e, 32'h4146893e} /* (20, 5, 10) {real, imag} */,
  {32'hc105d81a, 32'hc18468f1} /* (20, 5, 9) {real, imag} */,
  {32'h411aa1d9, 32'h411c5f98} /* (20, 5, 8) {real, imag} */,
  {32'h4010dc34, 32'h41730297} /* (20, 5, 7) {real, imag} */,
  {32'h41b4610c, 32'hc067c73b} /* (20, 5, 6) {real, imag} */,
  {32'hc1255955, 32'hc13c26ca} /* (20, 5, 5) {real, imag} */,
  {32'h41bd3304, 32'h406b6e60} /* (20, 5, 4) {real, imag} */,
  {32'h418625f8, 32'h411b65bc} /* (20, 5, 3) {real, imag} */,
  {32'hc1e0b282, 32'hc2499bde} /* (20, 5, 2) {real, imag} */,
  {32'h421a6ddc, 32'h42b178a3} /* (20, 5, 1) {real, imag} */,
  {32'h424aa5ed, 32'h428a429f} /* (20, 5, 0) {real, imag} */,
  {32'hc1fc09eb, 32'hc300e973} /* (20, 4, 31) {real, imag} */,
  {32'h42815489, 32'h428ed1b3} /* (20, 4, 30) {real, imag} */,
  {32'hc01be250, 32'h4093553a} /* (20, 4, 29) {real, imag} */,
  {32'hc1d5c348, 32'hbeea1da8} /* (20, 4, 28) {real, imag} */,
  {32'h41b765e3, 32'hc1ce5344} /* (20, 4, 27) {real, imag} */,
  {32'hc1d7da59, 32'hc1e7de52} /* (20, 4, 26) {real, imag} */,
  {32'h40df4006, 32'h41740a7e} /* (20, 4, 25) {real, imag} */,
  {32'h41ce0c7c, 32'hc0b95d3c} /* (20, 4, 24) {real, imag} */,
  {32'hc1071c90, 32'hc0d9c3c8} /* (20, 4, 23) {real, imag} */,
  {32'h41172054, 32'hbfbe34d6} /* (20, 4, 22) {real, imag} */,
  {32'h4145f0c8, 32'hc1385300} /* (20, 4, 21) {real, imag} */,
  {32'hc09231e4, 32'h40edc38c} /* (20, 4, 20) {real, imag} */,
  {32'h4164f95c, 32'hc1710963} /* (20, 4, 19) {real, imag} */,
  {32'hc107f912, 32'h40a17f4c} /* (20, 4, 18) {real, imag} */,
  {32'hc114ea90, 32'h41422195} /* (20, 4, 17) {real, imag} */,
  {32'h40357c39, 32'h40cb8f34} /* (20, 4, 16) {real, imag} */,
  {32'hc061d383, 32'hc11fb0e2} /* (20, 4, 15) {real, imag} */,
  {32'hc080aefa, 32'h41415543} /* (20, 4, 14) {real, imag} */,
  {32'h40e9202a, 32'hbe901850} /* (20, 4, 13) {real, imag} */,
  {32'hc117bc6a, 32'h4181bf96} /* (20, 4, 12) {real, imag} */,
  {32'hc17686de, 32'h40f8d113} /* (20, 4, 11) {real, imag} */,
  {32'hc1038bb5, 32'hc08a5a56} /* (20, 4, 10) {real, imag} */,
  {32'hbeffff20, 32'hc12ed022} /* (20, 4, 9) {real, imag} */,
  {32'h3ffb73e3, 32'h3e7df100} /* (20, 4, 8) {real, imag} */,
  {32'hc093965c, 32'hc1e34184} /* (20, 4, 7) {real, imag} */,
  {32'hc1857b17, 32'h4195999a} /* (20, 4, 6) {real, imag} */,
  {32'h41bea895, 32'h41e192d6} /* (20, 4, 5) {real, imag} */,
  {32'h400116ac, 32'hc189d6f4} /* (20, 4, 4) {real, imag} */,
  {32'hc1d8ac38, 32'hc22305c0} /* (20, 4, 3) {real, imag} */,
  {32'h430011c4, 32'h42a10ec4} /* (20, 4, 2) {real, imag} */,
  {32'hc3066ec0, 32'hc2790c92} /* (20, 4, 1) {real, imag} */,
  {32'hc2868616, 32'hc095598b} /* (20, 4, 0) {real, imag} */,
  {32'h42e8e9b9, 32'hc2de163e} /* (20, 3, 31) {real, imag} */,
  {32'hc286b455, 32'h43049385} /* (20, 3, 30) {real, imag} */,
  {32'hc1a9dbc1, 32'hc087c5f6} /* (20, 3, 29) {real, imag} */,
  {32'hc1dd0ef2, 32'hc214668c} /* (20, 3, 28) {real, imag} */,
  {32'hc058f320, 32'hc11bab82} /* (20, 3, 27) {real, imag} */,
  {32'hbf166be4, 32'hc0709e5c} /* (20, 3, 26) {real, imag} */,
  {32'hc1c28a8f, 32'h40bb0f46} /* (20, 3, 25) {real, imag} */,
  {32'hc0da3a72, 32'hc0560d08} /* (20, 3, 24) {real, imag} */,
  {32'hbfeb2830, 32'hc14616a7} /* (20, 3, 23) {real, imag} */,
  {32'hc03df5ce, 32'hc0ac98f4} /* (20, 3, 22) {real, imag} */,
  {32'hc0f01982, 32'h40a2894e} /* (20, 3, 21) {real, imag} */,
  {32'h40a34a6a, 32'h4077d575} /* (20, 3, 20) {real, imag} */,
  {32'hc112c8d0, 32'h40908d64} /* (20, 3, 19) {real, imag} */,
  {32'hc061520e, 32'h4036ab12} /* (20, 3, 18) {real, imag} */,
  {32'hbf32d772, 32'hc06fcf01} /* (20, 3, 17) {real, imag} */,
  {32'hbec7b3fa, 32'hc02fec0c} /* (20, 3, 16) {real, imag} */,
  {32'hc10762ae, 32'h3ef098e0} /* (20, 3, 15) {real, imag} */,
  {32'h40c6d120, 32'hbf036050} /* (20, 3, 14) {real, imag} */,
  {32'hc01e7d7e, 32'h411596ec} /* (20, 3, 13) {real, imag} */,
  {32'h414e70ba, 32'h4044cb48} /* (20, 3, 12) {real, imag} */,
  {32'hc03e104c, 32'h408d39ee} /* (20, 3, 11) {real, imag} */,
  {32'h416c316a, 32'h4102bb29} /* (20, 3, 10) {real, imag} */,
  {32'hc17f68e8, 32'hc0e5a600} /* (20, 3, 9) {real, imag} */,
  {32'hc101bb3a, 32'h418aabef} /* (20, 3, 8) {real, imag} */,
  {32'h419d71f9, 32'h3fdd5c38} /* (20, 3, 7) {real, imag} */,
  {32'h3ebfbb60, 32'hc11544ba} /* (20, 3, 6) {real, imag} */,
  {32'hc1a14155, 32'hbf62f0e0} /* (20, 3, 5) {real, imag} */,
  {32'h4218e171, 32'hc1058c4c} /* (20, 3, 4) {real, imag} */,
  {32'h421f48b2, 32'h4188b819} /* (20, 3, 3) {real, imag} */,
  {32'h41c8b5de, 32'h4309d2aa} /* (20, 3, 2) {real, imag} */,
  {32'hc318e2c7, 32'hc2a891b5} /* (20, 3, 1) {real, imag} */,
  {32'h412447d1, 32'h4174ecd2} /* (20, 3, 0) {real, imag} */,
  {32'h44a0d4b0, 32'h40993e6e} /* (20, 2, 31) {real, imag} */,
  {32'hc417a590, 32'h4357c390} /* (20, 2, 30) {real, imag} */,
  {32'h42124ba8, 32'hc16193bb} /* (20, 2, 29) {real, imag} */,
  {32'h41aa320d, 32'hc24b2e18} /* (20, 2, 28) {real, imag} */,
  {32'hc26226ad, 32'h40161cf0} /* (20, 2, 27) {real, imag} */,
  {32'h4194ceed, 32'h41411471} /* (20, 2, 26) {real, imag} */,
  {32'h4181bcec, 32'hc1af8576} /* (20, 2, 25) {real, imag} */,
  {32'hc1200584, 32'h42243d57} /* (20, 2, 24) {real, imag} */,
  {32'h3f9ca65c, 32'hc0c8728b} /* (20, 2, 23) {real, imag} */,
  {32'hc18ec44e, 32'hc156af92} /* (20, 2, 22) {real, imag} */,
  {32'h3f491000, 32'h4168af79} /* (20, 2, 21) {real, imag} */,
  {32'h40f9e3a8, 32'hc0543d10} /* (20, 2, 20) {real, imag} */,
  {32'hc109cf30, 32'h3f4c6fc4} /* (20, 2, 19) {real, imag} */,
  {32'hbef16b12, 32'hc0bbe3d3} /* (20, 2, 18) {real, imag} */,
  {32'hc0fb4408, 32'hc14f9bee} /* (20, 2, 17) {real, imag} */,
  {32'hbf7aeb0e, 32'hc0a2dc2a} /* (20, 2, 16) {real, imag} */,
  {32'h413014c1, 32'hc0ed1a6a} /* (20, 2, 15) {real, imag} */,
  {32'hc16530b4, 32'hc008d8ac} /* (20, 2, 14) {real, imag} */,
  {32'hc104a2fa, 32'hc0d52e63} /* (20, 2, 13) {real, imag} */,
  {32'h3fd586a4, 32'h402b00d8} /* (20, 2, 12) {real, imag} */,
  {32'h4126570a, 32'hc12930d0} /* (20, 2, 11) {real, imag} */,
  {32'h4157d422, 32'h413ee3ac} /* (20, 2, 10) {real, imag} */,
  {32'hbf8ac0e0, 32'h412d17b2} /* (20, 2, 9) {real, imag} */,
  {32'hc1d65898, 32'hc21925f4} /* (20, 2, 8) {real, imag} */,
  {32'h411e8ae0, 32'h40930a32} /* (20, 2, 7) {real, imag} */,
  {32'hc10ce8cd, 32'hc15d3819} /* (20, 2, 6) {real, imag} */,
  {32'hc2a03008, 32'hc2b1db17} /* (20, 2, 5) {real, imag} */,
  {32'h42ff0aeb, 32'h40d426f8} /* (20, 2, 4) {real, imag} */,
  {32'h411c25e9, 32'hc04395a6} /* (20, 2, 3) {real, imag} */,
  {32'hc3d0d7c1, 32'h42ace058} /* (20, 2, 2) {real, imag} */,
  {32'h44448726, 32'hc2ee840f} /* (20, 2, 1) {real, imag} */,
  {32'h44275dce, 32'h42ecb550} /* (20, 2, 0) {real, imag} */,
  {32'hc4db3350, 32'h43f56ab8} /* (20, 1, 31) {real, imag} */,
  {32'h43edbc2f, 32'h419f65a7} /* (20, 1, 30) {real, imag} */,
  {32'hc1e0731e, 32'hc1e59471} /* (20, 1, 29) {real, imag} */,
  {32'hc2934257, 32'hc2b8bb86} /* (20, 1, 28) {real, imag} */,
  {32'h4307550d, 32'h41116d18} /* (20, 1, 27) {real, imag} */,
  {32'h41d5c249, 32'hc1239f03} /* (20, 1, 26) {real, imag} */,
  {32'hc1738d96, 32'h418c1ed6} /* (20, 1, 25) {real, imag} */,
  {32'hc109d17b, 32'hc1c2817c} /* (20, 1, 24) {real, imag} */,
  {32'h3e57de40, 32'hc01a6e88} /* (20, 1, 23) {real, imag} */,
  {32'h40a23ff6, 32'hc16f6e2e} /* (20, 1, 22) {real, imag} */,
  {32'h412b1f1e, 32'h408791f8} /* (20, 1, 21) {real, imag} */,
  {32'hc0dddfab, 32'h409de5f7} /* (20, 1, 20) {real, imag} */,
  {32'h3fd45798, 32'hbfadc170} /* (20, 1, 19) {real, imag} */,
  {32'h40a3aa64, 32'hc17a716a} /* (20, 1, 18) {real, imag} */,
  {32'hc0cdefa8, 32'hc0b69388} /* (20, 1, 17) {real, imag} */,
  {32'hbec2fef8, 32'hc0851dc0} /* (20, 1, 16) {real, imag} */,
  {32'h40fe1e08, 32'hc08d20ab} /* (20, 1, 15) {real, imag} */,
  {32'h3fc87e42, 32'h4158a142} /* (20, 1, 14) {real, imag} */,
  {32'hc0884d52, 32'h4100f278} /* (20, 1, 13) {real, imag} */,
  {32'hc10e1ace, 32'h40d7b255} /* (20, 1, 12) {real, imag} */,
  {32'hc08c7bdc, 32'h41bdf1d7} /* (20, 1, 11) {real, imag} */,
  {32'h41b470f4, 32'h408a0fe3} /* (20, 1, 10) {real, imag} */,
  {32'h404cb25f, 32'hbee3c4f0} /* (20, 1, 9) {real, imag} */,
  {32'h418a1dde, 32'h41e990b1} /* (20, 1, 8) {real, imag} */,
  {32'hc21a6639, 32'hc18c1a32} /* (20, 1, 7) {real, imag} */,
  {32'h3fc6d2f0, 32'h40bbc3fa} /* (20, 1, 6) {real, imag} */,
  {32'h4270ad2f, 32'h4245485f} /* (20, 1, 5) {real, imag} */,
  {32'hc1c7bd5a, 32'hc2a4b38c} /* (20, 1, 4) {real, imag} */,
  {32'h426e8cc4, 32'h41cb97e1} /* (20, 1, 3) {real, imag} */,
  {32'h440b9b13, 32'h4414fd1c} /* (20, 1, 2) {real, imag} */,
  {32'hc51b5d9d, 32'hc4a444ab} /* (20, 1, 1) {real, imag} */,
  {32'hc5057347, 32'hc3a791d7} /* (20, 1, 0) {real, imag} */,
  {32'hc4c0efc0, 32'h44946c9f} /* (20, 0, 31) {real, imag} */,
  {32'h434cd765, 32'hc3a11e89} /* (20, 0, 30) {real, imag} */,
  {32'h413ec3b8, 32'hc1881810} /* (20, 0, 29) {real, imag} */,
  {32'hc106c05e, 32'hc2493621} /* (20, 0, 28) {real, imag} */,
  {32'h428202fd, 32'h419238cb} /* (20, 0, 27) {real, imag} */,
  {32'h3f3142a0, 32'hc1c40874} /* (20, 0, 26) {real, imag} */,
  {32'hbf0cb324, 32'h40c4b2b8} /* (20, 0, 25) {real, imag} */,
  {32'hc13dc6d5, 32'hc165ec6d} /* (20, 0, 24) {real, imag} */,
  {32'hc1029b1c, 32'h4199dd94} /* (20, 0, 23) {real, imag} */,
  {32'hc13d798e, 32'hc14a37b4} /* (20, 0, 22) {real, imag} */,
  {32'h4144a080, 32'h40b30d8c} /* (20, 0, 21) {real, imag} */,
  {32'h3e3d4480, 32'hc0fe0af6} /* (20, 0, 20) {real, imag} */,
  {32'hc08a194e, 32'hc112fc40} /* (20, 0, 19) {real, imag} */,
  {32'h40fae526, 32'h400c5816} /* (20, 0, 18) {real, imag} */,
  {32'hc022c801, 32'hc02f9340} /* (20, 0, 17) {real, imag} */,
  {32'hc0f23924, 32'h00000000} /* (20, 0, 16) {real, imag} */,
  {32'hc022c801, 32'h402f9340} /* (20, 0, 15) {real, imag} */,
  {32'h40fae526, 32'hc00c5816} /* (20, 0, 14) {real, imag} */,
  {32'hc08a194e, 32'h4112fc40} /* (20, 0, 13) {real, imag} */,
  {32'h3e3d4480, 32'h40fe0af6} /* (20, 0, 12) {real, imag} */,
  {32'h4144a080, 32'hc0b30d8c} /* (20, 0, 11) {real, imag} */,
  {32'hc13d798e, 32'h414a37b4} /* (20, 0, 10) {real, imag} */,
  {32'hc1029b1c, 32'hc199dd94} /* (20, 0, 9) {real, imag} */,
  {32'hc13dc6d5, 32'h4165ec6d} /* (20, 0, 8) {real, imag} */,
  {32'hbf0cb324, 32'hc0c4b2b8} /* (20, 0, 7) {real, imag} */,
  {32'h3f3142a0, 32'h41c40874} /* (20, 0, 6) {real, imag} */,
  {32'h428202fd, 32'hc19238cb} /* (20, 0, 5) {real, imag} */,
  {32'hc106c05e, 32'h42493621} /* (20, 0, 4) {real, imag} */,
  {32'h413ec3b8, 32'h41881810} /* (20, 0, 3) {real, imag} */,
  {32'h434cd765, 32'h43a11e89} /* (20, 0, 2) {real, imag} */,
  {32'hc4c0efc0, 32'hc4946c9f} /* (20, 0, 1) {real, imag} */,
  {32'hc50dc6b6, 32'h00000000} /* (20, 0, 0) {real, imag} */,
  {32'hc50d96c0, 32'h44926cb8} /* (19, 31, 31) {real, imag} */,
  {32'h440653f0, 32'hc4149d4d} /* (19, 31, 30) {real, imag} */,
  {32'h4227ab86, 32'h3efca780} /* (19, 31, 29) {real, imag} */,
  {32'hc25ac26a, 32'h42789b00} /* (19, 31, 28) {real, imag} */,
  {32'h425c707a, 32'hc2174044} /* (19, 31, 27) {real, imag} */,
  {32'h410db760, 32'hc039a8d8} /* (19, 31, 26) {real, imag} */,
  {32'hc17e6a95, 32'h409779ab} /* (19, 31, 25) {real, imag} */,
  {32'h41b8fbac, 32'hc1a399dc} /* (19, 31, 24) {real, imag} */,
  {32'hc1ea3b3f, 32'hbfba1744} /* (19, 31, 23) {real, imag} */,
  {32'h4187e204, 32'hbfa71c4a} /* (19, 31, 22) {real, imag} */,
  {32'h41c6c586, 32'hc15ba026} /* (19, 31, 21) {real, imag} */,
  {32'hc07a8334, 32'hc08d6764} /* (19, 31, 20) {real, imag} */,
  {32'hbfe172eb, 32'hc06be5f8} /* (19, 31, 19) {real, imag} */,
  {32'hc0899036, 32'hc14c92ce} /* (19, 31, 18) {real, imag} */,
  {32'h40c8eaea, 32'h3ffc2fa4} /* (19, 31, 17) {real, imag} */,
  {32'hc0552879, 32'h3c811980} /* (19, 31, 16) {real, imag} */,
  {32'hc0fe3945, 32'hbfaf1cfc} /* (19, 31, 15) {real, imag} */,
  {32'h4137e1e0, 32'h41b3eae0} /* (19, 31, 14) {real, imag} */,
  {32'h413263bc, 32'hbfeb920c} /* (19, 31, 13) {real, imag} */,
  {32'hbf9cf1f2, 32'hc11e022b} /* (19, 31, 12) {real, imag} */,
  {32'h412aef27, 32'h41c98c38} /* (19, 31, 11) {real, imag} */,
  {32'h40a7127e, 32'hc1295a08} /* (19, 31, 10) {real, imag} */,
  {32'h41cfccd1, 32'h40ea1754} /* (19, 31, 9) {real, imag} */,
  {32'h402c82e0, 32'h415e57fb} /* (19, 31, 8) {real, imag} */,
  {32'hc142ad45, 32'hc1f63974} /* (19, 31, 7) {real, imag} */,
  {32'h41e15250, 32'h4210711c} /* (19, 31, 6) {real, imag} */,
  {32'h42f8108b, 32'hc192529f} /* (19, 31, 5) {real, imag} */,
  {32'hc2989234, 32'h42996fae} /* (19, 31, 4) {real, imag} */,
  {32'hc1a1674d, 32'h422e63c3} /* (19, 31, 3) {real, imag} */,
  {32'h43d45f5f, 32'hc1a2f934} /* (19, 31, 2) {real, imag} */,
  {32'hc4c755b8, 32'hc3cef1e9} /* (19, 31, 1) {real, imag} */,
  {32'hc4f06f6a, 32'h439e44bc} /* (19, 31, 0) {real, imag} */,
  {32'h44341a12, 32'h430a4c11} /* (19, 30, 31) {real, imag} */,
  {32'hc3da912f, 32'hc2ef188a} /* (19, 30, 30) {real, imag} */,
  {32'h41946dcd, 32'hc1a50ed3} /* (19, 30, 29) {real, imag} */,
  {32'h42e8a60e, 32'h410d23c2} /* (19, 30, 28) {real, imag} */,
  {32'hc297ab95, 32'h42a2e8c7} /* (19, 30, 27) {real, imag} */,
  {32'h4102c26a, 32'h4039af58} /* (19, 30, 26) {real, imag} */,
  {32'h40ecdc44, 32'h413b3f66} /* (19, 30, 25) {real, imag} */,
  {32'hc0c86bd4, 32'h4244d424} /* (19, 30, 24) {real, imag} */,
  {32'h410f7533, 32'hc12b22eb} /* (19, 30, 23) {real, imag} */,
  {32'hbfe6ad3e, 32'hc10125ef} /* (19, 30, 22) {real, imag} */,
  {32'hc153d6a8, 32'h41ce17d4} /* (19, 30, 21) {real, imag} */,
  {32'hc134704e, 32'hbf7e7e2c} /* (19, 30, 20) {real, imag} */,
  {32'h3f938489, 32'hc13d4e69} /* (19, 30, 19) {real, imag} */,
  {32'h40614566, 32'h40b25b9e} /* (19, 30, 18) {real, imag} */,
  {32'h3fb426c4, 32'hbf96e272} /* (19, 30, 17) {real, imag} */,
  {32'h4110cbfe, 32'hbf5516bc} /* (19, 30, 16) {real, imag} */,
  {32'h3eccef60, 32'h413b548b} /* (19, 30, 15) {real, imag} */,
  {32'h40dbca44, 32'hbf73fe7c} /* (19, 30, 14) {real, imag} */,
  {32'hc11aa231, 32'hbff1d848} /* (19, 30, 13) {real, imag} */,
  {32'h414f24ed, 32'h411fc726} /* (19, 30, 12) {real, imag} */,
  {32'hc1bcb7f9, 32'hc1d04bce} /* (19, 30, 11) {real, imag} */,
  {32'h3f739674, 32'h410c3be0} /* (19, 30, 10) {real, imag} */,
  {32'hc124df02, 32'h4193f618} /* (19, 30, 9) {real, imag} */,
  {32'hc04e87c0, 32'hc1e6da45} /* (19, 30, 8) {real, imag} */,
  {32'h41543815, 32'h42131c38} /* (19, 30, 7) {real, imag} */,
  {32'hc107fc44, 32'hc175a83e} /* (19, 30, 6) {real, imag} */,
  {32'hc21d8382, 32'hc11546e2} /* (19, 30, 5) {real, imag} */,
  {32'h429139d3, 32'h42a5bd74} /* (19, 30, 4) {real, imag} */,
  {32'h4264ebc4, 32'hc11d3bea} /* (19, 30, 3) {real, imag} */,
  {32'hc4200bf6, 32'hc31783a5} /* (19, 30, 2) {real, imag} */,
  {32'h44983966, 32'h41ee873e} /* (19, 30, 1) {real, imag} */,
  {32'h4422870c, 32'hc2d27fe6} /* (19, 30, 0) {real, imag} */,
  {32'hc2f87158, 32'h42ffa6a3} /* (19, 29, 31) {real, imag} */,
  {32'h4290e6d0, 32'hc3044652} /* (19, 29, 30) {real, imag} */,
  {32'h421b4812, 32'h40bd9077} /* (19, 29, 29) {real, imag} */,
  {32'h41f03abd, 32'hc101f997} /* (19, 29, 28) {real, imag} */,
  {32'hc166997b, 32'hbf0d14a0} /* (19, 29, 27) {real, imag} */,
  {32'h41432411, 32'h3fa2c94e} /* (19, 29, 26) {real, imag} */,
  {32'hc1810248, 32'h40a7daac} /* (19, 29, 25) {real, imag} */,
  {32'h3fbf5a18, 32'hc0d37ff8} /* (19, 29, 24) {real, imag} */,
  {32'h41035da2, 32'h419bf923} /* (19, 29, 23) {real, imag} */,
  {32'h411baff1, 32'hc1213286} /* (19, 29, 22) {real, imag} */,
  {32'hc174f227, 32'h4119d71f} /* (19, 29, 21) {real, imag} */,
  {32'h41a7e896, 32'h3f9a2588} /* (19, 29, 20) {real, imag} */,
  {32'hc0f7d880, 32'hc0fbecfa} /* (19, 29, 19) {real, imag} */,
  {32'hc1072c9f, 32'hc08b7e99} /* (19, 29, 18) {real, imag} */,
  {32'hc11571a9, 32'h4062bc94} /* (19, 29, 17) {real, imag} */,
  {32'hc02d0c22, 32'h409b5293} /* (19, 29, 16) {real, imag} */,
  {32'h404b5068, 32'hc0ac92ba} /* (19, 29, 15) {real, imag} */,
  {32'h41855cd6, 32'h40e3d4e6} /* (19, 29, 14) {real, imag} */,
  {32'hc11ef57c, 32'hc192f3f4} /* (19, 29, 13) {real, imag} */,
  {32'h411ec64f, 32'h415e5611} /* (19, 29, 12) {real, imag} */,
  {32'h4096ccc1, 32'h3fc63cec} /* (19, 29, 11) {real, imag} */,
  {32'hc20aa34c, 32'h41d4624a} /* (19, 29, 10) {real, imag} */,
  {32'h40b1fb91, 32'hc1789852} /* (19, 29, 9) {real, imag} */,
  {32'h4134f57c, 32'h3f876960} /* (19, 29, 8) {real, imag} */,
  {32'hc1b02a8e, 32'hc1f556e4} /* (19, 29, 7) {real, imag} */,
  {32'h41047d8a, 32'h40df2cc2} /* (19, 29, 6) {real, imag} */,
  {32'hc064b90c, 32'h41e43918} /* (19, 29, 5) {real, imag} */,
  {32'hc1b73c64, 32'h413a94d5} /* (19, 29, 4) {real, imag} */,
  {32'hc20c2a7e, 32'h40cbd342} /* (19, 29, 3) {real, imag} */,
  {32'hc28324c7, 32'hc340b34e} /* (19, 29, 2) {real, imag} */,
  {32'h42ed1552, 32'h42ff18b3} /* (19, 29, 1) {real, imag} */,
  {32'hc1aa1f56, 32'hc212d83e} /* (19, 29, 0) {real, imag} */,
  {32'hc320ee6b, 32'h4295057c} /* (19, 28, 31) {real, imag} */,
  {32'h42db3682, 32'hc28b5a9b} /* (19, 28, 30) {real, imag} */,
  {32'hc20c1000, 32'h41de74b8} /* (19, 28, 29) {real, imag} */,
  {32'h41542306, 32'h4155c51a} /* (19, 28, 28) {real, imag} */,
  {32'hbff0d1aa, 32'hc1eb6441} /* (19, 28, 27) {real, imag} */,
  {32'hc113bf44, 32'hc0e3ede6} /* (19, 28, 26) {real, imag} */,
  {32'hc0cd0f69, 32'h4052922e} /* (19, 28, 25) {real, imag} */,
  {32'h408a7c58, 32'hc1157658} /* (19, 28, 24) {real, imag} */,
  {32'h3e7547a0, 32'h413f77df} /* (19, 28, 23) {real, imag} */,
  {32'hc126453a, 32'hbdf4a2c0} /* (19, 28, 22) {real, imag} */,
  {32'hc1331862, 32'hc0fc18d2} /* (19, 28, 21) {real, imag} */,
  {32'hc041d393, 32'h3f41d5e0} /* (19, 28, 20) {real, imag} */,
  {32'h41834280, 32'hc060beea} /* (19, 28, 19) {real, imag} */,
  {32'hc0cb3354, 32'hc15ff7bb} /* (19, 28, 18) {real, imag} */,
  {32'hbf8834a0, 32'h416555d2} /* (19, 28, 17) {real, imag} */,
  {32'hc112da76, 32'hc01e26ea} /* (19, 28, 16) {real, imag} */,
  {32'h404861d9, 32'h40b32eac} /* (19, 28, 15) {real, imag} */,
  {32'hc12641d6, 32'h3ee7a820} /* (19, 28, 14) {real, imag} */,
  {32'hc0d72b2e, 32'h41d38093} /* (19, 28, 13) {real, imag} */,
  {32'hc1a636ce, 32'h4105043f} /* (19, 28, 12) {real, imag} */,
  {32'h419d38f9, 32'hc00b214c} /* (19, 28, 11) {real, imag} */,
  {32'hbf155dc4, 32'hbf86a6a4} /* (19, 28, 10) {real, imag} */,
  {32'h3f3b57d0, 32'hc077d6aa} /* (19, 28, 9) {real, imag} */,
  {32'h41849765, 32'h402f96cc} /* (19, 28, 8) {real, imag} */,
  {32'h4104e112, 32'hc1a4b92a} /* (19, 28, 7) {real, imag} */,
  {32'hc214282e, 32'h41983514} /* (19, 28, 6) {real, imag} */,
  {32'h424071c9, 32'h42006161} /* (19, 28, 5) {real, imag} */,
  {32'hc22cd552, 32'h413024ae} /* (19, 28, 4) {real, imag} */,
  {32'hc18e63e5, 32'h40484d1e} /* (19, 28, 3) {real, imag} */,
  {32'h426dd8de, 32'hc26ca51b} /* (19, 28, 2) {real, imag} */,
  {32'hc226b5c0, 32'h42eefdb4} /* (19, 28, 1) {real, imag} */,
  {32'hc2919f9c, 32'h41a71882} /* (19, 28, 0) {real, imag} */,
  {32'h42826cc2, 32'hc29ceb15} /* (19, 27, 31) {real, imag} */,
  {32'hc21a71aa, 32'h4218a112} /* (19, 27, 30) {real, imag} */,
  {32'h40c11250, 32'hc0b1ee9b} /* (19, 27, 29) {real, imag} */,
  {32'h41b8956d, 32'hc07ae328} /* (19, 27, 28) {real, imag} */,
  {32'hc22977b9, 32'hc0636958} /* (19, 27, 27) {real, imag} */,
  {32'hc09c9743, 32'h4196bcec} /* (19, 27, 26) {real, imag} */,
  {32'h422b8570, 32'h408b872d} /* (19, 27, 25) {real, imag} */,
  {32'hc108b8a8, 32'h40939f89} /* (19, 27, 24) {real, imag} */,
  {32'hc0b53ed3, 32'hc19724c7} /* (19, 27, 23) {real, imag} */,
  {32'hc10855ff, 32'hc16b3dec} /* (19, 27, 22) {real, imag} */,
  {32'h40c65874, 32'h40b832c1} /* (19, 27, 21) {real, imag} */,
  {32'h41587bc4, 32'hc0261588} /* (19, 27, 20) {real, imag} */,
  {32'hc04ea606, 32'hbde2ff40} /* (19, 27, 19) {real, imag} */,
  {32'hbc8b9d60, 32'h40a88c9d} /* (19, 27, 18) {real, imag} */,
  {32'h410973a9, 32'h40cc8f5a} /* (19, 27, 17) {real, imag} */,
  {32'hc080d748, 32'hc11e8bc0} /* (19, 27, 16) {real, imag} */,
  {32'h419c751e, 32'hc0929ff2} /* (19, 27, 15) {real, imag} */,
  {32'h4116676a, 32'hc1733c61} /* (19, 27, 14) {real, imag} */,
  {32'hc0c6b7c4, 32'hc048c093} /* (19, 27, 13) {real, imag} */,
  {32'hc0e5bf52, 32'h3f4f7918} /* (19, 27, 12) {real, imag} */,
  {32'hc0ce5fbe, 32'hc114128f} /* (19, 27, 11) {real, imag} */,
  {32'h3f835870, 32'hc18c5db3} /* (19, 27, 10) {real, imag} */,
  {32'hc08496bc, 32'hc15fb443} /* (19, 27, 9) {real, imag} */,
  {32'hc133fd88, 32'h41908162} /* (19, 27, 8) {real, imag} */,
  {32'h4110cc68, 32'hc11f1b4e} /* (19, 27, 7) {real, imag} */,
  {32'h40dcde93, 32'hc181fbd1} /* (19, 27, 6) {real, imag} */,
  {32'hc1545832, 32'h41161d6b} /* (19, 27, 5) {real, imag} */,
  {32'hc18d3c62, 32'h4091bd70} /* (19, 27, 4) {real, imag} */,
  {32'h418f7300, 32'hc2072e5d} /* (19, 27, 3) {real, imag} */,
  {32'hc245716e, 32'hc0db76a2} /* (19, 27, 2) {real, imag} */,
  {32'h42d27f34, 32'h413bb466} /* (19, 27, 1) {real, imag} */,
  {32'h42335bde, 32'hc226520e} /* (19, 27, 0) {real, imag} */,
  {32'hc120fc08, 32'h3f487840} /* (19, 26, 31) {real, imag} */,
  {32'hc1082679, 32'h414602e8} /* (19, 26, 30) {real, imag} */,
  {32'h41e09a3d, 32'h418d7073} /* (19, 26, 29) {real, imag} */,
  {32'hc0d9d17a, 32'hc1d601fe} /* (19, 26, 28) {real, imag} */,
  {32'hc172708c, 32'h4186b3a2} /* (19, 26, 27) {real, imag} */,
  {32'h41f4b90e, 32'h411c5459} /* (19, 26, 26) {real, imag} */,
  {32'h403f0f70, 32'hbf1d3310} /* (19, 26, 25) {real, imag} */,
  {32'hc1871d73, 32'hc1bf1688} /* (19, 26, 24) {real, imag} */,
  {32'hc2037597, 32'h409db860} /* (19, 26, 23) {real, imag} */,
  {32'h40f52360, 32'h4080ff0c} /* (19, 26, 22) {real, imag} */,
  {32'hbfe3397c, 32'hc092e3d2} /* (19, 26, 21) {real, imag} */,
  {32'h405af764, 32'hbdadd860} /* (19, 26, 20) {real, imag} */,
  {32'h4066c008, 32'hc0e76597} /* (19, 26, 19) {real, imag} */,
  {32'h40bcbb34, 32'h41d0c56e} /* (19, 26, 18) {real, imag} */,
  {32'hc0f08ee4, 32'hc15aa2e1} /* (19, 26, 17) {real, imag} */,
  {32'hbfe3e088, 32'hbfebac5c} /* (19, 26, 16) {real, imag} */,
  {32'hbfddfaa6, 32'h41088d8c} /* (19, 26, 15) {real, imag} */,
  {32'hc14dbfe4, 32'h418c723a} /* (19, 26, 14) {real, imag} */,
  {32'h409c54c4, 32'hbf86321c} /* (19, 26, 13) {real, imag} */,
  {32'hbfa4e76d, 32'h407b9ce0} /* (19, 26, 12) {real, imag} */,
  {32'hc0b8b133, 32'hc08e468d} /* (19, 26, 11) {real, imag} */,
  {32'h41dc604b, 32'hc0637ecc} /* (19, 26, 10) {real, imag} */,
  {32'hc084bc76, 32'hc14f28f3} /* (19, 26, 9) {real, imag} */,
  {32'hc17eb02c, 32'h41ad7a0a} /* (19, 26, 8) {real, imag} */,
  {32'hc0bd4447, 32'h40392c38} /* (19, 26, 7) {real, imag} */,
  {32'hc0691fc0, 32'h40f0c93a} /* (19, 26, 6) {real, imag} */,
  {32'hc1105c0d, 32'h410a4c61} /* (19, 26, 5) {real, imag} */,
  {32'h40eeb21e, 32'hc11007f9} /* (19, 26, 4) {real, imag} */,
  {32'hc1b5c7ff, 32'hc0de49fc} /* (19, 26, 3) {real, imag} */,
  {32'hc0f2464c, 32'hc022b9f8} /* (19, 26, 2) {real, imag} */,
  {32'hc0fefcf3, 32'h4024e73e} /* (19, 26, 1) {real, imag} */,
  {32'hc030cfbc, 32'hc148823a} /* (19, 26, 0) {real, imag} */,
  {32'hbc5e3400, 32'h41b658aa} /* (19, 25, 31) {real, imag} */,
  {32'h412e4796, 32'hbee9cb20} /* (19, 25, 30) {real, imag} */,
  {32'h41a4558c, 32'hc10649d7} /* (19, 25, 29) {real, imag} */,
  {32'h4109e116, 32'h4073b504} /* (19, 25, 28) {real, imag} */,
  {32'h402a3790, 32'h403a3962} /* (19, 25, 27) {real, imag} */,
  {32'h4123b9dc, 32'h4123cba5} /* (19, 25, 26) {real, imag} */,
  {32'hc1b63d96, 32'hc0278ce7} /* (19, 25, 25) {real, imag} */,
  {32'hbf90fbc0, 32'hc0eac096} /* (19, 25, 24) {real, imag} */,
  {32'h414accc2, 32'h40885364} /* (19, 25, 23) {real, imag} */,
  {32'hc12b28ca, 32'h409dd2fa} /* (19, 25, 22) {real, imag} */,
  {32'hc0b2ef24, 32'hc04ecb51} /* (19, 25, 21) {real, imag} */,
  {32'hbf82c1f8, 32'hbf60e020} /* (19, 25, 20) {real, imag} */,
  {32'h41457595, 32'hc0d9b97a} /* (19, 25, 19) {real, imag} */,
  {32'hc0128e4e, 32'h40c91ca8} /* (19, 25, 18) {real, imag} */,
  {32'hc03e668a, 32'hc130bbc6} /* (19, 25, 17) {real, imag} */,
  {32'h410e8ce2, 32'h41590632} /* (19, 25, 16) {real, imag} */,
  {32'h40d42d9d, 32'hc0e50067} /* (19, 25, 15) {real, imag} */,
  {32'h4036562e, 32'h40ee3590} /* (19, 25, 14) {real, imag} */,
  {32'h3e606de0, 32'h40c839f4} /* (19, 25, 13) {real, imag} */,
  {32'hc04d48fc, 32'hc111f961} /* (19, 25, 12) {real, imag} */,
  {32'h413b2285, 32'hbfb64ee0} /* (19, 25, 11) {real, imag} */,
  {32'h40901794, 32'hbf820dd0} /* (19, 25, 10) {real, imag} */,
  {32'h3e2c7680, 32'hc1e03940} /* (19, 25, 9) {real, imag} */,
  {32'h402d9db2, 32'h41285522} /* (19, 25, 8) {real, imag} */,
  {32'hc10228bb, 32'h405179f6} /* (19, 25, 7) {real, imag} */,
  {32'hc102eae2, 32'h41b10672} /* (19, 25, 6) {real, imag} */,
  {32'h41b74788, 32'hc173e716} /* (19, 25, 5) {real, imag} */,
  {32'h40b6d0a4, 32'hc113d83a} /* (19, 25, 4) {real, imag} */,
  {32'hc11991c4, 32'h3f421b70} /* (19, 25, 3) {real, imag} */,
  {32'h404fc71f, 32'hc024536e} /* (19, 25, 2) {real, imag} */,
  {32'hc1eb5acd, 32'h4181bdf6} /* (19, 25, 1) {real, imag} */,
  {32'hbefb8bd0, 32'h41dd3b81} /* (19, 25, 0) {real, imag} */,
  {32'h418e2444, 32'hc20255e2} /* (19, 24, 31) {real, imag} */,
  {32'hc2082f95, 32'h418ed096} /* (19, 24, 30) {real, imag} */,
  {32'hc0b83e9a, 32'hc10fd540} /* (19, 24, 29) {real, imag} */,
  {32'h418efa06, 32'hc13d6898} /* (19, 24, 28) {real, imag} */,
  {32'h4118e6b8, 32'h42032d05} /* (19, 24, 27) {real, imag} */,
  {32'h41bf9aa8, 32'h415a923e} /* (19, 24, 26) {real, imag} */,
  {32'hc162a11d, 32'hbdd03fa0} /* (19, 24, 25) {real, imag} */,
  {32'hc1bb8c2a, 32'hc120f158} /* (19, 24, 24) {real, imag} */,
  {32'hc083ac35, 32'h413711f3} /* (19, 24, 23) {real, imag} */,
  {32'hc0df8de7, 32'hc0710b67} /* (19, 24, 22) {real, imag} */,
  {32'h4129bcd4, 32'hc13fcb1f} /* (19, 24, 21) {real, imag} */,
  {32'h4090a3c2, 32'h40f96b16} /* (19, 24, 20) {real, imag} */,
  {32'h3fd997f6, 32'h41a4acdd} /* (19, 24, 19) {real, imag} */,
  {32'h40ca2d5c, 32'hc12a7baa} /* (19, 24, 18) {real, imag} */,
  {32'h412ad4a5, 32'h40c31586} /* (19, 24, 17) {real, imag} */,
  {32'h40dacbba, 32'hc082309a} /* (19, 24, 16) {real, imag} */,
  {32'hc158cf56, 32'h409c29ca} /* (19, 24, 15) {real, imag} */,
  {32'hbfc710e4, 32'hc09a98fe} /* (19, 24, 14) {real, imag} */,
  {32'hc109fffc, 32'h40c104a2} /* (19, 24, 13) {real, imag} */,
  {32'hc0991e02, 32'h3fd0f430} /* (19, 24, 12) {real, imag} */,
  {32'h40af03c4, 32'h40d2aca8} /* (19, 24, 11) {real, imag} */,
  {32'hc0f85b2e, 32'h401dc874} /* (19, 24, 10) {real, imag} */,
  {32'hc15ce57a, 32'hc15ac673} /* (19, 24, 9) {real, imag} */,
  {32'hc136478e, 32'h40e4f9fc} /* (19, 24, 8) {real, imag} */,
  {32'h40de8cba, 32'hc0312ed8} /* (19, 24, 7) {real, imag} */,
  {32'hc160f108, 32'h409a4e03} /* (19, 24, 6) {real, imag} */,
  {32'hc192b746, 32'hc029de03} /* (19, 24, 5) {real, imag} */,
  {32'hc182e730, 32'hc1deaad3} /* (19, 24, 4) {real, imag} */,
  {32'h3e9d9940, 32'h41ad1e17} /* (19, 24, 3) {real, imag} */,
  {32'hc1b7d7d7, 32'hc1083db0} /* (19, 24, 2) {real, imag} */,
  {32'h420fd2ad, 32'hc200de7d} /* (19, 24, 1) {real, imag} */,
  {32'h41b75556, 32'hc185c36d} /* (19, 24, 0) {real, imag} */,
  {32'h3fa2150c, 32'h41cf3c73} /* (19, 23, 31) {real, imag} */,
  {32'hc092671b, 32'hc1d122ed} /* (19, 23, 30) {real, imag} */,
  {32'hbf9e958a, 32'h41c63506} /* (19, 23, 29) {real, imag} */,
  {32'hc10bd3ae, 32'h410d9e7a} /* (19, 23, 28) {real, imag} */,
  {32'h40c07476, 32'hc1a4fd1e} /* (19, 23, 27) {real, imag} */,
  {32'hbdd83880, 32'hc040b226} /* (19, 23, 26) {real, imag} */,
  {32'h3fb3125a, 32'hc081d186} /* (19, 23, 25) {real, imag} */,
  {32'hc15f6d73, 32'h413da109} /* (19, 23, 24) {real, imag} */,
  {32'h3f8b709c, 32'hc10bd287} /* (19, 23, 23) {real, imag} */,
  {32'h414ed0bc, 32'h40c6b75f} /* (19, 23, 22) {real, imag} */,
  {32'h40c91ae4, 32'hc10cbd70} /* (19, 23, 21) {real, imag} */,
  {32'hc08bc99b, 32'h40db371a} /* (19, 23, 20) {real, imag} */,
  {32'hbfe9368b, 32'h415f3e17} /* (19, 23, 19) {real, imag} */,
  {32'h40984ac4, 32'hc18e23a2} /* (19, 23, 18) {real, imag} */,
  {32'h410b6aa5, 32'h4169c7f0} /* (19, 23, 17) {real, imag} */,
  {32'hbf1c2870, 32'hbcfbc500} /* (19, 23, 16) {real, imag} */,
  {32'h4194be80, 32'hbfdb16d0} /* (19, 23, 15) {real, imag} */,
  {32'h3f7a4d00, 32'h410b650e} /* (19, 23, 14) {real, imag} */,
  {32'h4102fed6, 32'hc1ac3f02} /* (19, 23, 13) {real, imag} */,
  {32'hc01b5161, 32'hc05f0c02} /* (19, 23, 12) {real, imag} */,
  {32'hc1497cb8, 32'hc03e4d07} /* (19, 23, 11) {real, imag} */,
  {32'h4105b66a, 32'hc0de516d} /* (19, 23, 10) {real, imag} */,
  {32'hc1353168, 32'hc0e8211a} /* (19, 23, 9) {real, imag} */,
  {32'h401b55b6, 32'hc11fa0e4} /* (19, 23, 8) {real, imag} */,
  {32'h40ca7542, 32'hc0aa42b0} /* (19, 23, 7) {real, imag} */,
  {32'hc1df7430, 32'h408778e4} /* (19, 23, 6) {real, imag} */,
  {32'h408beff2, 32'h41ee5048} /* (19, 23, 5) {real, imag} */,
  {32'hc12e0c91, 32'h4149a753} /* (19, 23, 4) {real, imag} */,
  {32'h41bacf45, 32'hc0d119b8} /* (19, 23, 3) {real, imag} */,
  {32'hc17692ab, 32'hc22a495c} /* (19, 23, 2) {real, imag} */,
  {32'h4090293b, 32'hc18540ae} /* (19, 23, 1) {real, imag} */,
  {32'hbfa6ea9e, 32'h40117f98} /* (19, 23, 0) {real, imag} */,
  {32'hc113c848, 32'h418630c8} /* (19, 22, 31) {real, imag} */,
  {32'h41c464da, 32'hc148e6c6} /* (19, 22, 30) {real, imag} */,
  {32'hc169cde8, 32'hc0d72f88} /* (19, 22, 29) {real, imag} */,
  {32'hc1103e9c, 32'h40d88846} /* (19, 22, 28) {real, imag} */,
  {32'hc1621516, 32'hc0f4c836} /* (19, 22, 27) {real, imag} */,
  {32'hc1bbf721, 32'h41331880} /* (19, 22, 26) {real, imag} */,
  {32'hc14d1e7e, 32'h3f5c1a44} /* (19, 22, 25) {real, imag} */,
  {32'hc093a8c0, 32'hc1e31878} /* (19, 22, 24) {real, imag} */,
  {32'hc1b0ae04, 32'hc0e1269a} /* (19, 22, 23) {real, imag} */,
  {32'h3f932238, 32'h4096dc3c} /* (19, 22, 22) {real, imag} */,
  {32'h40dafb14, 32'h4106175c} /* (19, 22, 21) {real, imag} */,
  {32'hc16f9ab0, 32'hbffef1d2} /* (19, 22, 20) {real, imag} */,
  {32'h403a5e96, 32'h4088427f} /* (19, 22, 19) {real, imag} */,
  {32'h411c551c, 32'hc10002b2} /* (19, 22, 18) {real, imag} */,
  {32'hbf93924a, 32'h3d2e1100} /* (19, 22, 17) {real, imag} */,
  {32'hc1260e08, 32'h41adfa22} /* (19, 22, 16) {real, imag} */,
  {32'hc0eb27d0, 32'h41261bdd} /* (19, 22, 15) {real, imag} */,
  {32'h4108a17a, 32'hbfd410aa} /* (19, 22, 14) {real, imag} */,
  {32'h407042b0, 32'h4078cc50} /* (19, 22, 13) {real, imag} */,
  {32'h41202b04, 32'h40897b70} /* (19, 22, 12) {real, imag} */,
  {32'h3ffad38c, 32'hc1337604} /* (19, 22, 11) {real, imag} */,
  {32'hc0fdce1b, 32'hc0d1e272} /* (19, 22, 10) {real, imag} */,
  {32'h3ee24598, 32'h40ce695e} /* (19, 22, 9) {real, imag} */,
  {32'hc16fbf22, 32'hc1653d36} /* (19, 22, 8) {real, imag} */,
  {32'h419a9af9, 32'h417ff782} /* (19, 22, 7) {real, imag} */,
  {32'hc0f40fc9, 32'hc0d017c7} /* (19, 22, 6) {real, imag} */,
  {32'h40af24ce, 32'hbf765330} /* (19, 22, 5) {real, imag} */,
  {32'h4153451c, 32'hc1421426} /* (19, 22, 4) {real, imag} */,
  {32'hc15dab3e, 32'h40f96596} /* (19, 22, 3) {real, imag} */,
  {32'h406d9b02, 32'h41c5759b} /* (19, 22, 2) {real, imag} */,
  {32'h3fcb0c1e, 32'h4114554b} /* (19, 22, 1) {real, imag} */,
  {32'hc0d53874, 32'hbddc6040} /* (19, 22, 0) {real, imag} */,
  {32'h3ec5b620, 32'hc18eeb9d} /* (19, 21, 31) {real, imag} */,
  {32'h40d0a15e, 32'h4180ffda} /* (19, 21, 30) {real, imag} */,
  {32'hc115948f, 32'hbecb1660} /* (19, 21, 29) {real, imag} */,
  {32'h41085c22, 32'h415b53cd} /* (19, 21, 28) {real, imag} */,
  {32'hc0ab207c, 32'h40ca96d3} /* (19, 21, 27) {real, imag} */,
  {32'hc0405a93, 32'h4103153a} /* (19, 21, 26) {real, imag} */,
  {32'hc1781009, 32'hc11ebf7a} /* (19, 21, 25) {real, imag} */,
  {32'hc11934e6, 32'hc07375c9} /* (19, 21, 24) {real, imag} */,
  {32'hc0f8aba4, 32'h3f43a260} /* (19, 21, 23) {real, imag} */,
  {32'hc14f4687, 32'h410ae2ba} /* (19, 21, 22) {real, imag} */,
  {32'h409ea468, 32'h410b0e46} /* (19, 21, 21) {real, imag} */,
  {32'hc12c722d, 32'hc16bb1d0} /* (19, 21, 20) {real, imag} */,
  {32'h415f15b9, 32'h40c70dc6} /* (19, 21, 19) {real, imag} */,
  {32'hc124eb35, 32'hc0d9ae24} /* (19, 21, 18) {real, imag} */,
  {32'hc0fef14d, 32'hc0301e43} /* (19, 21, 17) {real, imag} */,
  {32'h40fba3b2, 32'h40bc76c0} /* (19, 21, 16) {real, imag} */,
  {32'h40022cc6, 32'hbf148f30} /* (19, 21, 15) {real, imag} */,
  {32'h411d989d, 32'h40fd79bb} /* (19, 21, 14) {real, imag} */,
  {32'h40a3408c, 32'h40ea76a5} /* (19, 21, 13) {real, imag} */,
  {32'h4042a75a, 32'h3fabf698} /* (19, 21, 12) {real, imag} */,
  {32'h417910c4, 32'hc1594d54} /* (19, 21, 11) {real, imag} */,
  {32'hc1154bfb, 32'hc153250b} /* (19, 21, 10) {real, imag} */,
  {32'h41018724, 32'hc058510e} /* (19, 21, 9) {real, imag} */,
  {32'hc1a92de6, 32'hc034740c} /* (19, 21, 8) {real, imag} */,
  {32'h4102406f, 32'h411c57a1} /* (19, 21, 7) {real, imag} */,
  {32'hc0e9b0ae, 32'h408ec48e} /* (19, 21, 6) {real, imag} */,
  {32'hc074f630, 32'hc12cb6a4} /* (19, 21, 5) {real, imag} */,
  {32'hc0886e32, 32'h412d8b2a} /* (19, 21, 4) {real, imag} */,
  {32'h41296676, 32'h400f6bca} /* (19, 21, 3) {real, imag} */,
  {32'hbffb843c, 32'h417d4829} /* (19, 21, 2) {real, imag} */,
  {32'h419c2b15, 32'h4000c507} /* (19, 21, 1) {real, imag} */,
  {32'h4202f94f, 32'hc143a0b4} /* (19, 21, 0) {real, imag} */,
  {32'h413f7ec1, 32'hc1235db8} /* (19, 20, 31) {real, imag} */,
  {32'hbf87ed54, 32'hc0a077ee} /* (19, 20, 30) {real, imag} */,
  {32'hc1029364, 32'h3b53a000} /* (19, 20, 29) {real, imag} */,
  {32'h4015eb6a, 32'h3ff2ab98} /* (19, 20, 28) {real, imag} */,
  {32'hc0b80d84, 32'hc12b46f3} /* (19, 20, 27) {real, imag} */,
  {32'hc0e25868, 32'h406f186a} /* (19, 20, 26) {real, imag} */,
  {32'hc10a6874, 32'h41261034} /* (19, 20, 25) {real, imag} */,
  {32'h418247a4, 32'h4113a01f} /* (19, 20, 24) {real, imag} */,
  {32'h41d7366f, 32'hc17d28d4} /* (19, 20, 23) {real, imag} */,
  {32'hc156247a, 32'hc1c70862} /* (19, 20, 22) {real, imag} */,
  {32'h410c9a4b, 32'hc0c95302} /* (19, 20, 21) {real, imag} */,
  {32'h3fdc6560, 32'h41871036} /* (19, 20, 20) {real, imag} */,
  {32'hc1aac912, 32'hbf0183b0} /* (19, 20, 19) {real, imag} */,
  {32'h4180672c, 32'hc003813c} /* (19, 20, 18) {real, imag} */,
  {32'h3fed7f40, 32'hc00e19b7} /* (19, 20, 17) {real, imag} */,
  {32'h410edefb, 32'h3e3cc500} /* (19, 20, 16) {real, imag} */,
  {32'h414c618e, 32'hc0cadde0} /* (19, 20, 15) {real, imag} */,
  {32'hc1808b60, 32'hc13a3ac0} /* (19, 20, 14) {real, imag} */,
  {32'hc09e240a, 32'h419e8a29} /* (19, 20, 13) {real, imag} */,
  {32'hc0888e42, 32'h4085edf6} /* (19, 20, 12) {real, imag} */,
  {32'hc1c77b87, 32'hc19dc757} /* (19, 20, 11) {real, imag} */,
  {32'hc0cc6f88, 32'hc0bda914} /* (19, 20, 10) {real, imag} */,
  {32'hbf8fdcf4, 32'h4117167d} /* (19, 20, 9) {real, imag} */,
  {32'hc0b92cf4, 32'hc0d46292} /* (19, 20, 8) {real, imag} */,
  {32'hc0c5851e, 32'h418e0760} /* (19, 20, 7) {real, imag} */,
  {32'h4199a17b, 32'hc1450c56} /* (19, 20, 6) {real, imag} */,
  {32'hc10fc47e, 32'hc0f0278f} /* (19, 20, 5) {real, imag} */,
  {32'hc194e264, 32'h4128cfbc} /* (19, 20, 4) {real, imag} */,
  {32'h40c5de43, 32'hc0bfcbcd} /* (19, 20, 3) {real, imag} */,
  {32'h4092902c, 32'h414c86b2} /* (19, 20, 2) {real, imag} */,
  {32'h40bcbe93, 32'h40e2f348} /* (19, 20, 1) {real, imag} */,
  {32'h41126f9b, 32'h3e0b3dc0} /* (19, 20, 0) {real, imag} */,
  {32'hc174069e, 32'h40576d11} /* (19, 19, 31) {real, imag} */,
  {32'hc0cd7ffc, 32'h40ef10de} /* (19, 19, 30) {real, imag} */,
  {32'h4169f39f, 32'hc0c1722a} /* (19, 19, 29) {real, imag} */,
  {32'hc1339fa4, 32'h4140c668} /* (19, 19, 28) {real, imag} */,
  {32'h4148ef50, 32'h41265b3f} /* (19, 19, 27) {real, imag} */,
  {32'h4199d886, 32'h3ed8c64e} /* (19, 19, 26) {real, imag} */,
  {32'hbff61604, 32'h40d213ca} /* (19, 19, 25) {real, imag} */,
  {32'h40e9bb28, 32'h4013d4eb} /* (19, 19, 24) {real, imag} */,
  {32'hc0760be2, 32'hc133f26b} /* (19, 19, 23) {real, imag} */,
  {32'h41a3fbe8, 32'h40e778da} /* (19, 19, 22) {real, imag} */,
  {32'hc029fcf6, 32'hc1f11246} /* (19, 19, 21) {real, imag} */,
  {32'h4157234c, 32'hc0e79836} /* (19, 19, 20) {real, imag} */,
  {32'hc136eeb0, 32'h41771af0} /* (19, 19, 19) {real, imag} */,
  {32'hc14705fc, 32'h41f5cff7} /* (19, 19, 18) {real, imag} */,
  {32'h4106cb08, 32'hc14e5517} /* (19, 19, 17) {real, imag} */,
  {32'h408f7d66, 32'hc006aa52} /* (19, 19, 16) {real, imag} */,
  {32'hc0eea98c, 32'h40b653ea} /* (19, 19, 15) {real, imag} */,
  {32'hbfff933f, 32'h41443bd1} /* (19, 19, 14) {real, imag} */,
  {32'h41101b56, 32'hc11aa538} /* (19, 19, 13) {real, imag} */,
  {32'hc07d495e, 32'h40e0e038} /* (19, 19, 12) {real, imag} */,
  {32'h40b1dbc8, 32'hc06da332} /* (19, 19, 11) {real, imag} */,
  {32'h40e6ecc3, 32'hc140c643} /* (19, 19, 10) {real, imag} */,
  {32'hc11551e1, 32'hbf97b210} /* (19, 19, 9) {real, imag} */,
  {32'hc1074d72, 32'h408ddad0} /* (19, 19, 8) {real, imag} */,
  {32'h40e14886, 32'hbfe561ac} /* (19, 19, 7) {real, imag} */,
  {32'hbfbf44ae, 32'hc10731d8} /* (19, 19, 6) {real, imag} */,
  {32'hc15d52f0, 32'hc0bfde90} /* (19, 19, 5) {real, imag} */,
  {32'hbebb3d08, 32'h41253688} /* (19, 19, 4) {real, imag} */,
  {32'hc1b069ae, 32'h416b45ca} /* (19, 19, 3) {real, imag} */,
  {32'hc0bf7f7d, 32'hc0d80e9a} /* (19, 19, 2) {real, imag} */,
  {32'h412c7cee, 32'hc045dff3} /* (19, 19, 1) {real, imag} */,
  {32'h409a0125, 32'h4003fafd} /* (19, 19, 0) {real, imag} */,
  {32'hc1357247, 32'hbfb04d28} /* (19, 18, 31) {real, imag} */,
  {32'h401843d8, 32'hbef34b48} /* (19, 18, 30) {real, imag} */,
  {32'hbfa3ae4b, 32'h3feed308} /* (19, 18, 29) {real, imag} */,
  {32'h40c8f3aa, 32'h404aa9fc} /* (19, 18, 28) {real, imag} */,
  {32'hc0ee3b2d, 32'h40d9e419} /* (19, 18, 27) {real, imag} */,
  {32'hc0daf0d6, 32'h4112f4e4} /* (19, 18, 26) {real, imag} */,
  {32'h41199d62, 32'h3fe6bb97} /* (19, 18, 25) {real, imag} */,
  {32'h406e1f74, 32'hc0abb1ab} /* (19, 18, 24) {real, imag} */,
  {32'hc1608d97, 32'hc02df0c3} /* (19, 18, 23) {real, imag} */,
  {32'h4116bcbe, 32'hc03c2b37} /* (19, 18, 22) {real, imag} */,
  {32'h3fe8795f, 32'h40d8fa54} /* (19, 18, 21) {real, imag} */,
  {32'h405e2570, 32'h408b5eeb} /* (19, 18, 20) {real, imag} */,
  {32'hc0813f30, 32'hc041b21f} /* (19, 18, 19) {real, imag} */,
  {32'h40cf743b, 32'h400d81b6} /* (19, 18, 18) {real, imag} */,
  {32'h410cbdbc, 32'hbfd4fcae} /* (19, 18, 17) {real, imag} */,
  {32'hc0f22b6a, 32'hc0f1c34c} /* (19, 18, 16) {real, imag} */,
  {32'hc0a7455c, 32'hc00d88f6} /* (19, 18, 15) {real, imag} */,
  {32'hc1325591, 32'h3fbff004} /* (19, 18, 14) {real, imag} */,
  {32'h40c212f8, 32'hc0e4065a} /* (19, 18, 13) {real, imag} */,
  {32'h409cb895, 32'hc1380ae4} /* (19, 18, 12) {real, imag} */,
  {32'h412856d8, 32'hbed3d1a0} /* (19, 18, 11) {real, imag} */,
  {32'h417521f8, 32'h41120d88} /* (19, 18, 10) {real, imag} */,
  {32'h41363802, 32'h40e430e2} /* (19, 18, 9) {real, imag} */,
  {32'h402f73e6, 32'hc09df35e} /* (19, 18, 8) {real, imag} */,
  {32'hc030162c, 32'hc09c3e66} /* (19, 18, 7) {real, imag} */,
  {32'h3f0fb6c8, 32'hc0a93c5b} /* (19, 18, 6) {real, imag} */,
  {32'h3ea5df38, 32'h3fa9d734} /* (19, 18, 5) {real, imag} */,
  {32'h40a6146e, 32'hc1989c20} /* (19, 18, 4) {real, imag} */,
  {32'hc030dc3a, 32'h40f54b02} /* (19, 18, 3) {real, imag} */,
  {32'hbdfd4c00, 32'h411573d5} /* (19, 18, 2) {real, imag} */,
  {32'h41449c92, 32'hc1a31b12} /* (19, 18, 1) {real, imag} */,
  {32'hc0e7542b, 32'hbf312158} /* (19, 18, 0) {real, imag} */,
  {32'h3fb064fa, 32'h40878794} /* (19, 17, 31) {real, imag} */,
  {32'h40278f08, 32'hc0973695} /* (19, 17, 30) {real, imag} */,
  {32'h3f81b110, 32'hbfde3349} /* (19, 17, 29) {real, imag} */,
  {32'h40abaa5a, 32'h40d1f4e8} /* (19, 17, 28) {real, imag} */,
  {32'h40c20878, 32'hc03998e2} /* (19, 17, 27) {real, imag} */,
  {32'h4161ea51, 32'h41957bf0} /* (19, 17, 26) {real, imag} */,
  {32'hbfbba038, 32'hc190edf4} /* (19, 17, 25) {real, imag} */,
  {32'h403ed2ff, 32'hc0944502} /* (19, 17, 24) {real, imag} */,
  {32'h40de79a4, 32'hbf7c9c0c} /* (19, 17, 23) {real, imag} */,
  {32'hbfb5f49c, 32'h415d87d8} /* (19, 17, 22) {real, imag} */,
  {32'h409b3052, 32'hc0a219ff} /* (19, 17, 21) {real, imag} */,
  {32'h400fd86c, 32'h40c25aef} /* (19, 17, 20) {real, imag} */,
  {32'hbfe423ac, 32'h3f818b88} /* (19, 17, 19) {real, imag} */,
  {32'hc0fe841e, 32'hc1635da4} /* (19, 17, 18) {real, imag} */,
  {32'h4095fe80, 32'hc1178ccc} /* (19, 17, 17) {real, imag} */,
  {32'h412f5a5c, 32'hc02c2f82} /* (19, 17, 16) {real, imag} */,
  {32'h403d99cc, 32'hc0bc8a48} /* (19, 17, 15) {real, imag} */,
  {32'h4109c8f8, 32'h3fdad057} /* (19, 17, 14) {real, imag} */,
  {32'h415bd79a, 32'h40ba56e6} /* (19, 17, 13) {real, imag} */,
  {32'hbf3bd7f2, 32'h401dddc4} /* (19, 17, 12) {real, imag} */,
  {32'h406c1814, 32'h40b50942} /* (19, 17, 11) {real, imag} */,
  {32'hc0a20322, 32'hc0ea4a74} /* (19, 17, 10) {real, imag} */,
  {32'hc108a09a, 32'hc0e832e6} /* (19, 17, 9) {real, imag} */,
  {32'hbf855962, 32'hc18daf75} /* (19, 17, 8) {real, imag} */,
  {32'h40bf5a72, 32'hc1234bd8} /* (19, 17, 7) {real, imag} */,
  {32'hc08468b2, 32'h40a37b84} /* (19, 17, 6) {real, imag} */,
  {32'hc172a6ff, 32'hc0e8368a} /* (19, 17, 5) {real, imag} */,
  {32'h4014dcd7, 32'h41870ced} /* (19, 17, 4) {real, imag} */,
  {32'hbf95748d, 32'hbfb924f0} /* (19, 17, 3) {real, imag} */,
  {32'h40ce91d1, 32'hbea3f680} /* (19, 17, 2) {real, imag} */,
  {32'h408547af, 32'hbf844619} /* (19, 17, 1) {real, imag} */,
  {32'h41267450, 32'h41052775} /* (19, 17, 0) {real, imag} */,
  {32'hbf8a387c, 32'hbf926228} /* (19, 16, 31) {real, imag} */,
  {32'hc0a760ba, 32'h41199406} /* (19, 16, 30) {real, imag} */,
  {32'h404df51e, 32'h4068e6dc} /* (19, 16, 29) {real, imag} */,
  {32'h3f174d75, 32'hc08ce4a0} /* (19, 16, 28) {real, imag} */,
  {32'hbf92f174, 32'hc09793c6} /* (19, 16, 27) {real, imag} */,
  {32'hbff8a327, 32'hc14903ac} /* (19, 16, 26) {real, imag} */,
  {32'h40a6d7d3, 32'h40ae8fda} /* (19, 16, 25) {real, imag} */,
  {32'hc1118ea6, 32'h406b9f25} /* (19, 16, 24) {real, imag} */,
  {32'hc00b0f53, 32'hc121f3cb} /* (19, 16, 23) {real, imag} */,
  {32'h408c08e6, 32'hc0a925d5} /* (19, 16, 22) {real, imag} */,
  {32'hc1113fc5, 32'h4005a732} /* (19, 16, 21) {real, imag} */,
  {32'hc0008007, 32'h40252550} /* (19, 16, 20) {real, imag} */,
  {32'hc11777f4, 32'hc0cfd009} /* (19, 16, 19) {real, imag} */,
  {32'h40af2db4, 32'hc0d22232} /* (19, 16, 18) {real, imag} */,
  {32'hc1112631, 32'hbf7403fa} /* (19, 16, 17) {real, imag} */,
  {32'hc0a9cc10, 32'h00000000} /* (19, 16, 16) {real, imag} */,
  {32'hc1112631, 32'h3f7403fa} /* (19, 16, 15) {real, imag} */,
  {32'h40af2db4, 32'h40d22232} /* (19, 16, 14) {real, imag} */,
  {32'hc11777f4, 32'h40cfd009} /* (19, 16, 13) {real, imag} */,
  {32'hc0008007, 32'hc0252550} /* (19, 16, 12) {real, imag} */,
  {32'hc1113fc5, 32'hc005a732} /* (19, 16, 11) {real, imag} */,
  {32'h408c08e6, 32'h40a925d5} /* (19, 16, 10) {real, imag} */,
  {32'hc00b0f53, 32'h4121f3cb} /* (19, 16, 9) {real, imag} */,
  {32'hc1118ea6, 32'hc06b9f25} /* (19, 16, 8) {real, imag} */,
  {32'h40a6d7d3, 32'hc0ae8fda} /* (19, 16, 7) {real, imag} */,
  {32'hbff8a327, 32'h414903ac} /* (19, 16, 6) {real, imag} */,
  {32'hbf92f174, 32'h409793c6} /* (19, 16, 5) {real, imag} */,
  {32'h3f174d75, 32'h408ce4a0} /* (19, 16, 4) {real, imag} */,
  {32'h404df51e, 32'hc068e6dc} /* (19, 16, 3) {real, imag} */,
  {32'hc0a760ba, 32'hc1199406} /* (19, 16, 2) {real, imag} */,
  {32'hbf8a387c, 32'h3f926228} /* (19, 16, 1) {real, imag} */,
  {32'hc121e5d3, 32'h00000000} /* (19, 16, 0) {real, imag} */,
  {32'h408547af, 32'h3f844619} /* (19, 15, 31) {real, imag} */,
  {32'h40ce91d1, 32'h3ea3f680} /* (19, 15, 30) {real, imag} */,
  {32'hbf95748d, 32'h3fb924f0} /* (19, 15, 29) {real, imag} */,
  {32'h4014dcd7, 32'hc1870ced} /* (19, 15, 28) {real, imag} */,
  {32'hc172a6ff, 32'h40e8368a} /* (19, 15, 27) {real, imag} */,
  {32'hc08468b2, 32'hc0a37b84} /* (19, 15, 26) {real, imag} */,
  {32'h40bf5a72, 32'h41234bd8} /* (19, 15, 25) {real, imag} */,
  {32'hbf855962, 32'h418daf75} /* (19, 15, 24) {real, imag} */,
  {32'hc108a09a, 32'h40e832e6} /* (19, 15, 23) {real, imag} */,
  {32'hc0a20322, 32'h40ea4a74} /* (19, 15, 22) {real, imag} */,
  {32'h406c1814, 32'hc0b50942} /* (19, 15, 21) {real, imag} */,
  {32'hbf3bd7f2, 32'hc01dddc4} /* (19, 15, 20) {real, imag} */,
  {32'h415bd79a, 32'hc0ba56e6} /* (19, 15, 19) {real, imag} */,
  {32'h4109c8f8, 32'hbfdad057} /* (19, 15, 18) {real, imag} */,
  {32'h403d99cc, 32'h40bc8a48} /* (19, 15, 17) {real, imag} */,
  {32'h412f5a5c, 32'h402c2f82} /* (19, 15, 16) {real, imag} */,
  {32'h4095fe80, 32'h41178ccc} /* (19, 15, 15) {real, imag} */,
  {32'hc0fe841e, 32'h41635da4} /* (19, 15, 14) {real, imag} */,
  {32'hbfe423ac, 32'hbf818b88} /* (19, 15, 13) {real, imag} */,
  {32'h400fd86c, 32'hc0c25aef} /* (19, 15, 12) {real, imag} */,
  {32'h409b3052, 32'h40a219ff} /* (19, 15, 11) {real, imag} */,
  {32'hbfb5f49c, 32'hc15d87d8} /* (19, 15, 10) {real, imag} */,
  {32'h40de79a4, 32'h3f7c9c0c} /* (19, 15, 9) {real, imag} */,
  {32'h403ed2ff, 32'h40944502} /* (19, 15, 8) {real, imag} */,
  {32'hbfbba038, 32'h4190edf4} /* (19, 15, 7) {real, imag} */,
  {32'h4161ea51, 32'hc1957bf0} /* (19, 15, 6) {real, imag} */,
  {32'h40c20878, 32'h403998e2} /* (19, 15, 5) {real, imag} */,
  {32'h40abaa5a, 32'hc0d1f4e8} /* (19, 15, 4) {real, imag} */,
  {32'h3f81b110, 32'h3fde3349} /* (19, 15, 3) {real, imag} */,
  {32'h40278f08, 32'h40973695} /* (19, 15, 2) {real, imag} */,
  {32'h3fb064fa, 32'hc0878794} /* (19, 15, 1) {real, imag} */,
  {32'h41267450, 32'hc1052775} /* (19, 15, 0) {real, imag} */,
  {32'h41449c92, 32'h41a31b12} /* (19, 14, 31) {real, imag} */,
  {32'hbdfd4c00, 32'hc11573d5} /* (19, 14, 30) {real, imag} */,
  {32'hc030dc3a, 32'hc0f54b02} /* (19, 14, 29) {real, imag} */,
  {32'h40a6146e, 32'h41989c20} /* (19, 14, 28) {real, imag} */,
  {32'h3ea5df38, 32'hbfa9d734} /* (19, 14, 27) {real, imag} */,
  {32'h3f0fb6c8, 32'h40a93c5b} /* (19, 14, 26) {real, imag} */,
  {32'hc030162c, 32'h409c3e66} /* (19, 14, 25) {real, imag} */,
  {32'h402f73e6, 32'h409df35e} /* (19, 14, 24) {real, imag} */,
  {32'h41363802, 32'hc0e430e2} /* (19, 14, 23) {real, imag} */,
  {32'h417521f8, 32'hc1120d88} /* (19, 14, 22) {real, imag} */,
  {32'h412856d8, 32'h3ed3d1a0} /* (19, 14, 21) {real, imag} */,
  {32'h409cb895, 32'h41380ae4} /* (19, 14, 20) {real, imag} */,
  {32'h40c212f8, 32'h40e4065a} /* (19, 14, 19) {real, imag} */,
  {32'hc1325591, 32'hbfbff004} /* (19, 14, 18) {real, imag} */,
  {32'hc0a7455c, 32'h400d88f6} /* (19, 14, 17) {real, imag} */,
  {32'hc0f22b6a, 32'h40f1c34c} /* (19, 14, 16) {real, imag} */,
  {32'h410cbdbc, 32'h3fd4fcae} /* (19, 14, 15) {real, imag} */,
  {32'h40cf743b, 32'hc00d81b6} /* (19, 14, 14) {real, imag} */,
  {32'hc0813f30, 32'h4041b21f} /* (19, 14, 13) {real, imag} */,
  {32'h405e2570, 32'hc08b5eeb} /* (19, 14, 12) {real, imag} */,
  {32'h3fe8795f, 32'hc0d8fa54} /* (19, 14, 11) {real, imag} */,
  {32'h4116bcbe, 32'h403c2b37} /* (19, 14, 10) {real, imag} */,
  {32'hc1608d97, 32'h402df0c3} /* (19, 14, 9) {real, imag} */,
  {32'h406e1f74, 32'h40abb1ab} /* (19, 14, 8) {real, imag} */,
  {32'h41199d62, 32'hbfe6bb97} /* (19, 14, 7) {real, imag} */,
  {32'hc0daf0d6, 32'hc112f4e4} /* (19, 14, 6) {real, imag} */,
  {32'hc0ee3b2d, 32'hc0d9e419} /* (19, 14, 5) {real, imag} */,
  {32'h40c8f3aa, 32'hc04aa9fc} /* (19, 14, 4) {real, imag} */,
  {32'hbfa3ae4b, 32'hbfeed308} /* (19, 14, 3) {real, imag} */,
  {32'h401843d8, 32'h3ef34b48} /* (19, 14, 2) {real, imag} */,
  {32'hc1357247, 32'h3fb04d28} /* (19, 14, 1) {real, imag} */,
  {32'hc0e7542b, 32'h3f312158} /* (19, 14, 0) {real, imag} */,
  {32'h412c7cee, 32'h4045dff3} /* (19, 13, 31) {real, imag} */,
  {32'hc0bf7f7d, 32'h40d80e9a} /* (19, 13, 30) {real, imag} */,
  {32'hc1b069ae, 32'hc16b45ca} /* (19, 13, 29) {real, imag} */,
  {32'hbebb3d08, 32'hc1253688} /* (19, 13, 28) {real, imag} */,
  {32'hc15d52f0, 32'h40bfde90} /* (19, 13, 27) {real, imag} */,
  {32'hbfbf44ae, 32'h410731d8} /* (19, 13, 26) {real, imag} */,
  {32'h40e14886, 32'h3fe561ac} /* (19, 13, 25) {real, imag} */,
  {32'hc1074d72, 32'hc08ddad0} /* (19, 13, 24) {real, imag} */,
  {32'hc11551e1, 32'h3f97b210} /* (19, 13, 23) {real, imag} */,
  {32'h40e6ecc3, 32'h4140c643} /* (19, 13, 22) {real, imag} */,
  {32'h40b1dbc8, 32'h406da332} /* (19, 13, 21) {real, imag} */,
  {32'hc07d495e, 32'hc0e0e038} /* (19, 13, 20) {real, imag} */,
  {32'h41101b56, 32'h411aa538} /* (19, 13, 19) {real, imag} */,
  {32'hbfff933f, 32'hc1443bd1} /* (19, 13, 18) {real, imag} */,
  {32'hc0eea98c, 32'hc0b653ea} /* (19, 13, 17) {real, imag} */,
  {32'h408f7d66, 32'h4006aa52} /* (19, 13, 16) {real, imag} */,
  {32'h4106cb08, 32'h414e5517} /* (19, 13, 15) {real, imag} */,
  {32'hc14705fc, 32'hc1f5cff7} /* (19, 13, 14) {real, imag} */,
  {32'hc136eeb0, 32'hc1771af0} /* (19, 13, 13) {real, imag} */,
  {32'h4157234c, 32'h40e79836} /* (19, 13, 12) {real, imag} */,
  {32'hc029fcf6, 32'h41f11246} /* (19, 13, 11) {real, imag} */,
  {32'h41a3fbe8, 32'hc0e778da} /* (19, 13, 10) {real, imag} */,
  {32'hc0760be2, 32'h4133f26b} /* (19, 13, 9) {real, imag} */,
  {32'h40e9bb28, 32'hc013d4eb} /* (19, 13, 8) {real, imag} */,
  {32'hbff61604, 32'hc0d213ca} /* (19, 13, 7) {real, imag} */,
  {32'h4199d886, 32'hbed8c64e} /* (19, 13, 6) {real, imag} */,
  {32'h4148ef50, 32'hc1265b3f} /* (19, 13, 5) {real, imag} */,
  {32'hc1339fa4, 32'hc140c668} /* (19, 13, 4) {real, imag} */,
  {32'h4169f39f, 32'h40c1722a} /* (19, 13, 3) {real, imag} */,
  {32'hc0cd7ffc, 32'hc0ef10de} /* (19, 13, 2) {real, imag} */,
  {32'hc174069e, 32'hc0576d11} /* (19, 13, 1) {real, imag} */,
  {32'h409a0125, 32'hc003fafd} /* (19, 13, 0) {real, imag} */,
  {32'h40bcbe93, 32'hc0e2f348} /* (19, 12, 31) {real, imag} */,
  {32'h4092902c, 32'hc14c86b2} /* (19, 12, 30) {real, imag} */,
  {32'h40c5de43, 32'h40bfcbcd} /* (19, 12, 29) {real, imag} */,
  {32'hc194e264, 32'hc128cfbc} /* (19, 12, 28) {real, imag} */,
  {32'hc10fc47e, 32'h40f0278f} /* (19, 12, 27) {real, imag} */,
  {32'h4199a17b, 32'h41450c56} /* (19, 12, 26) {real, imag} */,
  {32'hc0c5851e, 32'hc18e0760} /* (19, 12, 25) {real, imag} */,
  {32'hc0b92cf4, 32'h40d46292} /* (19, 12, 24) {real, imag} */,
  {32'hbf8fdcf4, 32'hc117167d} /* (19, 12, 23) {real, imag} */,
  {32'hc0cc6f88, 32'h40bda914} /* (19, 12, 22) {real, imag} */,
  {32'hc1c77b87, 32'h419dc757} /* (19, 12, 21) {real, imag} */,
  {32'hc0888e42, 32'hc085edf6} /* (19, 12, 20) {real, imag} */,
  {32'hc09e240a, 32'hc19e8a29} /* (19, 12, 19) {real, imag} */,
  {32'hc1808b60, 32'h413a3ac0} /* (19, 12, 18) {real, imag} */,
  {32'h414c618e, 32'h40cadde0} /* (19, 12, 17) {real, imag} */,
  {32'h410edefb, 32'hbe3cc500} /* (19, 12, 16) {real, imag} */,
  {32'h3fed7f40, 32'h400e19b7} /* (19, 12, 15) {real, imag} */,
  {32'h4180672c, 32'h4003813c} /* (19, 12, 14) {real, imag} */,
  {32'hc1aac912, 32'h3f0183b0} /* (19, 12, 13) {real, imag} */,
  {32'h3fdc6560, 32'hc1871036} /* (19, 12, 12) {real, imag} */,
  {32'h410c9a4b, 32'h40c95302} /* (19, 12, 11) {real, imag} */,
  {32'hc156247a, 32'h41c70862} /* (19, 12, 10) {real, imag} */,
  {32'h41d7366f, 32'h417d28d4} /* (19, 12, 9) {real, imag} */,
  {32'h418247a4, 32'hc113a01f} /* (19, 12, 8) {real, imag} */,
  {32'hc10a6874, 32'hc1261034} /* (19, 12, 7) {real, imag} */,
  {32'hc0e25868, 32'hc06f186a} /* (19, 12, 6) {real, imag} */,
  {32'hc0b80d84, 32'h412b46f3} /* (19, 12, 5) {real, imag} */,
  {32'h4015eb6a, 32'hbff2ab98} /* (19, 12, 4) {real, imag} */,
  {32'hc1029364, 32'hbb53a000} /* (19, 12, 3) {real, imag} */,
  {32'hbf87ed54, 32'h40a077ee} /* (19, 12, 2) {real, imag} */,
  {32'h413f7ec1, 32'h41235db8} /* (19, 12, 1) {real, imag} */,
  {32'h41126f9b, 32'hbe0b3dc0} /* (19, 12, 0) {real, imag} */,
  {32'h419c2b15, 32'hc000c507} /* (19, 11, 31) {real, imag} */,
  {32'hbffb843c, 32'hc17d4829} /* (19, 11, 30) {real, imag} */,
  {32'h41296676, 32'hc00f6bca} /* (19, 11, 29) {real, imag} */,
  {32'hc0886e32, 32'hc12d8b2a} /* (19, 11, 28) {real, imag} */,
  {32'hc074f630, 32'h412cb6a4} /* (19, 11, 27) {real, imag} */,
  {32'hc0e9b0ae, 32'hc08ec48e} /* (19, 11, 26) {real, imag} */,
  {32'h4102406f, 32'hc11c57a1} /* (19, 11, 25) {real, imag} */,
  {32'hc1a92de6, 32'h4034740c} /* (19, 11, 24) {real, imag} */,
  {32'h41018724, 32'h4058510e} /* (19, 11, 23) {real, imag} */,
  {32'hc1154bfb, 32'h4153250b} /* (19, 11, 22) {real, imag} */,
  {32'h417910c4, 32'h41594d54} /* (19, 11, 21) {real, imag} */,
  {32'h4042a75a, 32'hbfabf698} /* (19, 11, 20) {real, imag} */,
  {32'h40a3408c, 32'hc0ea76a5} /* (19, 11, 19) {real, imag} */,
  {32'h411d989d, 32'hc0fd79bb} /* (19, 11, 18) {real, imag} */,
  {32'h40022cc6, 32'h3f148f30} /* (19, 11, 17) {real, imag} */,
  {32'h40fba3b2, 32'hc0bc76c0} /* (19, 11, 16) {real, imag} */,
  {32'hc0fef14d, 32'h40301e43} /* (19, 11, 15) {real, imag} */,
  {32'hc124eb35, 32'h40d9ae24} /* (19, 11, 14) {real, imag} */,
  {32'h415f15b9, 32'hc0c70dc6} /* (19, 11, 13) {real, imag} */,
  {32'hc12c722d, 32'h416bb1d0} /* (19, 11, 12) {real, imag} */,
  {32'h409ea468, 32'hc10b0e46} /* (19, 11, 11) {real, imag} */,
  {32'hc14f4687, 32'hc10ae2ba} /* (19, 11, 10) {real, imag} */,
  {32'hc0f8aba4, 32'hbf43a260} /* (19, 11, 9) {real, imag} */,
  {32'hc11934e6, 32'h407375c9} /* (19, 11, 8) {real, imag} */,
  {32'hc1781009, 32'h411ebf7a} /* (19, 11, 7) {real, imag} */,
  {32'hc0405a93, 32'hc103153a} /* (19, 11, 6) {real, imag} */,
  {32'hc0ab207c, 32'hc0ca96d3} /* (19, 11, 5) {real, imag} */,
  {32'h41085c22, 32'hc15b53cd} /* (19, 11, 4) {real, imag} */,
  {32'hc115948f, 32'h3ecb1660} /* (19, 11, 3) {real, imag} */,
  {32'h40d0a15e, 32'hc180ffda} /* (19, 11, 2) {real, imag} */,
  {32'h3ec5b620, 32'h418eeb9d} /* (19, 11, 1) {real, imag} */,
  {32'h4202f94f, 32'h4143a0b4} /* (19, 11, 0) {real, imag} */,
  {32'h3fcb0c1e, 32'hc114554b} /* (19, 10, 31) {real, imag} */,
  {32'h406d9b02, 32'hc1c5759b} /* (19, 10, 30) {real, imag} */,
  {32'hc15dab3e, 32'hc0f96596} /* (19, 10, 29) {real, imag} */,
  {32'h4153451c, 32'h41421426} /* (19, 10, 28) {real, imag} */,
  {32'h40af24ce, 32'h3f765330} /* (19, 10, 27) {real, imag} */,
  {32'hc0f40fc9, 32'h40d017c7} /* (19, 10, 26) {real, imag} */,
  {32'h419a9af9, 32'hc17ff782} /* (19, 10, 25) {real, imag} */,
  {32'hc16fbf22, 32'h41653d36} /* (19, 10, 24) {real, imag} */,
  {32'h3ee24598, 32'hc0ce695e} /* (19, 10, 23) {real, imag} */,
  {32'hc0fdce1b, 32'h40d1e272} /* (19, 10, 22) {real, imag} */,
  {32'h3ffad38c, 32'h41337604} /* (19, 10, 21) {real, imag} */,
  {32'h41202b04, 32'hc0897b70} /* (19, 10, 20) {real, imag} */,
  {32'h407042b0, 32'hc078cc50} /* (19, 10, 19) {real, imag} */,
  {32'h4108a17a, 32'h3fd410aa} /* (19, 10, 18) {real, imag} */,
  {32'hc0eb27d0, 32'hc1261bdd} /* (19, 10, 17) {real, imag} */,
  {32'hc1260e08, 32'hc1adfa22} /* (19, 10, 16) {real, imag} */,
  {32'hbf93924a, 32'hbd2e1100} /* (19, 10, 15) {real, imag} */,
  {32'h411c551c, 32'h410002b2} /* (19, 10, 14) {real, imag} */,
  {32'h403a5e96, 32'hc088427f} /* (19, 10, 13) {real, imag} */,
  {32'hc16f9ab0, 32'h3ffef1d2} /* (19, 10, 12) {real, imag} */,
  {32'h40dafb14, 32'hc106175c} /* (19, 10, 11) {real, imag} */,
  {32'h3f932238, 32'hc096dc3c} /* (19, 10, 10) {real, imag} */,
  {32'hc1b0ae04, 32'h40e1269a} /* (19, 10, 9) {real, imag} */,
  {32'hc093a8c0, 32'h41e31878} /* (19, 10, 8) {real, imag} */,
  {32'hc14d1e7e, 32'hbf5c1a44} /* (19, 10, 7) {real, imag} */,
  {32'hc1bbf721, 32'hc1331880} /* (19, 10, 6) {real, imag} */,
  {32'hc1621516, 32'h40f4c836} /* (19, 10, 5) {real, imag} */,
  {32'hc1103e9c, 32'hc0d88846} /* (19, 10, 4) {real, imag} */,
  {32'hc169cde8, 32'h40d72f88} /* (19, 10, 3) {real, imag} */,
  {32'h41c464da, 32'h4148e6c6} /* (19, 10, 2) {real, imag} */,
  {32'hc113c848, 32'hc18630c8} /* (19, 10, 1) {real, imag} */,
  {32'hc0d53874, 32'h3ddc6040} /* (19, 10, 0) {real, imag} */,
  {32'h4090293b, 32'h418540ae} /* (19, 9, 31) {real, imag} */,
  {32'hc17692ab, 32'h422a495c} /* (19, 9, 30) {real, imag} */,
  {32'h41bacf45, 32'h40d119b8} /* (19, 9, 29) {real, imag} */,
  {32'hc12e0c91, 32'hc149a753} /* (19, 9, 28) {real, imag} */,
  {32'h408beff2, 32'hc1ee5048} /* (19, 9, 27) {real, imag} */,
  {32'hc1df7430, 32'hc08778e4} /* (19, 9, 26) {real, imag} */,
  {32'h40ca7542, 32'h40aa42b0} /* (19, 9, 25) {real, imag} */,
  {32'h401b55b6, 32'h411fa0e4} /* (19, 9, 24) {real, imag} */,
  {32'hc1353168, 32'h40e8211a} /* (19, 9, 23) {real, imag} */,
  {32'h4105b66a, 32'h40de516d} /* (19, 9, 22) {real, imag} */,
  {32'hc1497cb8, 32'h403e4d07} /* (19, 9, 21) {real, imag} */,
  {32'hc01b5161, 32'h405f0c02} /* (19, 9, 20) {real, imag} */,
  {32'h4102fed6, 32'h41ac3f02} /* (19, 9, 19) {real, imag} */,
  {32'h3f7a4d00, 32'hc10b650e} /* (19, 9, 18) {real, imag} */,
  {32'h4194be80, 32'h3fdb16d0} /* (19, 9, 17) {real, imag} */,
  {32'hbf1c2870, 32'h3cfbc500} /* (19, 9, 16) {real, imag} */,
  {32'h410b6aa5, 32'hc169c7f0} /* (19, 9, 15) {real, imag} */,
  {32'h40984ac4, 32'h418e23a2} /* (19, 9, 14) {real, imag} */,
  {32'hbfe9368b, 32'hc15f3e17} /* (19, 9, 13) {real, imag} */,
  {32'hc08bc99b, 32'hc0db371a} /* (19, 9, 12) {real, imag} */,
  {32'h40c91ae4, 32'h410cbd70} /* (19, 9, 11) {real, imag} */,
  {32'h414ed0bc, 32'hc0c6b75f} /* (19, 9, 10) {real, imag} */,
  {32'h3f8b709c, 32'h410bd287} /* (19, 9, 9) {real, imag} */,
  {32'hc15f6d73, 32'hc13da109} /* (19, 9, 8) {real, imag} */,
  {32'h3fb3125a, 32'h4081d186} /* (19, 9, 7) {real, imag} */,
  {32'hbdd83880, 32'h4040b226} /* (19, 9, 6) {real, imag} */,
  {32'h40c07476, 32'h41a4fd1e} /* (19, 9, 5) {real, imag} */,
  {32'hc10bd3ae, 32'hc10d9e7a} /* (19, 9, 4) {real, imag} */,
  {32'hbf9e958a, 32'hc1c63506} /* (19, 9, 3) {real, imag} */,
  {32'hc092671b, 32'h41d122ed} /* (19, 9, 2) {real, imag} */,
  {32'h3fa2150c, 32'hc1cf3c73} /* (19, 9, 1) {real, imag} */,
  {32'hbfa6ea9e, 32'hc0117f98} /* (19, 9, 0) {real, imag} */,
  {32'h420fd2ad, 32'h4200de7d} /* (19, 8, 31) {real, imag} */,
  {32'hc1b7d7d7, 32'h41083db0} /* (19, 8, 30) {real, imag} */,
  {32'h3e9d9940, 32'hc1ad1e17} /* (19, 8, 29) {real, imag} */,
  {32'hc182e730, 32'h41deaad3} /* (19, 8, 28) {real, imag} */,
  {32'hc192b746, 32'h4029de03} /* (19, 8, 27) {real, imag} */,
  {32'hc160f108, 32'hc09a4e03} /* (19, 8, 26) {real, imag} */,
  {32'h40de8cba, 32'h40312ed8} /* (19, 8, 25) {real, imag} */,
  {32'hc136478e, 32'hc0e4f9fc} /* (19, 8, 24) {real, imag} */,
  {32'hc15ce57a, 32'h415ac673} /* (19, 8, 23) {real, imag} */,
  {32'hc0f85b2e, 32'hc01dc874} /* (19, 8, 22) {real, imag} */,
  {32'h40af03c4, 32'hc0d2aca8} /* (19, 8, 21) {real, imag} */,
  {32'hc0991e02, 32'hbfd0f430} /* (19, 8, 20) {real, imag} */,
  {32'hc109fffc, 32'hc0c104a2} /* (19, 8, 19) {real, imag} */,
  {32'hbfc710e4, 32'h409a98fe} /* (19, 8, 18) {real, imag} */,
  {32'hc158cf56, 32'hc09c29ca} /* (19, 8, 17) {real, imag} */,
  {32'h40dacbba, 32'h4082309a} /* (19, 8, 16) {real, imag} */,
  {32'h412ad4a5, 32'hc0c31586} /* (19, 8, 15) {real, imag} */,
  {32'h40ca2d5c, 32'h412a7baa} /* (19, 8, 14) {real, imag} */,
  {32'h3fd997f6, 32'hc1a4acdd} /* (19, 8, 13) {real, imag} */,
  {32'h4090a3c2, 32'hc0f96b16} /* (19, 8, 12) {real, imag} */,
  {32'h4129bcd4, 32'h413fcb1f} /* (19, 8, 11) {real, imag} */,
  {32'hc0df8de7, 32'h40710b67} /* (19, 8, 10) {real, imag} */,
  {32'hc083ac35, 32'hc13711f3} /* (19, 8, 9) {real, imag} */,
  {32'hc1bb8c2a, 32'h4120f158} /* (19, 8, 8) {real, imag} */,
  {32'hc162a11d, 32'h3dd03fa0} /* (19, 8, 7) {real, imag} */,
  {32'h41bf9aa8, 32'hc15a923e} /* (19, 8, 6) {real, imag} */,
  {32'h4118e6b8, 32'hc2032d05} /* (19, 8, 5) {real, imag} */,
  {32'h418efa06, 32'h413d6898} /* (19, 8, 4) {real, imag} */,
  {32'hc0b83e9a, 32'h410fd540} /* (19, 8, 3) {real, imag} */,
  {32'hc2082f95, 32'hc18ed096} /* (19, 8, 2) {real, imag} */,
  {32'h418e2444, 32'h420255e2} /* (19, 8, 1) {real, imag} */,
  {32'h41b75556, 32'h4185c36d} /* (19, 8, 0) {real, imag} */,
  {32'hc1eb5acd, 32'hc181bdf6} /* (19, 7, 31) {real, imag} */,
  {32'h404fc71f, 32'h4024536e} /* (19, 7, 30) {real, imag} */,
  {32'hc11991c4, 32'hbf421b70} /* (19, 7, 29) {real, imag} */,
  {32'h40b6d0a4, 32'h4113d83a} /* (19, 7, 28) {real, imag} */,
  {32'h41b74788, 32'h4173e716} /* (19, 7, 27) {real, imag} */,
  {32'hc102eae2, 32'hc1b10672} /* (19, 7, 26) {real, imag} */,
  {32'hc10228bb, 32'hc05179f6} /* (19, 7, 25) {real, imag} */,
  {32'h402d9db2, 32'hc1285522} /* (19, 7, 24) {real, imag} */,
  {32'h3e2c7680, 32'h41e03940} /* (19, 7, 23) {real, imag} */,
  {32'h40901794, 32'h3f820dd0} /* (19, 7, 22) {real, imag} */,
  {32'h413b2285, 32'h3fb64ee0} /* (19, 7, 21) {real, imag} */,
  {32'hc04d48fc, 32'h4111f961} /* (19, 7, 20) {real, imag} */,
  {32'h3e606de0, 32'hc0c839f4} /* (19, 7, 19) {real, imag} */,
  {32'h4036562e, 32'hc0ee3590} /* (19, 7, 18) {real, imag} */,
  {32'h40d42d9d, 32'h40e50067} /* (19, 7, 17) {real, imag} */,
  {32'h410e8ce2, 32'hc1590632} /* (19, 7, 16) {real, imag} */,
  {32'hc03e668a, 32'h4130bbc6} /* (19, 7, 15) {real, imag} */,
  {32'hc0128e4e, 32'hc0c91ca8} /* (19, 7, 14) {real, imag} */,
  {32'h41457595, 32'h40d9b97a} /* (19, 7, 13) {real, imag} */,
  {32'hbf82c1f8, 32'h3f60e020} /* (19, 7, 12) {real, imag} */,
  {32'hc0b2ef24, 32'h404ecb51} /* (19, 7, 11) {real, imag} */,
  {32'hc12b28ca, 32'hc09dd2fa} /* (19, 7, 10) {real, imag} */,
  {32'h414accc2, 32'hc0885364} /* (19, 7, 9) {real, imag} */,
  {32'hbf90fbc0, 32'h40eac096} /* (19, 7, 8) {real, imag} */,
  {32'hc1b63d96, 32'h40278ce7} /* (19, 7, 7) {real, imag} */,
  {32'h4123b9dc, 32'hc123cba5} /* (19, 7, 6) {real, imag} */,
  {32'h402a3790, 32'hc03a3962} /* (19, 7, 5) {real, imag} */,
  {32'h4109e116, 32'hc073b504} /* (19, 7, 4) {real, imag} */,
  {32'h41a4558c, 32'h410649d7} /* (19, 7, 3) {real, imag} */,
  {32'h412e4796, 32'h3ee9cb20} /* (19, 7, 2) {real, imag} */,
  {32'hbc5e3400, 32'hc1b658aa} /* (19, 7, 1) {real, imag} */,
  {32'hbefb8bd0, 32'hc1dd3b81} /* (19, 7, 0) {real, imag} */,
  {32'hc0fefcf3, 32'hc024e73e} /* (19, 6, 31) {real, imag} */,
  {32'hc0f2464c, 32'h4022b9f8} /* (19, 6, 30) {real, imag} */,
  {32'hc1b5c7ff, 32'h40de49fc} /* (19, 6, 29) {real, imag} */,
  {32'h40eeb21e, 32'h411007f9} /* (19, 6, 28) {real, imag} */,
  {32'hc1105c0d, 32'hc10a4c61} /* (19, 6, 27) {real, imag} */,
  {32'hc0691fc0, 32'hc0f0c93a} /* (19, 6, 26) {real, imag} */,
  {32'hc0bd4447, 32'hc0392c38} /* (19, 6, 25) {real, imag} */,
  {32'hc17eb02c, 32'hc1ad7a0a} /* (19, 6, 24) {real, imag} */,
  {32'hc084bc76, 32'h414f28f3} /* (19, 6, 23) {real, imag} */,
  {32'h41dc604b, 32'h40637ecc} /* (19, 6, 22) {real, imag} */,
  {32'hc0b8b133, 32'h408e468d} /* (19, 6, 21) {real, imag} */,
  {32'hbfa4e76d, 32'hc07b9ce0} /* (19, 6, 20) {real, imag} */,
  {32'h409c54c4, 32'h3f86321c} /* (19, 6, 19) {real, imag} */,
  {32'hc14dbfe4, 32'hc18c723a} /* (19, 6, 18) {real, imag} */,
  {32'hbfddfaa6, 32'hc1088d8c} /* (19, 6, 17) {real, imag} */,
  {32'hbfe3e088, 32'h3febac5c} /* (19, 6, 16) {real, imag} */,
  {32'hc0f08ee4, 32'h415aa2e1} /* (19, 6, 15) {real, imag} */,
  {32'h40bcbb34, 32'hc1d0c56e} /* (19, 6, 14) {real, imag} */,
  {32'h4066c008, 32'h40e76597} /* (19, 6, 13) {real, imag} */,
  {32'h405af764, 32'h3dadd860} /* (19, 6, 12) {real, imag} */,
  {32'hbfe3397c, 32'h4092e3d2} /* (19, 6, 11) {real, imag} */,
  {32'h40f52360, 32'hc080ff0c} /* (19, 6, 10) {real, imag} */,
  {32'hc2037597, 32'hc09db860} /* (19, 6, 9) {real, imag} */,
  {32'hc1871d73, 32'h41bf1688} /* (19, 6, 8) {real, imag} */,
  {32'h403f0f70, 32'h3f1d3310} /* (19, 6, 7) {real, imag} */,
  {32'h41f4b90e, 32'hc11c5459} /* (19, 6, 6) {real, imag} */,
  {32'hc172708c, 32'hc186b3a2} /* (19, 6, 5) {real, imag} */,
  {32'hc0d9d17a, 32'h41d601fe} /* (19, 6, 4) {real, imag} */,
  {32'h41e09a3d, 32'hc18d7073} /* (19, 6, 3) {real, imag} */,
  {32'hc1082679, 32'hc14602e8} /* (19, 6, 2) {real, imag} */,
  {32'hc120fc08, 32'hbf487840} /* (19, 6, 1) {real, imag} */,
  {32'hc030cfbc, 32'h4148823a} /* (19, 6, 0) {real, imag} */,
  {32'h42d27f34, 32'hc13bb466} /* (19, 5, 31) {real, imag} */,
  {32'hc245716e, 32'h40db76a2} /* (19, 5, 30) {real, imag} */,
  {32'h418f7300, 32'h42072e5d} /* (19, 5, 29) {real, imag} */,
  {32'hc18d3c62, 32'hc091bd70} /* (19, 5, 28) {real, imag} */,
  {32'hc1545832, 32'hc1161d6b} /* (19, 5, 27) {real, imag} */,
  {32'h40dcde93, 32'h4181fbd1} /* (19, 5, 26) {real, imag} */,
  {32'h4110cc68, 32'h411f1b4e} /* (19, 5, 25) {real, imag} */,
  {32'hc133fd88, 32'hc1908162} /* (19, 5, 24) {real, imag} */,
  {32'hc08496bc, 32'h415fb443} /* (19, 5, 23) {real, imag} */,
  {32'h3f835870, 32'h418c5db3} /* (19, 5, 22) {real, imag} */,
  {32'hc0ce5fbe, 32'h4114128f} /* (19, 5, 21) {real, imag} */,
  {32'hc0e5bf52, 32'hbf4f7918} /* (19, 5, 20) {real, imag} */,
  {32'hc0c6b7c4, 32'h4048c093} /* (19, 5, 19) {real, imag} */,
  {32'h4116676a, 32'h41733c61} /* (19, 5, 18) {real, imag} */,
  {32'h419c751e, 32'h40929ff2} /* (19, 5, 17) {real, imag} */,
  {32'hc080d748, 32'h411e8bc0} /* (19, 5, 16) {real, imag} */,
  {32'h410973a9, 32'hc0cc8f5a} /* (19, 5, 15) {real, imag} */,
  {32'hbc8b9d60, 32'hc0a88c9d} /* (19, 5, 14) {real, imag} */,
  {32'hc04ea606, 32'h3de2ff40} /* (19, 5, 13) {real, imag} */,
  {32'h41587bc4, 32'h40261588} /* (19, 5, 12) {real, imag} */,
  {32'h40c65874, 32'hc0b832c1} /* (19, 5, 11) {real, imag} */,
  {32'hc10855ff, 32'h416b3dec} /* (19, 5, 10) {real, imag} */,
  {32'hc0b53ed3, 32'h419724c7} /* (19, 5, 9) {real, imag} */,
  {32'hc108b8a8, 32'hc0939f89} /* (19, 5, 8) {real, imag} */,
  {32'h422b8570, 32'hc08b872d} /* (19, 5, 7) {real, imag} */,
  {32'hc09c9743, 32'hc196bcec} /* (19, 5, 6) {real, imag} */,
  {32'hc22977b9, 32'h40636958} /* (19, 5, 5) {real, imag} */,
  {32'h41b8956d, 32'h407ae328} /* (19, 5, 4) {real, imag} */,
  {32'h40c11250, 32'h40b1ee9b} /* (19, 5, 3) {real, imag} */,
  {32'hc21a71aa, 32'hc218a112} /* (19, 5, 2) {real, imag} */,
  {32'h42826cc2, 32'h429ceb15} /* (19, 5, 1) {real, imag} */,
  {32'h42335bde, 32'h4226520e} /* (19, 5, 0) {real, imag} */,
  {32'hc226b5c0, 32'hc2eefdb4} /* (19, 4, 31) {real, imag} */,
  {32'h426dd8de, 32'h426ca51b} /* (19, 4, 30) {real, imag} */,
  {32'hc18e63e5, 32'hc0484d1e} /* (19, 4, 29) {real, imag} */,
  {32'hc22cd552, 32'hc13024ae} /* (19, 4, 28) {real, imag} */,
  {32'h424071c9, 32'hc2006161} /* (19, 4, 27) {real, imag} */,
  {32'hc214282e, 32'hc1983514} /* (19, 4, 26) {real, imag} */,
  {32'h4104e112, 32'h41a4b92a} /* (19, 4, 25) {real, imag} */,
  {32'h41849765, 32'hc02f96cc} /* (19, 4, 24) {real, imag} */,
  {32'h3f3b57d0, 32'h4077d6aa} /* (19, 4, 23) {real, imag} */,
  {32'hbf155dc4, 32'h3f86a6a4} /* (19, 4, 22) {real, imag} */,
  {32'h419d38f9, 32'h400b214c} /* (19, 4, 21) {real, imag} */,
  {32'hc1a636ce, 32'hc105043f} /* (19, 4, 20) {real, imag} */,
  {32'hc0d72b2e, 32'hc1d38093} /* (19, 4, 19) {real, imag} */,
  {32'hc12641d6, 32'hbee7a820} /* (19, 4, 18) {real, imag} */,
  {32'h404861d9, 32'hc0b32eac} /* (19, 4, 17) {real, imag} */,
  {32'hc112da76, 32'h401e26ea} /* (19, 4, 16) {real, imag} */,
  {32'hbf8834a0, 32'hc16555d2} /* (19, 4, 15) {real, imag} */,
  {32'hc0cb3354, 32'h415ff7bb} /* (19, 4, 14) {real, imag} */,
  {32'h41834280, 32'h4060beea} /* (19, 4, 13) {real, imag} */,
  {32'hc041d393, 32'hbf41d5e0} /* (19, 4, 12) {real, imag} */,
  {32'hc1331862, 32'h40fc18d2} /* (19, 4, 11) {real, imag} */,
  {32'hc126453a, 32'h3df4a2c0} /* (19, 4, 10) {real, imag} */,
  {32'h3e7547a0, 32'hc13f77df} /* (19, 4, 9) {real, imag} */,
  {32'h408a7c58, 32'h41157658} /* (19, 4, 8) {real, imag} */,
  {32'hc0cd0f69, 32'hc052922e} /* (19, 4, 7) {real, imag} */,
  {32'hc113bf44, 32'h40e3ede6} /* (19, 4, 6) {real, imag} */,
  {32'hbff0d1aa, 32'h41eb6441} /* (19, 4, 5) {real, imag} */,
  {32'h41542306, 32'hc155c51a} /* (19, 4, 4) {real, imag} */,
  {32'hc20c1000, 32'hc1de74b8} /* (19, 4, 3) {real, imag} */,
  {32'h42db3682, 32'h428b5a9b} /* (19, 4, 2) {real, imag} */,
  {32'hc320ee6b, 32'hc295057c} /* (19, 4, 1) {real, imag} */,
  {32'hc2919f9c, 32'hc1a71882} /* (19, 4, 0) {real, imag} */,
  {32'h42ed1552, 32'hc2ff18b3} /* (19, 3, 31) {real, imag} */,
  {32'hc28324c7, 32'h4340b34e} /* (19, 3, 30) {real, imag} */,
  {32'hc20c2a7e, 32'hc0cbd342} /* (19, 3, 29) {real, imag} */,
  {32'hc1b73c64, 32'hc13a94d5} /* (19, 3, 28) {real, imag} */,
  {32'hc064b90c, 32'hc1e43918} /* (19, 3, 27) {real, imag} */,
  {32'h41047d8a, 32'hc0df2cc2} /* (19, 3, 26) {real, imag} */,
  {32'hc1b02a8e, 32'h41f556e4} /* (19, 3, 25) {real, imag} */,
  {32'h4134f57c, 32'hbf876960} /* (19, 3, 24) {real, imag} */,
  {32'h40b1fb91, 32'h41789852} /* (19, 3, 23) {real, imag} */,
  {32'hc20aa34c, 32'hc1d4624a} /* (19, 3, 22) {real, imag} */,
  {32'h4096ccc1, 32'hbfc63cec} /* (19, 3, 21) {real, imag} */,
  {32'h411ec64f, 32'hc15e5611} /* (19, 3, 20) {real, imag} */,
  {32'hc11ef57c, 32'h4192f3f4} /* (19, 3, 19) {real, imag} */,
  {32'h41855cd6, 32'hc0e3d4e6} /* (19, 3, 18) {real, imag} */,
  {32'h404b5068, 32'h40ac92ba} /* (19, 3, 17) {real, imag} */,
  {32'hc02d0c22, 32'hc09b5293} /* (19, 3, 16) {real, imag} */,
  {32'hc11571a9, 32'hc062bc94} /* (19, 3, 15) {real, imag} */,
  {32'hc1072c9f, 32'h408b7e99} /* (19, 3, 14) {real, imag} */,
  {32'hc0f7d880, 32'h40fbecfa} /* (19, 3, 13) {real, imag} */,
  {32'h41a7e896, 32'hbf9a2588} /* (19, 3, 12) {real, imag} */,
  {32'hc174f227, 32'hc119d71f} /* (19, 3, 11) {real, imag} */,
  {32'h411baff1, 32'h41213286} /* (19, 3, 10) {real, imag} */,
  {32'h41035da2, 32'hc19bf923} /* (19, 3, 9) {real, imag} */,
  {32'h3fbf5a18, 32'h40d37ff8} /* (19, 3, 8) {real, imag} */,
  {32'hc1810248, 32'hc0a7daac} /* (19, 3, 7) {real, imag} */,
  {32'h41432411, 32'hbfa2c94e} /* (19, 3, 6) {real, imag} */,
  {32'hc166997b, 32'h3f0d14a0} /* (19, 3, 5) {real, imag} */,
  {32'h41f03abd, 32'h4101f997} /* (19, 3, 4) {real, imag} */,
  {32'h421b4812, 32'hc0bd9077} /* (19, 3, 3) {real, imag} */,
  {32'h4290e6d0, 32'h43044652} /* (19, 3, 2) {real, imag} */,
  {32'hc2f87158, 32'hc2ffa6a3} /* (19, 3, 1) {real, imag} */,
  {32'hc1aa1f56, 32'h4212d83e} /* (19, 3, 0) {real, imag} */,
  {32'h44983966, 32'hc1ee873e} /* (19, 2, 31) {real, imag} */,
  {32'hc4200bf6, 32'h431783a5} /* (19, 2, 30) {real, imag} */,
  {32'h4264ebc4, 32'h411d3bea} /* (19, 2, 29) {real, imag} */,
  {32'h429139d3, 32'hc2a5bd74} /* (19, 2, 28) {real, imag} */,
  {32'hc21d8382, 32'h411546e2} /* (19, 2, 27) {real, imag} */,
  {32'hc107fc44, 32'h4175a83e} /* (19, 2, 26) {real, imag} */,
  {32'h41543815, 32'hc2131c38} /* (19, 2, 25) {real, imag} */,
  {32'hc04e87c0, 32'h41e6da45} /* (19, 2, 24) {real, imag} */,
  {32'hc124df02, 32'hc193f618} /* (19, 2, 23) {real, imag} */,
  {32'h3f739674, 32'hc10c3be0} /* (19, 2, 22) {real, imag} */,
  {32'hc1bcb7f9, 32'h41d04bce} /* (19, 2, 21) {real, imag} */,
  {32'h414f24ed, 32'hc11fc726} /* (19, 2, 20) {real, imag} */,
  {32'hc11aa231, 32'h3ff1d848} /* (19, 2, 19) {real, imag} */,
  {32'h40dbca44, 32'h3f73fe7c} /* (19, 2, 18) {real, imag} */,
  {32'h3eccef60, 32'hc13b548b} /* (19, 2, 17) {real, imag} */,
  {32'h4110cbfe, 32'h3f5516bc} /* (19, 2, 16) {real, imag} */,
  {32'h3fb426c4, 32'h3f96e272} /* (19, 2, 15) {real, imag} */,
  {32'h40614566, 32'hc0b25b9e} /* (19, 2, 14) {real, imag} */,
  {32'h3f938489, 32'h413d4e69} /* (19, 2, 13) {real, imag} */,
  {32'hc134704e, 32'h3f7e7e2c} /* (19, 2, 12) {real, imag} */,
  {32'hc153d6a8, 32'hc1ce17d4} /* (19, 2, 11) {real, imag} */,
  {32'hbfe6ad3e, 32'h410125ef} /* (19, 2, 10) {real, imag} */,
  {32'h410f7533, 32'h412b22eb} /* (19, 2, 9) {real, imag} */,
  {32'hc0c86bd4, 32'hc244d424} /* (19, 2, 8) {real, imag} */,
  {32'h40ecdc44, 32'hc13b3f66} /* (19, 2, 7) {real, imag} */,
  {32'h4102c26a, 32'hc039af58} /* (19, 2, 6) {real, imag} */,
  {32'hc297ab95, 32'hc2a2e8c7} /* (19, 2, 5) {real, imag} */,
  {32'h42e8a60e, 32'hc10d23c2} /* (19, 2, 4) {real, imag} */,
  {32'h41946dcd, 32'h41a50ed3} /* (19, 2, 3) {real, imag} */,
  {32'hc3da912f, 32'h42ef188a} /* (19, 2, 2) {real, imag} */,
  {32'h44341a12, 32'hc30a4c11} /* (19, 2, 1) {real, imag} */,
  {32'h4422870c, 32'h42d27fe6} /* (19, 2, 0) {real, imag} */,
  {32'hc4c755b8, 32'h43cef1e9} /* (19, 1, 31) {real, imag} */,
  {32'h43d45f5f, 32'h41a2f934} /* (19, 1, 30) {real, imag} */,
  {32'hc1a1674d, 32'hc22e63c3} /* (19, 1, 29) {real, imag} */,
  {32'hc2989234, 32'hc2996fae} /* (19, 1, 28) {real, imag} */,
  {32'h42f8108b, 32'h4192529f} /* (19, 1, 27) {real, imag} */,
  {32'h41e15250, 32'hc210711c} /* (19, 1, 26) {real, imag} */,
  {32'hc142ad45, 32'h41f63974} /* (19, 1, 25) {real, imag} */,
  {32'h402c82e0, 32'hc15e57fb} /* (19, 1, 24) {real, imag} */,
  {32'h41cfccd1, 32'hc0ea1754} /* (19, 1, 23) {real, imag} */,
  {32'h40a7127e, 32'h41295a08} /* (19, 1, 22) {real, imag} */,
  {32'h412aef27, 32'hc1c98c38} /* (19, 1, 21) {real, imag} */,
  {32'hbf9cf1f2, 32'h411e022b} /* (19, 1, 20) {real, imag} */,
  {32'h413263bc, 32'h3feb920c} /* (19, 1, 19) {real, imag} */,
  {32'h4137e1e0, 32'hc1b3eae0} /* (19, 1, 18) {real, imag} */,
  {32'hc0fe3945, 32'h3faf1cfc} /* (19, 1, 17) {real, imag} */,
  {32'hc0552879, 32'hbc811980} /* (19, 1, 16) {real, imag} */,
  {32'h40c8eaea, 32'hbffc2fa4} /* (19, 1, 15) {real, imag} */,
  {32'hc0899036, 32'h414c92ce} /* (19, 1, 14) {real, imag} */,
  {32'hbfe172eb, 32'h406be5f8} /* (19, 1, 13) {real, imag} */,
  {32'hc07a8334, 32'h408d6764} /* (19, 1, 12) {real, imag} */,
  {32'h41c6c586, 32'h415ba026} /* (19, 1, 11) {real, imag} */,
  {32'h4187e204, 32'h3fa71c4a} /* (19, 1, 10) {real, imag} */,
  {32'hc1ea3b3f, 32'h3fba1744} /* (19, 1, 9) {real, imag} */,
  {32'h41b8fbac, 32'h41a399dc} /* (19, 1, 8) {real, imag} */,
  {32'hc17e6a95, 32'hc09779ab} /* (19, 1, 7) {real, imag} */,
  {32'h410db760, 32'h4039a8d8} /* (19, 1, 6) {real, imag} */,
  {32'h425c707a, 32'h42174044} /* (19, 1, 5) {real, imag} */,
  {32'hc25ac26a, 32'hc2789b00} /* (19, 1, 4) {real, imag} */,
  {32'h4227ab86, 32'hbefca780} /* (19, 1, 3) {real, imag} */,
  {32'h440653f0, 32'h44149d4d} /* (19, 1, 2) {real, imag} */,
  {32'hc50d96c0, 32'hc4926cb8} /* (19, 1, 1) {real, imag} */,
  {32'hc4f06f6a, 32'hc39e44bc} /* (19, 1, 0) {real, imag} */,
  {32'hc4b4955a, 32'h44871047} /* (19, 0, 31) {real, imag} */,
  {32'h432469c7, 32'hc39d60a3} /* (19, 0, 30) {real, imag} */,
  {32'hc14b3016, 32'hc21247de} /* (19, 0, 29) {real, imag} */,
  {32'hc1392829, 32'hc202596a} /* (19, 0, 28) {real, imag} */,
  {32'h4267ff0e, 32'h41e86c4d} /* (19, 0, 27) {real, imag} */,
  {32'h416c0766, 32'hc1b951c8} /* (19, 0, 26) {real, imag} */,
  {32'hc12ce883, 32'h40ef5ebe} /* (19, 0, 25) {real, imag} */,
  {32'h409f3d16, 32'hc196d38e} /* (19, 0, 24) {real, imag} */,
  {32'h42054f34, 32'hc167621a} /* (19, 0, 23) {real, imag} */,
  {32'hc0c5dd6c, 32'hc141b8fc} /* (19, 0, 22) {real, imag} */,
  {32'h4088e23c, 32'hc08f130f} /* (19, 0, 21) {real, imag} */,
  {32'h408a0bc8, 32'h3ff13f6e} /* (19, 0, 20) {real, imag} */,
  {32'h41435fa0, 32'h403f9ba4} /* (19, 0, 19) {real, imag} */,
  {32'h4125f34e, 32'hc073fffa} /* (19, 0, 18) {real, imag} */,
  {32'hbfcfa002, 32'hbff072d8} /* (19, 0, 17) {real, imag} */,
  {32'h41d4992e, 32'h00000000} /* (19, 0, 16) {real, imag} */,
  {32'hbfcfa002, 32'h3ff072d8} /* (19, 0, 15) {real, imag} */,
  {32'h4125f34e, 32'h4073fffa} /* (19, 0, 14) {real, imag} */,
  {32'h41435fa0, 32'hc03f9ba4} /* (19, 0, 13) {real, imag} */,
  {32'h408a0bc8, 32'hbff13f6e} /* (19, 0, 12) {real, imag} */,
  {32'h4088e23c, 32'h408f130f} /* (19, 0, 11) {real, imag} */,
  {32'hc0c5dd6c, 32'h4141b8fc} /* (19, 0, 10) {real, imag} */,
  {32'h42054f34, 32'h4167621a} /* (19, 0, 9) {real, imag} */,
  {32'h409f3d16, 32'h4196d38e} /* (19, 0, 8) {real, imag} */,
  {32'hc12ce883, 32'hc0ef5ebe} /* (19, 0, 7) {real, imag} */,
  {32'h416c0766, 32'h41b951c8} /* (19, 0, 6) {real, imag} */,
  {32'h4267ff0e, 32'hc1e86c4d} /* (19, 0, 5) {real, imag} */,
  {32'hc1392829, 32'h4202596a} /* (19, 0, 4) {real, imag} */,
  {32'hc14b3016, 32'h421247de} /* (19, 0, 3) {real, imag} */,
  {32'h432469c7, 32'h439d60a3} /* (19, 0, 2) {real, imag} */,
  {32'hc4b4955a, 32'hc4871047} /* (19, 0, 1) {real, imag} */,
  {32'hc502a720, 32'h00000000} /* (19, 0, 0) {real, imag} */,
  {32'hc4ee823b, 32'h44700eda} /* (18, 31, 31) {real, imag} */,
  {32'h43ea29e0, 32'hc4066126} /* (18, 31, 30) {real, imag} */,
  {32'hc1002ec0, 32'h42326612} /* (18, 31, 29) {real, imag} */,
  {32'hc28ec0fb, 32'h41f3042b} /* (18, 31, 28) {real, imag} */,
  {32'h4270565c, 32'hc226304d} /* (18, 31, 27) {real, imag} */,
  {32'h413d99f9, 32'h413b9e74} /* (18, 31, 26) {real, imag} */,
  {32'h41133642, 32'h413e826c} /* (18, 31, 25) {real, imag} */,
  {32'h41d59114, 32'hc225812a} /* (18, 31, 24) {real, imag} */,
  {32'h3ff7aa80, 32'hc020195d} /* (18, 31, 23) {real, imag} */,
  {32'hc04c2398, 32'hc12c2ff1} /* (18, 31, 22) {real, imag} */,
  {32'hc0c6b422, 32'hc1797b76} /* (18, 31, 21) {real, imag} */,
  {32'h417d21e6, 32'hc0aad8a0} /* (18, 31, 20) {real, imag} */,
  {32'hc04d6980, 32'hc042d80e} /* (18, 31, 19) {real, imag} */,
  {32'h40553931, 32'hc1aeca0a} /* (18, 31, 18) {real, imag} */,
  {32'hc128bc65, 32'h401fcaa5} /* (18, 31, 17) {real, imag} */,
  {32'h4119ee35, 32'hbf578718} /* (18, 31, 16) {real, imag} */,
  {32'h413162c4, 32'hc04f189d} /* (18, 31, 15) {real, imag} */,
  {32'h40834555, 32'hc01f2735} /* (18, 31, 14) {real, imag} */,
  {32'h41811eda, 32'h402fd45c} /* (18, 31, 13) {real, imag} */,
  {32'hc1e3cc12, 32'hc0b8bb6e} /* (18, 31, 12) {real, imag} */,
  {32'h41dbea6d, 32'h41bb826a} /* (18, 31, 11) {real, imag} */,
  {32'hbfd8b9ca, 32'hc139152c} /* (18, 31, 10) {real, imag} */,
  {32'hc086d7d4, 32'h41e51a0b} /* (18, 31, 9) {real, imag} */,
  {32'h416afe8a, 32'h41706d21} /* (18, 31, 8) {real, imag} */,
  {32'hc1343e0d, 32'hc1fa1f54} /* (18, 31, 7) {real, imag} */,
  {32'h423f9e19, 32'h420297ce} /* (18, 31, 6) {real, imag} */,
  {32'h42f4b350, 32'h41188ef4} /* (18, 31, 5) {real, imag} */,
  {32'hc29c0b24, 32'h42634bbd} /* (18, 31, 4) {real, imag} */,
  {32'hc12bd25c, 32'hc04813e0} /* (18, 31, 3) {real, imag} */,
  {32'h43b0f2ea, 32'h4248d7d4} /* (18, 31, 2) {real, imag} */,
  {32'hc4a59ac8, 32'hc396bdb0} /* (18, 31, 1) {real, imag} */,
  {32'hc4c974b6, 32'h438889b4} /* (18, 31, 0) {real, imag} */,
  {32'h441ef118, 32'h43063630} /* (18, 30, 31) {real, imag} */,
  {32'hc3bfb06a, 32'hc2e0251e} /* (18, 30, 30) {real, imag} */,
  {32'h421f44af, 32'hc1be5dcc} /* (18, 30, 29) {real, imag} */,
  {32'h42c76c6e, 32'h421b6e10} /* (18, 30, 28) {real, imag} */,
  {32'hc279d368, 32'h42acbb2f} /* (18, 30, 27) {real, imag} */,
  {32'h41b3f47c, 32'hc1bc609f} /* (18, 30, 26) {real, imag} */,
  {32'h41955588, 32'h4102905a} /* (18, 30, 25) {real, imag} */,
  {32'hc14253be, 32'h42234232} /* (18, 30, 24) {real, imag} */,
  {32'h418eae98, 32'h3eb4d750} /* (18, 30, 23) {real, imag} */,
  {32'hc078c564, 32'h407a6448} /* (18, 30, 22) {real, imag} */,
  {32'hc19b09f2, 32'h41c21458} /* (18, 30, 21) {real, imag} */,
  {32'h40d2f316, 32'hc1018188} /* (18, 30, 20) {real, imag} */,
  {32'h3fb0d500, 32'h40eb0c05} /* (18, 30, 19) {real, imag} */,
  {32'hc0361690, 32'h403c9606} /* (18, 30, 18) {real, imag} */,
  {32'h40d4502c, 32'h4093f18a} /* (18, 30, 17) {real, imag} */,
  {32'hbff10c6a, 32'h4053ddd4} /* (18, 30, 16) {real, imag} */,
  {32'h40e2e486, 32'h40887311} /* (18, 30, 15) {real, imag} */,
  {32'hc016983f, 32'hc15174bd} /* (18, 30, 14) {real, imag} */,
  {32'hc1146b9f, 32'hc03d1d20} /* (18, 30, 13) {real, imag} */,
  {32'h3f9b9b18, 32'h41068819} /* (18, 30, 12) {real, imag} */,
  {32'hc024dd75, 32'hc1b2dc6b} /* (18, 30, 11) {real, imag} */,
  {32'hbf97b9c4, 32'hc10d62d1} /* (18, 30, 10) {real, imag} */,
  {32'h408cdc66, 32'hbfcfaa3c} /* (18, 30, 9) {real, imag} */,
  {32'hc1613b0a, 32'hc158ef14} /* (18, 30, 8) {real, imag} */,
  {32'h41a1c464, 32'h41823f05} /* (18, 30, 7) {real, imag} */,
  {32'hc1330a2d, 32'hc14e353d} /* (18, 30, 6) {real, imag} */,
  {32'hc249ea44, 32'hc21c15e2} /* (18, 30, 5) {real, imag} */,
  {32'h42915d30, 32'h42a01cde} /* (18, 30, 4) {real, imag} */,
  {32'h420b143d, 32'hc1fe5615} /* (18, 30, 3) {real, imag} */,
  {32'hc4075d3a, 32'hc2e86d00} /* (18, 30, 2) {real, imag} */,
  {32'h4485513a, 32'h412712a0} /* (18, 30, 1) {real, imag} */,
  {32'h440dcf57, 32'hc2c25e41} /* (18, 30, 0) {real, imag} */,
  {32'hc2b48fa7, 32'h43260828} /* (18, 29, 31) {real, imag} */,
  {32'h42320704, 32'hc2c1a831} /* (18, 29, 30) {real, imag} */,
  {32'h41e00ead, 32'h424026d7} /* (18, 29, 29) {real, imag} */,
  {32'h41aea328, 32'hc203dfa6} /* (18, 29, 28) {real, imag} */,
  {32'hc04e3ad8, 32'hbfb32a90} /* (18, 29, 27) {real, imag} */,
  {32'h4187f5fd, 32'h40d99b5c} /* (18, 29, 26) {real, imag} */,
  {32'hc19fffc0, 32'hc1567e7a} /* (18, 29, 25) {real, imag} */,
  {32'hc19246d0, 32'h41952422} /* (18, 29, 24) {real, imag} */,
  {32'h41313a2d, 32'h40052554} /* (18, 29, 23) {real, imag} */,
  {32'h4180f45e, 32'h40d74fba} /* (18, 29, 22) {real, imag} */,
  {32'hc10973dc, 32'h405d9b4a} /* (18, 29, 21) {real, imag} */,
  {32'hc17e97ae, 32'hbfdf5a00} /* (18, 29, 20) {real, imag} */,
  {32'h40c9e798, 32'h418954a7} /* (18, 29, 19) {real, imag} */,
  {32'hc0ff1c46, 32'hbd9e5300} /* (18, 29, 18) {real, imag} */,
  {32'h40ad0e2a, 32'hc0696407} /* (18, 29, 17) {real, imag} */,
  {32'hc03bc42b, 32'h40377460} /* (18, 29, 16) {real, imag} */,
  {32'h3fcabcba, 32'h410934a2} /* (18, 29, 15) {real, imag} */,
  {32'h40432a18, 32'hc1109a89} /* (18, 29, 14) {real, imag} */,
  {32'h411cdb5d, 32'h3db19480} /* (18, 29, 13) {real, imag} */,
  {32'hc048c2fe, 32'h4158738c} /* (18, 29, 12) {real, imag} */,
  {32'h40a25c72, 32'h41b862d6} /* (18, 29, 11) {real, imag} */,
  {32'hc09011e6, 32'h41d9080b} /* (18, 29, 10) {real, imag} */,
  {32'h40bd12dc, 32'hc0977c17} /* (18, 29, 9) {real, imag} */,
  {32'h41aa120c, 32'h40593a4e} /* (18, 29, 8) {real, imag} */,
  {32'hc10b909a, 32'hc18302ce} /* (18, 29, 7) {real, imag} */,
  {32'hc1aac12a, 32'h41958560} /* (18, 29, 6) {real, imag} */,
  {32'h41d1bb1e, 32'h42170d95} /* (18, 29, 5) {real, imag} */,
  {32'hc1e4befe, 32'h3ea05de0} /* (18, 29, 4) {real, imag} */,
  {32'hc20aa8e9, 32'hc165ffcf} /* (18, 29, 3) {real, imag} */,
  {32'hc26e0f18, 32'hc3474fde} /* (18, 29, 2) {real, imag} */,
  {32'h42ca9d42, 32'h42fedc80} /* (18, 29, 1) {real, imag} */,
  {32'hbf3a5bc0, 32'h41026d97} /* (18, 29, 0) {real, imag} */,
  {32'hc2ffc6c7, 32'h42310953} /* (18, 28, 31) {real, imag} */,
  {32'h42d7928a, 32'hc267c8c7} /* (18, 28, 30) {real, imag} */,
  {32'hc01b8cb8, 32'h41818fab} /* (18, 28, 29) {real, imag} */,
  {32'h4198c316, 32'hc0865ea4} /* (18, 28, 28) {real, imag} */,
  {32'hc111795a, 32'hc1e3db25} /* (18, 28, 27) {real, imag} */,
  {32'hc1177314, 32'hc21ae2a6} /* (18, 28, 26) {real, imag} */,
  {32'hc062813a, 32'h400ff1f4} /* (18, 28, 25) {real, imag} */,
  {32'h4123e1be, 32'hc14f356b} /* (18, 28, 24) {real, imag} */,
  {32'h408f3ca8, 32'h40de4f87} /* (18, 28, 23) {real, imag} */,
  {32'h4199d7af, 32'h4190b966} /* (18, 28, 22) {real, imag} */,
  {32'h412c9bbe, 32'h3fbbda16} /* (18, 28, 21) {real, imag} */,
  {32'h406f3f67, 32'h41a31d7a} /* (18, 28, 20) {real, imag} */,
  {32'hc061f4be, 32'hc1434b59} /* (18, 28, 19) {real, imag} */,
  {32'h40081b3e, 32'hbfb0f1d0} /* (18, 28, 18) {real, imag} */,
  {32'h40b70e60, 32'h3fb275e0} /* (18, 28, 17) {real, imag} */,
  {32'hc1337658, 32'h40ad2a68} /* (18, 28, 16) {real, imag} */,
  {32'hc0815f50, 32'h3fec8440} /* (18, 28, 15) {real, imag} */,
  {32'hc0c3cd48, 32'h412c2125} /* (18, 28, 14) {real, imag} */,
  {32'hbf449070, 32'hc13d046b} /* (18, 28, 13) {real, imag} */,
  {32'h415ac598, 32'hbf80cf73} /* (18, 28, 12) {real, imag} */,
  {32'h3e2cb390, 32'h40e3109e} /* (18, 28, 11) {real, imag} */,
  {32'hc124f1a0, 32'hc18bb399} /* (18, 28, 10) {real, imag} */,
  {32'hc0df0bd2, 32'hc0e70ad4} /* (18, 28, 9) {real, imag} */,
  {32'h4074bd7e, 32'h3ee48ba8} /* (18, 28, 8) {real, imag} */,
  {32'hc086c778, 32'hc12a01ba} /* (18, 28, 7) {real, imag} */,
  {32'hc0dc34f6, 32'hc108da1c} /* (18, 28, 6) {real, imag} */,
  {32'h41baaf6e, 32'h419bf6e0} /* (18, 28, 5) {real, imag} */,
  {32'hc26caaf3, 32'h41c335ad} /* (18, 28, 4) {real, imag} */,
  {32'h403908ea, 32'h40dff103} /* (18, 28, 3) {real, imag} */,
  {32'h4185754b, 32'hc26609b9} /* (18, 28, 2) {real, imag} */,
  {32'hc2484ff7, 32'h4303b242} /* (18, 28, 1) {real, imag} */,
  {32'hc2818090, 32'h41c9ca12} /* (18, 28, 0) {real, imag} */,
  {32'h42681686, 32'hc290e72e} /* (18, 27, 31) {real, imag} */,
  {32'hc1ce6b93, 32'h4238f374} /* (18, 27, 30) {real, imag} */,
  {32'hc02d2e56, 32'hc0fe8db4} /* (18, 27, 29) {real, imag} */,
  {32'hc0725112, 32'hc18b0a0d} /* (18, 27, 28) {real, imag} */,
  {32'hc1d85a34, 32'hc11973f2} /* (18, 27, 27) {real, imag} */,
  {32'hc1aa97f4, 32'h41122791} /* (18, 27, 26) {real, imag} */,
  {32'h42151339, 32'hc1036c77} /* (18, 27, 25) {real, imag} */,
  {32'h41a26e57, 32'hc1579de6} /* (18, 27, 24) {real, imag} */,
  {32'h3e02aa08, 32'h41bec104} /* (18, 27, 23) {real, imag} */,
  {32'h4011fe8f, 32'h40a3906a} /* (18, 27, 22) {real, imag} */,
  {32'hc0ca4efa, 32'h41dc728b} /* (18, 27, 21) {real, imag} */,
  {32'h3e40e900, 32'h418f6592} /* (18, 27, 20) {real, imag} */,
  {32'h4156e875, 32'hc112d87e} /* (18, 27, 19) {real, imag} */,
  {32'h40a35792, 32'hc0e92dcb} /* (18, 27, 18) {real, imag} */,
  {32'h3f2b2268, 32'h3ef2d4d0} /* (18, 27, 17) {real, imag} */,
  {32'h40d15a50, 32'h40672d15} /* (18, 27, 16) {real, imag} */,
  {32'h3f3c89f6, 32'hc15f9d38} /* (18, 27, 15) {real, imag} */,
  {32'hc0ad566b, 32'hc1a14a7d} /* (18, 27, 14) {real, imag} */,
  {32'hc012765a, 32'h3f74d978} /* (18, 27, 13) {real, imag} */,
  {32'hc12f27a1, 32'h4049164c} /* (18, 27, 12) {real, imag} */,
  {32'hc174a2a4, 32'h4088ed37} /* (18, 27, 11) {real, imag} */,
  {32'h40f8e11f, 32'h40bc4a4f} /* (18, 27, 10) {real, imag} */,
  {32'h41331538, 32'h3fb42315} /* (18, 27, 9) {real, imag} */,
  {32'h3f126c1e, 32'h4191838e} /* (18, 27, 8) {real, imag} */,
  {32'h406cad1c, 32'hc11a1fc5} /* (18, 27, 7) {real, imag} */,
  {32'hc0a002d5, 32'hc1668fd7} /* (18, 27, 6) {real, imag} */,
  {32'h405dbc1c, 32'hc0cb5269} /* (18, 27, 5) {real, imag} */,
  {32'hc0bacc79, 32'h410a7920} /* (18, 27, 4) {real, imag} */,
  {32'h418f9346, 32'h40364c78} /* (18, 27, 3) {real, imag} */,
  {32'hc23c1b42, 32'hc17efceb} /* (18, 27, 2) {real, imag} */,
  {32'h42a9d441, 32'hc1e86370} /* (18, 27, 1) {real, imag} */,
  {32'h4226e5e7, 32'hc241347b} /* (18, 27, 0) {real, imag} */,
  {32'h4066e11c, 32'h40ffd4f3} /* (18, 26, 31) {real, imag} */,
  {32'h412298d6, 32'hc13c2be4} /* (18, 26, 30) {real, imag} */,
  {32'h40f251d8, 32'hc1121351} /* (18, 26, 29) {real, imag} */,
  {32'h408373e5, 32'hbf89fb8c} /* (18, 26, 28) {real, imag} */,
  {32'hc1702ad4, 32'hc0ef7bb1} /* (18, 26, 27) {real, imag} */,
  {32'h40fec143, 32'h41332e32} /* (18, 26, 26) {real, imag} */,
  {32'h41bf3470, 32'hc10dacb0} /* (18, 26, 25) {real, imag} */,
  {32'hc11717f0, 32'h3eae02a0} /* (18, 26, 24) {real, imag} */,
  {32'hc002bc54, 32'hc1016721} /* (18, 26, 23) {real, imag} */,
  {32'hc0ab5943, 32'hc02cfa27} /* (18, 26, 22) {real, imag} */,
  {32'hc0243448, 32'h419c3c45} /* (18, 26, 21) {real, imag} */,
  {32'h411896b4, 32'hc09ecee4} /* (18, 26, 20) {real, imag} */,
  {32'hc154feee, 32'hc0b3c034} /* (18, 26, 19) {real, imag} */,
  {32'h402e67ae, 32'hc02f15df} /* (18, 26, 18) {real, imag} */,
  {32'h4098106e, 32'hc0f758b0} /* (18, 26, 17) {real, imag} */,
  {32'h4038221c, 32'hc0cca0a8} /* (18, 26, 16) {real, imag} */,
  {32'h4015121b, 32'h403e7b92} /* (18, 26, 15) {real, imag} */,
  {32'hbfb4dcfc, 32'hc0d702ce} /* (18, 26, 14) {real, imag} */,
  {32'h40a6c33e, 32'h403c9148} /* (18, 26, 13) {real, imag} */,
  {32'h41285615, 32'hc095f74e} /* (18, 26, 12) {real, imag} */,
  {32'hbfdd5c6d, 32'h409d9944} /* (18, 26, 11) {real, imag} */,
  {32'h411a3e71, 32'hc116a9f1} /* (18, 26, 10) {real, imag} */,
  {32'h417c95d0, 32'h40ced53d} /* (18, 26, 9) {real, imag} */,
  {32'hc00431c4, 32'hbf8d5e38} /* (18, 26, 8) {real, imag} */,
  {32'hc0a7696a, 32'h4144d52e} /* (18, 26, 7) {real, imag} */,
  {32'h3f452a8c, 32'h40e64c6c} /* (18, 26, 6) {real, imag} */,
  {32'hc183ae76, 32'hc0962556} /* (18, 26, 5) {real, imag} */,
  {32'hc10bdb60, 32'hc022d910} /* (18, 26, 4) {real, imag} */,
  {32'hc1f947a8, 32'hc09bfaea} /* (18, 26, 3) {real, imag} */,
  {32'hc147e3fb, 32'h41b4bcdb} /* (18, 26, 2) {real, imag} */,
  {32'h41168407, 32'h40ca0da9} /* (18, 26, 1) {real, imag} */,
  {32'hc09ea980, 32'h41167201} /* (18, 26, 0) {real, imag} */,
  {32'hc1089c61, 32'h415efa54} /* (18, 25, 31) {real, imag} */,
  {32'h4119782c, 32'hc1cac280} /* (18, 25, 30) {real, imag} */,
  {32'h40274128, 32'hc040ae17} /* (18, 25, 29) {real, imag} */,
  {32'h41815c3c, 32'hc189f8f7} /* (18, 25, 28) {real, imag} */,
  {32'hc15e64c0, 32'h4110fce9} /* (18, 25, 27) {real, imag} */,
  {32'h41094ff2, 32'hc0337177} /* (18, 25, 26) {real, imag} */,
  {32'hc17f0cb9, 32'hc1832600} /* (18, 25, 25) {real, imag} */,
  {32'hc166ffde, 32'h41c397ce} /* (18, 25, 24) {real, imag} */,
  {32'hc196f172, 32'hc0bd4130} /* (18, 25, 23) {real, imag} */,
  {32'hc15b5c64, 32'hbeaf7600} /* (18, 25, 22) {real, imag} */,
  {32'h40adf2c6, 32'hc12fe1f8} /* (18, 25, 21) {real, imag} */,
  {32'h411c2a00, 32'hbff769c0} /* (18, 25, 20) {real, imag} */,
  {32'hc0f52dd1, 32'h406b7948} /* (18, 25, 19) {real, imag} */,
  {32'h3ec47380, 32'hc1924975} /* (18, 25, 18) {real, imag} */,
  {32'hc08cf666, 32'h40c38f80} /* (18, 25, 17) {real, imag} */,
  {32'hc06ee27a, 32'hbf8887fc} /* (18, 25, 16) {real, imag} */,
  {32'hc02f4798, 32'h4130e194} /* (18, 25, 15) {real, imag} */,
  {32'h411cc670, 32'hc1657840} /* (18, 25, 14) {real, imag} */,
  {32'hc160bc04, 32'h40354315} /* (18, 25, 13) {real, imag} */,
  {32'h40f6a654, 32'hbfff5270} /* (18, 25, 12) {real, imag} */,
  {32'hc0c61a6a, 32'hc1312c68} /* (18, 25, 11) {real, imag} */,
  {32'hc1553b6e, 32'h3fcd63ab} /* (18, 25, 10) {real, imag} */,
  {32'h41269425, 32'hc15f2b09} /* (18, 25, 9) {real, imag} */,
  {32'hbfa6c28c, 32'h40aa817a} /* (18, 25, 8) {real, imag} */,
  {32'hc1aa3959, 32'h41c0d96e} /* (18, 25, 7) {real, imag} */,
  {32'h414a1bd6, 32'h412e77c7} /* (18, 25, 6) {real, imag} */,
  {32'h4191ff38, 32'hc06129e4} /* (18, 25, 5) {real, imag} */,
  {32'h413ce270, 32'hc0d76006} /* (18, 25, 4) {real, imag} */,
  {32'hc11937b0, 32'h40e5547d} /* (18, 25, 3) {real, imag} */,
  {32'h41c26626, 32'h40572550} /* (18, 25, 2) {real, imag} */,
  {32'hc0c4742c, 32'h4193fe1e} /* (18, 25, 1) {real, imag} */,
  {32'hc1065c86, 32'h4168a097} /* (18, 25, 0) {real, imag} */,
  {32'h41a4a274, 32'hc1bbd90e} /* (18, 24, 31) {real, imag} */,
  {32'hc1ae4f33, 32'h41a79fd2} /* (18, 24, 30) {real, imag} */,
  {32'hc02844fa, 32'hbf9fa0ba} /* (18, 24, 29) {real, imag} */,
  {32'h409db65a, 32'hc01c4b41} /* (18, 24, 28) {real, imag} */,
  {32'h40095815, 32'h3fb82808} /* (18, 24, 27) {real, imag} */,
  {32'h40f23594, 32'h40b69b9d} /* (18, 24, 26) {real, imag} */,
  {32'hbf2587d0, 32'h3d417440} /* (18, 24, 25) {real, imag} */,
  {32'hc0e7807a, 32'hc1017f57} /* (18, 24, 24) {real, imag} */,
  {32'h4085f377, 32'h40a4cfda} /* (18, 24, 23) {real, imag} */,
  {32'h40b09488, 32'h4199dc28} /* (18, 24, 22) {real, imag} */,
  {32'h418360e8, 32'hbfc73e58} /* (18, 24, 21) {real, imag} */,
  {32'h4108072e, 32'hbf5ab0d0} /* (18, 24, 20) {real, imag} */,
  {32'hc13787b9, 32'h40fc9629} /* (18, 24, 19) {real, imag} */,
  {32'h4086e7fa, 32'h3ffc4b12} /* (18, 24, 18) {real, imag} */,
  {32'hc06d8e70, 32'hbf267500} /* (18, 24, 17) {real, imag} */,
  {32'hc0e93a5a, 32'hc080ea24} /* (18, 24, 16) {real, imag} */,
  {32'hc0be9580, 32'h408e6074} /* (18, 24, 15) {real, imag} */,
  {32'h40caa6c5, 32'h401e00e6} /* (18, 24, 14) {real, imag} */,
  {32'h4183e79c, 32'hc084c6cd} /* (18, 24, 13) {real, imag} */,
  {32'h411f8ebc, 32'h413f807a} /* (18, 24, 12) {real, imag} */,
  {32'hc182fa47, 32'hc0ac5295} /* (18, 24, 11) {real, imag} */,
  {32'hc1abd018, 32'hc02dbc82} /* (18, 24, 10) {real, imag} */,
  {32'hc15357be, 32'hc13dadf3} /* (18, 24, 9) {real, imag} */,
  {32'hc070c720, 32'h410e75bc} /* (18, 24, 8) {real, imag} */,
  {32'h4174a263, 32'h4121575e} /* (18, 24, 7) {real, imag} */,
  {32'hc0c28a4a, 32'h410ef21a} /* (18, 24, 6) {real, imag} */,
  {32'hc158047c, 32'h4033f9b5} /* (18, 24, 5) {real, imag} */,
  {32'h40c66a80, 32'hc19a2a99} /* (18, 24, 4) {real, imag} */,
  {32'h3f0ac2b0, 32'h40f9037a} /* (18, 24, 3) {real, imag} */,
  {32'hc21f0f48, 32'hc08cdccf} /* (18, 24, 2) {real, imag} */,
  {32'h424cb150, 32'hc20c0d71} /* (18, 24, 1) {real, imag} */,
  {32'h418bae06, 32'hc20b0557} /* (18, 24, 0) {real, imag} */,
  {32'hbf8c24c0, 32'h4142a79b} /* (18, 23, 31) {real, imag} */,
  {32'hc03f16a6, 32'hc177edee} /* (18, 23, 30) {real, imag} */,
  {32'hc0ccf12d, 32'hc0765444} /* (18, 23, 29) {real, imag} */,
  {32'h40073d34, 32'h41d3ee12} /* (18, 23, 28) {real, imag} */,
  {32'hc135dedb, 32'hc0aeca4a} /* (18, 23, 27) {real, imag} */,
  {32'h40fad470, 32'h40e7c5b1} /* (18, 23, 26) {real, imag} */,
  {32'hc1229d3d, 32'hbf007ea0} /* (18, 23, 25) {real, imag} */,
  {32'hc0f0c392, 32'h3fdada28} /* (18, 23, 24) {real, imag} */,
  {32'hc14f78c0, 32'h419289ae} /* (18, 23, 23) {real, imag} */,
  {32'h3f3a56f8, 32'hc1a8a20a} /* (18, 23, 22) {real, imag} */,
  {32'hc1e23c80, 32'hc19eb781} /* (18, 23, 21) {real, imag} */,
  {32'hc1257953, 32'h4082c6f6} /* (18, 23, 20) {real, imag} */,
  {32'h40947e26, 32'hc158895c} /* (18, 23, 19) {real, imag} */,
  {32'hc0b27778, 32'hc0021d5f} /* (18, 23, 18) {real, imag} */,
  {32'h3faf3662, 32'hc09891d4} /* (18, 23, 17) {real, imag} */,
  {32'h41709a9a, 32'h40b3cd96} /* (18, 23, 16) {real, imag} */,
  {32'h4082275e, 32'hc19f6ffe} /* (18, 23, 15) {real, imag} */,
  {32'h40cd74d0, 32'h41629c12} /* (18, 23, 14) {real, imag} */,
  {32'hc0ce54b8, 32'h4106b5ed} /* (18, 23, 13) {real, imag} */,
  {32'hc0e0aa19, 32'hc17d1e83} /* (18, 23, 12) {real, imag} */,
  {32'h413a3d79, 32'hc0ca3648} /* (18, 23, 11) {real, imag} */,
  {32'h416022a2, 32'h41b2e552} /* (18, 23, 10) {real, imag} */,
  {32'hc0dfe69c, 32'hc1a127d8} /* (18, 23, 9) {real, imag} */,
  {32'h4187a1f6, 32'h4127810c} /* (18, 23, 8) {real, imag} */,
  {32'hc14ea782, 32'hc1a8d47c} /* (18, 23, 7) {real, imag} */,
  {32'hc09638e5, 32'h41970567} /* (18, 23, 6) {real, imag} */,
  {32'h40aed934, 32'h415c8344} /* (18, 23, 5) {real, imag} */,
  {32'hc1868147, 32'h412a71f0} /* (18, 23, 4) {real, imag} */,
  {32'h418dcb36, 32'hc01c2207} /* (18, 23, 3) {real, imag} */,
  {32'hbe686ec0, 32'hc21fe30a} /* (18, 23, 2) {real, imag} */,
  {32'h40c78cdb, 32'h40dd63b0} /* (18, 23, 1) {real, imag} */,
  {32'h40db0059, 32'h40455da4} /* (18, 23, 0) {real, imag} */,
  {32'hc1915382, 32'h412a47fe} /* (18, 22, 31) {real, imag} */,
  {32'h41823b0a, 32'hc1d8cadc} /* (18, 22, 30) {real, imag} */,
  {32'hc1f8cd7c, 32'h410b0f55} /* (18, 22, 29) {real, imag} */,
  {32'hc15135be, 32'h418c9a5a} /* (18, 22, 28) {real, imag} */,
  {32'hc15c4ef8, 32'hc127c67e} /* (18, 22, 27) {real, imag} */,
  {32'hc189c652, 32'h4170b666} /* (18, 22, 26) {real, imag} */,
  {32'hbeb373b0, 32'hbe0b2b70} /* (18, 22, 25) {real, imag} */,
  {32'h40000aec, 32'hc0684340} /* (18, 22, 24) {real, imag} */,
  {32'hc09a4fbf, 32'hbf8395a0} /* (18, 22, 23) {real, imag} */,
  {32'h4089aa15, 32'hc174da06} /* (18, 22, 22) {real, imag} */,
  {32'h4184e3d5, 32'hc13afa88} /* (18, 22, 21) {real, imag} */,
  {32'h410fedc9, 32'h402b1f58} /* (18, 22, 20) {real, imag} */,
  {32'hc1567cb2, 32'hc08aca7a} /* (18, 22, 19) {real, imag} */,
  {32'h40d90ee0, 32'h41094de2} /* (18, 22, 18) {real, imag} */,
  {32'hc0b7933e, 32'h4150bcde} /* (18, 22, 17) {real, imag} */,
  {32'h3f951248, 32'hc0741b0d} /* (18, 22, 16) {real, imag} */,
  {32'hc00d049e, 32'h409d2cdc} /* (18, 22, 15) {real, imag} */,
  {32'hc005bf93, 32'h4117de0c} /* (18, 22, 14) {real, imag} */,
  {32'h404b12f6, 32'h40f9e3d5} /* (18, 22, 13) {real, imag} */,
  {32'hc0116647, 32'h40f18d64} /* (18, 22, 12) {real, imag} */,
  {32'hc08763cf, 32'h40114954} /* (18, 22, 11) {real, imag} */,
  {32'hc09e4ee4, 32'h41946131} /* (18, 22, 10) {real, imag} */,
  {32'hc10687d9, 32'hc1a81e12} /* (18, 22, 9) {real, imag} */,
  {32'hc0d0b588, 32'h3f8f53dc} /* (18, 22, 8) {real, imag} */,
  {32'hbefaac60, 32'h401c2600} /* (18, 22, 7) {real, imag} */,
  {32'h401aabf8, 32'hbff6384c} /* (18, 22, 6) {real, imag} */,
  {32'h40a71518, 32'hc03ddb87} /* (18, 22, 5) {real, imag} */,
  {32'hbffea7b0, 32'hc089e608} /* (18, 22, 4) {real, imag} */,
  {32'hc0da7cd1, 32'h4119c3af} /* (18, 22, 3) {real, imag} */,
  {32'h40e2a9d2, 32'h4154acbc} /* (18, 22, 2) {real, imag} */,
  {32'h3fa17b12, 32'hbd79db00} /* (18, 22, 1) {real, imag} */,
  {32'h41851758, 32'hbf90f790} /* (18, 22, 0) {real, imag} */,
  {32'hbf775106, 32'hc1e16006} /* (18, 21, 31) {real, imag} */,
  {32'h3fd68bd0, 32'h41401b0b} /* (18, 21, 30) {real, imag} */,
  {32'hc173c868, 32'hc1b43d52} /* (18, 21, 29) {real, imag} */,
  {32'hbfcc9dab, 32'hc18aad2d} /* (18, 21, 28) {real, imag} */,
  {32'h40665f6a, 32'h41d4a1aa} /* (18, 21, 27) {real, imag} */,
  {32'h41112699, 32'hc10ea340} /* (18, 21, 26) {real, imag} */,
  {32'h41242938, 32'h40dce20e} /* (18, 21, 25) {real, imag} */,
  {32'h41a83fa8, 32'hbfb0e27a} /* (18, 21, 24) {real, imag} */,
  {32'hc0b8f910, 32'h3e4ff0e0} /* (18, 21, 23) {real, imag} */,
  {32'h41166274, 32'h4043d304} /* (18, 21, 22) {real, imag} */,
  {32'h41b83316, 32'h40da4636} /* (18, 21, 21) {real, imag} */,
  {32'hc17453a6, 32'h40eb7c6a} /* (18, 21, 20) {real, imag} */,
  {32'hc11898c2, 32'h41202b0a} /* (18, 21, 19) {real, imag} */,
  {32'h40318192, 32'h41455b0f} /* (18, 21, 18) {real, imag} */,
  {32'hc195541a, 32'hc12a9232} /* (18, 21, 17) {real, imag} */,
  {32'hc084fb12, 32'hc0ff6a4e} /* (18, 21, 16) {real, imag} */,
  {32'h40977e5a, 32'h4033235f} /* (18, 21, 15) {real, imag} */,
  {32'h40432bd9, 32'h4046f8c0} /* (18, 21, 14) {real, imag} */,
  {32'h41411eba, 32'h407c059d} /* (18, 21, 13) {real, imag} */,
  {32'h3f24a95c, 32'h414b7288} /* (18, 21, 12) {real, imag} */,
  {32'hc1110e78, 32'h40df91bc} /* (18, 21, 11) {real, imag} */,
  {32'h41975be4, 32'hc004661f} /* (18, 21, 10) {real, imag} */,
  {32'hc1486ea6, 32'h419eb80c} /* (18, 21, 9) {real, imag} */,
  {32'hc0d67d52, 32'h4135009c} /* (18, 21, 8) {real, imag} */,
  {32'h41ceef9f, 32'h40bfd62d} /* (18, 21, 7) {real, imag} */,
  {32'h41688b53, 32'hc135c210} /* (18, 21, 6) {real, imag} */,
  {32'h40fdd55c, 32'hbf730590} /* (18, 21, 5) {real, imag} */,
  {32'h3dbe9a60, 32'hc0a240e0} /* (18, 21, 4) {real, imag} */,
  {32'hc12242b6, 32'h41670ba4} /* (18, 21, 3) {real, imag} */,
  {32'hc1654173, 32'h413051e9} /* (18, 21, 2) {real, imag} */,
  {32'h40a7949a, 32'hc032d392} /* (18, 21, 1) {real, imag} */,
  {32'h41120752, 32'hc15cedeb} /* (18, 21, 0) {real, imag} */,
  {32'hc0471fb0, 32'hc1329c2f} /* (18, 20, 31) {real, imag} */,
  {32'hc19ab664, 32'hbfc94cb4} /* (18, 20, 30) {real, imag} */,
  {32'hc08ff586, 32'h410bad8c} /* (18, 20, 29) {real, imag} */,
  {32'h401091fa, 32'h40a2173d} /* (18, 20, 28) {real, imag} */,
  {32'h4068e0ec, 32'hbee4886c} /* (18, 20, 27) {real, imag} */,
  {32'hc1262a54, 32'h403508e0} /* (18, 20, 26) {real, imag} */,
  {32'hc1024209, 32'h41aa681b} /* (18, 20, 25) {real, imag} */,
  {32'h3e65a7a0, 32'h41597184} /* (18, 20, 24) {real, imag} */,
  {32'hc0f3b0b3, 32'hc09bdef0} /* (18, 20, 23) {real, imag} */,
  {32'hbf3d1448, 32'hc037bd7e} /* (18, 20, 22) {real, imag} */,
  {32'hc0bd57c4, 32'hc0021a76} /* (18, 20, 21) {real, imag} */,
  {32'h410646c0, 32'hc1713927} /* (18, 20, 20) {real, imag} */,
  {32'h3f195ed2, 32'h406b5256} /* (18, 20, 19) {real, imag} */,
  {32'hc14c83f8, 32'h4120a826} /* (18, 20, 18) {real, imag} */,
  {32'h41332505, 32'hc09bcb72} /* (18, 20, 17) {real, imag} */,
  {32'hc0e976dd, 32'h40785484} /* (18, 20, 16) {real, imag} */,
  {32'hc0d4ca73, 32'h4062dc40} /* (18, 20, 15) {real, imag} */,
  {32'h40c24968, 32'h3e6d0740} /* (18, 20, 14) {real, imag} */,
  {32'hc143d6e6, 32'h40dff217} /* (18, 20, 13) {real, imag} */,
  {32'h41b8c16e, 32'hc08f9ed5} /* (18, 20, 12) {real, imag} */,
  {32'hc11adb9e, 32'hc119041b} /* (18, 20, 11) {real, imag} */,
  {32'hc1aa1811, 32'h40f5b4d7} /* (18, 20, 10) {real, imag} */,
  {32'hc0d8aa39, 32'hc0087955} /* (18, 20, 9) {real, imag} */,
  {32'hbf946d18, 32'hc19e2ac6} /* (18, 20, 8) {real, imag} */,
  {32'h403a321f, 32'hc0e459f0} /* (18, 20, 7) {real, imag} */,
  {32'hc114985f, 32'hc092654c} /* (18, 20, 6) {real, imag} */,
  {32'hc0711a41, 32'h40eb947e} /* (18, 20, 5) {real, imag} */,
  {32'h3feba57a, 32'h404f0cfa} /* (18, 20, 4) {real, imag} */,
  {32'h400ae748, 32'hc0f336c7} /* (18, 20, 3) {real, imag} */,
  {32'hc0f81319, 32'h40efbd08} /* (18, 20, 2) {real, imag} */,
  {32'h3ff8cbd0, 32'hc11b588f} /* (18, 20, 1) {real, imag} */,
  {32'h417bc074, 32'h4152bdb5} /* (18, 20, 0) {real, imag} */,
  {32'hc083c684, 32'hc08e70d8} /* (18, 19, 31) {real, imag} */,
  {32'h413084b8, 32'h410921ad} /* (18, 19, 30) {real, imag} */,
  {32'hc07f4f14, 32'h4131926f} /* (18, 19, 29) {real, imag} */,
  {32'hc02b3816, 32'hc122c0ce} /* (18, 19, 28) {real, imag} */,
  {32'h415f3f63, 32'h41740757} /* (18, 19, 27) {real, imag} */,
  {32'hc11c215b, 32'hc13ebe92} /* (18, 19, 26) {real, imag} */,
  {32'hc119f602, 32'h3f854184} /* (18, 19, 25) {real, imag} */,
  {32'h40d074e3, 32'h414f0f0c} /* (18, 19, 24) {real, imag} */,
  {32'hc0eb9820, 32'hc0f2172a} /* (18, 19, 23) {real, imag} */,
  {32'hc12436ca, 32'hc0c8202a} /* (18, 19, 22) {real, imag} */,
  {32'hbf332020, 32'hc0c8243f} /* (18, 19, 21) {real, imag} */,
  {32'hc0aafaee, 32'hc0d53c9d} /* (18, 19, 20) {real, imag} */,
  {32'h41275bd6, 32'h40941bd3} /* (18, 19, 19) {real, imag} */,
  {32'hc1113be8, 32'h3fae6a68} /* (18, 19, 18) {real, imag} */,
  {32'h406fe730, 32'hc001d07a} /* (18, 19, 17) {real, imag} */,
  {32'h40993c56, 32'hc0c86cae} /* (18, 19, 16) {real, imag} */,
  {32'h40a69095, 32'hc081ee48} /* (18, 19, 15) {real, imag} */,
  {32'h41aafe95, 32'hc0ce76b1} /* (18, 19, 14) {real, imag} */,
  {32'h41cf8df6, 32'h3f846b88} /* (18, 19, 13) {real, imag} */,
  {32'h4192a5e3, 32'hbfe2fe00} /* (18, 19, 12) {real, imag} */,
  {32'h4032cf65, 32'h404e84bc} /* (18, 19, 11) {real, imag} */,
  {32'h416394e4, 32'hc12617c9} /* (18, 19, 10) {real, imag} */,
  {32'h417cd9a4, 32'h4110f20f} /* (18, 19, 9) {real, imag} */,
  {32'h4020dfe9, 32'h4152fd32} /* (18, 19, 8) {real, imag} */,
  {32'hbfd60818, 32'h405782c8} /* (18, 19, 7) {real, imag} */,
  {32'hc1dca231, 32'h410aa398} /* (18, 19, 6) {real, imag} */,
  {32'hc0c95cec, 32'h414dfaf8} /* (18, 19, 5) {real, imag} */,
  {32'hc103f294, 32'hbfa0c7d2} /* (18, 19, 4) {real, imag} */,
  {32'h4010c27f, 32'hbf8a0c3e} /* (18, 19, 3) {real, imag} */,
  {32'h4033000b, 32'hc1a8271a} /* (18, 19, 2) {real, imag} */,
  {32'h40f85c80, 32'h3dd9b580} /* (18, 19, 1) {real, imag} */,
  {32'h3f823ba0, 32'h40e707f2} /* (18, 19, 0) {real, imag} */,
  {32'hc1114320, 32'hc08db4d8} /* (18, 18, 31) {real, imag} */,
  {32'h402740c4, 32'h40bfd1aa} /* (18, 18, 30) {real, imag} */,
  {32'hbf197858, 32'hc0daba38} /* (18, 18, 29) {real, imag} */,
  {32'h4095b7ab, 32'hc16a5468} /* (18, 18, 28) {real, imag} */,
  {32'hc0d47126, 32'hc02b1363} /* (18, 18, 27) {real, imag} */,
  {32'h3f6de2a0, 32'h41102074} /* (18, 18, 26) {real, imag} */,
  {32'hbf5527f8, 32'hbb87a800} /* (18, 18, 25) {real, imag} */,
  {32'hc0103bba, 32'hbf571880} /* (18, 18, 24) {real, imag} */,
  {32'hc0747b00, 32'h40f27f1e} /* (18, 18, 23) {real, imag} */,
  {32'hc0546084, 32'hc1410882} /* (18, 18, 22) {real, imag} */,
  {32'h403b5c68, 32'hc0b28fdc} /* (18, 18, 21) {real, imag} */,
  {32'h408c9a88, 32'h411b8521} /* (18, 18, 20) {real, imag} */,
  {32'h412f04f0, 32'hc08fe660} /* (18, 18, 19) {real, imag} */,
  {32'hc07cbbf8, 32'h41548273} /* (18, 18, 18) {real, imag} */,
  {32'hbfdd1d06, 32'hc0549b76} /* (18, 18, 17) {real, imag} */,
  {32'hc0afcc62, 32'hbefc52a0} /* (18, 18, 16) {real, imag} */,
  {32'h409c0bea, 32'h3e89dd08} /* (18, 18, 15) {real, imag} */,
  {32'h40993e0e, 32'hbfda3282} /* (18, 18, 14) {real, imag} */,
  {32'h417118d8, 32'hc12488ee} /* (18, 18, 13) {real, imag} */,
  {32'hbdee5fa0, 32'h418146bb} /* (18, 18, 12) {real, imag} */,
  {32'hbfb7d1c4, 32'h41b0feae} /* (18, 18, 11) {real, imag} */,
  {32'h40cbe98c, 32'h401e1ef2} /* (18, 18, 10) {real, imag} */,
  {32'hbf176348, 32'hc114b996} /* (18, 18, 9) {real, imag} */,
  {32'h3fbf8f1c, 32'h414a5870} /* (18, 18, 8) {real, imag} */,
  {32'hc169c87e, 32'h3e89d020} /* (18, 18, 7) {real, imag} */,
  {32'hc141ed54, 32'hbf323ae6} /* (18, 18, 6) {real, imag} */,
  {32'hc0cc7bb3, 32'h413a3adc} /* (18, 18, 5) {real, imag} */,
  {32'hc0c818e0, 32'hc0d83ee0} /* (18, 18, 4) {real, imag} */,
  {32'h410229c5, 32'hbf85c548} /* (18, 18, 3) {real, imag} */,
  {32'hc05b84a6, 32'h4097f9b6} /* (18, 18, 2) {real, imag} */,
  {32'h40f468b1, 32'hc14f1a22} /* (18, 18, 1) {real, imag} */,
  {32'h41572fe8, 32'hc12fd0ac} /* (18, 18, 0) {real, imag} */,
  {32'hc010ab79, 32'h41847832} /* (18, 17, 31) {real, imag} */,
  {32'hc0018330, 32'h40d37c10} /* (18, 17, 30) {real, imag} */,
  {32'hc0df6b56, 32'hbf9f5236} /* (18, 17, 29) {real, imag} */,
  {32'hbfa438ee, 32'h4039b613} /* (18, 17, 28) {real, imag} */,
  {32'h40f77f08, 32'hc16bef3c} /* (18, 17, 27) {real, imag} */,
  {32'hbfa89141, 32'h40875d0a} /* (18, 17, 26) {real, imag} */,
  {32'h4131ab08, 32'hbeba9880} /* (18, 17, 25) {real, imag} */,
  {32'h409d44fa, 32'hc185dc2f} /* (18, 17, 24) {real, imag} */,
  {32'h408a41d4, 32'h3f8c85e4} /* (18, 17, 23) {real, imag} */,
  {32'hbfc317b0, 32'hc14b2fed} /* (18, 17, 22) {real, imag} */,
  {32'hc0cb8611, 32'h402b6fa6} /* (18, 17, 21) {real, imag} */,
  {32'h41113122, 32'hbd95dac0} /* (18, 17, 20) {real, imag} */,
  {32'hbf8f7988, 32'h41215de0} /* (18, 17, 19) {real, imag} */,
  {32'h3f181a3a, 32'h411b3cef} /* (18, 17, 18) {real, imag} */,
  {32'h3f84c8a2, 32'h40c35e68} /* (18, 17, 17) {real, imag} */,
  {32'hbe633367, 32'hc0a36c66} /* (18, 17, 16) {real, imag} */,
  {32'hc08d5c5a, 32'h4056d4d2} /* (18, 17, 15) {real, imag} */,
  {32'h40fe5e06, 32'h40c747d7} /* (18, 17, 14) {real, imag} */,
  {32'h414ca010, 32'hc10f3f06} /* (18, 17, 13) {real, imag} */,
  {32'hc1240fc0, 32'h410b41c7} /* (18, 17, 12) {real, imag} */,
  {32'h4028f351, 32'hc0558d10} /* (18, 17, 11) {real, imag} */,
  {32'h413f876f, 32'hbf5a6edc} /* (18, 17, 10) {real, imag} */,
  {32'h4162d4c5, 32'h3fd1513c} /* (18, 17, 9) {real, imag} */,
  {32'hc015a1db, 32'h40641724} /* (18, 17, 8) {real, imag} */,
  {32'hc0bf6779, 32'hc10c2d3c} /* (18, 17, 7) {real, imag} */,
  {32'hc0f8e602, 32'hc098da7c} /* (18, 17, 6) {real, imag} */,
  {32'h3fb6a354, 32'hc0d30de6} /* (18, 17, 5) {real, imag} */,
  {32'h3f52481e, 32'hc0ba9d16} /* (18, 17, 4) {real, imag} */,
  {32'hc04f0e2a, 32'hc0a95ce9} /* (18, 17, 3) {real, imag} */,
  {32'h3f631588, 32'h3f828b10} /* (18, 17, 2) {real, imag} */,
  {32'hc07217f4, 32'hbf9854ee} /* (18, 17, 1) {real, imag} */,
  {32'h4089569a, 32'h3f4ed984} /* (18, 17, 0) {real, imag} */,
  {32'hc01f8ef4, 32'h409d9620} /* (18, 16, 31) {real, imag} */,
  {32'hc106bc9f, 32'hc0e2ce3a} /* (18, 16, 30) {real, imag} */,
  {32'hbe848458, 32'hc0247f48} /* (18, 16, 29) {real, imag} */,
  {32'h4161b9ed, 32'h40e4aa08} /* (18, 16, 28) {real, imag} */,
  {32'h401608c0, 32'h4092739a} /* (18, 16, 27) {real, imag} */,
  {32'hc0a5423e, 32'hc11d1af2} /* (18, 16, 26) {real, imag} */,
  {32'hbfaa88e6, 32'hc1523414} /* (18, 16, 25) {real, imag} */,
  {32'hbf3464c8, 32'h3fec91d0} /* (18, 16, 24) {real, imag} */,
  {32'h4036db4e, 32'h409fccb9} /* (18, 16, 23) {real, imag} */,
  {32'hc081086b, 32'h411766cc} /* (18, 16, 22) {real, imag} */,
  {32'h3ff01a48, 32'hc0dd3282} /* (18, 16, 21) {real, imag} */,
  {32'h3fda77be, 32'h40e240a3} /* (18, 16, 20) {real, imag} */,
  {32'h40c0f6eb, 32'h3f8cc7a8} /* (18, 16, 19) {real, imag} */,
  {32'hc02c5b1f, 32'h3ed52300} /* (18, 16, 18) {real, imag} */,
  {32'hc0015bff, 32'hc0c456f6} /* (18, 16, 17) {real, imag} */,
  {32'hc1361599, 32'h00000000} /* (18, 16, 16) {real, imag} */,
  {32'hc0015bff, 32'h40c456f6} /* (18, 16, 15) {real, imag} */,
  {32'hc02c5b1f, 32'hbed52300} /* (18, 16, 14) {real, imag} */,
  {32'h40c0f6eb, 32'hbf8cc7a8} /* (18, 16, 13) {real, imag} */,
  {32'h3fda77be, 32'hc0e240a3} /* (18, 16, 12) {real, imag} */,
  {32'h3ff01a48, 32'h40dd3282} /* (18, 16, 11) {real, imag} */,
  {32'hc081086b, 32'hc11766cc} /* (18, 16, 10) {real, imag} */,
  {32'h4036db4e, 32'hc09fccb9} /* (18, 16, 9) {real, imag} */,
  {32'hbf3464c8, 32'hbfec91d0} /* (18, 16, 8) {real, imag} */,
  {32'hbfaa88e6, 32'h41523414} /* (18, 16, 7) {real, imag} */,
  {32'hc0a5423e, 32'h411d1af2} /* (18, 16, 6) {real, imag} */,
  {32'h401608c0, 32'hc092739a} /* (18, 16, 5) {real, imag} */,
  {32'h4161b9ed, 32'hc0e4aa08} /* (18, 16, 4) {real, imag} */,
  {32'hbe848458, 32'h40247f48} /* (18, 16, 3) {real, imag} */,
  {32'hc106bc9f, 32'h40e2ce3a} /* (18, 16, 2) {real, imag} */,
  {32'hc01f8ef4, 32'hc09d9620} /* (18, 16, 1) {real, imag} */,
  {32'hc0090c88, 32'h00000000} /* (18, 16, 0) {real, imag} */,
  {32'hc07217f4, 32'h3f9854ee} /* (18, 15, 31) {real, imag} */,
  {32'h3f631588, 32'hbf828b10} /* (18, 15, 30) {real, imag} */,
  {32'hc04f0e2a, 32'h40a95ce9} /* (18, 15, 29) {real, imag} */,
  {32'h3f52481e, 32'h40ba9d16} /* (18, 15, 28) {real, imag} */,
  {32'h3fb6a354, 32'h40d30de6} /* (18, 15, 27) {real, imag} */,
  {32'hc0f8e602, 32'h4098da7c} /* (18, 15, 26) {real, imag} */,
  {32'hc0bf6779, 32'h410c2d3c} /* (18, 15, 25) {real, imag} */,
  {32'hc015a1db, 32'hc0641724} /* (18, 15, 24) {real, imag} */,
  {32'h4162d4c5, 32'hbfd1513c} /* (18, 15, 23) {real, imag} */,
  {32'h413f876f, 32'h3f5a6edc} /* (18, 15, 22) {real, imag} */,
  {32'h4028f351, 32'h40558d10} /* (18, 15, 21) {real, imag} */,
  {32'hc1240fc0, 32'hc10b41c7} /* (18, 15, 20) {real, imag} */,
  {32'h414ca010, 32'h410f3f06} /* (18, 15, 19) {real, imag} */,
  {32'h40fe5e06, 32'hc0c747d7} /* (18, 15, 18) {real, imag} */,
  {32'hc08d5c5a, 32'hc056d4d2} /* (18, 15, 17) {real, imag} */,
  {32'hbe633367, 32'h40a36c66} /* (18, 15, 16) {real, imag} */,
  {32'h3f84c8a2, 32'hc0c35e68} /* (18, 15, 15) {real, imag} */,
  {32'h3f181a3a, 32'hc11b3cef} /* (18, 15, 14) {real, imag} */,
  {32'hbf8f7988, 32'hc1215de0} /* (18, 15, 13) {real, imag} */,
  {32'h41113122, 32'h3d95dac0} /* (18, 15, 12) {real, imag} */,
  {32'hc0cb8611, 32'hc02b6fa6} /* (18, 15, 11) {real, imag} */,
  {32'hbfc317b0, 32'h414b2fed} /* (18, 15, 10) {real, imag} */,
  {32'h408a41d4, 32'hbf8c85e4} /* (18, 15, 9) {real, imag} */,
  {32'h409d44fa, 32'h4185dc2f} /* (18, 15, 8) {real, imag} */,
  {32'h4131ab08, 32'h3eba9880} /* (18, 15, 7) {real, imag} */,
  {32'hbfa89141, 32'hc0875d0a} /* (18, 15, 6) {real, imag} */,
  {32'h40f77f08, 32'h416bef3c} /* (18, 15, 5) {real, imag} */,
  {32'hbfa438ee, 32'hc039b613} /* (18, 15, 4) {real, imag} */,
  {32'hc0df6b56, 32'h3f9f5236} /* (18, 15, 3) {real, imag} */,
  {32'hc0018330, 32'hc0d37c10} /* (18, 15, 2) {real, imag} */,
  {32'hc010ab79, 32'hc1847832} /* (18, 15, 1) {real, imag} */,
  {32'h4089569a, 32'hbf4ed984} /* (18, 15, 0) {real, imag} */,
  {32'h40f468b1, 32'h414f1a22} /* (18, 14, 31) {real, imag} */,
  {32'hc05b84a6, 32'hc097f9b6} /* (18, 14, 30) {real, imag} */,
  {32'h410229c5, 32'h3f85c548} /* (18, 14, 29) {real, imag} */,
  {32'hc0c818e0, 32'h40d83ee0} /* (18, 14, 28) {real, imag} */,
  {32'hc0cc7bb3, 32'hc13a3adc} /* (18, 14, 27) {real, imag} */,
  {32'hc141ed54, 32'h3f323ae6} /* (18, 14, 26) {real, imag} */,
  {32'hc169c87e, 32'hbe89d020} /* (18, 14, 25) {real, imag} */,
  {32'h3fbf8f1c, 32'hc14a5870} /* (18, 14, 24) {real, imag} */,
  {32'hbf176348, 32'h4114b996} /* (18, 14, 23) {real, imag} */,
  {32'h40cbe98c, 32'hc01e1ef2} /* (18, 14, 22) {real, imag} */,
  {32'hbfb7d1c4, 32'hc1b0feae} /* (18, 14, 21) {real, imag} */,
  {32'hbdee5fa0, 32'hc18146bb} /* (18, 14, 20) {real, imag} */,
  {32'h417118d8, 32'h412488ee} /* (18, 14, 19) {real, imag} */,
  {32'h40993e0e, 32'h3fda3282} /* (18, 14, 18) {real, imag} */,
  {32'h409c0bea, 32'hbe89dd08} /* (18, 14, 17) {real, imag} */,
  {32'hc0afcc62, 32'h3efc52a0} /* (18, 14, 16) {real, imag} */,
  {32'hbfdd1d06, 32'h40549b76} /* (18, 14, 15) {real, imag} */,
  {32'hc07cbbf8, 32'hc1548273} /* (18, 14, 14) {real, imag} */,
  {32'h412f04f0, 32'h408fe660} /* (18, 14, 13) {real, imag} */,
  {32'h408c9a88, 32'hc11b8521} /* (18, 14, 12) {real, imag} */,
  {32'h403b5c68, 32'h40b28fdc} /* (18, 14, 11) {real, imag} */,
  {32'hc0546084, 32'h41410882} /* (18, 14, 10) {real, imag} */,
  {32'hc0747b00, 32'hc0f27f1e} /* (18, 14, 9) {real, imag} */,
  {32'hc0103bba, 32'h3f571880} /* (18, 14, 8) {real, imag} */,
  {32'hbf5527f8, 32'h3b87a800} /* (18, 14, 7) {real, imag} */,
  {32'h3f6de2a0, 32'hc1102074} /* (18, 14, 6) {real, imag} */,
  {32'hc0d47126, 32'h402b1363} /* (18, 14, 5) {real, imag} */,
  {32'h4095b7ab, 32'h416a5468} /* (18, 14, 4) {real, imag} */,
  {32'hbf197858, 32'h40daba38} /* (18, 14, 3) {real, imag} */,
  {32'h402740c4, 32'hc0bfd1aa} /* (18, 14, 2) {real, imag} */,
  {32'hc1114320, 32'h408db4d8} /* (18, 14, 1) {real, imag} */,
  {32'h41572fe8, 32'h412fd0ac} /* (18, 14, 0) {real, imag} */,
  {32'h40f85c80, 32'hbdd9b580} /* (18, 13, 31) {real, imag} */,
  {32'h4033000b, 32'h41a8271a} /* (18, 13, 30) {real, imag} */,
  {32'h4010c27f, 32'h3f8a0c3e} /* (18, 13, 29) {real, imag} */,
  {32'hc103f294, 32'h3fa0c7d2} /* (18, 13, 28) {real, imag} */,
  {32'hc0c95cec, 32'hc14dfaf8} /* (18, 13, 27) {real, imag} */,
  {32'hc1dca231, 32'hc10aa398} /* (18, 13, 26) {real, imag} */,
  {32'hbfd60818, 32'hc05782c8} /* (18, 13, 25) {real, imag} */,
  {32'h4020dfe9, 32'hc152fd32} /* (18, 13, 24) {real, imag} */,
  {32'h417cd9a4, 32'hc110f20f} /* (18, 13, 23) {real, imag} */,
  {32'h416394e4, 32'h412617c9} /* (18, 13, 22) {real, imag} */,
  {32'h4032cf65, 32'hc04e84bc} /* (18, 13, 21) {real, imag} */,
  {32'h4192a5e3, 32'h3fe2fe00} /* (18, 13, 20) {real, imag} */,
  {32'h41cf8df6, 32'hbf846b88} /* (18, 13, 19) {real, imag} */,
  {32'h41aafe95, 32'h40ce76b1} /* (18, 13, 18) {real, imag} */,
  {32'h40a69095, 32'h4081ee48} /* (18, 13, 17) {real, imag} */,
  {32'h40993c56, 32'h40c86cae} /* (18, 13, 16) {real, imag} */,
  {32'h406fe730, 32'h4001d07a} /* (18, 13, 15) {real, imag} */,
  {32'hc1113be8, 32'hbfae6a68} /* (18, 13, 14) {real, imag} */,
  {32'h41275bd6, 32'hc0941bd3} /* (18, 13, 13) {real, imag} */,
  {32'hc0aafaee, 32'h40d53c9d} /* (18, 13, 12) {real, imag} */,
  {32'hbf332020, 32'h40c8243f} /* (18, 13, 11) {real, imag} */,
  {32'hc12436ca, 32'h40c8202a} /* (18, 13, 10) {real, imag} */,
  {32'hc0eb9820, 32'h40f2172a} /* (18, 13, 9) {real, imag} */,
  {32'h40d074e3, 32'hc14f0f0c} /* (18, 13, 8) {real, imag} */,
  {32'hc119f602, 32'hbf854184} /* (18, 13, 7) {real, imag} */,
  {32'hc11c215b, 32'h413ebe92} /* (18, 13, 6) {real, imag} */,
  {32'h415f3f63, 32'hc1740757} /* (18, 13, 5) {real, imag} */,
  {32'hc02b3816, 32'h4122c0ce} /* (18, 13, 4) {real, imag} */,
  {32'hc07f4f14, 32'hc131926f} /* (18, 13, 3) {real, imag} */,
  {32'h413084b8, 32'hc10921ad} /* (18, 13, 2) {real, imag} */,
  {32'hc083c684, 32'h408e70d8} /* (18, 13, 1) {real, imag} */,
  {32'h3f823ba0, 32'hc0e707f2} /* (18, 13, 0) {real, imag} */,
  {32'h3ff8cbd0, 32'h411b588f} /* (18, 12, 31) {real, imag} */,
  {32'hc0f81319, 32'hc0efbd08} /* (18, 12, 30) {real, imag} */,
  {32'h400ae748, 32'h40f336c7} /* (18, 12, 29) {real, imag} */,
  {32'h3feba57a, 32'hc04f0cfa} /* (18, 12, 28) {real, imag} */,
  {32'hc0711a41, 32'hc0eb947e} /* (18, 12, 27) {real, imag} */,
  {32'hc114985f, 32'h4092654c} /* (18, 12, 26) {real, imag} */,
  {32'h403a321f, 32'h40e459f0} /* (18, 12, 25) {real, imag} */,
  {32'hbf946d18, 32'h419e2ac6} /* (18, 12, 24) {real, imag} */,
  {32'hc0d8aa39, 32'h40087955} /* (18, 12, 23) {real, imag} */,
  {32'hc1aa1811, 32'hc0f5b4d7} /* (18, 12, 22) {real, imag} */,
  {32'hc11adb9e, 32'h4119041b} /* (18, 12, 21) {real, imag} */,
  {32'h41b8c16e, 32'h408f9ed5} /* (18, 12, 20) {real, imag} */,
  {32'hc143d6e6, 32'hc0dff217} /* (18, 12, 19) {real, imag} */,
  {32'h40c24968, 32'hbe6d0740} /* (18, 12, 18) {real, imag} */,
  {32'hc0d4ca73, 32'hc062dc40} /* (18, 12, 17) {real, imag} */,
  {32'hc0e976dd, 32'hc0785484} /* (18, 12, 16) {real, imag} */,
  {32'h41332505, 32'h409bcb72} /* (18, 12, 15) {real, imag} */,
  {32'hc14c83f8, 32'hc120a826} /* (18, 12, 14) {real, imag} */,
  {32'h3f195ed2, 32'hc06b5256} /* (18, 12, 13) {real, imag} */,
  {32'h410646c0, 32'h41713927} /* (18, 12, 12) {real, imag} */,
  {32'hc0bd57c4, 32'h40021a76} /* (18, 12, 11) {real, imag} */,
  {32'hbf3d1448, 32'h4037bd7e} /* (18, 12, 10) {real, imag} */,
  {32'hc0f3b0b3, 32'h409bdef0} /* (18, 12, 9) {real, imag} */,
  {32'h3e65a7a0, 32'hc1597184} /* (18, 12, 8) {real, imag} */,
  {32'hc1024209, 32'hc1aa681b} /* (18, 12, 7) {real, imag} */,
  {32'hc1262a54, 32'hc03508e0} /* (18, 12, 6) {real, imag} */,
  {32'h4068e0ec, 32'h3ee4886c} /* (18, 12, 5) {real, imag} */,
  {32'h401091fa, 32'hc0a2173d} /* (18, 12, 4) {real, imag} */,
  {32'hc08ff586, 32'hc10bad8c} /* (18, 12, 3) {real, imag} */,
  {32'hc19ab664, 32'h3fc94cb4} /* (18, 12, 2) {real, imag} */,
  {32'hc0471fb0, 32'h41329c2f} /* (18, 12, 1) {real, imag} */,
  {32'h417bc074, 32'hc152bdb5} /* (18, 12, 0) {real, imag} */,
  {32'h40a7949a, 32'h4032d392} /* (18, 11, 31) {real, imag} */,
  {32'hc1654173, 32'hc13051e9} /* (18, 11, 30) {real, imag} */,
  {32'hc12242b6, 32'hc1670ba4} /* (18, 11, 29) {real, imag} */,
  {32'h3dbe9a60, 32'h40a240e0} /* (18, 11, 28) {real, imag} */,
  {32'h40fdd55c, 32'h3f730590} /* (18, 11, 27) {real, imag} */,
  {32'h41688b53, 32'h4135c210} /* (18, 11, 26) {real, imag} */,
  {32'h41ceef9f, 32'hc0bfd62d} /* (18, 11, 25) {real, imag} */,
  {32'hc0d67d52, 32'hc135009c} /* (18, 11, 24) {real, imag} */,
  {32'hc1486ea6, 32'hc19eb80c} /* (18, 11, 23) {real, imag} */,
  {32'h41975be4, 32'h4004661f} /* (18, 11, 22) {real, imag} */,
  {32'hc1110e78, 32'hc0df91bc} /* (18, 11, 21) {real, imag} */,
  {32'h3f24a95c, 32'hc14b7288} /* (18, 11, 20) {real, imag} */,
  {32'h41411eba, 32'hc07c059d} /* (18, 11, 19) {real, imag} */,
  {32'h40432bd9, 32'hc046f8c0} /* (18, 11, 18) {real, imag} */,
  {32'h40977e5a, 32'hc033235f} /* (18, 11, 17) {real, imag} */,
  {32'hc084fb12, 32'h40ff6a4e} /* (18, 11, 16) {real, imag} */,
  {32'hc195541a, 32'h412a9232} /* (18, 11, 15) {real, imag} */,
  {32'h40318192, 32'hc1455b0f} /* (18, 11, 14) {real, imag} */,
  {32'hc11898c2, 32'hc1202b0a} /* (18, 11, 13) {real, imag} */,
  {32'hc17453a6, 32'hc0eb7c6a} /* (18, 11, 12) {real, imag} */,
  {32'h41b83316, 32'hc0da4636} /* (18, 11, 11) {real, imag} */,
  {32'h41166274, 32'hc043d304} /* (18, 11, 10) {real, imag} */,
  {32'hc0b8f910, 32'hbe4ff0e0} /* (18, 11, 9) {real, imag} */,
  {32'h41a83fa8, 32'h3fb0e27a} /* (18, 11, 8) {real, imag} */,
  {32'h41242938, 32'hc0dce20e} /* (18, 11, 7) {real, imag} */,
  {32'h41112699, 32'h410ea340} /* (18, 11, 6) {real, imag} */,
  {32'h40665f6a, 32'hc1d4a1aa} /* (18, 11, 5) {real, imag} */,
  {32'hbfcc9dab, 32'h418aad2d} /* (18, 11, 4) {real, imag} */,
  {32'hc173c868, 32'h41b43d52} /* (18, 11, 3) {real, imag} */,
  {32'h3fd68bd0, 32'hc1401b0b} /* (18, 11, 2) {real, imag} */,
  {32'hbf775106, 32'h41e16006} /* (18, 11, 1) {real, imag} */,
  {32'h41120752, 32'h415cedeb} /* (18, 11, 0) {real, imag} */,
  {32'h3fa17b12, 32'h3d79db00} /* (18, 10, 31) {real, imag} */,
  {32'h40e2a9d2, 32'hc154acbc} /* (18, 10, 30) {real, imag} */,
  {32'hc0da7cd1, 32'hc119c3af} /* (18, 10, 29) {real, imag} */,
  {32'hbffea7b0, 32'h4089e608} /* (18, 10, 28) {real, imag} */,
  {32'h40a71518, 32'h403ddb87} /* (18, 10, 27) {real, imag} */,
  {32'h401aabf8, 32'h3ff6384c} /* (18, 10, 26) {real, imag} */,
  {32'hbefaac60, 32'hc01c2600} /* (18, 10, 25) {real, imag} */,
  {32'hc0d0b588, 32'hbf8f53dc} /* (18, 10, 24) {real, imag} */,
  {32'hc10687d9, 32'h41a81e12} /* (18, 10, 23) {real, imag} */,
  {32'hc09e4ee4, 32'hc1946131} /* (18, 10, 22) {real, imag} */,
  {32'hc08763cf, 32'hc0114954} /* (18, 10, 21) {real, imag} */,
  {32'hc0116647, 32'hc0f18d64} /* (18, 10, 20) {real, imag} */,
  {32'h404b12f6, 32'hc0f9e3d5} /* (18, 10, 19) {real, imag} */,
  {32'hc005bf93, 32'hc117de0c} /* (18, 10, 18) {real, imag} */,
  {32'hc00d049e, 32'hc09d2cdc} /* (18, 10, 17) {real, imag} */,
  {32'h3f951248, 32'h40741b0d} /* (18, 10, 16) {real, imag} */,
  {32'hc0b7933e, 32'hc150bcde} /* (18, 10, 15) {real, imag} */,
  {32'h40d90ee0, 32'hc1094de2} /* (18, 10, 14) {real, imag} */,
  {32'hc1567cb2, 32'h408aca7a} /* (18, 10, 13) {real, imag} */,
  {32'h410fedc9, 32'hc02b1f58} /* (18, 10, 12) {real, imag} */,
  {32'h4184e3d5, 32'h413afa88} /* (18, 10, 11) {real, imag} */,
  {32'h4089aa15, 32'h4174da06} /* (18, 10, 10) {real, imag} */,
  {32'hc09a4fbf, 32'h3f8395a0} /* (18, 10, 9) {real, imag} */,
  {32'h40000aec, 32'h40684340} /* (18, 10, 8) {real, imag} */,
  {32'hbeb373b0, 32'h3e0b2b70} /* (18, 10, 7) {real, imag} */,
  {32'hc189c652, 32'hc170b666} /* (18, 10, 6) {real, imag} */,
  {32'hc15c4ef8, 32'h4127c67e} /* (18, 10, 5) {real, imag} */,
  {32'hc15135be, 32'hc18c9a5a} /* (18, 10, 4) {real, imag} */,
  {32'hc1f8cd7c, 32'hc10b0f55} /* (18, 10, 3) {real, imag} */,
  {32'h41823b0a, 32'h41d8cadc} /* (18, 10, 2) {real, imag} */,
  {32'hc1915382, 32'hc12a47fe} /* (18, 10, 1) {real, imag} */,
  {32'h41851758, 32'h3f90f790} /* (18, 10, 0) {real, imag} */,
  {32'h40c78cdb, 32'hc0dd63b0} /* (18, 9, 31) {real, imag} */,
  {32'hbe686ec0, 32'h421fe30a} /* (18, 9, 30) {real, imag} */,
  {32'h418dcb36, 32'h401c2207} /* (18, 9, 29) {real, imag} */,
  {32'hc1868147, 32'hc12a71f0} /* (18, 9, 28) {real, imag} */,
  {32'h40aed934, 32'hc15c8344} /* (18, 9, 27) {real, imag} */,
  {32'hc09638e5, 32'hc1970567} /* (18, 9, 26) {real, imag} */,
  {32'hc14ea782, 32'h41a8d47c} /* (18, 9, 25) {real, imag} */,
  {32'h4187a1f6, 32'hc127810c} /* (18, 9, 24) {real, imag} */,
  {32'hc0dfe69c, 32'h41a127d8} /* (18, 9, 23) {real, imag} */,
  {32'h416022a2, 32'hc1b2e552} /* (18, 9, 22) {real, imag} */,
  {32'h413a3d79, 32'h40ca3648} /* (18, 9, 21) {real, imag} */,
  {32'hc0e0aa19, 32'h417d1e83} /* (18, 9, 20) {real, imag} */,
  {32'hc0ce54b8, 32'hc106b5ed} /* (18, 9, 19) {real, imag} */,
  {32'h40cd74d0, 32'hc1629c12} /* (18, 9, 18) {real, imag} */,
  {32'h4082275e, 32'h419f6ffe} /* (18, 9, 17) {real, imag} */,
  {32'h41709a9a, 32'hc0b3cd96} /* (18, 9, 16) {real, imag} */,
  {32'h3faf3662, 32'h409891d4} /* (18, 9, 15) {real, imag} */,
  {32'hc0b27778, 32'h40021d5f} /* (18, 9, 14) {real, imag} */,
  {32'h40947e26, 32'h4158895c} /* (18, 9, 13) {real, imag} */,
  {32'hc1257953, 32'hc082c6f6} /* (18, 9, 12) {real, imag} */,
  {32'hc1e23c80, 32'h419eb781} /* (18, 9, 11) {real, imag} */,
  {32'h3f3a56f8, 32'h41a8a20a} /* (18, 9, 10) {real, imag} */,
  {32'hc14f78c0, 32'hc19289ae} /* (18, 9, 9) {real, imag} */,
  {32'hc0f0c392, 32'hbfdada28} /* (18, 9, 8) {real, imag} */,
  {32'hc1229d3d, 32'h3f007ea0} /* (18, 9, 7) {real, imag} */,
  {32'h40fad470, 32'hc0e7c5b1} /* (18, 9, 6) {real, imag} */,
  {32'hc135dedb, 32'h40aeca4a} /* (18, 9, 5) {real, imag} */,
  {32'h40073d34, 32'hc1d3ee12} /* (18, 9, 4) {real, imag} */,
  {32'hc0ccf12d, 32'h40765444} /* (18, 9, 3) {real, imag} */,
  {32'hc03f16a6, 32'h4177edee} /* (18, 9, 2) {real, imag} */,
  {32'hbf8c24c0, 32'hc142a79b} /* (18, 9, 1) {real, imag} */,
  {32'h40db0059, 32'hc0455da4} /* (18, 9, 0) {real, imag} */,
  {32'h424cb150, 32'h420c0d71} /* (18, 8, 31) {real, imag} */,
  {32'hc21f0f48, 32'h408cdccf} /* (18, 8, 30) {real, imag} */,
  {32'h3f0ac2b0, 32'hc0f9037a} /* (18, 8, 29) {real, imag} */,
  {32'h40c66a80, 32'h419a2a99} /* (18, 8, 28) {real, imag} */,
  {32'hc158047c, 32'hc033f9b5} /* (18, 8, 27) {real, imag} */,
  {32'hc0c28a4a, 32'hc10ef21a} /* (18, 8, 26) {real, imag} */,
  {32'h4174a263, 32'hc121575e} /* (18, 8, 25) {real, imag} */,
  {32'hc070c720, 32'hc10e75bc} /* (18, 8, 24) {real, imag} */,
  {32'hc15357be, 32'h413dadf3} /* (18, 8, 23) {real, imag} */,
  {32'hc1abd018, 32'h402dbc82} /* (18, 8, 22) {real, imag} */,
  {32'hc182fa47, 32'h40ac5295} /* (18, 8, 21) {real, imag} */,
  {32'h411f8ebc, 32'hc13f807a} /* (18, 8, 20) {real, imag} */,
  {32'h4183e79c, 32'h4084c6cd} /* (18, 8, 19) {real, imag} */,
  {32'h40caa6c5, 32'hc01e00e6} /* (18, 8, 18) {real, imag} */,
  {32'hc0be9580, 32'hc08e6074} /* (18, 8, 17) {real, imag} */,
  {32'hc0e93a5a, 32'h4080ea24} /* (18, 8, 16) {real, imag} */,
  {32'hc06d8e70, 32'h3f267500} /* (18, 8, 15) {real, imag} */,
  {32'h4086e7fa, 32'hbffc4b12} /* (18, 8, 14) {real, imag} */,
  {32'hc13787b9, 32'hc0fc9629} /* (18, 8, 13) {real, imag} */,
  {32'h4108072e, 32'h3f5ab0d0} /* (18, 8, 12) {real, imag} */,
  {32'h418360e8, 32'h3fc73e58} /* (18, 8, 11) {real, imag} */,
  {32'h40b09488, 32'hc199dc28} /* (18, 8, 10) {real, imag} */,
  {32'h4085f377, 32'hc0a4cfda} /* (18, 8, 9) {real, imag} */,
  {32'hc0e7807a, 32'h41017f57} /* (18, 8, 8) {real, imag} */,
  {32'hbf2587d0, 32'hbd417440} /* (18, 8, 7) {real, imag} */,
  {32'h40f23594, 32'hc0b69b9d} /* (18, 8, 6) {real, imag} */,
  {32'h40095815, 32'hbfb82808} /* (18, 8, 5) {real, imag} */,
  {32'h409db65a, 32'h401c4b41} /* (18, 8, 4) {real, imag} */,
  {32'hc02844fa, 32'h3f9fa0ba} /* (18, 8, 3) {real, imag} */,
  {32'hc1ae4f33, 32'hc1a79fd2} /* (18, 8, 2) {real, imag} */,
  {32'h41a4a274, 32'h41bbd90e} /* (18, 8, 1) {real, imag} */,
  {32'h418bae06, 32'h420b0557} /* (18, 8, 0) {real, imag} */,
  {32'hc0c4742c, 32'hc193fe1e} /* (18, 7, 31) {real, imag} */,
  {32'h41c26626, 32'hc0572550} /* (18, 7, 30) {real, imag} */,
  {32'hc11937b0, 32'hc0e5547d} /* (18, 7, 29) {real, imag} */,
  {32'h413ce270, 32'h40d76006} /* (18, 7, 28) {real, imag} */,
  {32'h4191ff38, 32'h406129e4} /* (18, 7, 27) {real, imag} */,
  {32'h414a1bd6, 32'hc12e77c7} /* (18, 7, 26) {real, imag} */,
  {32'hc1aa3959, 32'hc1c0d96e} /* (18, 7, 25) {real, imag} */,
  {32'hbfa6c28c, 32'hc0aa817a} /* (18, 7, 24) {real, imag} */,
  {32'h41269425, 32'h415f2b09} /* (18, 7, 23) {real, imag} */,
  {32'hc1553b6e, 32'hbfcd63ab} /* (18, 7, 22) {real, imag} */,
  {32'hc0c61a6a, 32'h41312c68} /* (18, 7, 21) {real, imag} */,
  {32'h40f6a654, 32'h3fff5270} /* (18, 7, 20) {real, imag} */,
  {32'hc160bc04, 32'hc0354315} /* (18, 7, 19) {real, imag} */,
  {32'h411cc670, 32'h41657840} /* (18, 7, 18) {real, imag} */,
  {32'hc02f4798, 32'hc130e194} /* (18, 7, 17) {real, imag} */,
  {32'hc06ee27a, 32'h3f8887fc} /* (18, 7, 16) {real, imag} */,
  {32'hc08cf666, 32'hc0c38f80} /* (18, 7, 15) {real, imag} */,
  {32'h3ec47380, 32'h41924975} /* (18, 7, 14) {real, imag} */,
  {32'hc0f52dd1, 32'hc06b7948} /* (18, 7, 13) {real, imag} */,
  {32'h411c2a00, 32'h3ff769c0} /* (18, 7, 12) {real, imag} */,
  {32'h40adf2c6, 32'h412fe1f8} /* (18, 7, 11) {real, imag} */,
  {32'hc15b5c64, 32'h3eaf7600} /* (18, 7, 10) {real, imag} */,
  {32'hc196f172, 32'h40bd4130} /* (18, 7, 9) {real, imag} */,
  {32'hc166ffde, 32'hc1c397ce} /* (18, 7, 8) {real, imag} */,
  {32'hc17f0cb9, 32'h41832600} /* (18, 7, 7) {real, imag} */,
  {32'h41094ff2, 32'h40337177} /* (18, 7, 6) {real, imag} */,
  {32'hc15e64c0, 32'hc110fce9} /* (18, 7, 5) {real, imag} */,
  {32'h41815c3c, 32'h4189f8f7} /* (18, 7, 4) {real, imag} */,
  {32'h40274128, 32'h4040ae17} /* (18, 7, 3) {real, imag} */,
  {32'h4119782c, 32'h41cac280} /* (18, 7, 2) {real, imag} */,
  {32'hc1089c61, 32'hc15efa54} /* (18, 7, 1) {real, imag} */,
  {32'hc1065c86, 32'hc168a097} /* (18, 7, 0) {real, imag} */,
  {32'h41168407, 32'hc0ca0da9} /* (18, 6, 31) {real, imag} */,
  {32'hc147e3fb, 32'hc1b4bcdb} /* (18, 6, 30) {real, imag} */,
  {32'hc1f947a8, 32'h409bfaea} /* (18, 6, 29) {real, imag} */,
  {32'hc10bdb60, 32'h4022d910} /* (18, 6, 28) {real, imag} */,
  {32'hc183ae76, 32'h40962556} /* (18, 6, 27) {real, imag} */,
  {32'h3f452a8c, 32'hc0e64c6c} /* (18, 6, 26) {real, imag} */,
  {32'hc0a7696a, 32'hc144d52e} /* (18, 6, 25) {real, imag} */,
  {32'hc00431c4, 32'h3f8d5e38} /* (18, 6, 24) {real, imag} */,
  {32'h417c95d0, 32'hc0ced53d} /* (18, 6, 23) {real, imag} */,
  {32'h411a3e71, 32'h4116a9f1} /* (18, 6, 22) {real, imag} */,
  {32'hbfdd5c6d, 32'hc09d9944} /* (18, 6, 21) {real, imag} */,
  {32'h41285615, 32'h4095f74e} /* (18, 6, 20) {real, imag} */,
  {32'h40a6c33e, 32'hc03c9148} /* (18, 6, 19) {real, imag} */,
  {32'hbfb4dcfc, 32'h40d702ce} /* (18, 6, 18) {real, imag} */,
  {32'h4015121b, 32'hc03e7b92} /* (18, 6, 17) {real, imag} */,
  {32'h4038221c, 32'h40cca0a8} /* (18, 6, 16) {real, imag} */,
  {32'h4098106e, 32'h40f758b0} /* (18, 6, 15) {real, imag} */,
  {32'h402e67ae, 32'h402f15df} /* (18, 6, 14) {real, imag} */,
  {32'hc154feee, 32'h40b3c034} /* (18, 6, 13) {real, imag} */,
  {32'h411896b4, 32'h409ecee4} /* (18, 6, 12) {real, imag} */,
  {32'hc0243448, 32'hc19c3c45} /* (18, 6, 11) {real, imag} */,
  {32'hc0ab5943, 32'h402cfa27} /* (18, 6, 10) {real, imag} */,
  {32'hc002bc54, 32'h41016721} /* (18, 6, 9) {real, imag} */,
  {32'hc11717f0, 32'hbeae02a0} /* (18, 6, 8) {real, imag} */,
  {32'h41bf3470, 32'h410dacb0} /* (18, 6, 7) {real, imag} */,
  {32'h40fec143, 32'hc1332e32} /* (18, 6, 6) {real, imag} */,
  {32'hc1702ad4, 32'h40ef7bb1} /* (18, 6, 5) {real, imag} */,
  {32'h408373e5, 32'h3f89fb8c} /* (18, 6, 4) {real, imag} */,
  {32'h40f251d8, 32'h41121351} /* (18, 6, 3) {real, imag} */,
  {32'h412298d6, 32'h413c2be4} /* (18, 6, 2) {real, imag} */,
  {32'h4066e11c, 32'hc0ffd4f3} /* (18, 6, 1) {real, imag} */,
  {32'hc09ea980, 32'hc1167201} /* (18, 6, 0) {real, imag} */,
  {32'h42a9d441, 32'h41e86370} /* (18, 5, 31) {real, imag} */,
  {32'hc23c1b42, 32'h417efceb} /* (18, 5, 30) {real, imag} */,
  {32'h418f9346, 32'hc0364c78} /* (18, 5, 29) {real, imag} */,
  {32'hc0bacc79, 32'hc10a7920} /* (18, 5, 28) {real, imag} */,
  {32'h405dbc1c, 32'h40cb5269} /* (18, 5, 27) {real, imag} */,
  {32'hc0a002d5, 32'h41668fd7} /* (18, 5, 26) {real, imag} */,
  {32'h406cad1c, 32'h411a1fc5} /* (18, 5, 25) {real, imag} */,
  {32'h3f126c1e, 32'hc191838e} /* (18, 5, 24) {real, imag} */,
  {32'h41331538, 32'hbfb42315} /* (18, 5, 23) {real, imag} */,
  {32'h40f8e11f, 32'hc0bc4a4f} /* (18, 5, 22) {real, imag} */,
  {32'hc174a2a4, 32'hc088ed37} /* (18, 5, 21) {real, imag} */,
  {32'hc12f27a1, 32'hc049164c} /* (18, 5, 20) {real, imag} */,
  {32'hc012765a, 32'hbf74d978} /* (18, 5, 19) {real, imag} */,
  {32'hc0ad566b, 32'h41a14a7d} /* (18, 5, 18) {real, imag} */,
  {32'h3f3c89f6, 32'h415f9d38} /* (18, 5, 17) {real, imag} */,
  {32'h40d15a50, 32'hc0672d15} /* (18, 5, 16) {real, imag} */,
  {32'h3f2b2268, 32'hbef2d4d0} /* (18, 5, 15) {real, imag} */,
  {32'h40a35792, 32'h40e92dcb} /* (18, 5, 14) {real, imag} */,
  {32'h4156e875, 32'h4112d87e} /* (18, 5, 13) {real, imag} */,
  {32'h3e40e900, 32'hc18f6592} /* (18, 5, 12) {real, imag} */,
  {32'hc0ca4efa, 32'hc1dc728b} /* (18, 5, 11) {real, imag} */,
  {32'h4011fe8f, 32'hc0a3906a} /* (18, 5, 10) {real, imag} */,
  {32'h3e02aa08, 32'hc1bec104} /* (18, 5, 9) {real, imag} */,
  {32'h41a26e57, 32'h41579de6} /* (18, 5, 8) {real, imag} */,
  {32'h42151339, 32'h41036c77} /* (18, 5, 7) {real, imag} */,
  {32'hc1aa97f4, 32'hc1122791} /* (18, 5, 6) {real, imag} */,
  {32'hc1d85a34, 32'h411973f2} /* (18, 5, 5) {real, imag} */,
  {32'hc0725112, 32'h418b0a0d} /* (18, 5, 4) {real, imag} */,
  {32'hc02d2e56, 32'h40fe8db4} /* (18, 5, 3) {real, imag} */,
  {32'hc1ce6b93, 32'hc238f374} /* (18, 5, 2) {real, imag} */,
  {32'h42681686, 32'h4290e72e} /* (18, 5, 1) {real, imag} */,
  {32'h4226e5e7, 32'h4241347b} /* (18, 5, 0) {real, imag} */,
  {32'hc2484ff7, 32'hc303b242} /* (18, 4, 31) {real, imag} */,
  {32'h4185754b, 32'h426609b9} /* (18, 4, 30) {real, imag} */,
  {32'h403908ea, 32'hc0dff103} /* (18, 4, 29) {real, imag} */,
  {32'hc26caaf3, 32'hc1c335ad} /* (18, 4, 28) {real, imag} */,
  {32'h41baaf6e, 32'hc19bf6e0} /* (18, 4, 27) {real, imag} */,
  {32'hc0dc34f6, 32'h4108da1c} /* (18, 4, 26) {real, imag} */,
  {32'hc086c778, 32'h412a01ba} /* (18, 4, 25) {real, imag} */,
  {32'h4074bd7e, 32'hbee48ba8} /* (18, 4, 24) {real, imag} */,
  {32'hc0df0bd2, 32'h40e70ad4} /* (18, 4, 23) {real, imag} */,
  {32'hc124f1a0, 32'h418bb399} /* (18, 4, 22) {real, imag} */,
  {32'h3e2cb390, 32'hc0e3109e} /* (18, 4, 21) {real, imag} */,
  {32'h415ac598, 32'h3f80cf73} /* (18, 4, 20) {real, imag} */,
  {32'hbf449070, 32'h413d046b} /* (18, 4, 19) {real, imag} */,
  {32'hc0c3cd48, 32'hc12c2125} /* (18, 4, 18) {real, imag} */,
  {32'hc0815f50, 32'hbfec8440} /* (18, 4, 17) {real, imag} */,
  {32'hc1337658, 32'hc0ad2a68} /* (18, 4, 16) {real, imag} */,
  {32'h40b70e60, 32'hbfb275e0} /* (18, 4, 15) {real, imag} */,
  {32'h40081b3e, 32'h3fb0f1d0} /* (18, 4, 14) {real, imag} */,
  {32'hc061f4be, 32'h41434b59} /* (18, 4, 13) {real, imag} */,
  {32'h406f3f67, 32'hc1a31d7a} /* (18, 4, 12) {real, imag} */,
  {32'h412c9bbe, 32'hbfbbda16} /* (18, 4, 11) {real, imag} */,
  {32'h4199d7af, 32'hc190b966} /* (18, 4, 10) {real, imag} */,
  {32'h408f3ca8, 32'hc0de4f87} /* (18, 4, 9) {real, imag} */,
  {32'h4123e1be, 32'h414f356b} /* (18, 4, 8) {real, imag} */,
  {32'hc062813a, 32'hc00ff1f4} /* (18, 4, 7) {real, imag} */,
  {32'hc1177314, 32'h421ae2a6} /* (18, 4, 6) {real, imag} */,
  {32'hc111795a, 32'h41e3db25} /* (18, 4, 5) {real, imag} */,
  {32'h4198c316, 32'h40865ea4} /* (18, 4, 4) {real, imag} */,
  {32'hc01b8cb8, 32'hc1818fab} /* (18, 4, 3) {real, imag} */,
  {32'h42d7928a, 32'h4267c8c7} /* (18, 4, 2) {real, imag} */,
  {32'hc2ffc6c7, 32'hc2310953} /* (18, 4, 1) {real, imag} */,
  {32'hc2818090, 32'hc1c9ca12} /* (18, 4, 0) {real, imag} */,
  {32'h42ca9d42, 32'hc2fedc80} /* (18, 3, 31) {real, imag} */,
  {32'hc26e0f18, 32'h43474fde} /* (18, 3, 30) {real, imag} */,
  {32'hc20aa8e9, 32'h4165ffcf} /* (18, 3, 29) {real, imag} */,
  {32'hc1e4befe, 32'hbea05de0} /* (18, 3, 28) {real, imag} */,
  {32'h41d1bb1e, 32'hc2170d95} /* (18, 3, 27) {real, imag} */,
  {32'hc1aac12a, 32'hc1958560} /* (18, 3, 26) {real, imag} */,
  {32'hc10b909a, 32'h418302ce} /* (18, 3, 25) {real, imag} */,
  {32'h41aa120c, 32'hc0593a4e} /* (18, 3, 24) {real, imag} */,
  {32'h40bd12dc, 32'h40977c17} /* (18, 3, 23) {real, imag} */,
  {32'hc09011e6, 32'hc1d9080b} /* (18, 3, 22) {real, imag} */,
  {32'h40a25c72, 32'hc1b862d6} /* (18, 3, 21) {real, imag} */,
  {32'hc048c2fe, 32'hc158738c} /* (18, 3, 20) {real, imag} */,
  {32'h411cdb5d, 32'hbdb19480} /* (18, 3, 19) {real, imag} */,
  {32'h40432a18, 32'h41109a89} /* (18, 3, 18) {real, imag} */,
  {32'h3fcabcba, 32'hc10934a2} /* (18, 3, 17) {real, imag} */,
  {32'hc03bc42b, 32'hc0377460} /* (18, 3, 16) {real, imag} */,
  {32'h40ad0e2a, 32'h40696407} /* (18, 3, 15) {real, imag} */,
  {32'hc0ff1c46, 32'h3d9e5300} /* (18, 3, 14) {real, imag} */,
  {32'h40c9e798, 32'hc18954a7} /* (18, 3, 13) {real, imag} */,
  {32'hc17e97ae, 32'h3fdf5a00} /* (18, 3, 12) {real, imag} */,
  {32'hc10973dc, 32'hc05d9b4a} /* (18, 3, 11) {real, imag} */,
  {32'h4180f45e, 32'hc0d74fba} /* (18, 3, 10) {real, imag} */,
  {32'h41313a2d, 32'hc0052554} /* (18, 3, 9) {real, imag} */,
  {32'hc19246d0, 32'hc1952422} /* (18, 3, 8) {real, imag} */,
  {32'hc19fffc0, 32'h41567e7a} /* (18, 3, 7) {real, imag} */,
  {32'h4187f5fd, 32'hc0d99b5c} /* (18, 3, 6) {real, imag} */,
  {32'hc04e3ad8, 32'h3fb32a90} /* (18, 3, 5) {real, imag} */,
  {32'h41aea328, 32'h4203dfa6} /* (18, 3, 4) {real, imag} */,
  {32'h41e00ead, 32'hc24026d7} /* (18, 3, 3) {real, imag} */,
  {32'h42320704, 32'h42c1a831} /* (18, 3, 2) {real, imag} */,
  {32'hc2b48fa7, 32'hc3260828} /* (18, 3, 1) {real, imag} */,
  {32'hbf3a5bc0, 32'hc1026d97} /* (18, 3, 0) {real, imag} */,
  {32'h4485513a, 32'hc12712a0} /* (18, 2, 31) {real, imag} */,
  {32'hc4075d3a, 32'h42e86d00} /* (18, 2, 30) {real, imag} */,
  {32'h420b143d, 32'h41fe5615} /* (18, 2, 29) {real, imag} */,
  {32'h42915d30, 32'hc2a01cde} /* (18, 2, 28) {real, imag} */,
  {32'hc249ea44, 32'h421c15e2} /* (18, 2, 27) {real, imag} */,
  {32'hc1330a2d, 32'h414e353d} /* (18, 2, 26) {real, imag} */,
  {32'h41a1c464, 32'hc1823f05} /* (18, 2, 25) {real, imag} */,
  {32'hc1613b0a, 32'h4158ef14} /* (18, 2, 24) {real, imag} */,
  {32'h408cdc66, 32'h3fcfaa3c} /* (18, 2, 23) {real, imag} */,
  {32'hbf97b9c4, 32'h410d62d1} /* (18, 2, 22) {real, imag} */,
  {32'hc024dd75, 32'h41b2dc6b} /* (18, 2, 21) {real, imag} */,
  {32'h3f9b9b18, 32'hc1068819} /* (18, 2, 20) {real, imag} */,
  {32'hc1146b9f, 32'h403d1d20} /* (18, 2, 19) {real, imag} */,
  {32'hc016983f, 32'h415174bd} /* (18, 2, 18) {real, imag} */,
  {32'h40e2e486, 32'hc0887311} /* (18, 2, 17) {real, imag} */,
  {32'hbff10c6a, 32'hc053ddd4} /* (18, 2, 16) {real, imag} */,
  {32'h40d4502c, 32'hc093f18a} /* (18, 2, 15) {real, imag} */,
  {32'hc0361690, 32'hc03c9606} /* (18, 2, 14) {real, imag} */,
  {32'h3fb0d500, 32'hc0eb0c05} /* (18, 2, 13) {real, imag} */,
  {32'h40d2f316, 32'h41018188} /* (18, 2, 12) {real, imag} */,
  {32'hc19b09f2, 32'hc1c21458} /* (18, 2, 11) {real, imag} */,
  {32'hc078c564, 32'hc07a6448} /* (18, 2, 10) {real, imag} */,
  {32'h418eae98, 32'hbeb4d750} /* (18, 2, 9) {real, imag} */,
  {32'hc14253be, 32'hc2234232} /* (18, 2, 8) {real, imag} */,
  {32'h41955588, 32'hc102905a} /* (18, 2, 7) {real, imag} */,
  {32'h41b3f47c, 32'h41bc609f} /* (18, 2, 6) {real, imag} */,
  {32'hc279d368, 32'hc2acbb2f} /* (18, 2, 5) {real, imag} */,
  {32'h42c76c6e, 32'hc21b6e10} /* (18, 2, 4) {real, imag} */,
  {32'h421f44af, 32'h41be5dcc} /* (18, 2, 3) {real, imag} */,
  {32'hc3bfb06a, 32'h42e0251e} /* (18, 2, 2) {real, imag} */,
  {32'h441ef118, 32'hc3063630} /* (18, 2, 1) {real, imag} */,
  {32'h440dcf57, 32'h42c25e41} /* (18, 2, 0) {real, imag} */,
  {32'hc4a59ac8, 32'h4396bdb0} /* (18, 1, 31) {real, imag} */,
  {32'h43b0f2ea, 32'hc248d7d4} /* (18, 1, 30) {real, imag} */,
  {32'hc12bd25c, 32'h404813e0} /* (18, 1, 29) {real, imag} */,
  {32'hc29c0b24, 32'hc2634bbd} /* (18, 1, 28) {real, imag} */,
  {32'h42f4b350, 32'hc1188ef4} /* (18, 1, 27) {real, imag} */,
  {32'h423f9e19, 32'hc20297ce} /* (18, 1, 26) {real, imag} */,
  {32'hc1343e0d, 32'h41fa1f54} /* (18, 1, 25) {real, imag} */,
  {32'h416afe8a, 32'hc1706d21} /* (18, 1, 24) {real, imag} */,
  {32'hc086d7d4, 32'hc1e51a0b} /* (18, 1, 23) {real, imag} */,
  {32'hbfd8b9ca, 32'h4139152c} /* (18, 1, 22) {real, imag} */,
  {32'h41dbea6d, 32'hc1bb826a} /* (18, 1, 21) {real, imag} */,
  {32'hc1e3cc12, 32'h40b8bb6e} /* (18, 1, 20) {real, imag} */,
  {32'h41811eda, 32'hc02fd45c} /* (18, 1, 19) {real, imag} */,
  {32'h40834555, 32'h401f2735} /* (18, 1, 18) {real, imag} */,
  {32'h413162c4, 32'h404f189d} /* (18, 1, 17) {real, imag} */,
  {32'h4119ee35, 32'h3f578718} /* (18, 1, 16) {real, imag} */,
  {32'hc128bc65, 32'hc01fcaa5} /* (18, 1, 15) {real, imag} */,
  {32'h40553931, 32'h41aeca0a} /* (18, 1, 14) {real, imag} */,
  {32'hc04d6980, 32'h4042d80e} /* (18, 1, 13) {real, imag} */,
  {32'h417d21e6, 32'h40aad8a0} /* (18, 1, 12) {real, imag} */,
  {32'hc0c6b422, 32'h41797b76} /* (18, 1, 11) {real, imag} */,
  {32'hc04c2398, 32'h412c2ff1} /* (18, 1, 10) {real, imag} */,
  {32'h3ff7aa80, 32'h4020195d} /* (18, 1, 9) {real, imag} */,
  {32'h41d59114, 32'h4225812a} /* (18, 1, 8) {real, imag} */,
  {32'h41133642, 32'hc13e826c} /* (18, 1, 7) {real, imag} */,
  {32'h413d99f9, 32'hc13b9e74} /* (18, 1, 6) {real, imag} */,
  {32'h4270565c, 32'h4226304d} /* (18, 1, 5) {real, imag} */,
  {32'hc28ec0fb, 32'hc1f3042b} /* (18, 1, 4) {real, imag} */,
  {32'hc1002ec0, 32'hc2326612} /* (18, 1, 3) {real, imag} */,
  {32'h43ea29e0, 32'h44066126} /* (18, 1, 2) {real, imag} */,
  {32'hc4ee823b, 32'hc4700eda} /* (18, 1, 1) {real, imag} */,
  {32'hc4c974b6, 32'hc38889b4} /* (18, 1, 0) {real, imag} */,
  {32'hc4997341, 32'h4462c249} /* (18, 0, 31) {real, imag} */,
  {32'h4304c9ac, 32'hc387f00f} /* (18, 0, 30) {real, imag} */,
  {32'h4219ebdc, 32'hc1a0da9c} /* (18, 0, 29) {real, imag} */,
  {32'h4190b979, 32'hc1fb6b00} /* (18, 0, 28) {real, imag} */,
  {32'h4219ae56, 32'h416c8ae2} /* (18, 0, 27) {real, imag} */,
  {32'h41592cee, 32'h41a169f5} /* (18, 0, 26) {real, imag} */,
  {32'hc043118a, 32'h407e040c} /* (18, 0, 25) {real, imag} */,
  {32'h41858355, 32'hc20d6550} /* (18, 0, 24) {real, imag} */,
  {32'hc0ab37da, 32'hc04f3dce} /* (18, 0, 23) {real, imag} */,
  {32'h3fa9c570, 32'hc10bfc0a} /* (18, 0, 22) {real, imag} */,
  {32'h40b8d772, 32'hbe2afda0} /* (18, 0, 21) {real, imag} */,
  {32'h3f944520, 32'hc081e762} /* (18, 0, 20) {real, imag} */,
  {32'h410f81ce, 32'h4095d0fc} /* (18, 0, 19) {real, imag} */,
  {32'hbf07fff0, 32'hc098d6d0} /* (18, 0, 18) {real, imag} */,
  {32'h40e45abb, 32'h4123f8e2} /* (18, 0, 17) {real, imag} */,
  {32'hbfa25886, 32'h00000000} /* (18, 0, 16) {real, imag} */,
  {32'h40e45abb, 32'hc123f8e2} /* (18, 0, 15) {real, imag} */,
  {32'hbf07fff0, 32'h4098d6d0} /* (18, 0, 14) {real, imag} */,
  {32'h410f81ce, 32'hc095d0fc} /* (18, 0, 13) {real, imag} */,
  {32'h3f944520, 32'h4081e762} /* (18, 0, 12) {real, imag} */,
  {32'h40b8d772, 32'h3e2afda0} /* (18, 0, 11) {real, imag} */,
  {32'h3fa9c570, 32'h410bfc0a} /* (18, 0, 10) {real, imag} */,
  {32'hc0ab37da, 32'h404f3dce} /* (18, 0, 9) {real, imag} */,
  {32'h41858355, 32'h420d6550} /* (18, 0, 8) {real, imag} */,
  {32'hc043118a, 32'hc07e040c} /* (18, 0, 7) {real, imag} */,
  {32'h41592cee, 32'hc1a169f5} /* (18, 0, 6) {real, imag} */,
  {32'h4219ae56, 32'hc16c8ae2} /* (18, 0, 5) {real, imag} */,
  {32'h4190b979, 32'h41fb6b00} /* (18, 0, 4) {real, imag} */,
  {32'h4219ebdc, 32'h41a0da9c} /* (18, 0, 3) {real, imag} */,
  {32'h4304c9ac, 32'h4387f00f} /* (18, 0, 2) {real, imag} */,
  {32'hc4997341, 32'hc462c249} /* (18, 0, 1) {real, imag} */,
  {32'hc4d63932, 32'h00000000} /* (18, 0, 0) {real, imag} */,
  {32'hc4aaf334, 32'h44250cfc} /* (17, 31, 31) {real, imag} */,
  {32'h43b119ae, 32'hc3da851f} /* (17, 31, 30) {real, imag} */,
  {32'hc22d1d2b, 32'h425736df} /* (17, 31, 29) {real, imag} */,
  {32'hc22d22e4, 32'h41fe4f6d} /* (17, 31, 28) {real, imag} */,
  {32'h426f34bc, 32'hc219facb} /* (17, 31, 27) {real, imag} */,
  {32'h412a8dda, 32'h40108c04} /* (17, 31, 26) {real, imag} */,
  {32'hc1082fea, 32'h412a350a} /* (17, 31, 25) {real, imag} */,
  {32'h41a50ad9, 32'hc28df75e} /* (17, 31, 24) {real, imag} */,
  {32'hc059dcbc, 32'h40943fb1} /* (17, 31, 23) {real, imag} */,
  {32'h40be94db, 32'h3f19d878} /* (17, 31, 22) {real, imag} */,
  {32'h3f7015e0, 32'hc1d25396} /* (17, 31, 21) {real, imag} */,
  {32'h4166d210, 32'h414e21ae} /* (17, 31, 20) {real, imag} */,
  {32'hc18a5661, 32'h40aad338} /* (17, 31, 19) {real, imag} */,
  {32'hc182c1b2, 32'h406b45f4} /* (17, 31, 18) {real, imag} */,
  {32'h4138029a, 32'hbfb1f370} /* (17, 31, 17) {real, imag} */,
  {32'hc1194d8e, 32'h4129aef1} /* (17, 31, 16) {real, imag} */,
  {32'h40be2cb7, 32'hc185e109} /* (17, 31, 15) {real, imag} */,
  {32'hbfa02454, 32'hc07379a5} /* (17, 31, 14) {real, imag} */,
  {32'hc0077376, 32'hc007e550} /* (17, 31, 13) {real, imag} */,
  {32'h413b49f7, 32'hc13e1108} /* (17, 31, 12) {real, imag} */,
  {32'hc03e8df6, 32'h41926f32} /* (17, 31, 11) {real, imag} */,
  {32'hc051f9b6, 32'h411254de} /* (17, 31, 10) {real, imag} */,
  {32'hbe8ac650, 32'h4126c95f} /* (17, 31, 9) {real, imag} */,
  {32'h419f9115, 32'h420c2e6e} /* (17, 31, 8) {real, imag} */,
  {32'hc15ea69c, 32'hc166a351} /* (17, 31, 7) {real, imag} */,
  {32'h423476a8, 32'hc0fd81b3} /* (17, 31, 6) {real, imag} */,
  {32'h431a21f0, 32'hc14962a4} /* (17, 31, 5) {real, imag} */,
  {32'hc2798756, 32'h428e2986} /* (17, 31, 4) {real, imag} */,
  {32'hbfd78d70, 32'hc1a9f710} /* (17, 31, 3) {real, imag} */,
  {32'h438723ca, 32'h42507471} /* (17, 31, 2) {real, imag} */,
  {32'hc46325b8, 32'hc3204e43} /* (17, 31, 1) {real, imag} */,
  {32'hc48ef3c0, 32'h437de829} /* (17, 31, 0) {real, imag} */,
  {32'h43e45dc9, 32'h430390fb} /* (17, 30, 31) {real, imag} */,
  {32'hc38e17b0, 32'hc2ccefe8} /* (17, 30, 30) {real, imag} */,
  {32'h4224a4b4, 32'h40c3785f} /* (17, 30, 29) {real, imag} */,
  {32'h42cdf940, 32'h422cdad9} /* (17, 30, 28) {real, imag} */,
  {32'hc2aa10a1, 32'h429e6237} /* (17, 30, 27) {real, imag} */,
  {32'hbe644850, 32'hc20a2d36} /* (17, 30, 26) {real, imag} */,
  {32'h3febc9e9, 32'h410136c6} /* (17, 30, 25) {real, imag} */,
  {32'hc12299bb, 32'h414456ab} /* (17, 30, 24) {real, imag} */,
  {32'hc0f37bc8, 32'hc0dd08d7} /* (17, 30, 23) {real, imag} */,
  {32'h41299585, 32'hc0cb4fe4} /* (17, 30, 22) {real, imag} */,
  {32'hc03d5ae1, 32'h3fde1358} /* (17, 30, 21) {real, imag} */,
  {32'h4033c1d0, 32'h40e82340} /* (17, 30, 20) {real, imag} */,
  {32'h3fa11f96, 32'h40035031} /* (17, 30, 19) {real, imag} */,
  {32'hc145a022, 32'h4113a118} /* (17, 30, 18) {real, imag} */,
  {32'h40834f7e, 32'hc08eedc6} /* (17, 30, 17) {real, imag} */,
  {32'h40d2c800, 32'h405e694c} /* (17, 30, 16) {real, imag} */,
  {32'h3f17f04c, 32'h414619fc} /* (17, 30, 15) {real, imag} */,
  {32'h40c93973, 32'hc12248c7} /* (17, 30, 14) {real, imag} */,
  {32'h3fedae26, 32'hc02ff8d8} /* (17, 30, 13) {real, imag} */,
  {32'h3e9d8ac0, 32'h4132476c} /* (17, 30, 12) {real, imag} */,
  {32'hc094a283, 32'hc15995c9} /* (17, 30, 11) {real, imag} */,
  {32'hc099dee0, 32'hc12b02f3} /* (17, 30, 10) {real, imag} */,
  {32'hc0c7ef9d, 32'hc0de6cc8} /* (17, 30, 9) {real, imag} */,
  {32'hc24ba448, 32'hc1a86196} /* (17, 30, 8) {real, imag} */,
  {32'h42028a66, 32'h414e0f40} /* (17, 30, 7) {real, imag} */,
  {32'hbe2a4e00, 32'h410a4aee} /* (17, 30, 6) {real, imag} */,
  {32'hc27acdea, 32'hc228e65a} /* (17, 30, 5) {real, imag} */,
  {32'h4219df6a, 32'h428263c2} /* (17, 30, 4) {real, imag} */,
  {32'h428fef67, 32'hc0001cd8} /* (17, 30, 3) {real, imag} */,
  {32'hc3bd1670, 32'hc2a34ecf} /* (17, 30, 2) {real, imag} */,
  {32'h4447915e, 32'hc119cbf4} /* (17, 30, 1) {real, imag} */,
  {32'h43d3456d, 32'hc2afd54d} /* (17, 30, 0) {real, imag} */,
  {32'hc2654387, 32'h4305d28e} /* (17, 29, 31) {real, imag} */,
  {32'h4230f8ea, 32'hc2ab433c} /* (17, 29, 30) {real, imag} */,
  {32'h41b50749, 32'h4277ab50} /* (17, 29, 29) {real, imag} */,
  {32'h41c1ccfe, 32'hc2130496} /* (17, 29, 28) {real, imag} */,
  {32'hc1a4350a, 32'hc1b986f0} /* (17, 29, 27) {real, imag} */,
  {32'h40f2105a, 32'hc149a48d} /* (17, 29, 26) {real, imag} */,
  {32'hc10c2bab, 32'hc0cfd531} /* (17, 29, 25) {real, imag} */,
  {32'h40f2efa9, 32'h411ce4fc} /* (17, 29, 24) {real, imag} */,
  {32'h40c23098, 32'h40d80a4e} /* (17, 29, 23) {real, imag} */,
  {32'hc03cd734, 32'hc12e8d2a} /* (17, 29, 22) {real, imag} */,
  {32'h410364bd, 32'h3f3cf810} /* (17, 29, 21) {real, imag} */,
  {32'hc0a5bd73, 32'h418432b4} /* (17, 29, 20) {real, imag} */,
  {32'h408c8fbc, 32'h3f0b82b0} /* (17, 29, 19) {real, imag} */,
  {32'h40568e6d, 32'h3d33d740} /* (17, 29, 18) {real, imag} */,
  {32'h3fc00922, 32'h409ff018} /* (17, 29, 17) {real, imag} */,
  {32'hc13a2fd4, 32'hc10eb359} /* (17, 29, 16) {real, imag} */,
  {32'h41262c02, 32'h4137b195} /* (17, 29, 15) {real, imag} */,
  {32'hc1918005, 32'hc1235f08} /* (17, 29, 14) {real, imag} */,
  {32'hbfe3a8d2, 32'hc11d670a} /* (17, 29, 13) {real, imag} */,
  {32'hc09537ba, 32'hc03317b0} /* (17, 29, 12) {real, imag} */,
  {32'hc17be565, 32'hc10eb270} /* (17, 29, 11) {real, imag} */,
  {32'hc04bfca9, 32'hc097cc30} /* (17, 29, 10) {real, imag} */,
  {32'hc169063c, 32'h410bc7a0} /* (17, 29, 9) {real, imag} */,
  {32'hc049598c, 32'hc0ab2d17} /* (17, 29, 8) {real, imag} */,
  {32'hc0a2b79c, 32'hc19ba0c9} /* (17, 29, 7) {real, imag} */,
  {32'hc1edb4db, 32'h40ff7a40} /* (17, 29, 6) {real, imag} */,
  {32'h42207314, 32'h414b5c9e} /* (17, 29, 5) {real, imag} */,
  {32'hc226d3fa, 32'h41c1aa41} /* (17, 29, 4) {real, imag} */,
  {32'h410b0521, 32'h40f32a60} /* (17, 29, 3) {real, imag} */,
  {32'hc2389607, 32'hc318522a} /* (17, 29, 2) {real, imag} */,
  {32'h4300dd57, 32'h42b579f5} /* (17, 29, 1) {real, imag} */,
  {32'h420341ba, 32'h40833f42} /* (17, 29, 0) {real, imag} */,
  {32'hc2c04ae0, 32'h421d6da8} /* (17, 28, 31) {real, imag} */,
  {32'h42a29447, 32'hc2a39302} /* (17, 28, 30) {real, imag} */,
  {32'hc1dbbaa7, 32'h41e96c84} /* (17, 28, 29) {real, imag} */,
  {32'h41b5a3fe, 32'hc0c31bfa} /* (17, 28, 28) {real, imag} */,
  {32'hc1cd42d7, 32'hc1a26184} /* (17, 28, 27) {real, imag} */,
  {32'hbfd80170, 32'hc1e88f71} /* (17, 28, 26) {real, imag} */,
  {32'hc190ec04, 32'h41a2e694} /* (17, 28, 25) {real, imag} */,
  {32'h41498354, 32'h404f3887} /* (17, 28, 24) {real, imag} */,
  {32'h40346804, 32'hc0d43eeb} /* (17, 28, 23) {real, imag} */,
  {32'h41336582, 32'h405ea772} /* (17, 28, 22) {real, imag} */,
  {32'h4121376b, 32'h412198e2} /* (17, 28, 21) {real, imag} */,
  {32'hc0edaac3, 32'h40518c38} /* (17, 28, 20) {real, imag} */,
  {32'h3e8c3c60, 32'hc184eb5d} /* (17, 28, 19) {real, imag} */,
  {32'h40a066c8, 32'hbf1062b8} /* (17, 28, 18) {real, imag} */,
  {32'h40a5e585, 32'hc0acc103} /* (17, 28, 17) {real, imag} */,
  {32'h4141e00c, 32'hc1002555} /* (17, 28, 16) {real, imag} */,
  {32'hc131be4a, 32'h4126acea} /* (17, 28, 15) {real, imag} */,
  {32'h414ba620, 32'h40a414c0} /* (17, 28, 14) {real, imag} */,
  {32'h4056db14, 32'h403a0161} /* (17, 28, 13) {real, imag} */,
  {32'h40e9525a, 32'h408ec5d9} /* (17, 28, 12) {real, imag} */,
  {32'hbf92ed97, 32'hc174f120} /* (17, 28, 11) {real, imag} */,
  {32'hc07e56e3, 32'hc14d006c} /* (17, 28, 10) {real, imag} */,
  {32'hc157e283, 32'hbf86e4ee} /* (17, 28, 9) {real, imag} */,
  {32'h41e7814d, 32'h41e7e69c} /* (17, 28, 8) {real, imag} */,
  {32'h4039665a, 32'hc10e25e2} /* (17, 28, 7) {real, imag} */,
  {32'hc1757136, 32'hc0d7b64c} /* (17, 28, 6) {real, imag} */,
  {32'h419ea620, 32'h3e3b7ad0} /* (17, 28, 5) {real, imag} */,
  {32'hc2715196, 32'h41d27f96} /* (17, 28, 4) {real, imag} */,
  {32'h41660558, 32'h41c89c82} /* (17, 28, 3) {real, imag} */,
  {32'h414ae830, 32'hc25911df} /* (17, 28, 2) {real, imag} */,
  {32'hc1c4f2d4, 32'h42d419ba} /* (17, 28, 1) {real, imag} */,
  {32'hc29cbe58, 32'h4273c19b} /* (17, 28, 0) {real, imag} */,
  {32'h4231115a, 32'hc2a15aad} /* (17, 27, 31) {real, imag} */,
  {32'h4108be06, 32'h4222e1ac} /* (17, 27, 30) {real, imag} */,
  {32'hc0252f50, 32'hc1550cb8} /* (17, 27, 29) {real, imag} */,
  {32'hc0b5fc26, 32'hc0e72f2d} /* (17, 27, 28) {real, imag} */,
  {32'hc1a65d44, 32'hc1b70752} /* (17, 27, 27) {real, imag} */,
  {32'h3f9257b0, 32'h420a1da8} /* (17, 27, 26) {real, imag} */,
  {32'hc1cbb574, 32'hc1d393a4} /* (17, 27, 25) {real, imag} */,
  {32'h4147e471, 32'h413bc81a} /* (17, 27, 24) {real, imag} */,
  {32'h41945d6e, 32'h41814249} /* (17, 27, 23) {real, imag} */,
  {32'h415e8afb, 32'h40727918} /* (17, 27, 22) {real, imag} */,
  {32'hc12de120, 32'hc0037aac} /* (17, 27, 21) {real, imag} */,
  {32'hbf05c15a, 32'h416acd4c} /* (17, 27, 20) {real, imag} */,
  {32'h41091c18, 32'hc158718e} /* (17, 27, 19) {real, imag} */,
  {32'h40c522ca, 32'hc0974341} /* (17, 27, 18) {real, imag} */,
  {32'h401578f2, 32'h40c60530} /* (17, 27, 17) {real, imag} */,
  {32'h411e0188, 32'h40620910} /* (17, 27, 16) {real, imag} */,
  {32'h40002650, 32'h40c6687d} /* (17, 27, 15) {real, imag} */,
  {32'h409ccafe, 32'h403c30ce} /* (17, 27, 14) {real, imag} */,
  {32'hc05eed69, 32'h3f19238c} /* (17, 27, 13) {real, imag} */,
  {32'h41678729, 32'h41276fc6} /* (17, 27, 12) {real, imag} */,
  {32'hc0a357ce, 32'hc08fc2e4} /* (17, 27, 11) {real, imag} */,
  {32'hc1933d1e, 32'h4177daf8} /* (17, 27, 10) {real, imag} */,
  {32'hbf678388, 32'h40a7a49a} /* (17, 27, 9) {real, imag} */,
  {32'hc0fa2238, 32'hc1039ad4} /* (17, 27, 8) {real, imag} */,
  {32'h41075cea, 32'hc09e30c0} /* (17, 27, 7) {real, imag} */,
  {32'h3f086558, 32'hc1684462} /* (17, 27, 6) {real, imag} */,
  {32'h4103344e, 32'hc02aacb8} /* (17, 27, 5) {real, imag} */,
  {32'hc18c3c2e, 32'hc1006192} /* (17, 27, 4) {real, imag} */,
  {32'h40e9ee35, 32'hc09f5d45} /* (17, 27, 3) {real, imag} */,
  {32'hc21b94ba, 32'h40984324} /* (17, 27, 2) {real, imag} */,
  {32'h42bc336d, 32'hc1fa391f} /* (17, 27, 1) {real, imag} */,
  {32'h41ecaa0f, 32'hc2353dfb} /* (17, 27, 0) {real, imag} */,
  {32'h419c0ad1, 32'h3fcc1b98} /* (17, 26, 31) {real, imag} */,
  {32'h40d750d2, 32'h400beeda} /* (17, 26, 30) {real, imag} */,
  {32'hc1701db7, 32'h409f5cb3} /* (17, 26, 29) {real, imag} */,
  {32'h410975f8, 32'hc0e55a7e} /* (17, 26, 28) {real, imag} */,
  {32'hbed71f40, 32'hc0a76230} /* (17, 26, 27) {real, imag} */,
  {32'hc082fb68, 32'hbfc0043c} /* (17, 26, 26) {real, imag} */,
  {32'h41c61766, 32'hc0231105} /* (17, 26, 25) {real, imag} */,
  {32'hc2076142, 32'h40a9f186} /* (17, 26, 24) {real, imag} */,
  {32'h41943509, 32'h41589656} /* (17, 26, 23) {real, imag} */,
  {32'hc1b5e78a, 32'h40eab484} /* (17, 26, 22) {real, imag} */,
  {32'h40a57003, 32'hc109045d} /* (17, 26, 21) {real, imag} */,
  {32'h412c306e, 32'h40c64b40} /* (17, 26, 20) {real, imag} */,
  {32'h405797f8, 32'h416f3ecf} /* (17, 26, 19) {real, imag} */,
  {32'hbfec8da4, 32'h418a70fb} /* (17, 26, 18) {real, imag} */,
  {32'hc13017bf, 32'h40d6c220} /* (17, 26, 17) {real, imag} */,
  {32'hbf1d27c0, 32'h40ca5d24} /* (17, 26, 16) {real, imag} */,
  {32'hbf35d0c0, 32'hc11a1159} /* (17, 26, 15) {real, imag} */,
  {32'h411a0c3a, 32'hc17cdda0} /* (17, 26, 14) {real, imag} */,
  {32'hc02a7715, 32'h407e474b} /* (17, 26, 13) {real, imag} */,
  {32'h3f6f84b0, 32'hbf81144f} /* (17, 26, 12) {real, imag} */,
  {32'h40e69aeb, 32'h3fa19564} /* (17, 26, 11) {real, imag} */,
  {32'hc16a9c85, 32'hc11d64d6} /* (17, 26, 10) {real, imag} */,
  {32'h41189e84, 32'h40f1d3dc} /* (17, 26, 9) {real, imag} */,
  {32'hc13bb20f, 32'h40564e42} /* (17, 26, 8) {real, imag} */,
  {32'h412cca39, 32'hc14b0fe8} /* (17, 26, 7) {real, imag} */,
  {32'h418258de, 32'hc021d861} /* (17, 26, 6) {real, imag} */,
  {32'hc0c61f40, 32'h414ab8e0} /* (17, 26, 5) {real, imag} */,
  {32'hc089a4bb, 32'hc1799f9f} /* (17, 26, 4) {real, imag} */,
  {32'hbe4afc70, 32'h420252a7} /* (17, 26, 3) {real, imag} */,
  {32'hc1c0960e, 32'h40d70cfb} /* (17, 26, 2) {real, imag} */,
  {32'h41d47d58, 32'hc0af9170} /* (17, 26, 1) {real, imag} */,
  {32'hc148770f, 32'h40a44bb6} /* (17, 26, 0) {real, imag} */,
  {32'hc0a21d4c, 32'h40cea690} /* (17, 25, 31) {real, imag} */,
  {32'hc10ebeae, 32'hc0b16189} /* (17, 25, 30) {real, imag} */,
  {32'hc1597566, 32'h3ef6a980} /* (17, 25, 29) {real, imag} */,
  {32'h41c1ce0c, 32'hc0b50339} /* (17, 25, 28) {real, imag} */,
  {32'hc13fece6, 32'h410e8190} /* (17, 25, 27) {real, imag} */,
  {32'h3fbbdd50, 32'h41e220a0} /* (17, 25, 26) {real, imag} */,
  {32'h4048af70, 32'hbe6f15e0} /* (17, 25, 25) {real, imag} */,
  {32'hc09af406, 32'h41168f58} /* (17, 25, 24) {real, imag} */,
  {32'h4078df06, 32'hc1991d74} /* (17, 25, 23) {real, imag} */,
  {32'hc0d8cdf1, 32'h40d4c8af} /* (17, 25, 22) {real, imag} */,
  {32'h4107033d, 32'h409d59a7} /* (17, 25, 21) {real, imag} */,
  {32'h3f63693f, 32'hc1184337} /* (17, 25, 20) {real, imag} */,
  {32'hc072bbff, 32'h410825d2} /* (17, 25, 19) {real, imag} */,
  {32'hc12ba945, 32'hc043fee1} /* (17, 25, 18) {real, imag} */,
  {32'h40e334c6, 32'h3f16d614} /* (17, 25, 17) {real, imag} */,
  {32'h413b7d54, 32'hc175c08d} /* (17, 25, 16) {real, imag} */,
  {32'hc084ceb0, 32'h41290fe5} /* (17, 25, 15) {real, imag} */,
  {32'hbe72a660, 32'h411f8c56} /* (17, 25, 14) {real, imag} */,
  {32'h40b4fda5, 32'hc0ac22c6} /* (17, 25, 13) {real, imag} */,
  {32'h408c5b15, 32'h40222e3d} /* (17, 25, 12) {real, imag} */,
  {32'h417ef63c, 32'hc15c15f4} /* (17, 25, 11) {real, imag} */,
  {32'h4180cf70, 32'hc120d1c0} /* (17, 25, 10) {real, imag} */,
  {32'hbfb8e294, 32'hc14162b1} /* (17, 25, 9) {real, imag} */,
  {32'hbfad47c4, 32'hbfec9560} /* (17, 25, 8) {real, imag} */,
  {32'hbfe4f840, 32'h4168819b} /* (17, 25, 7) {real, imag} */,
  {32'hc1a202aa, 32'h408be56c} /* (17, 25, 6) {real, imag} */,
  {32'hc17ce140, 32'h40f574e4} /* (17, 25, 5) {real, imag} */,
  {32'hc0ce81b4, 32'hc1b440e0} /* (17, 25, 4) {real, imag} */,
  {32'hc081af26, 32'hc02c7d13} /* (17, 25, 3) {real, imag} */,
  {32'h42128712, 32'h4138a2b3} /* (17, 25, 2) {real, imag} */,
  {32'hc0c306d4, 32'hc05d9518} /* (17, 25, 1) {real, imag} */,
  {32'hc128a444, 32'hc1adcd86} /* (17, 25, 0) {real, imag} */,
  {32'h414dd8a0, 32'hc15cee6c} /* (17, 24, 31) {real, imag} */,
  {32'hc1aa00ee, 32'h418a558c} /* (17, 24, 30) {real, imag} */,
  {32'hc0a060ec, 32'hc1cd3f04} /* (17, 24, 29) {real, imag} */,
  {32'h420c2766, 32'hc08dfe6b} /* (17, 24, 28) {real, imag} */,
  {32'hbfd84030, 32'hc1669dc0} /* (17, 24, 27) {real, imag} */,
  {32'hc0e67990, 32'hc0567dc8} /* (17, 24, 26) {real, imag} */,
  {32'hc119ae6f, 32'hc15e18c8} /* (17, 24, 25) {real, imag} */,
  {32'h40bb8bc0, 32'h417a636e} /* (17, 24, 24) {real, imag} */,
  {32'h413b2c56, 32'hc07ca8a8} /* (17, 24, 23) {real, imag} */,
  {32'hc030ee0c, 32'hc0af83d2} /* (17, 24, 22) {real, imag} */,
  {32'h4102b87e, 32'hbf0a9212} /* (17, 24, 21) {real, imag} */,
  {32'h41810d72, 32'hc150abe0} /* (17, 24, 20) {real, imag} */,
  {32'hc1022c74, 32'hc0cfe76a} /* (17, 24, 19) {real, imag} */,
  {32'h40004c33, 32'h4113c6d4} /* (17, 24, 18) {real, imag} */,
  {32'hc06c6594, 32'h3d74cac0} /* (17, 24, 17) {real, imag} */,
  {32'h411e2791, 32'h407bcc8e} /* (17, 24, 16) {real, imag} */,
  {32'hc08e1725, 32'hc0b18f24} /* (17, 24, 15) {real, imag} */,
  {32'h4041a8ad, 32'hc10ea972} /* (17, 24, 14) {real, imag} */,
  {32'hbf96165c, 32'h3fa933ea} /* (17, 24, 13) {real, imag} */,
  {32'h4013278c, 32'hc1035490} /* (17, 24, 12) {real, imag} */,
  {32'hc12855cd, 32'hc100491f} /* (17, 24, 11) {real, imag} */,
  {32'hc0899b3c, 32'h4180d8d6} /* (17, 24, 10) {real, imag} */,
  {32'h40dac23a, 32'hc0fc370a} /* (17, 24, 9) {real, imag} */,
  {32'hc200aa9b, 32'hc0b80978} /* (17, 24, 8) {real, imag} */,
  {32'h40868c50, 32'hc0c993a6} /* (17, 24, 7) {real, imag} */,
  {32'hc1266aad, 32'h3f8f2d20} /* (17, 24, 6) {real, imag} */,
  {32'h407dc456, 32'h4102f736} /* (17, 24, 5) {real, imag} */,
  {32'h413bb5cf, 32'hc0879bc4} /* (17, 24, 4) {real, imag} */,
  {32'hbf97a4b8, 32'h413f32e1} /* (17, 24, 3) {real, imag} */,
  {32'hc214bc10, 32'hc198df3c} /* (17, 24, 2) {real, imag} */,
  {32'h420d1468, 32'hc1d34360} /* (17, 24, 1) {real, imag} */,
  {32'h41773b30, 32'hc1044b34} /* (17, 24, 0) {real, imag} */,
  {32'h4198da5b, 32'h42281a51} /* (17, 23, 31) {real, imag} */,
  {32'hc08d153b, 32'hc0a54723} /* (17, 23, 30) {real, imag} */,
  {32'hc189cd7c, 32'h3f3d12b8} /* (17, 23, 29) {real, imag} */,
  {32'h402e1ac0, 32'h418eff12} /* (17, 23, 28) {real, imag} */,
  {32'hc14210fb, 32'h40585528} /* (17, 23, 27) {real, imag} */,
  {32'hbf0e1b20, 32'hc0ec2828} /* (17, 23, 26) {real, imag} */,
  {32'h402d7d54, 32'h3b65d000} /* (17, 23, 25) {real, imag} */,
  {32'hc0c4eec0, 32'hc0b0efe3} /* (17, 23, 24) {real, imag} */,
  {32'h41799966, 32'hbf991808} /* (17, 23, 23) {real, imag} */,
  {32'hc0b09bec, 32'hc00d69c6} /* (17, 23, 22) {real, imag} */,
  {32'hc199ec52, 32'h4114cfab} /* (17, 23, 21) {real, imag} */,
  {32'hc14ce0ae, 32'h4040ada8} /* (17, 23, 20) {real, imag} */,
  {32'h40bd236a, 32'hc1a863c0} /* (17, 23, 19) {real, imag} */,
  {32'h40388cda, 32'h4155a87f} /* (17, 23, 18) {real, imag} */,
  {32'hc032a35c, 32'hc18435f1} /* (17, 23, 17) {real, imag} */,
  {32'hc09918e8, 32'hc0197d02} /* (17, 23, 16) {real, imag} */,
  {32'hc0f19f4c, 32'hc10ddd42} /* (17, 23, 15) {real, imag} */,
  {32'h40ed8a8b, 32'h41566c2f} /* (17, 23, 14) {real, imag} */,
  {32'hc112c012, 32'hc0978e79} /* (17, 23, 13) {real, imag} */,
  {32'h402a86de, 32'h41adf0fa} /* (17, 23, 12) {real, imag} */,
  {32'h4196fe56, 32'h40533273} /* (17, 23, 11) {real, imag} */,
  {32'hbf813480, 32'h41788e89} /* (17, 23, 10) {real, imag} */,
  {32'hbf836b64, 32'hc10b2c9b} /* (17, 23, 9) {real, imag} */,
  {32'h4138baf2, 32'hc2078aeb} /* (17, 23, 8) {real, imag} */,
  {32'hc0f3f890, 32'hc0b14db8} /* (17, 23, 7) {real, imag} */,
  {32'h3feb3690, 32'hc1c2f3c1} /* (17, 23, 6) {real, imag} */,
  {32'h40e50ac4, 32'hc0cd9ea1} /* (17, 23, 5) {real, imag} */,
  {32'hc17de05c, 32'h4136d576} /* (17, 23, 4) {real, imag} */,
  {32'h41002016, 32'hc10e551f} /* (17, 23, 3) {real, imag} */,
  {32'hc0cc6edd, 32'hc0ad3992} /* (17, 23, 2) {real, imag} */,
  {32'hc0cceeb8, 32'h40ae5b4b} /* (17, 23, 1) {real, imag} */,
  {32'h412f1767, 32'hc053ac8f} /* (17, 23, 0) {real, imag} */,
  {32'hc18fa6c2, 32'hbfacf8a4} /* (17, 22, 31) {real, imag} */,
  {32'h40388076, 32'hc0a547a2} /* (17, 22, 30) {real, imag} */,
  {32'h40cb7de6, 32'h40fb7685} /* (17, 22, 29) {real, imag} */,
  {32'h3fb95c30, 32'h4094ce7c} /* (17, 22, 28) {real, imag} */,
  {32'h40e9b0a4, 32'h40f6a8a3} /* (17, 22, 27) {real, imag} */,
  {32'h40baa6a7, 32'hc00e9be2} /* (17, 22, 26) {real, imag} */,
  {32'hc0cd2042, 32'h3f81d4d8} /* (17, 22, 25) {real, imag} */,
  {32'h3ff3ce9b, 32'hc0ebe44e} /* (17, 22, 24) {real, imag} */,
  {32'h40acb65c, 32'h4105ca6f} /* (17, 22, 23) {real, imag} */,
  {32'hc0859ff2, 32'hc0cb940c} /* (17, 22, 22) {real, imag} */,
  {32'hc1af96b2, 32'hc116a26e} /* (17, 22, 21) {real, imag} */,
  {32'hc1277e70, 32'h40adb817} /* (17, 22, 20) {real, imag} */,
  {32'hbfa91a20, 32'h40d343b5} /* (17, 22, 19) {real, imag} */,
  {32'hc0d5f370, 32'h3fe5c40c} /* (17, 22, 18) {real, imag} */,
  {32'hc1811be2, 32'h3fc07cd4} /* (17, 22, 17) {real, imag} */,
  {32'h40ea7ebf, 32'h40d8a490} /* (17, 22, 16) {real, imag} */,
  {32'h4119d7ec, 32'hbff5f7a1} /* (17, 22, 15) {real, imag} */,
  {32'h411cdc65, 32'hbf8a3280} /* (17, 22, 14) {real, imag} */,
  {32'hbfaad272, 32'h3f625340} /* (17, 22, 13) {real, imag} */,
  {32'hc01a3807, 32'h3f3962f0} /* (17, 22, 12) {real, imag} */,
  {32'h4158b25c, 32'hc12f70b3} /* (17, 22, 11) {real, imag} */,
  {32'hc125bba4, 32'hc15f96c4} /* (17, 22, 10) {real, imag} */,
  {32'hc00a0ac0, 32'h3ff13bf8} /* (17, 22, 9) {real, imag} */,
  {32'h412ee91c, 32'h412caccb} /* (17, 22, 8) {real, imag} */,
  {32'h3ed00878, 32'h406ed1b3} /* (17, 22, 7) {real, imag} */,
  {32'h410f5a86, 32'hc059e5d8} /* (17, 22, 6) {real, imag} */,
  {32'h40f7faf8, 32'h41487f2c} /* (17, 22, 5) {real, imag} */,
  {32'hc0caaec9, 32'hc0b2594e} /* (17, 22, 4) {real, imag} */,
  {32'hc07e838d, 32'h408178df} /* (17, 22, 3) {real, imag} */,
  {32'hbff8e098, 32'hc0b06d2b} /* (17, 22, 2) {real, imag} */,
  {32'hc1110f01, 32'h4087f32a} /* (17, 22, 1) {real, imag} */,
  {32'hbff2ea9c, 32'hc14a36b5} /* (17, 22, 0) {real, imag} */,
  {32'hbff2801e, 32'hc154d49a} /* (17, 21, 31) {real, imag} */,
  {32'h41324fb6, 32'h417599c8} /* (17, 21, 30) {real, imag} */,
  {32'hc09f4d2b, 32'hbee32680} /* (17, 21, 29) {real, imag} */,
  {32'hc1328e41, 32'hc0d4dd6a} /* (17, 21, 28) {real, imag} */,
  {32'hc0b10a90, 32'h419c3618} /* (17, 21, 27) {real, imag} */,
  {32'h3e782a00, 32'hc1a63c00} /* (17, 21, 26) {real, imag} */,
  {32'h40ad3175, 32'h413747b5} /* (17, 21, 25) {real, imag} */,
  {32'hc1447703, 32'h4190c22a} /* (17, 21, 24) {real, imag} */,
  {32'hc13a246c, 32'hc12f0e9e} /* (17, 21, 23) {real, imag} */,
  {32'h418e55f2, 32'hbec5ab98} /* (17, 21, 22) {real, imag} */,
  {32'hc00f27de, 32'h40a0fe62} /* (17, 21, 21) {real, imag} */,
  {32'hc0f9b023, 32'hc0d8a404} /* (17, 21, 20) {real, imag} */,
  {32'h408d9400, 32'h40e268e3} /* (17, 21, 19) {real, imag} */,
  {32'hbf5f3688, 32'h400e6000} /* (17, 21, 18) {real, imag} */,
  {32'h408bebf4, 32'hc14a09c8} /* (17, 21, 17) {real, imag} */,
  {32'hc10a8dcb, 32'h414d4039} /* (17, 21, 16) {real, imag} */,
  {32'h3f99d877, 32'h3eadedd0} /* (17, 21, 15) {real, imag} */,
  {32'hc13f9209, 32'h4066121e} /* (17, 21, 14) {real, imag} */,
  {32'h3f3f65d8, 32'h40dc9527} /* (17, 21, 13) {real, imag} */,
  {32'hc0d4670d, 32'h3fba9a28} /* (17, 21, 12) {real, imag} */,
  {32'hc1a1fd78, 32'h402264ec} /* (17, 21, 11) {real, imag} */,
  {32'hc0b9becc, 32'h3fa95646} /* (17, 21, 10) {real, imag} */,
  {32'hc1540c5d, 32'h414decb1} /* (17, 21, 9) {real, imag} */,
  {32'hc180efde, 32'h40b5cbc5} /* (17, 21, 8) {real, imag} */,
  {32'h3fbd3ca4, 32'h4020099c} /* (17, 21, 7) {real, imag} */,
  {32'hc1299cd2, 32'hc0d27574} /* (17, 21, 6) {real, imag} */,
  {32'hc0602a24, 32'h41900bb5} /* (17, 21, 5) {real, imag} */,
  {32'h41acadd4, 32'hc0e89f4e} /* (17, 21, 4) {real, imag} */,
  {32'hc01afcd4, 32'hc14d3cc9} /* (17, 21, 3) {real, imag} */,
  {32'h4149ad6c, 32'h3fc81ba4} /* (17, 21, 2) {real, imag} */,
  {32'h4100dc11, 32'hc1a8e124} /* (17, 21, 1) {real, imag} */,
  {32'h418f4503, 32'hc15e391e} /* (17, 21, 0) {real, imag} */,
  {32'h408c9bd3, 32'h3f5abd40} /* (17, 20, 31) {real, imag} */,
  {32'h414e66cb, 32'h40cdc575} /* (17, 20, 30) {real, imag} */,
  {32'hc0974c49, 32'hbf486100} /* (17, 20, 29) {real, imag} */,
  {32'hc1581e80, 32'h40ea5f77} /* (17, 20, 28) {real, imag} */,
  {32'hc0044804, 32'h405c6832} /* (17, 20, 27) {real, imag} */,
  {32'h40cfcb68, 32'h40eb6705} /* (17, 20, 26) {real, imag} */,
  {32'hc0ac0e33, 32'h408b3d4e} /* (17, 20, 25) {real, imag} */,
  {32'h41d4b99d, 32'h4111c7c4} /* (17, 20, 24) {real, imag} */,
  {32'hc1515e18, 32'h4101ad04} /* (17, 20, 23) {real, imag} */,
  {32'hc0778612, 32'h40bb4604} /* (17, 20, 22) {real, imag} */,
  {32'h41afcb32, 32'hc00b2c34} /* (17, 20, 21) {real, imag} */,
  {32'hc097f504, 32'h411b02ba} /* (17, 20, 20) {real, imag} */,
  {32'hc0578119, 32'h40da9e42} /* (17, 20, 19) {real, imag} */,
  {32'h412050d4, 32'hc0df58a6} /* (17, 20, 18) {real, imag} */,
  {32'hc087cd1a, 32'hbfcb69da} /* (17, 20, 17) {real, imag} */,
  {32'hc15b3e13, 32'hc082220a} /* (17, 20, 16) {real, imag} */,
  {32'hc0f3db29, 32'h4010e2a4} /* (17, 20, 15) {real, imag} */,
  {32'h40e082ec, 32'h408bcb99} /* (17, 20, 14) {real, imag} */,
  {32'h40633af2, 32'h3f939b08} /* (17, 20, 13) {real, imag} */,
  {32'hc15cae30, 32'hbf72747c} /* (17, 20, 12) {real, imag} */,
  {32'hc0535182, 32'h41bbe6aa} /* (17, 20, 11) {real, imag} */,
  {32'h4166520b, 32'hc14e9606} /* (17, 20, 10) {real, imag} */,
  {32'h4045d9b2, 32'h4116ae00} /* (17, 20, 9) {real, imag} */,
  {32'h415816f0, 32'hc1463ce0} /* (17, 20, 8) {real, imag} */,
  {32'hc0e98e8f, 32'hc105bb29} /* (17, 20, 7) {real, imag} */,
  {32'h4127604a, 32'hc10c6d31} /* (17, 20, 6) {real, imag} */,
  {32'h40455e1d, 32'h40095ad8} /* (17, 20, 5) {real, imag} */,
  {32'h3fd33122, 32'hbde16880} /* (17, 20, 4) {real, imag} */,
  {32'hc11b1de2, 32'hc0fb5b28} /* (17, 20, 3) {real, imag} */,
  {32'h404ad6d8, 32'hbffebe30} /* (17, 20, 2) {real, imag} */,
  {32'hc109324e, 32'h40859769} /* (17, 20, 1) {real, imag} */,
  {32'hc16acf5f, 32'h406a3d4d} /* (17, 20, 0) {real, imag} */,
  {32'hc1be1052, 32'hbe617b00} /* (17, 19, 31) {real, imag} */,
  {32'hc0be6fd4, 32'hc134ef6e} /* (17, 19, 30) {real, imag} */,
  {32'h40b952c8, 32'h40cac8fc} /* (17, 19, 29) {real, imag} */,
  {32'h40c876d9, 32'h419909d6} /* (17, 19, 28) {real, imag} */,
  {32'hc16c1018, 32'hc12b8c44} /* (17, 19, 27) {real, imag} */,
  {32'h417bef96, 32'h410d9675} /* (17, 19, 26) {real, imag} */,
  {32'h3faa3b16, 32'hc0b0ba8d} /* (17, 19, 25) {real, imag} */,
  {32'h41169f2c, 32'hc0fc5f0a} /* (17, 19, 24) {real, imag} */,
  {32'hc1208dab, 32'hc0979400} /* (17, 19, 23) {real, imag} */,
  {32'h414313a0, 32'h3f1451d4} /* (17, 19, 22) {real, imag} */,
  {32'hc15633d4, 32'h41996611} /* (17, 19, 21) {real, imag} */,
  {32'h40a4d978, 32'h40d65c8a} /* (17, 19, 20) {real, imag} */,
  {32'h40a6db87, 32'h3f1d6fe8} /* (17, 19, 19) {real, imag} */,
  {32'hc1c451f6, 32'hbf8267c0} /* (17, 19, 18) {real, imag} */,
  {32'h4144cb66, 32'h409c3fe5} /* (17, 19, 17) {real, imag} */,
  {32'h4040acb6, 32'h416645cb} /* (17, 19, 16) {real, imag} */,
  {32'hbf048c84, 32'hc10f0438} /* (17, 19, 15) {real, imag} */,
  {32'h409aab95, 32'hc0d6ec5c} /* (17, 19, 14) {real, imag} */,
  {32'hc02f3610, 32'hc1368f5e} /* (17, 19, 13) {real, imag} */,
  {32'h405196dc, 32'hc033c7ee} /* (17, 19, 12) {real, imag} */,
  {32'h40684efd, 32'hc1670bc3} /* (17, 19, 11) {real, imag} */,
  {32'hc1104ffb, 32'h40d56177} /* (17, 19, 10) {real, imag} */,
  {32'h40804424, 32'hc0e4d601} /* (17, 19, 9) {real, imag} */,
  {32'hc0653648, 32'h40ecff59} /* (17, 19, 8) {real, imag} */,
  {32'hbf493148, 32'h413218cd} /* (17, 19, 7) {real, imag} */,
  {32'hc0cc7117, 32'h41118d62} /* (17, 19, 6) {real, imag} */,
  {32'h413b7ff4, 32'h416ad9cf} /* (17, 19, 5) {real, imag} */,
  {32'hc1248862, 32'hc0929fc4} /* (17, 19, 4) {real, imag} */,
  {32'hc0aa8b6c, 32'h40e2929f} /* (17, 19, 3) {real, imag} */,
  {32'hc102c924, 32'h40e12d4e} /* (17, 19, 2) {real, imag} */,
  {32'hbff82350, 32'hc1732dbc} /* (17, 19, 1) {real, imag} */,
  {32'h40a3d74e, 32'h40d82467} /* (17, 19, 0) {real, imag} */,
  {32'h40ed0667, 32'hc130c6c2} /* (17, 18, 31) {real, imag} */,
  {32'h40279a74, 32'h3f530870} /* (17, 18, 30) {real, imag} */,
  {32'hc15b4b0b, 32'h412c01ca} /* (17, 18, 29) {real, imag} */,
  {32'h41321590, 32'h41448864} /* (17, 18, 28) {real, imag} */,
  {32'h40ad6630, 32'hc080be6a} /* (17, 18, 27) {real, imag} */,
  {32'h40450325, 32'h40c91538} /* (17, 18, 26) {real, imag} */,
  {32'h41194eca, 32'h3fac8d20} /* (17, 18, 25) {real, imag} */,
  {32'h40f17687, 32'h40ca629f} /* (17, 18, 24) {real, imag} */,
  {32'h4154ea1e, 32'h413d6ff1} /* (17, 18, 23) {real, imag} */,
  {32'hc17088ef, 32'hbf8cfee0} /* (17, 18, 22) {real, imag} */,
  {32'hbf98b7e4, 32'hbe827688} /* (17, 18, 21) {real, imag} */,
  {32'hc026fda2, 32'h403064b0} /* (17, 18, 20) {real, imag} */,
  {32'hc102173a, 32'hbb20a000} /* (17, 18, 19) {real, imag} */,
  {32'h409ceb31, 32'hc18bcb12} /* (17, 18, 18) {real, imag} */,
  {32'hc0adfd30, 32'h41017bea} /* (17, 18, 17) {real, imag} */,
  {32'h40452e56, 32'hc04db3ee} /* (17, 18, 16) {real, imag} */,
  {32'h4007dc44, 32'hc0a0e004} /* (17, 18, 15) {real, imag} */,
  {32'h4138cbb6, 32'h3d8e5010} /* (17, 18, 14) {real, imag} */,
  {32'hc0fd348f, 32'hc0229696} /* (17, 18, 13) {real, imag} */,
  {32'hc0a25da8, 32'hc1126155} /* (17, 18, 12) {real, imag} */,
  {32'hbd71d3c0, 32'hc05afa8e} /* (17, 18, 11) {real, imag} */,
  {32'hbf258e6c, 32'hbf618e0c} /* (17, 18, 10) {real, imag} */,
  {32'h4158cdb4, 32'hbfa5252a} /* (17, 18, 9) {real, imag} */,
  {32'hc0229df6, 32'hbfb4ba26} /* (17, 18, 8) {real, imag} */,
  {32'hc107678e, 32'h3d06dc80} /* (17, 18, 7) {real, imag} */,
  {32'h41179b82, 32'hc08a4d0d} /* (17, 18, 6) {real, imag} */,
  {32'hc113475a, 32'h406a50e3} /* (17, 18, 5) {real, imag} */,
  {32'hbfac0ee4, 32'hc0bdc1bc} /* (17, 18, 4) {real, imag} */,
  {32'h418c9aa0, 32'h40f12a4a} /* (17, 18, 3) {real, imag} */,
  {32'hc113c92d, 32'hbfbaf65a} /* (17, 18, 2) {real, imag} */,
  {32'h410cad42, 32'hc05b3113} /* (17, 18, 1) {real, imag} */,
  {32'hbf2f4e0c, 32'hc1422354} /* (17, 18, 0) {real, imag} */,
  {32'hc0bca8e2, 32'h40fb5a8a} /* (17, 17, 31) {real, imag} */,
  {32'hbff80b84, 32'h410f7e34} /* (17, 17, 30) {real, imag} */,
  {32'h412f1d5a, 32'hc07c75e2} /* (17, 17, 29) {real, imag} */,
  {32'hc1045b82, 32'hbff9c2d8} /* (17, 17, 28) {real, imag} */,
  {32'h40ee596e, 32'hc018bfc0} /* (17, 17, 27) {real, imag} */,
  {32'hc0d07d69, 32'hc1ab83e0} /* (17, 17, 26) {real, imag} */,
  {32'h404d42b7, 32'h41468410} /* (17, 17, 25) {real, imag} */,
  {32'hc0db715d, 32'hc071bf78} /* (17, 17, 24) {real, imag} */,
  {32'hc094baaf, 32'h4151ab7b} /* (17, 17, 23) {real, imag} */,
  {32'hc05449b2, 32'hbffe1262} /* (17, 17, 22) {real, imag} */,
  {32'hc0433d74, 32'h41005223} /* (17, 17, 21) {real, imag} */,
  {32'h40dc69a2, 32'hc13b82b7} /* (17, 17, 20) {real, imag} */,
  {32'h413d5295, 32'hc04a6d2c} /* (17, 17, 19) {real, imag} */,
  {32'h40b19da0, 32'h40fbe7a8} /* (17, 17, 18) {real, imag} */,
  {32'h40bac9aa, 32'h4066cae8} /* (17, 17, 17) {real, imag} */,
  {32'hbba01700, 32'hc0b6763c} /* (17, 17, 16) {real, imag} */,
  {32'hc058f06e, 32'h41525fbe} /* (17, 17, 15) {real, imag} */,
  {32'h410ee659, 32'h3ea56da0} /* (17, 17, 14) {real, imag} */,
  {32'hc0a6f4e4, 32'hc100ddce} /* (17, 17, 13) {real, imag} */,
  {32'h419b78e5, 32'h3f8d6686} /* (17, 17, 12) {real, imag} */,
  {32'hc181ba7b, 32'h4182a412} /* (17, 17, 11) {real, imag} */,
  {32'h400c9224, 32'hc13c7caa} /* (17, 17, 10) {real, imag} */,
  {32'hc0a1f79f, 32'hc10a9d60} /* (17, 17, 9) {real, imag} */,
  {32'h4159017b, 32'hc0801d84} /* (17, 17, 8) {real, imag} */,
  {32'h4108ab06, 32'h3f9f537c} /* (17, 17, 7) {real, imag} */,
  {32'hc134ea22, 32'h40dcd3b6} /* (17, 17, 6) {real, imag} */,
  {32'h410d91c2, 32'hc0250d3a} /* (17, 17, 5) {real, imag} */,
  {32'hbfa15940, 32'h4085a064} /* (17, 17, 4) {real, imag} */,
  {32'hbfc0fdb0, 32'hc0318fbc} /* (17, 17, 3) {real, imag} */,
  {32'hc1085406, 32'hc1397d34} /* (17, 17, 2) {real, imag} */,
  {32'h40cac849, 32'h413d4283} /* (17, 17, 1) {real, imag} */,
  {32'h4142f7eb, 32'h4012f6a5} /* (17, 17, 0) {real, imag} */,
  {32'h40aed0ab, 32'hc129c1f9} /* (17, 16, 31) {real, imag} */,
  {32'hbf4ea908, 32'hc02040ec} /* (17, 16, 30) {real, imag} */,
  {32'hc085a32c, 32'hc09ff758} /* (17, 16, 29) {real, imag} */,
  {32'hbe07cbc0, 32'hc12b8cdd} /* (17, 16, 28) {real, imag} */,
  {32'hc052e95f, 32'hc0fa5344} /* (17, 16, 27) {real, imag} */,
  {32'h40cef036, 32'h4135d13c} /* (17, 16, 26) {real, imag} */,
  {32'hc0c40955, 32'h3f948c04} /* (17, 16, 25) {real, imag} */,
  {32'h404f15af, 32'hc0913aaa} /* (17, 16, 24) {real, imag} */,
  {32'hc090e126, 32'h3e819e30} /* (17, 16, 23) {real, imag} */,
  {32'h3ffa9095, 32'hc089bebc} /* (17, 16, 22) {real, imag} */,
  {32'hc0261b84, 32'h4115ba92} /* (17, 16, 21) {real, imag} */,
  {32'hbdfe10c0, 32'h413ae6a8} /* (17, 16, 20) {real, imag} */,
  {32'hc08fc8ee, 32'hbf3ecb1c} /* (17, 16, 19) {real, imag} */,
  {32'h402999f8, 32'hc0d3fba1} /* (17, 16, 18) {real, imag} */,
  {32'hc1611614, 32'h41080314} /* (17, 16, 17) {real, imag} */,
  {32'hc034025c, 32'h00000000} /* (17, 16, 16) {real, imag} */,
  {32'hc1611614, 32'hc1080314} /* (17, 16, 15) {real, imag} */,
  {32'h402999f8, 32'h40d3fba1} /* (17, 16, 14) {real, imag} */,
  {32'hc08fc8ee, 32'h3f3ecb1c} /* (17, 16, 13) {real, imag} */,
  {32'hbdfe10c0, 32'hc13ae6a8} /* (17, 16, 12) {real, imag} */,
  {32'hc0261b84, 32'hc115ba92} /* (17, 16, 11) {real, imag} */,
  {32'h3ffa9095, 32'h4089bebc} /* (17, 16, 10) {real, imag} */,
  {32'hc090e126, 32'hbe819e30} /* (17, 16, 9) {real, imag} */,
  {32'h404f15af, 32'h40913aaa} /* (17, 16, 8) {real, imag} */,
  {32'hc0c40955, 32'hbf948c04} /* (17, 16, 7) {real, imag} */,
  {32'h40cef036, 32'hc135d13c} /* (17, 16, 6) {real, imag} */,
  {32'hc052e95f, 32'h40fa5344} /* (17, 16, 5) {real, imag} */,
  {32'hbe07cbc0, 32'h412b8cdd} /* (17, 16, 4) {real, imag} */,
  {32'hc085a32c, 32'h409ff758} /* (17, 16, 3) {real, imag} */,
  {32'hbf4ea908, 32'h402040ec} /* (17, 16, 2) {real, imag} */,
  {32'h40aed0ab, 32'h4129c1f9} /* (17, 16, 1) {real, imag} */,
  {32'hc096b4c2, 32'h00000000} /* (17, 16, 0) {real, imag} */,
  {32'h40cac849, 32'hc13d4283} /* (17, 15, 31) {real, imag} */,
  {32'hc1085406, 32'h41397d34} /* (17, 15, 30) {real, imag} */,
  {32'hbfc0fdb0, 32'h40318fbc} /* (17, 15, 29) {real, imag} */,
  {32'hbfa15940, 32'hc085a064} /* (17, 15, 28) {real, imag} */,
  {32'h410d91c2, 32'h40250d3a} /* (17, 15, 27) {real, imag} */,
  {32'hc134ea22, 32'hc0dcd3b6} /* (17, 15, 26) {real, imag} */,
  {32'h4108ab06, 32'hbf9f537c} /* (17, 15, 25) {real, imag} */,
  {32'h4159017b, 32'h40801d84} /* (17, 15, 24) {real, imag} */,
  {32'hc0a1f79f, 32'h410a9d60} /* (17, 15, 23) {real, imag} */,
  {32'h400c9224, 32'h413c7caa} /* (17, 15, 22) {real, imag} */,
  {32'hc181ba7b, 32'hc182a412} /* (17, 15, 21) {real, imag} */,
  {32'h419b78e5, 32'hbf8d6686} /* (17, 15, 20) {real, imag} */,
  {32'hc0a6f4e4, 32'h4100ddce} /* (17, 15, 19) {real, imag} */,
  {32'h410ee659, 32'hbea56da0} /* (17, 15, 18) {real, imag} */,
  {32'hc058f06e, 32'hc1525fbe} /* (17, 15, 17) {real, imag} */,
  {32'hbba01700, 32'h40b6763c} /* (17, 15, 16) {real, imag} */,
  {32'h40bac9aa, 32'hc066cae8} /* (17, 15, 15) {real, imag} */,
  {32'h40b19da0, 32'hc0fbe7a8} /* (17, 15, 14) {real, imag} */,
  {32'h413d5295, 32'h404a6d2c} /* (17, 15, 13) {real, imag} */,
  {32'h40dc69a2, 32'h413b82b7} /* (17, 15, 12) {real, imag} */,
  {32'hc0433d74, 32'hc1005223} /* (17, 15, 11) {real, imag} */,
  {32'hc05449b2, 32'h3ffe1262} /* (17, 15, 10) {real, imag} */,
  {32'hc094baaf, 32'hc151ab7b} /* (17, 15, 9) {real, imag} */,
  {32'hc0db715d, 32'h4071bf78} /* (17, 15, 8) {real, imag} */,
  {32'h404d42b7, 32'hc1468410} /* (17, 15, 7) {real, imag} */,
  {32'hc0d07d69, 32'h41ab83e0} /* (17, 15, 6) {real, imag} */,
  {32'h40ee596e, 32'h4018bfc0} /* (17, 15, 5) {real, imag} */,
  {32'hc1045b82, 32'h3ff9c2d8} /* (17, 15, 4) {real, imag} */,
  {32'h412f1d5a, 32'h407c75e2} /* (17, 15, 3) {real, imag} */,
  {32'hbff80b84, 32'hc10f7e34} /* (17, 15, 2) {real, imag} */,
  {32'hc0bca8e2, 32'hc0fb5a8a} /* (17, 15, 1) {real, imag} */,
  {32'h4142f7eb, 32'hc012f6a5} /* (17, 15, 0) {real, imag} */,
  {32'h410cad42, 32'h405b3113} /* (17, 14, 31) {real, imag} */,
  {32'hc113c92d, 32'h3fbaf65a} /* (17, 14, 30) {real, imag} */,
  {32'h418c9aa0, 32'hc0f12a4a} /* (17, 14, 29) {real, imag} */,
  {32'hbfac0ee4, 32'h40bdc1bc} /* (17, 14, 28) {real, imag} */,
  {32'hc113475a, 32'hc06a50e3} /* (17, 14, 27) {real, imag} */,
  {32'h41179b82, 32'h408a4d0d} /* (17, 14, 26) {real, imag} */,
  {32'hc107678e, 32'hbd06dc80} /* (17, 14, 25) {real, imag} */,
  {32'hc0229df6, 32'h3fb4ba26} /* (17, 14, 24) {real, imag} */,
  {32'h4158cdb4, 32'h3fa5252a} /* (17, 14, 23) {real, imag} */,
  {32'hbf258e6c, 32'h3f618e0c} /* (17, 14, 22) {real, imag} */,
  {32'hbd71d3c0, 32'h405afa8e} /* (17, 14, 21) {real, imag} */,
  {32'hc0a25da8, 32'h41126155} /* (17, 14, 20) {real, imag} */,
  {32'hc0fd348f, 32'h40229696} /* (17, 14, 19) {real, imag} */,
  {32'h4138cbb6, 32'hbd8e5010} /* (17, 14, 18) {real, imag} */,
  {32'h4007dc44, 32'h40a0e004} /* (17, 14, 17) {real, imag} */,
  {32'h40452e56, 32'h404db3ee} /* (17, 14, 16) {real, imag} */,
  {32'hc0adfd30, 32'hc1017bea} /* (17, 14, 15) {real, imag} */,
  {32'h409ceb31, 32'h418bcb12} /* (17, 14, 14) {real, imag} */,
  {32'hc102173a, 32'h3b20a000} /* (17, 14, 13) {real, imag} */,
  {32'hc026fda2, 32'hc03064b0} /* (17, 14, 12) {real, imag} */,
  {32'hbf98b7e4, 32'h3e827688} /* (17, 14, 11) {real, imag} */,
  {32'hc17088ef, 32'h3f8cfee0} /* (17, 14, 10) {real, imag} */,
  {32'h4154ea1e, 32'hc13d6ff1} /* (17, 14, 9) {real, imag} */,
  {32'h40f17687, 32'hc0ca629f} /* (17, 14, 8) {real, imag} */,
  {32'h41194eca, 32'hbfac8d20} /* (17, 14, 7) {real, imag} */,
  {32'h40450325, 32'hc0c91538} /* (17, 14, 6) {real, imag} */,
  {32'h40ad6630, 32'h4080be6a} /* (17, 14, 5) {real, imag} */,
  {32'h41321590, 32'hc1448864} /* (17, 14, 4) {real, imag} */,
  {32'hc15b4b0b, 32'hc12c01ca} /* (17, 14, 3) {real, imag} */,
  {32'h40279a74, 32'hbf530870} /* (17, 14, 2) {real, imag} */,
  {32'h40ed0667, 32'h4130c6c2} /* (17, 14, 1) {real, imag} */,
  {32'hbf2f4e0c, 32'h41422354} /* (17, 14, 0) {real, imag} */,
  {32'hbff82350, 32'h41732dbc} /* (17, 13, 31) {real, imag} */,
  {32'hc102c924, 32'hc0e12d4e} /* (17, 13, 30) {real, imag} */,
  {32'hc0aa8b6c, 32'hc0e2929f} /* (17, 13, 29) {real, imag} */,
  {32'hc1248862, 32'h40929fc4} /* (17, 13, 28) {real, imag} */,
  {32'h413b7ff4, 32'hc16ad9cf} /* (17, 13, 27) {real, imag} */,
  {32'hc0cc7117, 32'hc1118d62} /* (17, 13, 26) {real, imag} */,
  {32'hbf493148, 32'hc13218cd} /* (17, 13, 25) {real, imag} */,
  {32'hc0653648, 32'hc0ecff59} /* (17, 13, 24) {real, imag} */,
  {32'h40804424, 32'h40e4d601} /* (17, 13, 23) {real, imag} */,
  {32'hc1104ffb, 32'hc0d56177} /* (17, 13, 22) {real, imag} */,
  {32'h40684efd, 32'h41670bc3} /* (17, 13, 21) {real, imag} */,
  {32'h405196dc, 32'h4033c7ee} /* (17, 13, 20) {real, imag} */,
  {32'hc02f3610, 32'h41368f5e} /* (17, 13, 19) {real, imag} */,
  {32'h409aab95, 32'h40d6ec5c} /* (17, 13, 18) {real, imag} */,
  {32'hbf048c84, 32'h410f0438} /* (17, 13, 17) {real, imag} */,
  {32'h4040acb6, 32'hc16645cb} /* (17, 13, 16) {real, imag} */,
  {32'h4144cb66, 32'hc09c3fe5} /* (17, 13, 15) {real, imag} */,
  {32'hc1c451f6, 32'h3f8267c0} /* (17, 13, 14) {real, imag} */,
  {32'h40a6db87, 32'hbf1d6fe8} /* (17, 13, 13) {real, imag} */,
  {32'h40a4d978, 32'hc0d65c8a} /* (17, 13, 12) {real, imag} */,
  {32'hc15633d4, 32'hc1996611} /* (17, 13, 11) {real, imag} */,
  {32'h414313a0, 32'hbf1451d4} /* (17, 13, 10) {real, imag} */,
  {32'hc1208dab, 32'h40979400} /* (17, 13, 9) {real, imag} */,
  {32'h41169f2c, 32'h40fc5f0a} /* (17, 13, 8) {real, imag} */,
  {32'h3faa3b16, 32'h40b0ba8d} /* (17, 13, 7) {real, imag} */,
  {32'h417bef96, 32'hc10d9675} /* (17, 13, 6) {real, imag} */,
  {32'hc16c1018, 32'h412b8c44} /* (17, 13, 5) {real, imag} */,
  {32'h40c876d9, 32'hc19909d6} /* (17, 13, 4) {real, imag} */,
  {32'h40b952c8, 32'hc0cac8fc} /* (17, 13, 3) {real, imag} */,
  {32'hc0be6fd4, 32'h4134ef6e} /* (17, 13, 2) {real, imag} */,
  {32'hc1be1052, 32'h3e617b00} /* (17, 13, 1) {real, imag} */,
  {32'h40a3d74e, 32'hc0d82467} /* (17, 13, 0) {real, imag} */,
  {32'hc109324e, 32'hc0859769} /* (17, 12, 31) {real, imag} */,
  {32'h404ad6d8, 32'h3ffebe30} /* (17, 12, 30) {real, imag} */,
  {32'hc11b1de2, 32'h40fb5b28} /* (17, 12, 29) {real, imag} */,
  {32'h3fd33122, 32'h3de16880} /* (17, 12, 28) {real, imag} */,
  {32'h40455e1d, 32'hc0095ad8} /* (17, 12, 27) {real, imag} */,
  {32'h4127604a, 32'h410c6d31} /* (17, 12, 26) {real, imag} */,
  {32'hc0e98e8f, 32'h4105bb29} /* (17, 12, 25) {real, imag} */,
  {32'h415816f0, 32'h41463ce0} /* (17, 12, 24) {real, imag} */,
  {32'h4045d9b2, 32'hc116ae00} /* (17, 12, 23) {real, imag} */,
  {32'h4166520b, 32'h414e9606} /* (17, 12, 22) {real, imag} */,
  {32'hc0535182, 32'hc1bbe6aa} /* (17, 12, 21) {real, imag} */,
  {32'hc15cae30, 32'h3f72747c} /* (17, 12, 20) {real, imag} */,
  {32'h40633af2, 32'hbf939b08} /* (17, 12, 19) {real, imag} */,
  {32'h40e082ec, 32'hc08bcb99} /* (17, 12, 18) {real, imag} */,
  {32'hc0f3db29, 32'hc010e2a4} /* (17, 12, 17) {real, imag} */,
  {32'hc15b3e13, 32'h4082220a} /* (17, 12, 16) {real, imag} */,
  {32'hc087cd1a, 32'h3fcb69da} /* (17, 12, 15) {real, imag} */,
  {32'h412050d4, 32'h40df58a6} /* (17, 12, 14) {real, imag} */,
  {32'hc0578119, 32'hc0da9e42} /* (17, 12, 13) {real, imag} */,
  {32'hc097f504, 32'hc11b02ba} /* (17, 12, 12) {real, imag} */,
  {32'h41afcb32, 32'h400b2c34} /* (17, 12, 11) {real, imag} */,
  {32'hc0778612, 32'hc0bb4604} /* (17, 12, 10) {real, imag} */,
  {32'hc1515e18, 32'hc101ad04} /* (17, 12, 9) {real, imag} */,
  {32'h41d4b99d, 32'hc111c7c4} /* (17, 12, 8) {real, imag} */,
  {32'hc0ac0e33, 32'hc08b3d4e} /* (17, 12, 7) {real, imag} */,
  {32'h40cfcb68, 32'hc0eb6705} /* (17, 12, 6) {real, imag} */,
  {32'hc0044804, 32'hc05c6832} /* (17, 12, 5) {real, imag} */,
  {32'hc1581e80, 32'hc0ea5f77} /* (17, 12, 4) {real, imag} */,
  {32'hc0974c49, 32'h3f486100} /* (17, 12, 3) {real, imag} */,
  {32'h414e66cb, 32'hc0cdc575} /* (17, 12, 2) {real, imag} */,
  {32'h408c9bd3, 32'hbf5abd40} /* (17, 12, 1) {real, imag} */,
  {32'hc16acf5f, 32'hc06a3d4d} /* (17, 12, 0) {real, imag} */,
  {32'h4100dc11, 32'h41a8e124} /* (17, 11, 31) {real, imag} */,
  {32'h4149ad6c, 32'hbfc81ba4} /* (17, 11, 30) {real, imag} */,
  {32'hc01afcd4, 32'h414d3cc9} /* (17, 11, 29) {real, imag} */,
  {32'h41acadd4, 32'h40e89f4e} /* (17, 11, 28) {real, imag} */,
  {32'hc0602a24, 32'hc1900bb5} /* (17, 11, 27) {real, imag} */,
  {32'hc1299cd2, 32'h40d27574} /* (17, 11, 26) {real, imag} */,
  {32'h3fbd3ca4, 32'hc020099c} /* (17, 11, 25) {real, imag} */,
  {32'hc180efde, 32'hc0b5cbc5} /* (17, 11, 24) {real, imag} */,
  {32'hc1540c5d, 32'hc14decb1} /* (17, 11, 23) {real, imag} */,
  {32'hc0b9becc, 32'hbfa95646} /* (17, 11, 22) {real, imag} */,
  {32'hc1a1fd78, 32'hc02264ec} /* (17, 11, 21) {real, imag} */,
  {32'hc0d4670d, 32'hbfba9a28} /* (17, 11, 20) {real, imag} */,
  {32'h3f3f65d8, 32'hc0dc9527} /* (17, 11, 19) {real, imag} */,
  {32'hc13f9209, 32'hc066121e} /* (17, 11, 18) {real, imag} */,
  {32'h3f99d877, 32'hbeadedd0} /* (17, 11, 17) {real, imag} */,
  {32'hc10a8dcb, 32'hc14d4039} /* (17, 11, 16) {real, imag} */,
  {32'h408bebf4, 32'h414a09c8} /* (17, 11, 15) {real, imag} */,
  {32'hbf5f3688, 32'hc00e6000} /* (17, 11, 14) {real, imag} */,
  {32'h408d9400, 32'hc0e268e3} /* (17, 11, 13) {real, imag} */,
  {32'hc0f9b023, 32'h40d8a404} /* (17, 11, 12) {real, imag} */,
  {32'hc00f27de, 32'hc0a0fe62} /* (17, 11, 11) {real, imag} */,
  {32'h418e55f2, 32'h3ec5ab98} /* (17, 11, 10) {real, imag} */,
  {32'hc13a246c, 32'h412f0e9e} /* (17, 11, 9) {real, imag} */,
  {32'hc1447703, 32'hc190c22a} /* (17, 11, 8) {real, imag} */,
  {32'h40ad3175, 32'hc13747b5} /* (17, 11, 7) {real, imag} */,
  {32'h3e782a00, 32'h41a63c00} /* (17, 11, 6) {real, imag} */,
  {32'hc0b10a90, 32'hc19c3618} /* (17, 11, 5) {real, imag} */,
  {32'hc1328e41, 32'h40d4dd6a} /* (17, 11, 4) {real, imag} */,
  {32'hc09f4d2b, 32'h3ee32680} /* (17, 11, 3) {real, imag} */,
  {32'h41324fb6, 32'hc17599c8} /* (17, 11, 2) {real, imag} */,
  {32'hbff2801e, 32'h4154d49a} /* (17, 11, 1) {real, imag} */,
  {32'h418f4503, 32'h415e391e} /* (17, 11, 0) {real, imag} */,
  {32'hc1110f01, 32'hc087f32a} /* (17, 10, 31) {real, imag} */,
  {32'hbff8e098, 32'h40b06d2b} /* (17, 10, 30) {real, imag} */,
  {32'hc07e838d, 32'hc08178df} /* (17, 10, 29) {real, imag} */,
  {32'hc0caaec9, 32'h40b2594e} /* (17, 10, 28) {real, imag} */,
  {32'h40f7faf8, 32'hc1487f2c} /* (17, 10, 27) {real, imag} */,
  {32'h410f5a86, 32'h4059e5d8} /* (17, 10, 26) {real, imag} */,
  {32'h3ed00878, 32'hc06ed1b3} /* (17, 10, 25) {real, imag} */,
  {32'h412ee91c, 32'hc12caccb} /* (17, 10, 24) {real, imag} */,
  {32'hc00a0ac0, 32'hbff13bf8} /* (17, 10, 23) {real, imag} */,
  {32'hc125bba4, 32'h415f96c4} /* (17, 10, 22) {real, imag} */,
  {32'h4158b25c, 32'h412f70b3} /* (17, 10, 21) {real, imag} */,
  {32'hc01a3807, 32'hbf3962f0} /* (17, 10, 20) {real, imag} */,
  {32'hbfaad272, 32'hbf625340} /* (17, 10, 19) {real, imag} */,
  {32'h411cdc65, 32'h3f8a3280} /* (17, 10, 18) {real, imag} */,
  {32'h4119d7ec, 32'h3ff5f7a1} /* (17, 10, 17) {real, imag} */,
  {32'h40ea7ebf, 32'hc0d8a490} /* (17, 10, 16) {real, imag} */,
  {32'hc1811be2, 32'hbfc07cd4} /* (17, 10, 15) {real, imag} */,
  {32'hc0d5f370, 32'hbfe5c40c} /* (17, 10, 14) {real, imag} */,
  {32'hbfa91a20, 32'hc0d343b5} /* (17, 10, 13) {real, imag} */,
  {32'hc1277e70, 32'hc0adb817} /* (17, 10, 12) {real, imag} */,
  {32'hc1af96b2, 32'h4116a26e} /* (17, 10, 11) {real, imag} */,
  {32'hc0859ff2, 32'h40cb940c} /* (17, 10, 10) {real, imag} */,
  {32'h40acb65c, 32'hc105ca6f} /* (17, 10, 9) {real, imag} */,
  {32'h3ff3ce9b, 32'h40ebe44e} /* (17, 10, 8) {real, imag} */,
  {32'hc0cd2042, 32'hbf81d4d8} /* (17, 10, 7) {real, imag} */,
  {32'h40baa6a7, 32'h400e9be2} /* (17, 10, 6) {real, imag} */,
  {32'h40e9b0a4, 32'hc0f6a8a3} /* (17, 10, 5) {real, imag} */,
  {32'h3fb95c30, 32'hc094ce7c} /* (17, 10, 4) {real, imag} */,
  {32'h40cb7de6, 32'hc0fb7685} /* (17, 10, 3) {real, imag} */,
  {32'h40388076, 32'h40a547a2} /* (17, 10, 2) {real, imag} */,
  {32'hc18fa6c2, 32'h3facf8a4} /* (17, 10, 1) {real, imag} */,
  {32'hbff2ea9c, 32'h414a36b5} /* (17, 10, 0) {real, imag} */,
  {32'hc0cceeb8, 32'hc0ae5b4b} /* (17, 9, 31) {real, imag} */,
  {32'hc0cc6edd, 32'h40ad3992} /* (17, 9, 30) {real, imag} */,
  {32'h41002016, 32'h410e551f} /* (17, 9, 29) {real, imag} */,
  {32'hc17de05c, 32'hc136d576} /* (17, 9, 28) {real, imag} */,
  {32'h40e50ac4, 32'h40cd9ea1} /* (17, 9, 27) {real, imag} */,
  {32'h3feb3690, 32'h41c2f3c1} /* (17, 9, 26) {real, imag} */,
  {32'hc0f3f890, 32'h40b14db8} /* (17, 9, 25) {real, imag} */,
  {32'h4138baf2, 32'h42078aeb} /* (17, 9, 24) {real, imag} */,
  {32'hbf836b64, 32'h410b2c9b} /* (17, 9, 23) {real, imag} */,
  {32'hbf813480, 32'hc1788e89} /* (17, 9, 22) {real, imag} */,
  {32'h4196fe56, 32'hc0533273} /* (17, 9, 21) {real, imag} */,
  {32'h402a86de, 32'hc1adf0fa} /* (17, 9, 20) {real, imag} */,
  {32'hc112c012, 32'h40978e79} /* (17, 9, 19) {real, imag} */,
  {32'h40ed8a8b, 32'hc1566c2f} /* (17, 9, 18) {real, imag} */,
  {32'hc0f19f4c, 32'h410ddd42} /* (17, 9, 17) {real, imag} */,
  {32'hc09918e8, 32'h40197d02} /* (17, 9, 16) {real, imag} */,
  {32'hc032a35c, 32'h418435f1} /* (17, 9, 15) {real, imag} */,
  {32'h40388cda, 32'hc155a87f} /* (17, 9, 14) {real, imag} */,
  {32'h40bd236a, 32'h41a863c0} /* (17, 9, 13) {real, imag} */,
  {32'hc14ce0ae, 32'hc040ada8} /* (17, 9, 12) {real, imag} */,
  {32'hc199ec52, 32'hc114cfab} /* (17, 9, 11) {real, imag} */,
  {32'hc0b09bec, 32'h400d69c6} /* (17, 9, 10) {real, imag} */,
  {32'h41799966, 32'h3f991808} /* (17, 9, 9) {real, imag} */,
  {32'hc0c4eec0, 32'h40b0efe3} /* (17, 9, 8) {real, imag} */,
  {32'h402d7d54, 32'hbb65d000} /* (17, 9, 7) {real, imag} */,
  {32'hbf0e1b20, 32'h40ec2828} /* (17, 9, 6) {real, imag} */,
  {32'hc14210fb, 32'hc0585528} /* (17, 9, 5) {real, imag} */,
  {32'h402e1ac0, 32'hc18eff12} /* (17, 9, 4) {real, imag} */,
  {32'hc189cd7c, 32'hbf3d12b8} /* (17, 9, 3) {real, imag} */,
  {32'hc08d153b, 32'h40a54723} /* (17, 9, 2) {real, imag} */,
  {32'h4198da5b, 32'hc2281a51} /* (17, 9, 1) {real, imag} */,
  {32'h412f1767, 32'h4053ac8f} /* (17, 9, 0) {real, imag} */,
  {32'h420d1468, 32'h41d34360} /* (17, 8, 31) {real, imag} */,
  {32'hc214bc10, 32'h4198df3c} /* (17, 8, 30) {real, imag} */,
  {32'hbf97a4b8, 32'hc13f32e1} /* (17, 8, 29) {real, imag} */,
  {32'h413bb5cf, 32'h40879bc4} /* (17, 8, 28) {real, imag} */,
  {32'h407dc456, 32'hc102f736} /* (17, 8, 27) {real, imag} */,
  {32'hc1266aad, 32'hbf8f2d20} /* (17, 8, 26) {real, imag} */,
  {32'h40868c50, 32'h40c993a6} /* (17, 8, 25) {real, imag} */,
  {32'hc200aa9b, 32'h40b80978} /* (17, 8, 24) {real, imag} */,
  {32'h40dac23a, 32'h40fc370a} /* (17, 8, 23) {real, imag} */,
  {32'hc0899b3c, 32'hc180d8d6} /* (17, 8, 22) {real, imag} */,
  {32'hc12855cd, 32'h4100491f} /* (17, 8, 21) {real, imag} */,
  {32'h4013278c, 32'h41035490} /* (17, 8, 20) {real, imag} */,
  {32'hbf96165c, 32'hbfa933ea} /* (17, 8, 19) {real, imag} */,
  {32'h4041a8ad, 32'h410ea972} /* (17, 8, 18) {real, imag} */,
  {32'hc08e1725, 32'h40b18f24} /* (17, 8, 17) {real, imag} */,
  {32'h411e2791, 32'hc07bcc8e} /* (17, 8, 16) {real, imag} */,
  {32'hc06c6594, 32'hbd74cac0} /* (17, 8, 15) {real, imag} */,
  {32'h40004c33, 32'hc113c6d4} /* (17, 8, 14) {real, imag} */,
  {32'hc1022c74, 32'h40cfe76a} /* (17, 8, 13) {real, imag} */,
  {32'h41810d72, 32'h4150abe0} /* (17, 8, 12) {real, imag} */,
  {32'h4102b87e, 32'h3f0a9212} /* (17, 8, 11) {real, imag} */,
  {32'hc030ee0c, 32'h40af83d2} /* (17, 8, 10) {real, imag} */,
  {32'h413b2c56, 32'h407ca8a8} /* (17, 8, 9) {real, imag} */,
  {32'h40bb8bc0, 32'hc17a636e} /* (17, 8, 8) {real, imag} */,
  {32'hc119ae6f, 32'h415e18c8} /* (17, 8, 7) {real, imag} */,
  {32'hc0e67990, 32'h40567dc8} /* (17, 8, 6) {real, imag} */,
  {32'hbfd84030, 32'h41669dc0} /* (17, 8, 5) {real, imag} */,
  {32'h420c2766, 32'h408dfe6b} /* (17, 8, 4) {real, imag} */,
  {32'hc0a060ec, 32'h41cd3f04} /* (17, 8, 3) {real, imag} */,
  {32'hc1aa00ee, 32'hc18a558c} /* (17, 8, 2) {real, imag} */,
  {32'h414dd8a0, 32'h415cee6c} /* (17, 8, 1) {real, imag} */,
  {32'h41773b30, 32'h41044b34} /* (17, 8, 0) {real, imag} */,
  {32'hc0c306d4, 32'h405d9518} /* (17, 7, 31) {real, imag} */,
  {32'h42128712, 32'hc138a2b3} /* (17, 7, 30) {real, imag} */,
  {32'hc081af26, 32'h402c7d13} /* (17, 7, 29) {real, imag} */,
  {32'hc0ce81b4, 32'h41b440e0} /* (17, 7, 28) {real, imag} */,
  {32'hc17ce140, 32'hc0f574e4} /* (17, 7, 27) {real, imag} */,
  {32'hc1a202aa, 32'hc08be56c} /* (17, 7, 26) {real, imag} */,
  {32'hbfe4f840, 32'hc168819b} /* (17, 7, 25) {real, imag} */,
  {32'hbfad47c4, 32'h3fec9560} /* (17, 7, 24) {real, imag} */,
  {32'hbfb8e294, 32'h414162b1} /* (17, 7, 23) {real, imag} */,
  {32'h4180cf70, 32'h4120d1c0} /* (17, 7, 22) {real, imag} */,
  {32'h417ef63c, 32'h415c15f4} /* (17, 7, 21) {real, imag} */,
  {32'h408c5b15, 32'hc0222e3d} /* (17, 7, 20) {real, imag} */,
  {32'h40b4fda5, 32'h40ac22c6} /* (17, 7, 19) {real, imag} */,
  {32'hbe72a660, 32'hc11f8c56} /* (17, 7, 18) {real, imag} */,
  {32'hc084ceb0, 32'hc1290fe5} /* (17, 7, 17) {real, imag} */,
  {32'h413b7d54, 32'h4175c08d} /* (17, 7, 16) {real, imag} */,
  {32'h40e334c6, 32'hbf16d614} /* (17, 7, 15) {real, imag} */,
  {32'hc12ba945, 32'h4043fee1} /* (17, 7, 14) {real, imag} */,
  {32'hc072bbff, 32'hc10825d2} /* (17, 7, 13) {real, imag} */,
  {32'h3f63693f, 32'h41184337} /* (17, 7, 12) {real, imag} */,
  {32'h4107033d, 32'hc09d59a7} /* (17, 7, 11) {real, imag} */,
  {32'hc0d8cdf1, 32'hc0d4c8af} /* (17, 7, 10) {real, imag} */,
  {32'h4078df06, 32'h41991d74} /* (17, 7, 9) {real, imag} */,
  {32'hc09af406, 32'hc1168f58} /* (17, 7, 8) {real, imag} */,
  {32'h4048af70, 32'h3e6f15e0} /* (17, 7, 7) {real, imag} */,
  {32'h3fbbdd50, 32'hc1e220a0} /* (17, 7, 6) {real, imag} */,
  {32'hc13fece6, 32'hc10e8190} /* (17, 7, 5) {real, imag} */,
  {32'h41c1ce0c, 32'h40b50339} /* (17, 7, 4) {real, imag} */,
  {32'hc1597566, 32'hbef6a980} /* (17, 7, 3) {real, imag} */,
  {32'hc10ebeae, 32'h40b16189} /* (17, 7, 2) {real, imag} */,
  {32'hc0a21d4c, 32'hc0cea690} /* (17, 7, 1) {real, imag} */,
  {32'hc128a444, 32'h41adcd86} /* (17, 7, 0) {real, imag} */,
  {32'h41d47d58, 32'h40af9170} /* (17, 6, 31) {real, imag} */,
  {32'hc1c0960e, 32'hc0d70cfb} /* (17, 6, 30) {real, imag} */,
  {32'hbe4afc70, 32'hc20252a7} /* (17, 6, 29) {real, imag} */,
  {32'hc089a4bb, 32'h41799f9f} /* (17, 6, 28) {real, imag} */,
  {32'hc0c61f40, 32'hc14ab8e0} /* (17, 6, 27) {real, imag} */,
  {32'h418258de, 32'h4021d861} /* (17, 6, 26) {real, imag} */,
  {32'h412cca39, 32'h414b0fe8} /* (17, 6, 25) {real, imag} */,
  {32'hc13bb20f, 32'hc0564e42} /* (17, 6, 24) {real, imag} */,
  {32'h41189e84, 32'hc0f1d3dc} /* (17, 6, 23) {real, imag} */,
  {32'hc16a9c85, 32'h411d64d6} /* (17, 6, 22) {real, imag} */,
  {32'h40e69aeb, 32'hbfa19564} /* (17, 6, 21) {real, imag} */,
  {32'h3f6f84b0, 32'h3f81144f} /* (17, 6, 20) {real, imag} */,
  {32'hc02a7715, 32'hc07e474b} /* (17, 6, 19) {real, imag} */,
  {32'h411a0c3a, 32'h417cdda0} /* (17, 6, 18) {real, imag} */,
  {32'hbf35d0c0, 32'h411a1159} /* (17, 6, 17) {real, imag} */,
  {32'hbf1d27c0, 32'hc0ca5d24} /* (17, 6, 16) {real, imag} */,
  {32'hc13017bf, 32'hc0d6c220} /* (17, 6, 15) {real, imag} */,
  {32'hbfec8da4, 32'hc18a70fb} /* (17, 6, 14) {real, imag} */,
  {32'h405797f8, 32'hc16f3ecf} /* (17, 6, 13) {real, imag} */,
  {32'h412c306e, 32'hc0c64b40} /* (17, 6, 12) {real, imag} */,
  {32'h40a57003, 32'h4109045d} /* (17, 6, 11) {real, imag} */,
  {32'hc1b5e78a, 32'hc0eab484} /* (17, 6, 10) {real, imag} */,
  {32'h41943509, 32'hc1589656} /* (17, 6, 9) {real, imag} */,
  {32'hc2076142, 32'hc0a9f186} /* (17, 6, 8) {real, imag} */,
  {32'h41c61766, 32'h40231105} /* (17, 6, 7) {real, imag} */,
  {32'hc082fb68, 32'h3fc0043c} /* (17, 6, 6) {real, imag} */,
  {32'hbed71f40, 32'h40a76230} /* (17, 6, 5) {real, imag} */,
  {32'h410975f8, 32'h40e55a7e} /* (17, 6, 4) {real, imag} */,
  {32'hc1701db7, 32'hc09f5cb3} /* (17, 6, 3) {real, imag} */,
  {32'h40d750d2, 32'hc00beeda} /* (17, 6, 2) {real, imag} */,
  {32'h419c0ad1, 32'hbfcc1b98} /* (17, 6, 1) {real, imag} */,
  {32'hc148770f, 32'hc0a44bb6} /* (17, 6, 0) {real, imag} */,
  {32'h42bc336d, 32'h41fa391f} /* (17, 5, 31) {real, imag} */,
  {32'hc21b94ba, 32'hc0984324} /* (17, 5, 30) {real, imag} */,
  {32'h40e9ee35, 32'h409f5d45} /* (17, 5, 29) {real, imag} */,
  {32'hc18c3c2e, 32'h41006192} /* (17, 5, 28) {real, imag} */,
  {32'h4103344e, 32'h402aacb8} /* (17, 5, 27) {real, imag} */,
  {32'h3f086558, 32'h41684462} /* (17, 5, 26) {real, imag} */,
  {32'h41075cea, 32'h409e30c0} /* (17, 5, 25) {real, imag} */,
  {32'hc0fa2238, 32'h41039ad4} /* (17, 5, 24) {real, imag} */,
  {32'hbf678388, 32'hc0a7a49a} /* (17, 5, 23) {real, imag} */,
  {32'hc1933d1e, 32'hc177daf8} /* (17, 5, 22) {real, imag} */,
  {32'hc0a357ce, 32'h408fc2e4} /* (17, 5, 21) {real, imag} */,
  {32'h41678729, 32'hc1276fc6} /* (17, 5, 20) {real, imag} */,
  {32'hc05eed69, 32'hbf19238c} /* (17, 5, 19) {real, imag} */,
  {32'h409ccafe, 32'hc03c30ce} /* (17, 5, 18) {real, imag} */,
  {32'h40002650, 32'hc0c6687d} /* (17, 5, 17) {real, imag} */,
  {32'h411e0188, 32'hc0620910} /* (17, 5, 16) {real, imag} */,
  {32'h401578f2, 32'hc0c60530} /* (17, 5, 15) {real, imag} */,
  {32'h40c522ca, 32'h40974341} /* (17, 5, 14) {real, imag} */,
  {32'h41091c18, 32'h4158718e} /* (17, 5, 13) {real, imag} */,
  {32'hbf05c15a, 32'hc16acd4c} /* (17, 5, 12) {real, imag} */,
  {32'hc12de120, 32'h40037aac} /* (17, 5, 11) {real, imag} */,
  {32'h415e8afb, 32'hc0727918} /* (17, 5, 10) {real, imag} */,
  {32'h41945d6e, 32'hc1814249} /* (17, 5, 9) {real, imag} */,
  {32'h4147e471, 32'hc13bc81a} /* (17, 5, 8) {real, imag} */,
  {32'hc1cbb574, 32'h41d393a4} /* (17, 5, 7) {real, imag} */,
  {32'h3f9257b0, 32'hc20a1da8} /* (17, 5, 6) {real, imag} */,
  {32'hc1a65d44, 32'h41b70752} /* (17, 5, 5) {real, imag} */,
  {32'hc0b5fc26, 32'h40e72f2d} /* (17, 5, 4) {real, imag} */,
  {32'hc0252f50, 32'h41550cb8} /* (17, 5, 3) {real, imag} */,
  {32'h4108be06, 32'hc222e1ac} /* (17, 5, 2) {real, imag} */,
  {32'h4231115a, 32'h42a15aad} /* (17, 5, 1) {real, imag} */,
  {32'h41ecaa0f, 32'h42353dfb} /* (17, 5, 0) {real, imag} */,
  {32'hc1c4f2d4, 32'hc2d419ba} /* (17, 4, 31) {real, imag} */,
  {32'h414ae830, 32'h425911df} /* (17, 4, 30) {real, imag} */,
  {32'h41660558, 32'hc1c89c82} /* (17, 4, 29) {real, imag} */,
  {32'hc2715196, 32'hc1d27f96} /* (17, 4, 28) {real, imag} */,
  {32'h419ea620, 32'hbe3b7ad0} /* (17, 4, 27) {real, imag} */,
  {32'hc1757136, 32'h40d7b64c} /* (17, 4, 26) {real, imag} */,
  {32'h4039665a, 32'h410e25e2} /* (17, 4, 25) {real, imag} */,
  {32'h41e7814d, 32'hc1e7e69c} /* (17, 4, 24) {real, imag} */,
  {32'hc157e283, 32'h3f86e4ee} /* (17, 4, 23) {real, imag} */,
  {32'hc07e56e3, 32'h414d006c} /* (17, 4, 22) {real, imag} */,
  {32'hbf92ed97, 32'h4174f120} /* (17, 4, 21) {real, imag} */,
  {32'h40e9525a, 32'hc08ec5d9} /* (17, 4, 20) {real, imag} */,
  {32'h4056db14, 32'hc03a0161} /* (17, 4, 19) {real, imag} */,
  {32'h414ba620, 32'hc0a414c0} /* (17, 4, 18) {real, imag} */,
  {32'hc131be4a, 32'hc126acea} /* (17, 4, 17) {real, imag} */,
  {32'h4141e00c, 32'h41002555} /* (17, 4, 16) {real, imag} */,
  {32'h40a5e585, 32'h40acc103} /* (17, 4, 15) {real, imag} */,
  {32'h40a066c8, 32'h3f1062b8} /* (17, 4, 14) {real, imag} */,
  {32'h3e8c3c60, 32'h4184eb5d} /* (17, 4, 13) {real, imag} */,
  {32'hc0edaac3, 32'hc0518c38} /* (17, 4, 12) {real, imag} */,
  {32'h4121376b, 32'hc12198e2} /* (17, 4, 11) {real, imag} */,
  {32'h41336582, 32'hc05ea772} /* (17, 4, 10) {real, imag} */,
  {32'h40346804, 32'h40d43eeb} /* (17, 4, 9) {real, imag} */,
  {32'h41498354, 32'hc04f3887} /* (17, 4, 8) {real, imag} */,
  {32'hc190ec04, 32'hc1a2e694} /* (17, 4, 7) {real, imag} */,
  {32'hbfd80170, 32'h41e88f71} /* (17, 4, 6) {real, imag} */,
  {32'hc1cd42d7, 32'h41a26184} /* (17, 4, 5) {real, imag} */,
  {32'h41b5a3fe, 32'h40c31bfa} /* (17, 4, 4) {real, imag} */,
  {32'hc1dbbaa7, 32'hc1e96c84} /* (17, 4, 3) {real, imag} */,
  {32'h42a29447, 32'h42a39302} /* (17, 4, 2) {real, imag} */,
  {32'hc2c04ae0, 32'hc21d6da8} /* (17, 4, 1) {real, imag} */,
  {32'hc29cbe58, 32'hc273c19b} /* (17, 4, 0) {real, imag} */,
  {32'h4300dd57, 32'hc2b579f5} /* (17, 3, 31) {real, imag} */,
  {32'hc2389607, 32'h4318522a} /* (17, 3, 30) {real, imag} */,
  {32'h410b0521, 32'hc0f32a60} /* (17, 3, 29) {real, imag} */,
  {32'hc226d3fa, 32'hc1c1aa41} /* (17, 3, 28) {real, imag} */,
  {32'h42207314, 32'hc14b5c9e} /* (17, 3, 27) {real, imag} */,
  {32'hc1edb4db, 32'hc0ff7a40} /* (17, 3, 26) {real, imag} */,
  {32'hc0a2b79c, 32'h419ba0c9} /* (17, 3, 25) {real, imag} */,
  {32'hc049598c, 32'h40ab2d17} /* (17, 3, 24) {real, imag} */,
  {32'hc169063c, 32'hc10bc7a0} /* (17, 3, 23) {real, imag} */,
  {32'hc04bfca9, 32'h4097cc30} /* (17, 3, 22) {real, imag} */,
  {32'hc17be565, 32'h410eb270} /* (17, 3, 21) {real, imag} */,
  {32'hc09537ba, 32'h403317b0} /* (17, 3, 20) {real, imag} */,
  {32'hbfe3a8d2, 32'h411d670a} /* (17, 3, 19) {real, imag} */,
  {32'hc1918005, 32'h41235f08} /* (17, 3, 18) {real, imag} */,
  {32'h41262c02, 32'hc137b195} /* (17, 3, 17) {real, imag} */,
  {32'hc13a2fd4, 32'h410eb359} /* (17, 3, 16) {real, imag} */,
  {32'h3fc00922, 32'hc09ff018} /* (17, 3, 15) {real, imag} */,
  {32'h40568e6d, 32'hbd33d740} /* (17, 3, 14) {real, imag} */,
  {32'h408c8fbc, 32'hbf0b82b0} /* (17, 3, 13) {real, imag} */,
  {32'hc0a5bd73, 32'hc18432b4} /* (17, 3, 12) {real, imag} */,
  {32'h410364bd, 32'hbf3cf810} /* (17, 3, 11) {real, imag} */,
  {32'hc03cd734, 32'h412e8d2a} /* (17, 3, 10) {real, imag} */,
  {32'h40c23098, 32'hc0d80a4e} /* (17, 3, 9) {real, imag} */,
  {32'h40f2efa9, 32'hc11ce4fc} /* (17, 3, 8) {real, imag} */,
  {32'hc10c2bab, 32'h40cfd531} /* (17, 3, 7) {real, imag} */,
  {32'h40f2105a, 32'h4149a48d} /* (17, 3, 6) {real, imag} */,
  {32'hc1a4350a, 32'h41b986f0} /* (17, 3, 5) {real, imag} */,
  {32'h41c1ccfe, 32'h42130496} /* (17, 3, 4) {real, imag} */,
  {32'h41b50749, 32'hc277ab50} /* (17, 3, 3) {real, imag} */,
  {32'h4230f8ea, 32'h42ab433c} /* (17, 3, 2) {real, imag} */,
  {32'hc2654387, 32'hc305d28e} /* (17, 3, 1) {real, imag} */,
  {32'h420341ba, 32'hc0833f42} /* (17, 3, 0) {real, imag} */,
  {32'h4447915e, 32'h4119cbf4} /* (17, 2, 31) {real, imag} */,
  {32'hc3bd1670, 32'h42a34ecf} /* (17, 2, 30) {real, imag} */,
  {32'h428fef67, 32'h40001cd8} /* (17, 2, 29) {real, imag} */,
  {32'h4219df6a, 32'hc28263c2} /* (17, 2, 28) {real, imag} */,
  {32'hc27acdea, 32'h4228e65a} /* (17, 2, 27) {real, imag} */,
  {32'hbe2a4e00, 32'hc10a4aee} /* (17, 2, 26) {real, imag} */,
  {32'h42028a66, 32'hc14e0f40} /* (17, 2, 25) {real, imag} */,
  {32'hc24ba448, 32'h41a86196} /* (17, 2, 24) {real, imag} */,
  {32'hc0c7ef9d, 32'h40de6cc8} /* (17, 2, 23) {real, imag} */,
  {32'hc099dee0, 32'h412b02f3} /* (17, 2, 22) {real, imag} */,
  {32'hc094a283, 32'h415995c9} /* (17, 2, 21) {real, imag} */,
  {32'h3e9d8ac0, 32'hc132476c} /* (17, 2, 20) {real, imag} */,
  {32'h3fedae26, 32'h402ff8d8} /* (17, 2, 19) {real, imag} */,
  {32'h40c93973, 32'h412248c7} /* (17, 2, 18) {real, imag} */,
  {32'h3f17f04c, 32'hc14619fc} /* (17, 2, 17) {real, imag} */,
  {32'h40d2c800, 32'hc05e694c} /* (17, 2, 16) {real, imag} */,
  {32'h40834f7e, 32'h408eedc6} /* (17, 2, 15) {real, imag} */,
  {32'hc145a022, 32'hc113a118} /* (17, 2, 14) {real, imag} */,
  {32'h3fa11f96, 32'hc0035031} /* (17, 2, 13) {real, imag} */,
  {32'h4033c1d0, 32'hc0e82340} /* (17, 2, 12) {real, imag} */,
  {32'hc03d5ae1, 32'hbfde1358} /* (17, 2, 11) {real, imag} */,
  {32'h41299585, 32'h40cb4fe4} /* (17, 2, 10) {real, imag} */,
  {32'hc0f37bc8, 32'h40dd08d7} /* (17, 2, 9) {real, imag} */,
  {32'hc12299bb, 32'hc14456ab} /* (17, 2, 8) {real, imag} */,
  {32'h3febc9e9, 32'hc10136c6} /* (17, 2, 7) {real, imag} */,
  {32'hbe644850, 32'h420a2d36} /* (17, 2, 6) {real, imag} */,
  {32'hc2aa10a1, 32'hc29e6237} /* (17, 2, 5) {real, imag} */,
  {32'h42cdf940, 32'hc22cdad9} /* (17, 2, 4) {real, imag} */,
  {32'h4224a4b4, 32'hc0c3785f} /* (17, 2, 3) {real, imag} */,
  {32'hc38e17b0, 32'h42ccefe8} /* (17, 2, 2) {real, imag} */,
  {32'h43e45dc9, 32'hc30390fb} /* (17, 2, 1) {real, imag} */,
  {32'h43d3456d, 32'h42afd54d} /* (17, 2, 0) {real, imag} */,
  {32'hc46325b8, 32'h43204e43} /* (17, 1, 31) {real, imag} */,
  {32'h438723ca, 32'hc2507471} /* (17, 1, 30) {real, imag} */,
  {32'hbfd78d70, 32'h41a9f710} /* (17, 1, 29) {real, imag} */,
  {32'hc2798756, 32'hc28e2986} /* (17, 1, 28) {real, imag} */,
  {32'h431a21f0, 32'h414962a4} /* (17, 1, 27) {real, imag} */,
  {32'h423476a8, 32'h40fd81b3} /* (17, 1, 26) {real, imag} */,
  {32'hc15ea69c, 32'h4166a351} /* (17, 1, 25) {real, imag} */,
  {32'h419f9115, 32'hc20c2e6e} /* (17, 1, 24) {real, imag} */,
  {32'hbe8ac650, 32'hc126c95f} /* (17, 1, 23) {real, imag} */,
  {32'hc051f9b6, 32'hc11254de} /* (17, 1, 22) {real, imag} */,
  {32'hc03e8df6, 32'hc1926f32} /* (17, 1, 21) {real, imag} */,
  {32'h413b49f7, 32'h413e1108} /* (17, 1, 20) {real, imag} */,
  {32'hc0077376, 32'h4007e550} /* (17, 1, 19) {real, imag} */,
  {32'hbfa02454, 32'h407379a5} /* (17, 1, 18) {real, imag} */,
  {32'h40be2cb7, 32'h4185e109} /* (17, 1, 17) {real, imag} */,
  {32'hc1194d8e, 32'hc129aef1} /* (17, 1, 16) {real, imag} */,
  {32'h4138029a, 32'h3fb1f370} /* (17, 1, 15) {real, imag} */,
  {32'hc182c1b2, 32'hc06b45f4} /* (17, 1, 14) {real, imag} */,
  {32'hc18a5661, 32'hc0aad338} /* (17, 1, 13) {real, imag} */,
  {32'h4166d210, 32'hc14e21ae} /* (17, 1, 12) {real, imag} */,
  {32'h3f7015e0, 32'h41d25396} /* (17, 1, 11) {real, imag} */,
  {32'h40be94db, 32'hbf19d878} /* (17, 1, 10) {real, imag} */,
  {32'hc059dcbc, 32'hc0943fb1} /* (17, 1, 9) {real, imag} */,
  {32'h41a50ad9, 32'h428df75e} /* (17, 1, 8) {real, imag} */,
  {32'hc1082fea, 32'hc12a350a} /* (17, 1, 7) {real, imag} */,
  {32'h412a8dda, 32'hc0108c04} /* (17, 1, 6) {real, imag} */,
  {32'h426f34bc, 32'h4219facb} /* (17, 1, 5) {real, imag} */,
  {32'hc22d22e4, 32'hc1fe4f6d} /* (17, 1, 4) {real, imag} */,
  {32'hc22d1d2b, 32'hc25736df} /* (17, 1, 3) {real, imag} */,
  {32'h43b119ae, 32'h43da851f} /* (17, 1, 2) {real, imag} */,
  {32'hc4aaf334, 32'hc4250cfc} /* (17, 1, 1) {real, imag} */,
  {32'hc48ef3c0, 32'hc37de829} /* (17, 1, 0) {real, imag} */,
  {32'hc4671599, 32'h4422213a} /* (17, 0, 31) {real, imag} */,
  {32'h42a5bd79, 32'hc363558b} /* (17, 0, 30) {real, imag} */,
  {32'h4271d857, 32'h41e52f40} /* (17, 0, 29) {real, imag} */,
  {32'h4113d84e, 32'hc1c8ef74} /* (17, 0, 28) {real, imag} */,
  {32'h41f4c91c, 32'h422b5e56} /* (17, 0, 27) {real, imag} */,
  {32'h3ff93b08, 32'hc0d95845} /* (17, 0, 26) {real, imag} */,
  {32'hc0faba63, 32'h417da962} /* (17, 0, 25) {real, imag} */,
  {32'h41fc9351, 32'hc13bb64e} /* (17, 0, 24) {real, imag} */,
  {32'h40aa1894, 32'hc16e5358} /* (17, 0, 23) {real, imag} */,
  {32'h40c2ac6e, 32'h408ee08e} /* (17, 0, 22) {real, imag} */,
  {32'h418b1072, 32'hc1b0c811} /* (17, 0, 21) {real, imag} */,
  {32'h401fcefa, 32'h409b7fb2} /* (17, 0, 20) {real, imag} */,
  {32'h4117bee2, 32'h41295176} /* (17, 0, 19) {real, imag} */,
  {32'hc128fa80, 32'hc0ec2939} /* (17, 0, 18) {real, imag} */,
  {32'hc033dc7f, 32'h4104f2a3} /* (17, 0, 17) {real, imag} */,
  {32'hc14448a2, 32'h00000000} /* (17, 0, 16) {real, imag} */,
  {32'hc033dc7f, 32'hc104f2a3} /* (17, 0, 15) {real, imag} */,
  {32'hc128fa80, 32'h40ec2939} /* (17, 0, 14) {real, imag} */,
  {32'h4117bee2, 32'hc1295176} /* (17, 0, 13) {real, imag} */,
  {32'h401fcefa, 32'hc09b7fb2} /* (17, 0, 12) {real, imag} */,
  {32'h418b1072, 32'h41b0c811} /* (17, 0, 11) {real, imag} */,
  {32'h40c2ac6e, 32'hc08ee08e} /* (17, 0, 10) {real, imag} */,
  {32'h40aa1894, 32'h416e5358} /* (17, 0, 9) {real, imag} */,
  {32'h41fc9351, 32'h413bb64e} /* (17, 0, 8) {real, imag} */,
  {32'hc0faba63, 32'hc17da962} /* (17, 0, 7) {real, imag} */,
  {32'h3ff93b08, 32'h40d95845} /* (17, 0, 6) {real, imag} */,
  {32'h41f4c91c, 32'hc22b5e56} /* (17, 0, 5) {real, imag} */,
  {32'h4113d84e, 32'h41c8ef74} /* (17, 0, 4) {real, imag} */,
  {32'h4271d857, 32'hc1e52f40} /* (17, 0, 3) {real, imag} */,
  {32'h42a5bd79, 32'h4363558b} /* (17, 0, 2) {real, imag} */,
  {32'hc4671599, 32'hc422213a} /* (17, 0, 1) {real, imag} */,
  {32'hc48c0ae0, 32'h00000000} /* (17, 0, 0) {real, imag} */,
  {32'hc416a040, 32'h4370ba5d} /* (16, 31, 31) {real, imag} */,
  {32'h43003086, 32'hc3542f73} /* (16, 31, 30) {real, imag} */,
  {32'hc1fee1ff, 32'hc13a5880} /* (16, 31, 29) {real, imag} */,
  {32'hc23a5c66, 32'h41249777} /* (16, 31, 28) {real, imag} */,
  {32'h427660e2, 32'hc1f518ce} /* (16, 31, 27) {real, imag} */,
  {32'hc090c21a, 32'hc19679ee} /* (16, 31, 26) {real, imag} */,
  {32'hc00f8e26, 32'h41a0ac28} /* (16, 31, 25) {real, imag} */,
  {32'h40fe7128, 32'hc1bd5189} /* (16, 31, 24) {real, imag} */,
  {32'h41128433, 32'hc0ffd64c} /* (16, 31, 23) {real, imag} */,
  {32'h40878c98, 32'hc061d634} /* (16, 31, 22) {real, imag} */,
  {32'h40754fc6, 32'hc1cf6f50} /* (16, 31, 21) {real, imag} */,
  {32'hc10bd5c4, 32'h41aa38c2} /* (16, 31, 20) {real, imag} */,
  {32'h3eba93a8, 32'hc057d8c8} /* (16, 31, 19) {real, imag} */,
  {32'hbf2c29cc, 32'hc0e4d42a} /* (16, 31, 18) {real, imag} */,
  {32'hbf38b92c, 32'hc0952676} /* (16, 31, 17) {real, imag} */,
  {32'hc0c43076, 32'hc13151b0} /* (16, 31, 16) {real, imag} */,
  {32'hc13d88f8, 32'h40659aef} /* (16, 31, 15) {real, imag} */,
  {32'h400488e8, 32'hc0c4c194} /* (16, 31, 14) {real, imag} */,
  {32'h3e571d80, 32'hc150cc18} /* (16, 31, 13) {real, imag} */,
  {32'h40c597a8, 32'h41496438} /* (16, 31, 12) {real, imag} */,
  {32'hbf805608, 32'h41b04976} /* (16, 31, 11) {real, imag} */,
  {32'hc095f084, 32'hc0d65155} /* (16, 31, 10) {real, imag} */,
  {32'hc147fb94, 32'hc161bd66} /* (16, 31, 9) {real, imag} */,
  {32'hbe9a22b0, 32'h414ca71f} /* (16, 31, 8) {real, imag} */,
  {32'hc122288c, 32'hc1317902} /* (16, 31, 7) {real, imag} */,
  {32'h421fb484, 32'h3f3e6d20} /* (16, 31, 6) {real, imag} */,
  {32'h42ac0bc7, 32'h406f9e22} /* (16, 31, 5) {real, imag} */,
  {32'hc1e7daa7, 32'h427fb5b5} /* (16, 31, 4) {real, imag} */,
  {32'hc0a62fb2, 32'hc2161134} /* (16, 31, 3) {real, imag} */,
  {32'h42ceb9cb, 32'h422d3df8} /* (16, 31, 2) {real, imag} */,
  {32'hc3a9e471, 32'hc1f7d62e} /* (16, 31, 1) {real, imag} */,
  {32'hc3dbf39e, 32'h4356e162} /* (16, 31, 0) {real, imag} */,
  {32'h43525d58, 32'h42874e32} /* (16, 30, 31) {real, imag} */,
  {32'hc3135ae8, 32'hc2557096} /* (16, 30, 30) {real, imag} */,
  {32'h424e23a5, 32'h4208953e} /* (16, 30, 29) {real, imag} */,
  {32'h428cd20f, 32'h427ba005} /* (16, 30, 28) {real, imag} */,
  {32'hc227d671, 32'h4205cc47} /* (16, 30, 27) {real, imag} */,
  {32'h41460f24, 32'hc2086788} /* (16, 30, 26) {real, imag} */,
  {32'h41015ed4, 32'h41a8dbae} /* (16, 30, 25) {real, imag} */,
  {32'hbf889ec0, 32'h419e9816} /* (16, 30, 24) {real, imag} */,
  {32'hc1375fee, 32'hc1413fc8} /* (16, 30, 23) {real, imag} */,
  {32'hc0e9d6d9, 32'hc11f7780} /* (16, 30, 22) {real, imag} */,
  {32'h3f6ce7e8, 32'h4133794e} /* (16, 30, 21) {real, imag} */,
  {32'hc1b2f796, 32'hc10b6330} /* (16, 30, 20) {real, imag} */,
  {32'h40883189, 32'hc1295024} /* (16, 30, 19) {real, imag} */,
  {32'hc100a7b6, 32'h41363e1f} /* (16, 30, 18) {real, imag} */,
  {32'hc142b1cf, 32'hc02eceec} /* (16, 30, 17) {real, imag} */,
  {32'hc032db5d, 32'hc0aae302} /* (16, 30, 16) {real, imag} */,
  {32'hc1054dc6, 32'h404b1777} /* (16, 30, 15) {real, imag} */,
  {32'hc029ca0b, 32'h3ec3d998} /* (16, 30, 14) {real, imag} */,
  {32'hc134a8cc, 32'h3f36c77e} /* (16, 30, 13) {real, imag} */,
  {32'h40b6fcaa, 32'h4087d80a} /* (16, 30, 12) {real, imag} */,
  {32'h3e024e20, 32'hc1c0d919} /* (16, 30, 11) {real, imag} */,
  {32'hc04edfa3, 32'h40ca6495} /* (16, 30, 10) {real, imag} */,
  {32'hc14c89d3, 32'hc18cc3a5} /* (16, 30, 9) {real, imag} */,
  {32'hc2085792, 32'hc1566ed8} /* (16, 30, 8) {real, imag} */,
  {32'h41d35b7e, 32'h42144c77} /* (16, 30, 7) {real, imag} */,
  {32'h408f1896, 32'hc164c2ed} /* (16, 30, 6) {real, imag} */,
  {32'hc1fd5c0e, 32'hc196de1c} /* (16, 30, 5) {real, imag} */,
  {32'h41c53ad6, 32'h41b337ce} /* (16, 30, 4) {real, imag} */,
  {32'h4290f9ee, 32'hc1a6bee2} /* (16, 30, 3) {real, imag} */,
  {32'hc32b9d67, 32'hc216c7cd} /* (16, 30, 2) {real, imag} */,
  {32'h43b5b55c, 32'h42082d55} /* (16, 30, 1) {real, imag} */,
  {32'h432463d3, 32'hc289471a} /* (16, 30, 0) {real, imag} */,
  {32'hc2026ac2, 32'h42a3f852} /* (16, 29, 31) {real, imag} */,
  {32'h42971188, 32'hc216f3d0} /* (16, 29, 30) {real, imag} */,
  {32'h410cfc1b, 32'h417dfa0d} /* (16, 29, 29) {real, imag} */,
  {32'h4190803e, 32'hc19d0864} /* (16, 29, 28) {real, imag} */,
  {32'hc18e1e02, 32'hc1002733} /* (16, 29, 27) {real, imag} */,
  {32'hc18005d0, 32'hc08311c2} /* (16, 29, 26) {real, imag} */,
  {32'hc0d0444c, 32'h411b23b6} /* (16, 29, 25) {real, imag} */,
  {32'h4002eb04, 32'h418226a3} /* (16, 29, 24) {real, imag} */,
  {32'hc18f8df1, 32'hc0e87389} /* (16, 29, 23) {real, imag} */,
  {32'h3eeacb50, 32'h4188e3c5} /* (16, 29, 22) {real, imag} */,
  {32'h4167c226, 32'h409fbefd} /* (16, 29, 21) {real, imag} */,
  {32'hc1316220, 32'h40fecc8b} /* (16, 29, 20) {real, imag} */,
  {32'hc14d823d, 32'h40ba483a} /* (16, 29, 19) {real, imag} */,
  {32'h414d49bd, 32'h3ffc036a} /* (16, 29, 18) {real, imag} */,
  {32'h4148a698, 32'hc12f8729} /* (16, 29, 17) {real, imag} */,
  {32'h4094aec2, 32'hc0d777d5} /* (16, 29, 16) {real, imag} */,
  {32'hc09ac3ce, 32'h403295e6} /* (16, 29, 15) {real, imag} */,
  {32'hbf35b548, 32'h40b23e14} /* (16, 29, 14) {real, imag} */,
  {32'hbfff8368, 32'h4101c5aa} /* (16, 29, 13) {real, imag} */,
  {32'hbea18910, 32'hc06ab9b7} /* (16, 29, 12) {real, imag} */,
  {32'h41502bdd, 32'hbf9431be} /* (16, 29, 11) {real, imag} */,
  {32'h3e96ec70, 32'h40c0ba5d} /* (16, 29, 10) {real, imag} */,
  {32'hc1512ec5, 32'hc0178b56} /* (16, 29, 9) {real, imag} */,
  {32'hc0dcea7a, 32'h3ff58794} /* (16, 29, 8) {real, imag} */,
  {32'hc1baa252, 32'hc1abb9e5} /* (16, 29, 7) {real, imag} */,
  {32'hc0188f58, 32'hbfa196b6} /* (16, 29, 6) {real, imag} */,
  {32'h416191b8, 32'hc0668ad4} /* (16, 29, 5) {real, imag} */,
  {32'hc146e227, 32'hbfbf4d74} /* (16, 29, 4) {real, imag} */,
  {32'hc1c8b58a, 32'hc1979098} /* (16, 29, 3) {real, imag} */,
  {32'h41ab2c82, 32'hc2a46962} /* (16, 29, 2) {real, imag} */,
  {32'h42d5e0dc, 32'h4250b5ec} /* (16, 29, 1) {real, imag} */,
  {32'h41905f7a, 32'hc1a4b14b} /* (16, 29, 0) {real, imag} */,
  {32'hc20ce2be, 32'h4215a388} /* (16, 28, 31) {real, imag} */,
  {32'h42176092, 32'hc278c2f9} /* (16, 28, 30) {real, imag} */,
  {32'hc17d33a6, 32'h408b24d8} /* (16, 28, 29) {real, imag} */,
  {32'hc103fc49, 32'h41d7fa27} /* (16, 28, 28) {real, imag} */,
  {32'hc18aae12, 32'hc10239a2} /* (16, 28, 27) {real, imag} */,
  {32'hc123d011, 32'h4124bb9c} /* (16, 28, 26) {real, imag} */,
  {32'hc1db095a, 32'h40960a48} /* (16, 28, 25) {real, imag} */,
  {32'h4191f692, 32'hc12d68be} /* (16, 28, 24) {real, imag} */,
  {32'hc11930da, 32'hc181ad64} /* (16, 28, 23) {real, imag} */,
  {32'h41a38449, 32'hc0094c7c} /* (16, 28, 22) {real, imag} */,
  {32'hc0cb16fe, 32'h411ec8b7} /* (16, 28, 21) {real, imag} */,
  {32'h40707691, 32'hc00a6a56} /* (16, 28, 20) {real, imag} */,
  {32'hc14b4da3, 32'hc105ef57} /* (16, 28, 19) {real, imag} */,
  {32'hc0a41c75, 32'hc0ce2ff2} /* (16, 28, 18) {real, imag} */,
  {32'h41146a74, 32'h404a939e} /* (16, 28, 17) {real, imag} */,
  {32'hc09e3c68, 32'h409ae6a6} /* (16, 28, 16) {real, imag} */,
  {32'hc10576e6, 32'hbf8c59a6} /* (16, 28, 15) {real, imag} */,
  {32'h4092e2e9, 32'hc027d58e} /* (16, 28, 14) {real, imag} */,
  {32'h3fa4c4b0, 32'hc064b6d6} /* (16, 28, 13) {real, imag} */,
  {32'hc0053f98, 32'hc0cc0c12} /* (16, 28, 12) {real, imag} */,
  {32'hbf64ad36, 32'h40baa582} /* (16, 28, 11) {real, imag} */,
  {32'h4061fc82, 32'hc085ff20} /* (16, 28, 10) {real, imag} */,
  {32'h402cfae6, 32'hbf69bf10} /* (16, 28, 9) {real, imag} */,
  {32'h42099a8e, 32'h41b8d4ff} /* (16, 28, 8) {real, imag} */,
  {32'hc19cb690, 32'hbd317400} /* (16, 28, 7) {real, imag} */,
  {32'hc1259ff8, 32'hc08d4d5f} /* (16, 28, 6) {real, imag} */,
  {32'h4194e39b, 32'hc0a89d65} /* (16, 28, 5) {real, imag} */,
  {32'hc21c27aa, 32'hc0fc8e5e} /* (16, 28, 4) {real, imag} */,
  {32'hc020bf02, 32'h421ae6e1} /* (16, 28, 3) {real, imag} */,
  {32'h420f346b, 32'hc1c7f420} /* (16, 28, 2) {real, imag} */,
  {32'hc0fef748, 32'h428e53ee} /* (16, 28, 1) {real, imag} */,
  {32'hc28acaa1, 32'h4296486a} /* (16, 28, 0) {real, imag} */,
  {32'h41a0dc8e, 32'hc25c1706} /* (16, 27, 31) {real, imag} */,
  {32'hc046f4b8, 32'h42366d87} /* (16, 27, 30) {real, imag} */,
  {32'hc12489dd, 32'h3fb24d8c} /* (16, 27, 29) {real, imag} */,
  {32'h4154b8f5, 32'hbf632e98} /* (16, 27, 28) {real, imag} */,
  {32'hc1e00008, 32'hc1dcbb5b} /* (16, 27, 27) {real, imag} */,
  {32'hc04f8582, 32'hc0cf2bf4} /* (16, 27, 26) {real, imag} */,
  {32'hbf9854b8, 32'hc186caac} /* (16, 27, 25) {real, imag} */,
  {32'h40ce175e, 32'hc11a4fe6} /* (16, 27, 24) {real, imag} */,
  {32'hc178c88c, 32'hc01e1b2a} /* (16, 27, 23) {real, imag} */,
  {32'hc1041c64, 32'h41c378ea} /* (16, 27, 22) {real, imag} */,
  {32'h418f13c0, 32'hc1018f4d} /* (16, 27, 21) {real, imag} */,
  {32'h416e77ad, 32'hc118a145} /* (16, 27, 20) {real, imag} */,
  {32'hc0051cda, 32'h406a0f04} /* (16, 27, 19) {real, imag} */,
  {32'h41093b1a, 32'h406ac28b} /* (16, 27, 18) {real, imag} */,
  {32'hc11c228f, 32'hc12bbf3b} /* (16, 27, 17) {real, imag} */,
  {32'hc12e3380, 32'hc10d46b1} /* (16, 27, 16) {real, imag} */,
  {32'h3fc84a76, 32'hbf80c8e1} /* (16, 27, 15) {real, imag} */,
  {32'h402f3984, 32'h3fab52b8} /* (16, 27, 14) {real, imag} */,
  {32'h3e7db080, 32'h4130760e} /* (16, 27, 13) {real, imag} */,
  {32'hc12b2d92, 32'hbf8b64e0} /* (16, 27, 12) {real, imag} */,
  {32'hc08bab9e, 32'h40d14531} /* (16, 27, 11) {real, imag} */,
  {32'h3f1b9680, 32'hc13b0653} /* (16, 27, 10) {real, imag} */,
  {32'hc103a542, 32'hbfd8a9e8} /* (16, 27, 9) {real, imag} */,
  {32'hc1b94790, 32'hc1429a9f} /* (16, 27, 8) {real, imag} */,
  {32'hc0d4e649, 32'h40c34098} /* (16, 27, 7) {real, imag} */,
  {32'hc06144db, 32'hc185ebf2} /* (16, 27, 6) {real, imag} */,
  {32'h405db322, 32'hc1a6a638} /* (16, 27, 5) {real, imag} */,
  {32'h401dce72, 32'hc15b7df2} /* (16, 27, 4) {real, imag} */,
  {32'h41318f0c, 32'hc1d2cc37} /* (16, 27, 3) {real, imag} */,
  {32'hc1dde820, 32'h41dae196} /* (16, 27, 2) {real, imag} */,
  {32'h425146f0, 32'hc1eab79a} /* (16, 27, 1) {real, imag} */,
  {32'h413619bc, 32'hc224ad66} /* (16, 27, 0) {real, imag} */,
  {32'h419c7b22, 32'hc03cc0b0} /* (16, 26, 31) {real, imag} */,
  {32'h4149149e, 32'h407bba58} /* (16, 26, 30) {real, imag} */,
  {32'h40960241, 32'hc0ee1746} /* (16, 26, 29) {real, imag} */,
  {32'h3fa327c0, 32'hc1b0f047} /* (16, 26, 28) {real, imag} */,
  {32'hc0350853, 32'h409c36f4} /* (16, 26, 27) {real, imag} */,
  {32'h4078c06a, 32'hbe09c6b0} /* (16, 26, 26) {real, imag} */,
  {32'h41af4862, 32'hbfe719f8} /* (16, 26, 25) {real, imag} */,
  {32'hc011c108, 32'h41803afc} /* (16, 26, 24) {real, imag} */,
  {32'h3e2c44e0, 32'h3fad4c3c} /* (16, 26, 23) {real, imag} */,
  {32'hc1a48c5d, 32'hc02dc1ac} /* (16, 26, 22) {real, imag} */,
  {32'hc15df51b, 32'hc118e706} /* (16, 26, 21) {real, imag} */,
  {32'h4143dae3, 32'h3eb15270} /* (16, 26, 20) {real, imag} */,
  {32'h413acf5e, 32'h41843cfb} /* (16, 26, 19) {real, imag} */,
  {32'h414f250a, 32'hc0ae7ffe} /* (16, 26, 18) {real, imag} */,
  {32'h40abb11d, 32'hc101672d} /* (16, 26, 17) {real, imag} */,
  {32'hc00b14c0, 32'h3ff03d4a} /* (16, 26, 16) {real, imag} */,
  {32'h40c7ac93, 32'hbf1e9f4a} /* (16, 26, 15) {real, imag} */,
  {32'hc0205ba6, 32'h41901716} /* (16, 26, 14) {real, imag} */,
  {32'h40f8964e, 32'hbfa533bf} /* (16, 26, 13) {real, imag} */,
  {32'hbfb5a018, 32'h41b85db2} /* (16, 26, 12) {real, imag} */,
  {32'hbeaf36b0, 32'hc08860fc} /* (16, 26, 11) {real, imag} */,
  {32'h40dc52dc, 32'h3ff3cbfc} /* (16, 26, 10) {real, imag} */,
  {32'hc0eb0490, 32'hbfb19bc0} /* (16, 26, 9) {real, imag} */,
  {32'h401fc3c1, 32'h416846a6} /* (16, 26, 8) {real, imag} */,
  {32'h405e029e, 32'hc18cbda7} /* (16, 26, 7) {real, imag} */,
  {32'hc01ebc74, 32'h40512764} /* (16, 26, 6) {real, imag} */,
  {32'hbc417c00, 32'hc06afc42} /* (16, 26, 5) {real, imag} */,
  {32'hc1039244, 32'hc13650b5} /* (16, 26, 4) {real, imag} */,
  {32'h3f6cebe4, 32'h41c6318b} /* (16, 26, 3) {real, imag} */,
  {32'hc1e34a9f, 32'hc0531000} /* (16, 26, 2) {real, imag} */,
  {32'h416a83e1, 32'hc00e69cc} /* (16, 26, 1) {real, imag} */,
  {32'hc164373a, 32'h41c7785a} /* (16, 26, 0) {real, imag} */,
  {32'hc20e2258, 32'hc1412336} /* (16, 25, 31) {real, imag} */,
  {32'h4115fb1a, 32'h41641866} /* (16, 25, 30) {real, imag} */,
  {32'hc025b60c, 32'h40697c23} /* (16, 25, 29) {real, imag} */,
  {32'h419a940c, 32'hc0be27ed} /* (16, 25, 28) {real, imag} */,
  {32'h40c54229, 32'hc107814e} /* (16, 25, 27) {real, imag} */,
  {32'hc0f4ca63, 32'h40f88243} /* (16, 25, 26) {real, imag} */,
  {32'h4038b28d, 32'h3fcc36d8} /* (16, 25, 25) {real, imag} */,
  {32'hc1481bec, 32'h3f9ca6bc} /* (16, 25, 24) {real, imag} */,
  {32'hc0b48c16, 32'h411f5a90} /* (16, 25, 23) {real, imag} */,
  {32'h3fe64f44, 32'hc146108e} /* (16, 25, 22) {real, imag} */,
  {32'h411cb243, 32'h416dec23} /* (16, 25, 21) {real, imag} */,
  {32'hc0e7da49, 32'h3f6be698} /* (16, 25, 20) {real, imag} */,
  {32'hc1167886, 32'h41572bce} /* (16, 25, 19) {real, imag} */,
  {32'h410f3f86, 32'hbfdf0ce2} /* (16, 25, 18) {real, imag} */,
  {32'hc177365a, 32'hc0f63554} /* (16, 25, 17) {real, imag} */,
  {32'h40e91d02, 32'h40a83555} /* (16, 25, 16) {real, imag} */,
  {32'hc0ea4d8c, 32'h40091450} /* (16, 25, 15) {real, imag} */,
  {32'hc0bcd34b, 32'h40dc146b} /* (16, 25, 14) {real, imag} */,
  {32'h408fc175, 32'h41bd2980} /* (16, 25, 13) {real, imag} */,
  {32'hc1ad22ab, 32'hc08904e0} /* (16, 25, 12) {real, imag} */,
  {32'h410dc0ac, 32'hc0b6abdc} /* (16, 25, 11) {real, imag} */,
  {32'h40cc6de2, 32'h40f47b89} /* (16, 25, 10) {real, imag} */,
  {32'h4173b8a2, 32'hc0ed1bb8} /* (16, 25, 9) {real, imag} */,
  {32'hc001e20f, 32'hbdacad80} /* (16, 25, 8) {real, imag} */,
  {32'hc0dda323, 32'h403ba25a} /* (16, 25, 7) {real, imag} */,
  {32'h409d4e34, 32'h408a75e8} /* (16, 25, 6) {real, imag} */,
  {32'hc02c55ef, 32'h3f42a76c} /* (16, 25, 5) {real, imag} */,
  {32'hc17ebc5e, 32'hc0e17932} /* (16, 25, 4) {real, imag} */,
  {32'hc1bd531a, 32'h3ef08240} /* (16, 25, 3) {real, imag} */,
  {32'h415938be, 32'h41bf75e4} /* (16, 25, 2) {real, imag} */,
  {32'h3ff3a648, 32'hc203c1b0} /* (16, 25, 1) {real, imag} */,
  {32'hc02b7490, 32'h41321a3c} /* (16, 25, 0) {real, imag} */,
  {32'h41bafc54, 32'hc1f19911} /* (16, 24, 31) {real, imag} */,
  {32'hc0e2054c, 32'hbfe75f36} /* (16, 24, 30) {real, imag} */,
  {32'hc1100690, 32'hc12a6a21} /* (16, 24, 29) {real, imag} */,
  {32'h3fc75044, 32'h41a0916d} /* (16, 24, 28) {real, imag} */,
  {32'h413de063, 32'h417b5a17} /* (16, 24, 27) {real, imag} */,
  {32'h416302e4, 32'h419518b9} /* (16, 24, 26) {real, imag} */,
  {32'hc1199166, 32'hc1881508} /* (16, 24, 25) {real, imag} */,
  {32'hc01cbd02, 32'h4170eb11} /* (16, 24, 24) {real, imag} */,
  {32'h4131c973, 32'hc021db98} /* (16, 24, 23) {real, imag} */,
  {32'hc1403fbe, 32'hc0c652de} /* (16, 24, 22) {real, imag} */,
  {32'hc15ff4e4, 32'hc13cdc1a} /* (16, 24, 21) {real, imag} */,
  {32'h4146f27e, 32'hc0093d4e} /* (16, 24, 20) {real, imag} */,
  {32'hc0abf8c2, 32'hbf4aca60} /* (16, 24, 19) {real, imag} */,
  {32'hc089583c, 32'hc119f0ed} /* (16, 24, 18) {real, imag} */,
  {32'h41636aee, 32'hc0b147ac} /* (16, 24, 17) {real, imag} */,
  {32'hbff5c088, 32'hc0e756d5} /* (16, 24, 16) {real, imag} */,
  {32'h40251ffb, 32'h3f416e2a} /* (16, 24, 15) {real, imag} */,
  {32'h40c9b438, 32'hc124083c} /* (16, 24, 14) {real, imag} */,
  {32'hc18f07fa, 32'h416f5374} /* (16, 24, 13) {real, imag} */,
  {32'hc06dd372, 32'hc07afdcc} /* (16, 24, 12) {real, imag} */,
  {32'h3e031f10, 32'hc10b4763} /* (16, 24, 11) {real, imag} */,
  {32'hc134f0c2, 32'h418589df} /* (16, 24, 10) {real, imag} */,
  {32'h41952c9a, 32'h4084102d} /* (16, 24, 9) {real, imag} */,
  {32'hc1bb4e97, 32'h3fe17ca0} /* (16, 24, 8) {real, imag} */,
  {32'h3e15fc60, 32'h4116bd29} /* (16, 24, 7) {real, imag} */,
  {32'hc208a4fb, 32'hc18385de} /* (16, 24, 6) {real, imag} */,
  {32'hc117b41f, 32'hbf2d34ac} /* (16, 24, 5) {real, imag} */,
  {32'h40df0298, 32'h4181a8fe} /* (16, 24, 4) {real, imag} */,
  {32'hc1685e3a, 32'h3ee9b080} /* (16, 24, 3) {real, imag} */,
  {32'hc1be68b2, 32'h416fd801} /* (16, 24, 2) {real, imag} */,
  {32'h40f92d32, 32'hc20e7938} /* (16, 24, 1) {real, imag} */,
  {32'h4174daed, 32'hc116a838} /* (16, 24, 0) {real, imag} */,
  {32'hc10f69c9, 32'h40e1725c} /* (16, 23, 31) {real, imag} */,
  {32'hc1595fe8, 32'hc1d94b4e} /* (16, 23, 30) {real, imag} */,
  {32'h401851d6, 32'h3e1e1d80} /* (16, 23, 29) {real, imag} */,
  {32'hc1293bb8, 32'hc12c3dab} /* (16, 23, 28) {real, imag} */,
  {32'h3fc9154b, 32'h3e894d40} /* (16, 23, 27) {real, imag} */,
  {32'h418ab3b2, 32'h41b89c90} /* (16, 23, 26) {real, imag} */,
  {32'h419af1cb, 32'hc0c793c6} /* (16, 23, 25) {real, imag} */,
  {32'hc13e5da1, 32'hc0a3af6b} /* (16, 23, 24) {real, imag} */,
  {32'h41343dc9, 32'hc14405ae} /* (16, 23, 23) {real, imag} */,
  {32'hc1a1ca96, 32'h41199872} /* (16, 23, 22) {real, imag} */,
  {32'h410ed7ec, 32'hc119cf89} /* (16, 23, 21) {real, imag} */,
  {32'h40ba1339, 32'hc0b4a265} /* (16, 23, 20) {real, imag} */,
  {32'hc0a33aa7, 32'hbf62496c} /* (16, 23, 19) {real, imag} */,
  {32'h40f95a54, 32'h3f759184} /* (16, 23, 18) {real, imag} */,
  {32'h40e01d24, 32'hc10dc252} /* (16, 23, 17) {real, imag} */,
  {32'hbf2eb338, 32'hc1113a07} /* (16, 23, 16) {real, imag} */,
  {32'h4112a36e, 32'hc1072ae6} /* (16, 23, 15) {real, imag} */,
  {32'h40fc7b59, 32'hc1381228} /* (16, 23, 14) {real, imag} */,
  {32'hbff7874a, 32'h40a0cb22} /* (16, 23, 13) {real, imag} */,
  {32'h40e9cf4b, 32'hc144b732} /* (16, 23, 12) {real, imag} */,
  {32'hc10d8e04, 32'h41173746} /* (16, 23, 11) {real, imag} */,
  {32'hc108ef1f, 32'hc15b6b3a} /* (16, 23, 10) {real, imag} */,
  {32'hc1381999, 32'hc16d484c} /* (16, 23, 9) {real, imag} */,
  {32'h3efe5800, 32'hc077aa8b} /* (16, 23, 8) {real, imag} */,
  {32'h3ffb3ede, 32'h4156a950} /* (16, 23, 7) {real, imag} */,
  {32'h41b22a8b, 32'hc107132c} /* (16, 23, 6) {real, imag} */,
  {32'h411325f2, 32'h40a3b785} /* (16, 23, 5) {real, imag} */,
  {32'hc10fdbb2, 32'hc03330c0} /* (16, 23, 4) {real, imag} */,
  {32'h4107e81b, 32'h4104da68} /* (16, 23, 3) {real, imag} */,
  {32'hc13af3aa, 32'hc0866a1b} /* (16, 23, 2) {real, imag} */,
  {32'hc0eced88, 32'hc1791898} /* (16, 23, 1) {real, imag} */,
  {32'h4101cf3d, 32'h4180fb34} /* (16, 23, 0) {real, imag} */,
  {32'h3f01f0b0, 32'h411a3298} /* (16, 22, 31) {real, imag} */,
  {32'h4121afc8, 32'h4082d55a} /* (16, 22, 30) {real, imag} */,
  {32'hc0b65c0e, 32'h40f121a2} /* (16, 22, 29) {real, imag} */,
  {32'h411b498c, 32'h41ca9b39} /* (16, 22, 28) {real, imag} */,
  {32'h40ef9d00, 32'hc0467517} /* (16, 22, 27) {real, imag} */,
  {32'h40461b26, 32'hc14c05a0} /* (16, 22, 26) {real, imag} */,
  {32'h404f9478, 32'h405f3462} /* (16, 22, 25) {real, imag} */,
  {32'hc11d4e97, 32'hc1323c9e} /* (16, 22, 24) {real, imag} */,
  {32'h40a40f4c, 32'hc030f870} /* (16, 22, 23) {real, imag} */,
  {32'h41925ae8, 32'hc090f0c3} /* (16, 22, 22) {real, imag} */,
  {32'h41194178, 32'hbdcb8a30} /* (16, 22, 21) {real, imag} */,
  {32'hc17410a0, 32'hc0bc72d6} /* (16, 22, 20) {real, imag} */,
  {32'h406387d8, 32'h416f5fb5} /* (16, 22, 19) {real, imag} */,
  {32'hc181e9fd, 32'hc15701d3} /* (16, 22, 18) {real, imag} */,
  {32'h40ce2324, 32'h40b528d7} /* (16, 22, 17) {real, imag} */,
  {32'hc135ff1a, 32'hc129d092} /* (16, 22, 16) {real, imag} */,
  {32'h3fd9e73a, 32'hc1bbc68c} /* (16, 22, 15) {real, imag} */,
  {32'h401cbb54, 32'hc04d690d} /* (16, 22, 14) {real, imag} */,
  {32'h41b5f964, 32'hc1213ff7} /* (16, 22, 13) {real, imag} */,
  {32'h416c0107, 32'h4182ad62} /* (16, 22, 12) {real, imag} */,
  {32'hc03e9554, 32'h41d67618} /* (16, 22, 11) {real, imag} */,
  {32'hc0c8a849, 32'hc13e0c27} /* (16, 22, 10) {real, imag} */,
  {32'h4150d99f, 32'h41044364} /* (16, 22, 9) {real, imag} */,
  {32'hc0ce1d87, 32'hc08491ee} /* (16, 22, 8) {real, imag} */,
  {32'hc17dbe89, 32'hc09fb19a} /* (16, 22, 7) {real, imag} */,
  {32'hc10ffbaa, 32'hc1805166} /* (16, 22, 6) {real, imag} */,
  {32'hc190de90, 32'hc09d5560} /* (16, 22, 5) {real, imag} */,
  {32'hc1861950, 32'h3fca81b8} /* (16, 22, 4) {real, imag} */,
  {32'hc111d38c, 32'hc068439f} /* (16, 22, 3) {real, imag} */,
  {32'h4183e306, 32'hc18dbfdc} /* (16, 22, 2) {real, imag} */,
  {32'h3f192688, 32'h4113b20e} /* (16, 22, 1) {real, imag} */,
  {32'hc08ae0e6, 32'h3ea43d30} /* (16, 22, 0) {real, imag} */,
  {32'h40f42859, 32'hc0fae46d} /* (16, 21, 31) {real, imag} */,
  {32'h4105a62b, 32'h412579a7} /* (16, 21, 30) {real, imag} */,
  {32'hc0d7c77b, 32'h41190f94} /* (16, 21, 29) {real, imag} */,
  {32'hc1475cd6, 32'h40720474} /* (16, 21, 28) {real, imag} */,
  {32'h3f61d300, 32'h4113e7ba} /* (16, 21, 27) {real, imag} */,
  {32'hc083fc47, 32'hc07c1e84} /* (16, 21, 26) {real, imag} */,
  {32'hc1ee11e8, 32'h3fcc8fc3} /* (16, 21, 25) {real, imag} */,
  {32'h4188b7f1, 32'hc1aeef45} /* (16, 21, 24) {real, imag} */,
  {32'hbfc309dc, 32'hc154321c} /* (16, 21, 23) {real, imag} */,
  {32'hc089cb2e, 32'h40099941} /* (16, 21, 22) {real, imag} */,
  {32'h4150d457, 32'h40fb1054} /* (16, 21, 21) {real, imag} */,
  {32'hc10a1ba6, 32'h40c2a748} /* (16, 21, 20) {real, imag} */,
  {32'hc1513d12, 32'hc16d0ef4} /* (16, 21, 19) {real, imag} */,
  {32'hc149ad96, 32'h3f89afc4} /* (16, 21, 18) {real, imag} */,
  {32'h4147d4fa, 32'hbb848200} /* (16, 21, 17) {real, imag} */,
  {32'hbdb92540, 32'hc1637ff1} /* (16, 21, 16) {real, imag} */,
  {32'hc0b7c2ca, 32'h409bbdef} /* (16, 21, 15) {real, imag} */,
  {32'h412eeffc, 32'hbff08ddc} /* (16, 21, 14) {real, imag} */,
  {32'hc0cb0ea8, 32'hbf64ab00} /* (16, 21, 13) {real, imag} */,
  {32'hc18e24ad, 32'hc1c82e02} /* (16, 21, 12) {real, imag} */,
  {32'hbf910e58, 32'h407a6f0c} /* (16, 21, 11) {real, imag} */,
  {32'h413a6004, 32'hc049f90c} /* (16, 21, 10) {real, imag} */,
  {32'h41ad8660, 32'h407c98f8} /* (16, 21, 9) {real, imag} */,
  {32'hbf3a0f00, 32'hc0092e5a} /* (16, 21, 8) {real, imag} */,
  {32'h400d3cc7, 32'hc1011628} /* (16, 21, 7) {real, imag} */,
  {32'h41531dfa, 32'h41d812b5} /* (16, 21, 6) {real, imag} */,
  {32'hc0d0c494, 32'h4197f5dc} /* (16, 21, 5) {real, imag} */,
  {32'h4114ca48, 32'hc12e70a4} /* (16, 21, 4) {real, imag} */,
  {32'h4191ae65, 32'h40b218b5} /* (16, 21, 3) {real, imag} */,
  {32'hc0132f28, 32'h3ec5c718} /* (16, 21, 2) {real, imag} */,
  {32'hbf2dca90, 32'h406b2840} /* (16, 21, 1) {real, imag} */,
  {32'h419acd5a, 32'hc121ac34} /* (16, 21, 0) {real, imag} */,
  {32'hbf8ca0dc, 32'hc0530146} /* (16, 20, 31) {real, imag} */,
  {32'hbe2d8900, 32'h401baf21} /* (16, 20, 30) {real, imag} */,
  {32'hc12a3deb, 32'hc114651a} /* (16, 20, 29) {real, imag} */,
  {32'hc06c15a6, 32'h40949879} /* (16, 20, 28) {real, imag} */,
  {32'hc0d7f7b3, 32'h409e2778} /* (16, 20, 27) {real, imag} */,
  {32'h40bec7d0, 32'h41130070} /* (16, 20, 26) {real, imag} */,
  {32'h40b749ad, 32'h3e5ddd20} /* (16, 20, 25) {real, imag} */,
  {32'hbf9d72a8, 32'hc18fad80} /* (16, 20, 24) {real, imag} */,
  {32'h4005e55c, 32'hbf9eed0c} /* (16, 20, 23) {real, imag} */,
  {32'h40e4edbe, 32'hc1410586} /* (16, 20, 22) {real, imag} */,
  {32'hc0caa815, 32'hc046dcb2} /* (16, 20, 21) {real, imag} */,
  {32'h40280910, 32'h4189a76c} /* (16, 20, 20) {real, imag} */,
  {32'hc0be43cf, 32'h4039cea8} /* (16, 20, 19) {real, imag} */,
  {32'hc10a1115, 32'h4125a04c} /* (16, 20, 18) {real, imag} */,
  {32'hbfd35114, 32'hc052ff1c} /* (16, 20, 17) {real, imag} */,
  {32'h3ecde2d4, 32'hbfb3ede2} /* (16, 20, 16) {real, imag} */,
  {32'hc0e543b2, 32'h419aa1a3} /* (16, 20, 15) {real, imag} */,
  {32'hc095ef9b, 32'hc1923193} /* (16, 20, 14) {real, imag} */,
  {32'h418b5523, 32'hc0030112} /* (16, 20, 13) {real, imag} */,
  {32'hc0c43a97, 32'h4084b8fa} /* (16, 20, 12) {real, imag} */,
  {32'hc18064a2, 32'h4103663b} /* (16, 20, 11) {real, imag} */,
  {32'hbff7669f, 32'hc18f40c2} /* (16, 20, 10) {real, imag} */,
  {32'hc129cab9, 32'hc0cde0b5} /* (16, 20, 9) {real, imag} */,
  {32'h40c091df, 32'h40a7a6a6} /* (16, 20, 8) {real, imag} */,
  {32'h3fe55f20, 32'hbeb20b78} /* (16, 20, 7) {real, imag} */,
  {32'h4075486d, 32'h41690f70} /* (16, 20, 6) {real, imag} */,
  {32'hc10237f4, 32'h408fa772} /* (16, 20, 5) {real, imag} */,
  {32'h3bc62200, 32'h3ee40a20} /* (16, 20, 4) {real, imag} */,
  {32'hc04d876b, 32'h41072dcc} /* (16, 20, 3) {real, imag} */,
  {32'h417a5444, 32'hc09e1ca2} /* (16, 20, 2) {real, imag} */,
  {32'hc127b835, 32'hbe5beec0} /* (16, 20, 1) {real, imag} */,
  {32'h40353da6, 32'h408e11fc} /* (16, 20, 0) {real, imag} */,
  {32'hc11735f4, 32'h41367d3e} /* (16, 19, 31) {real, imag} */,
  {32'hc0b53adb, 32'h3faebf2e} /* (16, 19, 30) {real, imag} */,
  {32'hc0603aec, 32'hc17da553} /* (16, 19, 29) {real, imag} */,
  {32'hbfe51d88, 32'h41346ff9} /* (16, 19, 28) {real, imag} */,
  {32'h3fa107b1, 32'h40bfe432} /* (16, 19, 27) {real, imag} */,
  {32'h3ff11356, 32'hc1db34e6} /* (16, 19, 26) {real, imag} */,
  {32'hc1414d4a, 32'h410f7559} /* (16, 19, 25) {real, imag} */,
  {32'h419d685c, 32'hbfe73930} /* (16, 19, 24) {real, imag} */,
  {32'hbd9de940, 32'hc1324954} /* (16, 19, 23) {real, imag} */,
  {32'h41895a34, 32'hc14cc114} /* (16, 19, 22) {real, imag} */,
  {32'hc0b3a8a6, 32'hc0ec4cc1} /* (16, 19, 21) {real, imag} */,
  {32'h40e5dda4, 32'h414e5280} /* (16, 19, 20) {real, imag} */,
  {32'hc062405c, 32'h3f8cb371} /* (16, 19, 19) {real, imag} */,
  {32'h40adba14, 32'hc02e1069} /* (16, 19, 18) {real, imag} */,
  {32'h412014d6, 32'h409e61aa} /* (16, 19, 17) {real, imag} */,
  {32'hc10de0fd, 32'h4102b515} /* (16, 19, 16) {real, imag} */,
  {32'h40182cd0, 32'hc07e1861} /* (16, 19, 15) {real, imag} */,
  {32'h4045b92c, 32'hbfb93ff4} /* (16, 19, 14) {real, imag} */,
  {32'h4112908a, 32'hc06599de} /* (16, 19, 13) {real, imag} */,
  {32'hc001eda8, 32'hc06ca543} /* (16, 19, 12) {real, imag} */,
  {32'h402edf42, 32'h401d035f} /* (16, 19, 11) {real, imag} */,
  {32'hbe59cc30, 32'h409a80e6} /* (16, 19, 10) {real, imag} */,
  {32'hc07d5580, 32'hc0200c42} /* (16, 19, 9) {real, imag} */,
  {32'hc182e43f, 32'h40f0c816} /* (16, 19, 8) {real, imag} */,
  {32'h3f7dd340, 32'hc184f1ee} /* (16, 19, 7) {real, imag} */,
  {32'hc181fd21, 32'hc11db568} /* (16, 19, 6) {real, imag} */,
  {32'h415bb36b, 32'hbfbe834c} /* (16, 19, 5) {real, imag} */,
  {32'hbc6ee680, 32'hc0787ed6} /* (16, 19, 4) {real, imag} */,
  {32'h40825cf3, 32'hc1273b38} /* (16, 19, 3) {real, imag} */,
  {32'h4088a2e3, 32'h40bdccd6} /* (16, 19, 2) {real, imag} */,
  {32'hbe4d4aa0, 32'h40489c7c} /* (16, 19, 1) {real, imag} */,
  {32'h4114ef5e, 32'h40d35019} /* (16, 19, 0) {real, imag} */,
  {32'h40ce0811, 32'hc01d3cce} /* (16, 18, 31) {real, imag} */,
  {32'hc08258b4, 32'h410b9474} /* (16, 18, 30) {real, imag} */,
  {32'h40bb583d, 32'h41264ab4} /* (16, 18, 29) {real, imag} */,
  {32'h40a7a766, 32'hc0dea23b} /* (16, 18, 28) {real, imag} */,
  {32'h3f18bf38, 32'h40926c6e} /* (16, 18, 27) {real, imag} */,
  {32'hc1300030, 32'h408ca6fa} /* (16, 18, 26) {real, imag} */,
  {32'hbf8c1a3c, 32'h4189a076} /* (16, 18, 25) {real, imag} */,
  {32'hc11262e9, 32'hc020357c} /* (16, 18, 24) {real, imag} */,
  {32'h3ee3f160, 32'h40b7537a} /* (16, 18, 23) {real, imag} */,
  {32'hbfc32a34, 32'h419cadaa} /* (16, 18, 22) {real, imag} */,
  {32'h406b5a4a, 32'h3f1b6af0} /* (16, 18, 21) {real, imag} */,
  {32'hc015d314, 32'hc1877534} /* (16, 18, 20) {real, imag} */,
  {32'h40ab97e1, 32'h410e0940} /* (16, 18, 19) {real, imag} */,
  {32'h3e722fe8, 32'hc127de98} /* (16, 18, 18) {real, imag} */,
  {32'h410966b6, 32'h3faaa1aa} /* (16, 18, 17) {real, imag} */,
  {32'hc134376f, 32'h3fd9a214} /* (16, 18, 16) {real, imag} */,
  {32'hc1112859, 32'hc15fe9f0} /* (16, 18, 15) {real, imag} */,
  {32'hc1115e02, 32'h3e4e7360} /* (16, 18, 14) {real, imag} */,
  {32'hc029e36c, 32'h4084f060} /* (16, 18, 13) {real, imag} */,
  {32'hc017e7e0, 32'hc0b4aeed} /* (16, 18, 12) {real, imag} */,
  {32'h41060fbe, 32'hc0498b72} /* (16, 18, 11) {real, imag} */,
  {32'hc12966ee, 32'h40e463ce} /* (16, 18, 10) {real, imag} */,
  {32'h3ffbe2ea, 32'h41915462} /* (16, 18, 9) {real, imag} */,
  {32'h4118d928, 32'h410de5a4} /* (16, 18, 8) {real, imag} */,
  {32'h40c580cf, 32'hc12c0560} /* (16, 18, 7) {real, imag} */,
  {32'h412c316c, 32'h408a96f7} /* (16, 18, 6) {real, imag} */,
  {32'h408d79e8, 32'hc1307d21} /* (16, 18, 5) {real, imag} */,
  {32'h41698586, 32'h410ef6af} /* (16, 18, 4) {real, imag} */,
  {32'h403fdb2b, 32'hbfd31278} /* (16, 18, 3) {real, imag} */,
  {32'h40968743, 32'h4032cf72} /* (16, 18, 2) {real, imag} */,
  {32'h40b2b50b, 32'hc134ad20} /* (16, 18, 1) {real, imag} */,
  {32'hc0eb84a3, 32'hc18a40de} /* (16, 18, 0) {real, imag} */,
  {32'hc0462245, 32'h410e5ac6} /* (16, 17, 31) {real, imag} */,
  {32'h408c0c53, 32'h3f09c638} /* (16, 17, 30) {real, imag} */,
  {32'h3fffac28, 32'hc13882e0} /* (16, 17, 29) {real, imag} */,
  {32'hbf263296, 32'hc0ace88e} /* (16, 17, 28) {real, imag} */,
  {32'hc0b2ce8a, 32'hbf6bbd3a} /* (16, 17, 27) {real, imag} */,
  {32'h3ed05840, 32'h412960f6} /* (16, 17, 26) {real, imag} */,
  {32'h3fca4774, 32'hc08dc8b8} /* (16, 17, 25) {real, imag} */,
  {32'hc07cc876, 32'h40cc1fb2} /* (16, 17, 24) {real, imag} */,
  {32'h412f9704, 32'h413012d3} /* (16, 17, 23) {real, imag} */,
  {32'hc0c944b3, 32'hc08e94a8} /* (16, 17, 22) {real, imag} */,
  {32'h40b99cd5, 32'h41af28b6} /* (16, 17, 21) {real, imag} */,
  {32'hc0443202, 32'h416906b5} /* (16, 17, 20) {real, imag} */,
  {32'h3e5cc100, 32'hc03a909b} /* (16, 17, 19) {real, imag} */,
  {32'hc110e5da, 32'h412e1f53} /* (16, 17, 18) {real, imag} */,
  {32'hc0088ea8, 32'h40f38a42} /* (16, 17, 17) {real, imag} */,
  {32'h3fb078d0, 32'hbdb92270} /* (16, 17, 16) {real, imag} */,
  {32'hbf22c0b8, 32'hc11075a8} /* (16, 17, 15) {real, imag} */,
  {32'h41394087, 32'hc0a7001b} /* (16, 17, 14) {real, imag} */,
  {32'hc0a6816c, 32'hc14575b7} /* (16, 17, 13) {real, imag} */,
  {32'hc078e5f0, 32'hc088d284} /* (16, 17, 12) {real, imag} */,
  {32'hc17bdc8f, 32'h40c0e90e} /* (16, 17, 11) {real, imag} */,
  {32'h4133e1bb, 32'h410b7ff0} /* (16, 17, 10) {real, imag} */,
  {32'h40e47389, 32'h4008c577} /* (16, 17, 9) {real, imag} */,
  {32'h40e63b2c, 32'hc002450b} /* (16, 17, 8) {real, imag} */,
  {32'h4100fd1a, 32'h41127b78} /* (16, 17, 7) {real, imag} */,
  {32'h40d1320d, 32'hc12fc0bc} /* (16, 17, 6) {real, imag} */,
  {32'hc09ccfb2, 32'h41244556} /* (16, 17, 5) {real, imag} */,
  {32'hbf2c2cdc, 32'h4077b260} /* (16, 17, 4) {real, imag} */,
  {32'h40f3a6d0, 32'h40bf046a} /* (16, 17, 3) {real, imag} */,
  {32'hc0f3aedc, 32'h3f3cb940} /* (16, 17, 2) {real, imag} */,
  {32'h409e6998, 32'hc06ee26a} /* (16, 17, 1) {real, imag} */,
  {32'h40016c62, 32'hc0618c12} /* (16, 17, 0) {real, imag} */,
  {32'h3e8f7344, 32'hc07d1b94} /* (16, 16, 31) {real, imag} */,
  {32'hbf108d80, 32'hc0d8f684} /* (16, 16, 30) {real, imag} */,
  {32'hc0ce884f, 32'h40795643} /* (16, 16, 29) {real, imag} */,
  {32'hbf9853d7, 32'hc1203216} /* (16, 16, 28) {real, imag} */,
  {32'hc0e7b5a0, 32'hc0c8bc34} /* (16, 16, 27) {real, imag} */,
  {32'hc0a17485, 32'h40af8b28} /* (16, 16, 26) {real, imag} */,
  {32'h410202a0, 32'h4105954a} /* (16, 16, 25) {real, imag} */,
  {32'hc1380873, 32'hc0a575bb} /* (16, 16, 24) {real, imag} */,
  {32'hc0a0b7f8, 32'hbe98c8c8} /* (16, 16, 23) {real, imag} */,
  {32'hc0a78fec, 32'h40c08f7a} /* (16, 16, 22) {real, imag} */,
  {32'h3ff5c469, 32'hc0a329dc} /* (16, 16, 21) {real, imag} */,
  {32'h414abf08, 32'hc125bf3a} /* (16, 16, 20) {real, imag} */,
  {32'hbe0c6f88, 32'h41124a00} /* (16, 16, 19) {real, imag} */,
  {32'h40823e92, 32'hc0e392b6} /* (16, 16, 18) {real, imag} */,
  {32'h401bc844, 32'h3c5e4e00} /* (16, 16, 17) {real, imag} */,
  {32'h4048067c, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h401bc844, 32'hbc5e4e00} /* (16, 16, 15) {real, imag} */,
  {32'h40823e92, 32'h40e392b6} /* (16, 16, 14) {real, imag} */,
  {32'hbe0c6f88, 32'hc1124a00} /* (16, 16, 13) {real, imag} */,
  {32'h414abf08, 32'h4125bf3a} /* (16, 16, 12) {real, imag} */,
  {32'h3ff5c469, 32'h40a329dc} /* (16, 16, 11) {real, imag} */,
  {32'hc0a78fec, 32'hc0c08f7a} /* (16, 16, 10) {real, imag} */,
  {32'hc0a0b7f8, 32'h3e98c8c8} /* (16, 16, 9) {real, imag} */,
  {32'hc1380873, 32'h40a575bb} /* (16, 16, 8) {real, imag} */,
  {32'h410202a0, 32'hc105954a} /* (16, 16, 7) {real, imag} */,
  {32'hc0a17485, 32'hc0af8b28} /* (16, 16, 6) {real, imag} */,
  {32'hc0e7b5a0, 32'h40c8bc34} /* (16, 16, 5) {real, imag} */,
  {32'hbf9853d7, 32'h41203216} /* (16, 16, 4) {real, imag} */,
  {32'hc0ce884f, 32'hc0795643} /* (16, 16, 3) {real, imag} */,
  {32'hbf108d80, 32'h40d8f684} /* (16, 16, 2) {real, imag} */,
  {32'h3e8f7344, 32'h407d1b94} /* (16, 16, 1) {real, imag} */,
  {32'hc09eef1f, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h409e6998, 32'h406ee26a} /* (16, 15, 31) {real, imag} */,
  {32'hc0f3aedc, 32'hbf3cb940} /* (16, 15, 30) {real, imag} */,
  {32'h40f3a6d0, 32'hc0bf046a} /* (16, 15, 29) {real, imag} */,
  {32'hbf2c2cdc, 32'hc077b260} /* (16, 15, 28) {real, imag} */,
  {32'hc09ccfb2, 32'hc1244556} /* (16, 15, 27) {real, imag} */,
  {32'h40d1320d, 32'h412fc0bc} /* (16, 15, 26) {real, imag} */,
  {32'h4100fd1a, 32'hc1127b78} /* (16, 15, 25) {real, imag} */,
  {32'h40e63b2c, 32'h4002450b} /* (16, 15, 24) {real, imag} */,
  {32'h40e47389, 32'hc008c577} /* (16, 15, 23) {real, imag} */,
  {32'h4133e1bb, 32'hc10b7ff0} /* (16, 15, 22) {real, imag} */,
  {32'hc17bdc8f, 32'hc0c0e90e} /* (16, 15, 21) {real, imag} */,
  {32'hc078e5f0, 32'h4088d284} /* (16, 15, 20) {real, imag} */,
  {32'hc0a6816c, 32'h414575b7} /* (16, 15, 19) {real, imag} */,
  {32'h41394087, 32'h40a7001b} /* (16, 15, 18) {real, imag} */,
  {32'hbf22c0b8, 32'h411075a8} /* (16, 15, 17) {real, imag} */,
  {32'h3fb078d0, 32'h3db92270} /* (16, 15, 16) {real, imag} */,
  {32'hc0088ea8, 32'hc0f38a42} /* (16, 15, 15) {real, imag} */,
  {32'hc110e5da, 32'hc12e1f53} /* (16, 15, 14) {real, imag} */,
  {32'h3e5cc100, 32'h403a909b} /* (16, 15, 13) {real, imag} */,
  {32'hc0443202, 32'hc16906b5} /* (16, 15, 12) {real, imag} */,
  {32'h40b99cd5, 32'hc1af28b6} /* (16, 15, 11) {real, imag} */,
  {32'hc0c944b3, 32'h408e94a8} /* (16, 15, 10) {real, imag} */,
  {32'h412f9704, 32'hc13012d3} /* (16, 15, 9) {real, imag} */,
  {32'hc07cc876, 32'hc0cc1fb2} /* (16, 15, 8) {real, imag} */,
  {32'h3fca4774, 32'h408dc8b8} /* (16, 15, 7) {real, imag} */,
  {32'h3ed05840, 32'hc12960f6} /* (16, 15, 6) {real, imag} */,
  {32'hc0b2ce8a, 32'h3f6bbd3a} /* (16, 15, 5) {real, imag} */,
  {32'hbf263296, 32'h40ace88e} /* (16, 15, 4) {real, imag} */,
  {32'h3fffac28, 32'h413882e0} /* (16, 15, 3) {real, imag} */,
  {32'h408c0c53, 32'hbf09c638} /* (16, 15, 2) {real, imag} */,
  {32'hc0462245, 32'hc10e5ac6} /* (16, 15, 1) {real, imag} */,
  {32'h40016c62, 32'h40618c12} /* (16, 15, 0) {real, imag} */,
  {32'h40b2b50b, 32'h4134ad20} /* (16, 14, 31) {real, imag} */,
  {32'h40968743, 32'hc032cf72} /* (16, 14, 30) {real, imag} */,
  {32'h403fdb2b, 32'h3fd31278} /* (16, 14, 29) {real, imag} */,
  {32'h41698586, 32'hc10ef6af} /* (16, 14, 28) {real, imag} */,
  {32'h408d79e8, 32'h41307d21} /* (16, 14, 27) {real, imag} */,
  {32'h412c316c, 32'hc08a96f7} /* (16, 14, 26) {real, imag} */,
  {32'h40c580cf, 32'h412c0560} /* (16, 14, 25) {real, imag} */,
  {32'h4118d928, 32'hc10de5a4} /* (16, 14, 24) {real, imag} */,
  {32'h3ffbe2ea, 32'hc1915462} /* (16, 14, 23) {real, imag} */,
  {32'hc12966ee, 32'hc0e463ce} /* (16, 14, 22) {real, imag} */,
  {32'h41060fbe, 32'h40498b72} /* (16, 14, 21) {real, imag} */,
  {32'hc017e7e0, 32'h40b4aeed} /* (16, 14, 20) {real, imag} */,
  {32'hc029e36c, 32'hc084f060} /* (16, 14, 19) {real, imag} */,
  {32'hc1115e02, 32'hbe4e7360} /* (16, 14, 18) {real, imag} */,
  {32'hc1112859, 32'h415fe9f0} /* (16, 14, 17) {real, imag} */,
  {32'hc134376f, 32'hbfd9a214} /* (16, 14, 16) {real, imag} */,
  {32'h410966b6, 32'hbfaaa1aa} /* (16, 14, 15) {real, imag} */,
  {32'h3e722fe8, 32'h4127de98} /* (16, 14, 14) {real, imag} */,
  {32'h40ab97e1, 32'hc10e0940} /* (16, 14, 13) {real, imag} */,
  {32'hc015d314, 32'h41877534} /* (16, 14, 12) {real, imag} */,
  {32'h406b5a4a, 32'hbf1b6af0} /* (16, 14, 11) {real, imag} */,
  {32'hbfc32a34, 32'hc19cadaa} /* (16, 14, 10) {real, imag} */,
  {32'h3ee3f160, 32'hc0b7537a} /* (16, 14, 9) {real, imag} */,
  {32'hc11262e9, 32'h4020357c} /* (16, 14, 8) {real, imag} */,
  {32'hbf8c1a3c, 32'hc189a076} /* (16, 14, 7) {real, imag} */,
  {32'hc1300030, 32'hc08ca6fa} /* (16, 14, 6) {real, imag} */,
  {32'h3f18bf38, 32'hc0926c6e} /* (16, 14, 5) {real, imag} */,
  {32'h40a7a766, 32'h40dea23b} /* (16, 14, 4) {real, imag} */,
  {32'h40bb583d, 32'hc1264ab4} /* (16, 14, 3) {real, imag} */,
  {32'hc08258b4, 32'hc10b9474} /* (16, 14, 2) {real, imag} */,
  {32'h40ce0811, 32'h401d3cce} /* (16, 14, 1) {real, imag} */,
  {32'hc0eb84a3, 32'h418a40de} /* (16, 14, 0) {real, imag} */,
  {32'hbe4d4aa0, 32'hc0489c7c} /* (16, 13, 31) {real, imag} */,
  {32'h4088a2e3, 32'hc0bdccd6} /* (16, 13, 30) {real, imag} */,
  {32'h40825cf3, 32'h41273b38} /* (16, 13, 29) {real, imag} */,
  {32'hbc6ee680, 32'h40787ed6} /* (16, 13, 28) {real, imag} */,
  {32'h415bb36b, 32'h3fbe834c} /* (16, 13, 27) {real, imag} */,
  {32'hc181fd21, 32'h411db568} /* (16, 13, 26) {real, imag} */,
  {32'h3f7dd340, 32'h4184f1ee} /* (16, 13, 25) {real, imag} */,
  {32'hc182e43f, 32'hc0f0c816} /* (16, 13, 24) {real, imag} */,
  {32'hc07d5580, 32'h40200c42} /* (16, 13, 23) {real, imag} */,
  {32'hbe59cc30, 32'hc09a80e6} /* (16, 13, 22) {real, imag} */,
  {32'h402edf42, 32'hc01d035f} /* (16, 13, 21) {real, imag} */,
  {32'hc001eda8, 32'h406ca543} /* (16, 13, 20) {real, imag} */,
  {32'h4112908a, 32'h406599de} /* (16, 13, 19) {real, imag} */,
  {32'h4045b92c, 32'h3fb93ff4} /* (16, 13, 18) {real, imag} */,
  {32'h40182cd0, 32'h407e1861} /* (16, 13, 17) {real, imag} */,
  {32'hc10de0fd, 32'hc102b515} /* (16, 13, 16) {real, imag} */,
  {32'h412014d6, 32'hc09e61aa} /* (16, 13, 15) {real, imag} */,
  {32'h40adba14, 32'h402e1069} /* (16, 13, 14) {real, imag} */,
  {32'hc062405c, 32'hbf8cb371} /* (16, 13, 13) {real, imag} */,
  {32'h40e5dda4, 32'hc14e5280} /* (16, 13, 12) {real, imag} */,
  {32'hc0b3a8a6, 32'h40ec4cc1} /* (16, 13, 11) {real, imag} */,
  {32'h41895a34, 32'h414cc114} /* (16, 13, 10) {real, imag} */,
  {32'hbd9de940, 32'h41324954} /* (16, 13, 9) {real, imag} */,
  {32'h419d685c, 32'h3fe73930} /* (16, 13, 8) {real, imag} */,
  {32'hc1414d4a, 32'hc10f7559} /* (16, 13, 7) {real, imag} */,
  {32'h3ff11356, 32'h41db34e6} /* (16, 13, 6) {real, imag} */,
  {32'h3fa107b1, 32'hc0bfe432} /* (16, 13, 5) {real, imag} */,
  {32'hbfe51d88, 32'hc1346ff9} /* (16, 13, 4) {real, imag} */,
  {32'hc0603aec, 32'h417da553} /* (16, 13, 3) {real, imag} */,
  {32'hc0b53adb, 32'hbfaebf2e} /* (16, 13, 2) {real, imag} */,
  {32'hc11735f4, 32'hc1367d3e} /* (16, 13, 1) {real, imag} */,
  {32'h4114ef5e, 32'hc0d35019} /* (16, 13, 0) {real, imag} */,
  {32'hc127b835, 32'h3e5beec0} /* (16, 12, 31) {real, imag} */,
  {32'h417a5444, 32'h409e1ca2} /* (16, 12, 30) {real, imag} */,
  {32'hc04d876b, 32'hc1072dcc} /* (16, 12, 29) {real, imag} */,
  {32'h3bc62200, 32'hbee40a20} /* (16, 12, 28) {real, imag} */,
  {32'hc10237f4, 32'hc08fa772} /* (16, 12, 27) {real, imag} */,
  {32'h4075486d, 32'hc1690f70} /* (16, 12, 26) {real, imag} */,
  {32'h3fe55f20, 32'h3eb20b78} /* (16, 12, 25) {real, imag} */,
  {32'h40c091df, 32'hc0a7a6a6} /* (16, 12, 24) {real, imag} */,
  {32'hc129cab9, 32'h40cde0b5} /* (16, 12, 23) {real, imag} */,
  {32'hbff7669f, 32'h418f40c2} /* (16, 12, 22) {real, imag} */,
  {32'hc18064a2, 32'hc103663b} /* (16, 12, 21) {real, imag} */,
  {32'hc0c43a97, 32'hc084b8fa} /* (16, 12, 20) {real, imag} */,
  {32'h418b5523, 32'h40030112} /* (16, 12, 19) {real, imag} */,
  {32'hc095ef9b, 32'h41923193} /* (16, 12, 18) {real, imag} */,
  {32'hc0e543b2, 32'hc19aa1a3} /* (16, 12, 17) {real, imag} */,
  {32'h3ecde2d4, 32'h3fb3ede2} /* (16, 12, 16) {real, imag} */,
  {32'hbfd35114, 32'h4052ff1c} /* (16, 12, 15) {real, imag} */,
  {32'hc10a1115, 32'hc125a04c} /* (16, 12, 14) {real, imag} */,
  {32'hc0be43cf, 32'hc039cea8} /* (16, 12, 13) {real, imag} */,
  {32'h40280910, 32'hc189a76c} /* (16, 12, 12) {real, imag} */,
  {32'hc0caa815, 32'h4046dcb2} /* (16, 12, 11) {real, imag} */,
  {32'h40e4edbe, 32'h41410586} /* (16, 12, 10) {real, imag} */,
  {32'h4005e55c, 32'h3f9eed0c} /* (16, 12, 9) {real, imag} */,
  {32'hbf9d72a8, 32'h418fad80} /* (16, 12, 8) {real, imag} */,
  {32'h40b749ad, 32'hbe5ddd20} /* (16, 12, 7) {real, imag} */,
  {32'h40bec7d0, 32'hc1130070} /* (16, 12, 6) {real, imag} */,
  {32'hc0d7f7b3, 32'hc09e2778} /* (16, 12, 5) {real, imag} */,
  {32'hc06c15a6, 32'hc0949879} /* (16, 12, 4) {real, imag} */,
  {32'hc12a3deb, 32'h4114651a} /* (16, 12, 3) {real, imag} */,
  {32'hbe2d8900, 32'hc01baf21} /* (16, 12, 2) {real, imag} */,
  {32'hbf8ca0dc, 32'h40530146} /* (16, 12, 1) {real, imag} */,
  {32'h40353da6, 32'hc08e11fc} /* (16, 12, 0) {real, imag} */,
  {32'hbf2dca90, 32'hc06b2840} /* (16, 11, 31) {real, imag} */,
  {32'hc0132f28, 32'hbec5c718} /* (16, 11, 30) {real, imag} */,
  {32'h4191ae65, 32'hc0b218b5} /* (16, 11, 29) {real, imag} */,
  {32'h4114ca48, 32'h412e70a4} /* (16, 11, 28) {real, imag} */,
  {32'hc0d0c494, 32'hc197f5dc} /* (16, 11, 27) {real, imag} */,
  {32'h41531dfa, 32'hc1d812b5} /* (16, 11, 26) {real, imag} */,
  {32'h400d3cc7, 32'h41011628} /* (16, 11, 25) {real, imag} */,
  {32'hbf3a0f00, 32'h40092e5a} /* (16, 11, 24) {real, imag} */,
  {32'h41ad8660, 32'hc07c98f8} /* (16, 11, 23) {real, imag} */,
  {32'h413a6004, 32'h4049f90c} /* (16, 11, 22) {real, imag} */,
  {32'hbf910e58, 32'hc07a6f0c} /* (16, 11, 21) {real, imag} */,
  {32'hc18e24ad, 32'h41c82e02} /* (16, 11, 20) {real, imag} */,
  {32'hc0cb0ea8, 32'h3f64ab00} /* (16, 11, 19) {real, imag} */,
  {32'h412eeffc, 32'h3ff08ddc} /* (16, 11, 18) {real, imag} */,
  {32'hc0b7c2ca, 32'hc09bbdef} /* (16, 11, 17) {real, imag} */,
  {32'hbdb92540, 32'h41637ff1} /* (16, 11, 16) {real, imag} */,
  {32'h4147d4fa, 32'h3b848200} /* (16, 11, 15) {real, imag} */,
  {32'hc149ad96, 32'hbf89afc4} /* (16, 11, 14) {real, imag} */,
  {32'hc1513d12, 32'h416d0ef4} /* (16, 11, 13) {real, imag} */,
  {32'hc10a1ba6, 32'hc0c2a748} /* (16, 11, 12) {real, imag} */,
  {32'h4150d457, 32'hc0fb1054} /* (16, 11, 11) {real, imag} */,
  {32'hc089cb2e, 32'hc0099941} /* (16, 11, 10) {real, imag} */,
  {32'hbfc309dc, 32'h4154321c} /* (16, 11, 9) {real, imag} */,
  {32'h4188b7f1, 32'h41aeef45} /* (16, 11, 8) {real, imag} */,
  {32'hc1ee11e8, 32'hbfcc8fc3} /* (16, 11, 7) {real, imag} */,
  {32'hc083fc47, 32'h407c1e84} /* (16, 11, 6) {real, imag} */,
  {32'h3f61d300, 32'hc113e7ba} /* (16, 11, 5) {real, imag} */,
  {32'hc1475cd6, 32'hc0720474} /* (16, 11, 4) {real, imag} */,
  {32'hc0d7c77b, 32'hc1190f94} /* (16, 11, 3) {real, imag} */,
  {32'h4105a62b, 32'hc12579a7} /* (16, 11, 2) {real, imag} */,
  {32'h40f42859, 32'h40fae46d} /* (16, 11, 1) {real, imag} */,
  {32'h419acd5a, 32'h4121ac34} /* (16, 11, 0) {real, imag} */,
  {32'h3f192688, 32'hc113b20e} /* (16, 10, 31) {real, imag} */,
  {32'h4183e306, 32'h418dbfdc} /* (16, 10, 30) {real, imag} */,
  {32'hc111d38c, 32'h4068439f} /* (16, 10, 29) {real, imag} */,
  {32'hc1861950, 32'hbfca81b8} /* (16, 10, 28) {real, imag} */,
  {32'hc190de90, 32'h409d5560} /* (16, 10, 27) {real, imag} */,
  {32'hc10ffbaa, 32'h41805166} /* (16, 10, 26) {real, imag} */,
  {32'hc17dbe89, 32'h409fb19a} /* (16, 10, 25) {real, imag} */,
  {32'hc0ce1d87, 32'h408491ee} /* (16, 10, 24) {real, imag} */,
  {32'h4150d99f, 32'hc1044364} /* (16, 10, 23) {real, imag} */,
  {32'hc0c8a849, 32'h413e0c27} /* (16, 10, 22) {real, imag} */,
  {32'hc03e9554, 32'hc1d67618} /* (16, 10, 21) {real, imag} */,
  {32'h416c0107, 32'hc182ad62} /* (16, 10, 20) {real, imag} */,
  {32'h41b5f964, 32'h41213ff7} /* (16, 10, 19) {real, imag} */,
  {32'h401cbb54, 32'h404d690d} /* (16, 10, 18) {real, imag} */,
  {32'h3fd9e73a, 32'h41bbc68c} /* (16, 10, 17) {real, imag} */,
  {32'hc135ff1a, 32'h4129d092} /* (16, 10, 16) {real, imag} */,
  {32'h40ce2324, 32'hc0b528d7} /* (16, 10, 15) {real, imag} */,
  {32'hc181e9fd, 32'h415701d3} /* (16, 10, 14) {real, imag} */,
  {32'h406387d8, 32'hc16f5fb5} /* (16, 10, 13) {real, imag} */,
  {32'hc17410a0, 32'h40bc72d6} /* (16, 10, 12) {real, imag} */,
  {32'h41194178, 32'h3dcb8a30} /* (16, 10, 11) {real, imag} */,
  {32'h41925ae8, 32'h4090f0c3} /* (16, 10, 10) {real, imag} */,
  {32'h40a40f4c, 32'h4030f870} /* (16, 10, 9) {real, imag} */,
  {32'hc11d4e97, 32'h41323c9e} /* (16, 10, 8) {real, imag} */,
  {32'h404f9478, 32'hc05f3462} /* (16, 10, 7) {real, imag} */,
  {32'h40461b26, 32'h414c05a0} /* (16, 10, 6) {real, imag} */,
  {32'h40ef9d00, 32'h40467517} /* (16, 10, 5) {real, imag} */,
  {32'h411b498c, 32'hc1ca9b39} /* (16, 10, 4) {real, imag} */,
  {32'hc0b65c0e, 32'hc0f121a2} /* (16, 10, 3) {real, imag} */,
  {32'h4121afc8, 32'hc082d55a} /* (16, 10, 2) {real, imag} */,
  {32'h3f01f0b0, 32'hc11a3298} /* (16, 10, 1) {real, imag} */,
  {32'hc08ae0e6, 32'hbea43d30} /* (16, 10, 0) {real, imag} */,
  {32'hc0eced88, 32'h41791898} /* (16, 9, 31) {real, imag} */,
  {32'hc13af3aa, 32'h40866a1b} /* (16, 9, 30) {real, imag} */,
  {32'h4107e81b, 32'hc104da68} /* (16, 9, 29) {real, imag} */,
  {32'hc10fdbb2, 32'h403330c0} /* (16, 9, 28) {real, imag} */,
  {32'h411325f2, 32'hc0a3b785} /* (16, 9, 27) {real, imag} */,
  {32'h41b22a8b, 32'h4107132c} /* (16, 9, 26) {real, imag} */,
  {32'h3ffb3ede, 32'hc156a950} /* (16, 9, 25) {real, imag} */,
  {32'h3efe5800, 32'h4077aa8b} /* (16, 9, 24) {real, imag} */,
  {32'hc1381999, 32'h416d484c} /* (16, 9, 23) {real, imag} */,
  {32'hc108ef1f, 32'h415b6b3a} /* (16, 9, 22) {real, imag} */,
  {32'hc10d8e04, 32'hc1173746} /* (16, 9, 21) {real, imag} */,
  {32'h40e9cf4b, 32'h4144b732} /* (16, 9, 20) {real, imag} */,
  {32'hbff7874a, 32'hc0a0cb22} /* (16, 9, 19) {real, imag} */,
  {32'h40fc7b59, 32'h41381228} /* (16, 9, 18) {real, imag} */,
  {32'h4112a36e, 32'h41072ae6} /* (16, 9, 17) {real, imag} */,
  {32'hbf2eb338, 32'h41113a07} /* (16, 9, 16) {real, imag} */,
  {32'h40e01d24, 32'h410dc252} /* (16, 9, 15) {real, imag} */,
  {32'h40f95a54, 32'hbf759184} /* (16, 9, 14) {real, imag} */,
  {32'hc0a33aa7, 32'h3f62496c} /* (16, 9, 13) {real, imag} */,
  {32'h40ba1339, 32'h40b4a265} /* (16, 9, 12) {real, imag} */,
  {32'h410ed7ec, 32'h4119cf89} /* (16, 9, 11) {real, imag} */,
  {32'hc1a1ca96, 32'hc1199872} /* (16, 9, 10) {real, imag} */,
  {32'h41343dc9, 32'h414405ae} /* (16, 9, 9) {real, imag} */,
  {32'hc13e5da1, 32'h40a3af6b} /* (16, 9, 8) {real, imag} */,
  {32'h419af1cb, 32'h40c793c6} /* (16, 9, 7) {real, imag} */,
  {32'h418ab3b2, 32'hc1b89c90} /* (16, 9, 6) {real, imag} */,
  {32'h3fc9154b, 32'hbe894d40} /* (16, 9, 5) {real, imag} */,
  {32'hc1293bb8, 32'h412c3dab} /* (16, 9, 4) {real, imag} */,
  {32'h401851d6, 32'hbe1e1d80} /* (16, 9, 3) {real, imag} */,
  {32'hc1595fe8, 32'h41d94b4e} /* (16, 9, 2) {real, imag} */,
  {32'hc10f69c9, 32'hc0e1725c} /* (16, 9, 1) {real, imag} */,
  {32'h4101cf3d, 32'hc180fb34} /* (16, 9, 0) {real, imag} */,
  {32'h40f92d32, 32'h420e7938} /* (16, 8, 31) {real, imag} */,
  {32'hc1be68b2, 32'hc16fd801} /* (16, 8, 30) {real, imag} */,
  {32'hc1685e3a, 32'hbee9b080} /* (16, 8, 29) {real, imag} */,
  {32'h40df0298, 32'hc181a8fe} /* (16, 8, 28) {real, imag} */,
  {32'hc117b41f, 32'h3f2d34ac} /* (16, 8, 27) {real, imag} */,
  {32'hc208a4fb, 32'h418385de} /* (16, 8, 26) {real, imag} */,
  {32'h3e15fc60, 32'hc116bd29} /* (16, 8, 25) {real, imag} */,
  {32'hc1bb4e97, 32'hbfe17ca0} /* (16, 8, 24) {real, imag} */,
  {32'h41952c9a, 32'hc084102d} /* (16, 8, 23) {real, imag} */,
  {32'hc134f0c2, 32'hc18589df} /* (16, 8, 22) {real, imag} */,
  {32'h3e031f10, 32'h410b4763} /* (16, 8, 21) {real, imag} */,
  {32'hc06dd372, 32'h407afdcc} /* (16, 8, 20) {real, imag} */,
  {32'hc18f07fa, 32'hc16f5374} /* (16, 8, 19) {real, imag} */,
  {32'h40c9b438, 32'h4124083c} /* (16, 8, 18) {real, imag} */,
  {32'h40251ffb, 32'hbf416e2a} /* (16, 8, 17) {real, imag} */,
  {32'hbff5c088, 32'h40e756d5} /* (16, 8, 16) {real, imag} */,
  {32'h41636aee, 32'h40b147ac} /* (16, 8, 15) {real, imag} */,
  {32'hc089583c, 32'h4119f0ed} /* (16, 8, 14) {real, imag} */,
  {32'hc0abf8c2, 32'h3f4aca60} /* (16, 8, 13) {real, imag} */,
  {32'h4146f27e, 32'h40093d4e} /* (16, 8, 12) {real, imag} */,
  {32'hc15ff4e4, 32'h413cdc1a} /* (16, 8, 11) {real, imag} */,
  {32'hc1403fbe, 32'h40c652de} /* (16, 8, 10) {real, imag} */,
  {32'h4131c973, 32'h4021db98} /* (16, 8, 9) {real, imag} */,
  {32'hc01cbd02, 32'hc170eb11} /* (16, 8, 8) {real, imag} */,
  {32'hc1199166, 32'h41881508} /* (16, 8, 7) {real, imag} */,
  {32'h416302e4, 32'hc19518b9} /* (16, 8, 6) {real, imag} */,
  {32'h413de063, 32'hc17b5a17} /* (16, 8, 5) {real, imag} */,
  {32'h3fc75044, 32'hc1a0916d} /* (16, 8, 4) {real, imag} */,
  {32'hc1100690, 32'h412a6a21} /* (16, 8, 3) {real, imag} */,
  {32'hc0e2054c, 32'h3fe75f36} /* (16, 8, 2) {real, imag} */,
  {32'h41bafc54, 32'h41f19911} /* (16, 8, 1) {real, imag} */,
  {32'h4174daed, 32'h4116a838} /* (16, 8, 0) {real, imag} */,
  {32'h3ff3a648, 32'h4203c1b0} /* (16, 7, 31) {real, imag} */,
  {32'h415938be, 32'hc1bf75e4} /* (16, 7, 30) {real, imag} */,
  {32'hc1bd531a, 32'hbef08240} /* (16, 7, 29) {real, imag} */,
  {32'hc17ebc5e, 32'h40e17932} /* (16, 7, 28) {real, imag} */,
  {32'hc02c55ef, 32'hbf42a76c} /* (16, 7, 27) {real, imag} */,
  {32'h409d4e34, 32'hc08a75e8} /* (16, 7, 26) {real, imag} */,
  {32'hc0dda323, 32'hc03ba25a} /* (16, 7, 25) {real, imag} */,
  {32'hc001e20f, 32'h3dacad80} /* (16, 7, 24) {real, imag} */,
  {32'h4173b8a2, 32'h40ed1bb8} /* (16, 7, 23) {real, imag} */,
  {32'h40cc6de2, 32'hc0f47b89} /* (16, 7, 22) {real, imag} */,
  {32'h410dc0ac, 32'h40b6abdc} /* (16, 7, 21) {real, imag} */,
  {32'hc1ad22ab, 32'h408904e0} /* (16, 7, 20) {real, imag} */,
  {32'h408fc175, 32'hc1bd2980} /* (16, 7, 19) {real, imag} */,
  {32'hc0bcd34b, 32'hc0dc146b} /* (16, 7, 18) {real, imag} */,
  {32'hc0ea4d8c, 32'hc0091450} /* (16, 7, 17) {real, imag} */,
  {32'h40e91d02, 32'hc0a83555} /* (16, 7, 16) {real, imag} */,
  {32'hc177365a, 32'h40f63554} /* (16, 7, 15) {real, imag} */,
  {32'h410f3f86, 32'h3fdf0ce2} /* (16, 7, 14) {real, imag} */,
  {32'hc1167886, 32'hc1572bce} /* (16, 7, 13) {real, imag} */,
  {32'hc0e7da49, 32'hbf6be698} /* (16, 7, 12) {real, imag} */,
  {32'h411cb243, 32'hc16dec23} /* (16, 7, 11) {real, imag} */,
  {32'h3fe64f44, 32'h4146108e} /* (16, 7, 10) {real, imag} */,
  {32'hc0b48c16, 32'hc11f5a90} /* (16, 7, 9) {real, imag} */,
  {32'hc1481bec, 32'hbf9ca6bc} /* (16, 7, 8) {real, imag} */,
  {32'h4038b28d, 32'hbfcc36d8} /* (16, 7, 7) {real, imag} */,
  {32'hc0f4ca63, 32'hc0f88243} /* (16, 7, 6) {real, imag} */,
  {32'h40c54229, 32'h4107814e} /* (16, 7, 5) {real, imag} */,
  {32'h419a940c, 32'h40be27ed} /* (16, 7, 4) {real, imag} */,
  {32'hc025b60c, 32'hc0697c23} /* (16, 7, 3) {real, imag} */,
  {32'h4115fb1a, 32'hc1641866} /* (16, 7, 2) {real, imag} */,
  {32'hc20e2258, 32'h41412336} /* (16, 7, 1) {real, imag} */,
  {32'hc02b7490, 32'hc1321a3c} /* (16, 7, 0) {real, imag} */,
  {32'h416a83e1, 32'h400e69cc} /* (16, 6, 31) {real, imag} */,
  {32'hc1e34a9f, 32'h40531000} /* (16, 6, 30) {real, imag} */,
  {32'h3f6cebe4, 32'hc1c6318b} /* (16, 6, 29) {real, imag} */,
  {32'hc1039244, 32'h413650b5} /* (16, 6, 28) {real, imag} */,
  {32'hbc417c00, 32'h406afc42} /* (16, 6, 27) {real, imag} */,
  {32'hc01ebc74, 32'hc0512764} /* (16, 6, 26) {real, imag} */,
  {32'h405e029e, 32'h418cbda7} /* (16, 6, 25) {real, imag} */,
  {32'h401fc3c1, 32'hc16846a6} /* (16, 6, 24) {real, imag} */,
  {32'hc0eb0490, 32'h3fb19bc0} /* (16, 6, 23) {real, imag} */,
  {32'h40dc52dc, 32'hbff3cbfc} /* (16, 6, 22) {real, imag} */,
  {32'hbeaf36b0, 32'h408860fc} /* (16, 6, 21) {real, imag} */,
  {32'hbfb5a018, 32'hc1b85db2} /* (16, 6, 20) {real, imag} */,
  {32'h40f8964e, 32'h3fa533bf} /* (16, 6, 19) {real, imag} */,
  {32'hc0205ba6, 32'hc1901716} /* (16, 6, 18) {real, imag} */,
  {32'h40c7ac93, 32'h3f1e9f4a} /* (16, 6, 17) {real, imag} */,
  {32'hc00b14c0, 32'hbff03d4a} /* (16, 6, 16) {real, imag} */,
  {32'h40abb11d, 32'h4101672d} /* (16, 6, 15) {real, imag} */,
  {32'h414f250a, 32'h40ae7ffe} /* (16, 6, 14) {real, imag} */,
  {32'h413acf5e, 32'hc1843cfb} /* (16, 6, 13) {real, imag} */,
  {32'h4143dae3, 32'hbeb15270} /* (16, 6, 12) {real, imag} */,
  {32'hc15df51b, 32'h4118e706} /* (16, 6, 11) {real, imag} */,
  {32'hc1a48c5d, 32'h402dc1ac} /* (16, 6, 10) {real, imag} */,
  {32'h3e2c44e0, 32'hbfad4c3c} /* (16, 6, 9) {real, imag} */,
  {32'hc011c108, 32'hc1803afc} /* (16, 6, 8) {real, imag} */,
  {32'h41af4862, 32'h3fe719f8} /* (16, 6, 7) {real, imag} */,
  {32'h4078c06a, 32'h3e09c6b0} /* (16, 6, 6) {real, imag} */,
  {32'hc0350853, 32'hc09c36f4} /* (16, 6, 5) {real, imag} */,
  {32'h3fa327c0, 32'h41b0f047} /* (16, 6, 4) {real, imag} */,
  {32'h40960241, 32'h40ee1746} /* (16, 6, 3) {real, imag} */,
  {32'h4149149e, 32'hc07bba58} /* (16, 6, 2) {real, imag} */,
  {32'h419c7b22, 32'h403cc0b0} /* (16, 6, 1) {real, imag} */,
  {32'hc164373a, 32'hc1c7785a} /* (16, 6, 0) {real, imag} */,
  {32'h425146f0, 32'h41eab79a} /* (16, 5, 31) {real, imag} */,
  {32'hc1dde820, 32'hc1dae196} /* (16, 5, 30) {real, imag} */,
  {32'h41318f0c, 32'h41d2cc37} /* (16, 5, 29) {real, imag} */,
  {32'h401dce72, 32'h415b7df2} /* (16, 5, 28) {real, imag} */,
  {32'h405db322, 32'h41a6a638} /* (16, 5, 27) {real, imag} */,
  {32'hc06144db, 32'h4185ebf2} /* (16, 5, 26) {real, imag} */,
  {32'hc0d4e649, 32'hc0c34098} /* (16, 5, 25) {real, imag} */,
  {32'hc1b94790, 32'h41429a9f} /* (16, 5, 24) {real, imag} */,
  {32'hc103a542, 32'h3fd8a9e8} /* (16, 5, 23) {real, imag} */,
  {32'h3f1b9680, 32'h413b0653} /* (16, 5, 22) {real, imag} */,
  {32'hc08bab9e, 32'hc0d14531} /* (16, 5, 21) {real, imag} */,
  {32'hc12b2d92, 32'h3f8b64e0} /* (16, 5, 20) {real, imag} */,
  {32'h3e7db080, 32'hc130760e} /* (16, 5, 19) {real, imag} */,
  {32'h402f3984, 32'hbfab52b8} /* (16, 5, 18) {real, imag} */,
  {32'h3fc84a76, 32'h3f80c8e1} /* (16, 5, 17) {real, imag} */,
  {32'hc12e3380, 32'h410d46b1} /* (16, 5, 16) {real, imag} */,
  {32'hc11c228f, 32'h412bbf3b} /* (16, 5, 15) {real, imag} */,
  {32'h41093b1a, 32'hc06ac28b} /* (16, 5, 14) {real, imag} */,
  {32'hc0051cda, 32'hc06a0f04} /* (16, 5, 13) {real, imag} */,
  {32'h416e77ad, 32'h4118a145} /* (16, 5, 12) {real, imag} */,
  {32'h418f13c0, 32'h41018f4d} /* (16, 5, 11) {real, imag} */,
  {32'hc1041c64, 32'hc1c378ea} /* (16, 5, 10) {real, imag} */,
  {32'hc178c88c, 32'h401e1b2a} /* (16, 5, 9) {real, imag} */,
  {32'h40ce175e, 32'h411a4fe6} /* (16, 5, 8) {real, imag} */,
  {32'hbf9854b8, 32'h4186caac} /* (16, 5, 7) {real, imag} */,
  {32'hc04f8582, 32'h40cf2bf4} /* (16, 5, 6) {real, imag} */,
  {32'hc1e00008, 32'h41dcbb5b} /* (16, 5, 5) {real, imag} */,
  {32'h4154b8f5, 32'h3f632e98} /* (16, 5, 4) {real, imag} */,
  {32'hc12489dd, 32'hbfb24d8c} /* (16, 5, 3) {real, imag} */,
  {32'hc046f4b8, 32'hc2366d87} /* (16, 5, 2) {real, imag} */,
  {32'h41a0dc8e, 32'h425c1706} /* (16, 5, 1) {real, imag} */,
  {32'h413619bc, 32'h4224ad66} /* (16, 5, 0) {real, imag} */,
  {32'hc0fef748, 32'hc28e53ee} /* (16, 4, 31) {real, imag} */,
  {32'h420f346b, 32'h41c7f420} /* (16, 4, 30) {real, imag} */,
  {32'hc020bf02, 32'hc21ae6e1} /* (16, 4, 29) {real, imag} */,
  {32'hc21c27aa, 32'h40fc8e5e} /* (16, 4, 28) {real, imag} */,
  {32'h4194e39b, 32'h40a89d65} /* (16, 4, 27) {real, imag} */,
  {32'hc1259ff8, 32'h408d4d5f} /* (16, 4, 26) {real, imag} */,
  {32'hc19cb690, 32'h3d317400} /* (16, 4, 25) {real, imag} */,
  {32'h42099a8e, 32'hc1b8d4ff} /* (16, 4, 24) {real, imag} */,
  {32'h402cfae6, 32'h3f69bf10} /* (16, 4, 23) {real, imag} */,
  {32'h4061fc82, 32'h4085ff20} /* (16, 4, 22) {real, imag} */,
  {32'hbf64ad36, 32'hc0baa582} /* (16, 4, 21) {real, imag} */,
  {32'hc0053f98, 32'h40cc0c12} /* (16, 4, 20) {real, imag} */,
  {32'h3fa4c4b0, 32'h4064b6d6} /* (16, 4, 19) {real, imag} */,
  {32'h4092e2e9, 32'h4027d58e} /* (16, 4, 18) {real, imag} */,
  {32'hc10576e6, 32'h3f8c59a6} /* (16, 4, 17) {real, imag} */,
  {32'hc09e3c68, 32'hc09ae6a6} /* (16, 4, 16) {real, imag} */,
  {32'h41146a74, 32'hc04a939e} /* (16, 4, 15) {real, imag} */,
  {32'hc0a41c75, 32'h40ce2ff2} /* (16, 4, 14) {real, imag} */,
  {32'hc14b4da3, 32'h4105ef57} /* (16, 4, 13) {real, imag} */,
  {32'h40707691, 32'h400a6a56} /* (16, 4, 12) {real, imag} */,
  {32'hc0cb16fe, 32'hc11ec8b7} /* (16, 4, 11) {real, imag} */,
  {32'h41a38449, 32'h40094c7c} /* (16, 4, 10) {real, imag} */,
  {32'hc11930da, 32'h4181ad64} /* (16, 4, 9) {real, imag} */,
  {32'h4191f692, 32'h412d68be} /* (16, 4, 8) {real, imag} */,
  {32'hc1db095a, 32'hc0960a48} /* (16, 4, 7) {real, imag} */,
  {32'hc123d011, 32'hc124bb9c} /* (16, 4, 6) {real, imag} */,
  {32'hc18aae12, 32'h410239a2} /* (16, 4, 5) {real, imag} */,
  {32'hc103fc49, 32'hc1d7fa27} /* (16, 4, 4) {real, imag} */,
  {32'hc17d33a6, 32'hc08b24d8} /* (16, 4, 3) {real, imag} */,
  {32'h42176092, 32'h4278c2f9} /* (16, 4, 2) {real, imag} */,
  {32'hc20ce2be, 32'hc215a388} /* (16, 4, 1) {real, imag} */,
  {32'hc28acaa1, 32'hc296486a} /* (16, 4, 0) {real, imag} */,
  {32'h42d5e0dc, 32'hc250b5ec} /* (16, 3, 31) {real, imag} */,
  {32'h41ab2c82, 32'h42a46962} /* (16, 3, 30) {real, imag} */,
  {32'hc1c8b58a, 32'h41979098} /* (16, 3, 29) {real, imag} */,
  {32'hc146e227, 32'h3fbf4d74} /* (16, 3, 28) {real, imag} */,
  {32'h416191b8, 32'h40668ad4} /* (16, 3, 27) {real, imag} */,
  {32'hc0188f58, 32'h3fa196b6} /* (16, 3, 26) {real, imag} */,
  {32'hc1baa252, 32'h41abb9e5} /* (16, 3, 25) {real, imag} */,
  {32'hc0dcea7a, 32'hbff58794} /* (16, 3, 24) {real, imag} */,
  {32'hc1512ec5, 32'h40178b56} /* (16, 3, 23) {real, imag} */,
  {32'h3e96ec70, 32'hc0c0ba5d} /* (16, 3, 22) {real, imag} */,
  {32'h41502bdd, 32'h3f9431be} /* (16, 3, 21) {real, imag} */,
  {32'hbea18910, 32'h406ab9b7} /* (16, 3, 20) {real, imag} */,
  {32'hbfff8368, 32'hc101c5aa} /* (16, 3, 19) {real, imag} */,
  {32'hbf35b548, 32'hc0b23e14} /* (16, 3, 18) {real, imag} */,
  {32'hc09ac3ce, 32'hc03295e6} /* (16, 3, 17) {real, imag} */,
  {32'h4094aec2, 32'h40d777d5} /* (16, 3, 16) {real, imag} */,
  {32'h4148a698, 32'h412f8729} /* (16, 3, 15) {real, imag} */,
  {32'h414d49bd, 32'hbffc036a} /* (16, 3, 14) {real, imag} */,
  {32'hc14d823d, 32'hc0ba483a} /* (16, 3, 13) {real, imag} */,
  {32'hc1316220, 32'hc0fecc8b} /* (16, 3, 12) {real, imag} */,
  {32'h4167c226, 32'hc09fbefd} /* (16, 3, 11) {real, imag} */,
  {32'h3eeacb50, 32'hc188e3c5} /* (16, 3, 10) {real, imag} */,
  {32'hc18f8df1, 32'h40e87389} /* (16, 3, 9) {real, imag} */,
  {32'h4002eb04, 32'hc18226a3} /* (16, 3, 8) {real, imag} */,
  {32'hc0d0444c, 32'hc11b23b6} /* (16, 3, 7) {real, imag} */,
  {32'hc18005d0, 32'h408311c2} /* (16, 3, 6) {real, imag} */,
  {32'hc18e1e02, 32'h41002733} /* (16, 3, 5) {real, imag} */,
  {32'h4190803e, 32'h419d0864} /* (16, 3, 4) {real, imag} */,
  {32'h410cfc1b, 32'hc17dfa0d} /* (16, 3, 3) {real, imag} */,
  {32'h42971188, 32'h4216f3d0} /* (16, 3, 2) {real, imag} */,
  {32'hc2026ac2, 32'hc2a3f852} /* (16, 3, 1) {real, imag} */,
  {32'h41905f7a, 32'h41a4b14b} /* (16, 3, 0) {real, imag} */,
  {32'h43b5b55c, 32'hc2082d55} /* (16, 2, 31) {real, imag} */,
  {32'hc32b9d67, 32'h4216c7cd} /* (16, 2, 30) {real, imag} */,
  {32'h4290f9ee, 32'h41a6bee2} /* (16, 2, 29) {real, imag} */,
  {32'h41c53ad6, 32'hc1b337ce} /* (16, 2, 28) {real, imag} */,
  {32'hc1fd5c0e, 32'h4196de1c} /* (16, 2, 27) {real, imag} */,
  {32'h408f1896, 32'h4164c2ed} /* (16, 2, 26) {real, imag} */,
  {32'h41d35b7e, 32'hc2144c77} /* (16, 2, 25) {real, imag} */,
  {32'hc2085792, 32'h41566ed8} /* (16, 2, 24) {real, imag} */,
  {32'hc14c89d3, 32'h418cc3a5} /* (16, 2, 23) {real, imag} */,
  {32'hc04edfa3, 32'hc0ca6495} /* (16, 2, 22) {real, imag} */,
  {32'h3e024e20, 32'h41c0d919} /* (16, 2, 21) {real, imag} */,
  {32'h40b6fcaa, 32'hc087d80a} /* (16, 2, 20) {real, imag} */,
  {32'hc134a8cc, 32'hbf36c77e} /* (16, 2, 19) {real, imag} */,
  {32'hc029ca0b, 32'hbec3d998} /* (16, 2, 18) {real, imag} */,
  {32'hc1054dc6, 32'hc04b1777} /* (16, 2, 17) {real, imag} */,
  {32'hc032db5d, 32'h40aae302} /* (16, 2, 16) {real, imag} */,
  {32'hc142b1cf, 32'h402eceec} /* (16, 2, 15) {real, imag} */,
  {32'hc100a7b6, 32'hc1363e1f} /* (16, 2, 14) {real, imag} */,
  {32'h40883189, 32'h41295024} /* (16, 2, 13) {real, imag} */,
  {32'hc1b2f796, 32'h410b6330} /* (16, 2, 12) {real, imag} */,
  {32'h3f6ce7e8, 32'hc133794e} /* (16, 2, 11) {real, imag} */,
  {32'hc0e9d6d9, 32'h411f7780} /* (16, 2, 10) {real, imag} */,
  {32'hc1375fee, 32'h41413fc8} /* (16, 2, 9) {real, imag} */,
  {32'hbf889ec0, 32'hc19e9816} /* (16, 2, 8) {real, imag} */,
  {32'h41015ed4, 32'hc1a8dbae} /* (16, 2, 7) {real, imag} */,
  {32'h41460f24, 32'h42086788} /* (16, 2, 6) {real, imag} */,
  {32'hc227d671, 32'hc205cc47} /* (16, 2, 5) {real, imag} */,
  {32'h428cd20f, 32'hc27ba005} /* (16, 2, 4) {real, imag} */,
  {32'h424e23a5, 32'hc208953e} /* (16, 2, 3) {real, imag} */,
  {32'hc3135ae8, 32'h42557096} /* (16, 2, 2) {real, imag} */,
  {32'h43525d58, 32'hc2874e32} /* (16, 2, 1) {real, imag} */,
  {32'h432463d3, 32'h4289471a} /* (16, 2, 0) {real, imag} */,
  {32'hc3a9e471, 32'h41f7d62e} /* (16, 1, 31) {real, imag} */,
  {32'h42ceb9cb, 32'hc22d3df8} /* (16, 1, 30) {real, imag} */,
  {32'hc0a62fb2, 32'h42161134} /* (16, 1, 29) {real, imag} */,
  {32'hc1e7daa7, 32'hc27fb5b5} /* (16, 1, 28) {real, imag} */,
  {32'h42ac0bc7, 32'hc06f9e22} /* (16, 1, 27) {real, imag} */,
  {32'h421fb484, 32'hbf3e6d20} /* (16, 1, 26) {real, imag} */,
  {32'hc122288c, 32'h41317902} /* (16, 1, 25) {real, imag} */,
  {32'hbe9a22b0, 32'hc14ca71f} /* (16, 1, 24) {real, imag} */,
  {32'hc147fb94, 32'h4161bd66} /* (16, 1, 23) {real, imag} */,
  {32'hc095f084, 32'h40d65155} /* (16, 1, 22) {real, imag} */,
  {32'hbf805608, 32'hc1b04976} /* (16, 1, 21) {real, imag} */,
  {32'h40c597a8, 32'hc1496438} /* (16, 1, 20) {real, imag} */,
  {32'h3e571d80, 32'h4150cc18} /* (16, 1, 19) {real, imag} */,
  {32'h400488e8, 32'h40c4c194} /* (16, 1, 18) {real, imag} */,
  {32'hc13d88f8, 32'hc0659aef} /* (16, 1, 17) {real, imag} */,
  {32'hc0c43076, 32'h413151b0} /* (16, 1, 16) {real, imag} */,
  {32'hbf38b92c, 32'h40952676} /* (16, 1, 15) {real, imag} */,
  {32'hbf2c29cc, 32'h40e4d42a} /* (16, 1, 14) {real, imag} */,
  {32'h3eba93a8, 32'h4057d8c8} /* (16, 1, 13) {real, imag} */,
  {32'hc10bd5c4, 32'hc1aa38c2} /* (16, 1, 12) {real, imag} */,
  {32'h40754fc6, 32'h41cf6f50} /* (16, 1, 11) {real, imag} */,
  {32'h40878c98, 32'h4061d634} /* (16, 1, 10) {real, imag} */,
  {32'h41128433, 32'h40ffd64c} /* (16, 1, 9) {real, imag} */,
  {32'h40fe7128, 32'h41bd5189} /* (16, 1, 8) {real, imag} */,
  {32'hc00f8e26, 32'hc1a0ac28} /* (16, 1, 7) {real, imag} */,
  {32'hc090c21a, 32'h419679ee} /* (16, 1, 6) {real, imag} */,
  {32'h427660e2, 32'h41f518ce} /* (16, 1, 5) {real, imag} */,
  {32'hc23a5c66, 32'hc1249777} /* (16, 1, 4) {real, imag} */,
  {32'hc1fee1ff, 32'h413a5880} /* (16, 1, 3) {real, imag} */,
  {32'h43003086, 32'h43542f73} /* (16, 1, 2) {real, imag} */,
  {32'hc416a040, 32'hc370ba5d} /* (16, 1, 1) {real, imag} */,
  {32'hc3dbf39e, 32'hc356e162} /* (16, 1, 0) {real, imag} */,
  {32'hc3e20ab6, 32'h4390a64a} /* (16, 0, 31) {real, imag} */,
  {32'h41f42fc5, 32'hc2c73f5d} /* (16, 0, 30) {real, imag} */,
  {32'h41fe0f7d, 32'h410ad063} /* (16, 0, 29) {real, imag} */,
  {32'hc1b7660c, 32'hc20cbb86} /* (16, 0, 28) {real, imag} */,
  {32'h4146f808, 32'h402514b8} /* (16, 0, 27) {real, imag} */,
  {32'h415da8ad, 32'hc1562bfb} /* (16, 0, 26) {real, imag} */,
  {32'h408ac698, 32'hc0db7eea} /* (16, 0, 25) {real, imag} */,
  {32'h40d52678, 32'hc0adb9b2} /* (16, 0, 24) {real, imag} */,
  {32'h41945767, 32'hc0c64972} /* (16, 0, 23) {real, imag} */,
  {32'hbf58ca10, 32'h3ef49bc0} /* (16, 0, 22) {real, imag} */,
  {32'h4000c83c, 32'hc0ccbe07} /* (16, 0, 21) {real, imag} */,
  {32'h40d5eba4, 32'h3edeb5b0} /* (16, 0, 20) {real, imag} */,
  {32'hc0845d26, 32'h3f863b3b} /* (16, 0, 19) {real, imag} */,
  {32'hc14611c8, 32'h3fbb0930} /* (16, 0, 18) {real, imag} */,
  {32'h40503e54, 32'hc0eab21c} /* (16, 0, 17) {real, imag} */,
  {32'hc00d19a7, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h40503e54, 32'h40eab21c} /* (16, 0, 15) {real, imag} */,
  {32'hc14611c8, 32'hbfbb0930} /* (16, 0, 14) {real, imag} */,
  {32'hc0845d26, 32'hbf863b3b} /* (16, 0, 13) {real, imag} */,
  {32'h40d5eba4, 32'hbedeb5b0} /* (16, 0, 12) {real, imag} */,
  {32'h4000c83c, 32'h40ccbe07} /* (16, 0, 11) {real, imag} */,
  {32'hbf58ca10, 32'hbef49bc0} /* (16, 0, 10) {real, imag} */,
  {32'h41945767, 32'h40c64972} /* (16, 0, 9) {real, imag} */,
  {32'h40d52678, 32'h40adb9b2} /* (16, 0, 8) {real, imag} */,
  {32'h408ac698, 32'h40db7eea} /* (16, 0, 7) {real, imag} */,
  {32'h415da8ad, 32'h41562bfb} /* (16, 0, 6) {real, imag} */,
  {32'h4146f808, 32'hc02514b8} /* (16, 0, 5) {real, imag} */,
  {32'hc1b7660c, 32'h420cbb86} /* (16, 0, 4) {real, imag} */,
  {32'h41fe0f7d, 32'hc10ad063} /* (16, 0, 3) {real, imag} */,
  {32'h41f42fc5, 32'h42c73f5d} /* (16, 0, 2) {real, imag} */,
  {32'hc3e20ab6, 32'hc390a64a} /* (16, 0, 1) {real, imag} */,
  {32'hc3c20fa8, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h43deba7e, 32'hc3a76652} /* (15, 31, 31) {real, imag} */,
  {32'hc3582234, 32'h43079866} /* (15, 31, 30) {real, imag} */,
  {32'hc27e0c61, 32'hc0ef4938} /* (15, 31, 29) {real, imag} */,
  {32'hc1c0ee98, 32'hc230abe2} /* (15, 31, 28) {real, imag} */,
  {32'hc1470a0a, 32'h41239f68} /* (15, 31, 27) {real, imag} */,
  {32'h415d400e, 32'h4177816f} /* (15, 31, 26) {real, imag} */,
  {32'h41e36749, 32'hc133a78e} /* (15, 31, 25) {real, imag} */,
  {32'hc19c2dfb, 32'h41a15b96} /* (15, 31, 24) {real, imag} */,
  {32'h3f2a78da, 32'hc0b2ed53} /* (15, 31, 23) {real, imag} */,
  {32'h400bcd7e, 32'h410aad7a} /* (15, 31, 22) {real, imag} */,
  {32'hc0f318b2, 32'h3f52feb0} /* (15, 31, 21) {real, imag} */,
  {32'hc1062490, 32'h41933f61} /* (15, 31, 20) {real, imag} */,
  {32'h4177cc9e, 32'h3f90055a} /* (15, 31, 19) {real, imag} */,
  {32'h413ef1c5, 32'h40ef4662} /* (15, 31, 18) {real, imag} */,
  {32'hc0fa9b04, 32'hc10faaf0} /* (15, 31, 17) {real, imag} */,
  {32'h40aa6adf, 32'h418bfdf0} /* (15, 31, 16) {real, imag} */,
  {32'h412a92c4, 32'h40562f48} /* (15, 31, 15) {real, imag} */,
  {32'hc0563de8, 32'hc10bc191} /* (15, 31, 14) {real, imag} */,
  {32'h40c26fe1, 32'hc1987dd0} /* (15, 31, 13) {real, imag} */,
  {32'h4160bff3, 32'h3fcbd704} /* (15, 31, 12) {real, imag} */,
  {32'hc1764074, 32'hc103b3d4} /* (15, 31, 11) {real, imag} */,
  {32'h4187daa9, 32'h40a7086c} /* (15, 31, 10) {real, imag} */,
  {32'hc143235a, 32'hc187b618} /* (15, 31, 9) {real, imag} */,
  {32'hc149a74e, 32'hc135d01a} /* (15, 31, 8) {real, imag} */,
  {32'hc010a002, 32'hc16a7351} /* (15, 31, 7) {real, imag} */,
  {32'h41d73571, 32'h417115ce} /* (15, 31, 6) {real, imag} */,
  {32'hc2310238, 32'hc1b4d6e6} /* (15, 31, 5) {real, imag} */,
  {32'h42458192, 32'h41999196} /* (15, 31, 4) {real, imag} */,
  {32'hc0c0fadc, 32'hc27f0978} /* (15, 31, 3) {real, imag} */,
  {32'hc3104efa, 32'h4218cc8b} /* (15, 31, 2) {real, imag} */,
  {32'h43d60f50, 32'h43086eb9} /* (15, 31, 1) {real, imag} */,
  {32'h43d4b47b, 32'h42ce2f16} /* (15, 31, 0) {real, imag} */,
  {32'hc31dbeae, 32'h41aa6c18} /* (15, 30, 31) {real, imag} */,
  {32'h42ec5e68, 32'h41312d1c} /* (15, 30, 30) {real, imag} */,
  {32'h41ab8b3f, 32'h410a9278} /* (15, 30, 29) {real, imag} */,
  {32'h40e9a620, 32'h427a85c9} /* (15, 30, 28) {real, imag} */,
  {32'h41bfdd0d, 32'hc2279d04} /* (15, 30, 27) {real, imag} */,
  {32'h4020a6df, 32'hc164eab7} /* (15, 30, 26) {real, imag} */,
  {32'hbe2ab738, 32'hc0d32c30} /* (15, 30, 25) {real, imag} */,
  {32'h41f18c62, 32'hbff18db0} /* (15, 30, 24) {real, imag} */,
  {32'hc10bf8c0, 32'hc1005efe} /* (15, 30, 23) {real, imag} */,
  {32'hc18bedac, 32'h41065a68} /* (15, 30, 22) {real, imag} */,
  {32'hc12d1c62, 32'hc110aedd} /* (15, 30, 21) {real, imag} */,
  {32'h408e462c, 32'hc1486628} /* (15, 30, 20) {real, imag} */,
  {32'h40940144, 32'h3fb0bfba} /* (15, 30, 19) {real, imag} */,
  {32'h40bc4161, 32'hc1796a64} /* (15, 30, 18) {real, imag} */,
  {32'h3ee3c278, 32'h408d37ae} /* (15, 30, 17) {real, imag} */,
  {32'hc0bb5706, 32'h40dd9872} /* (15, 30, 16) {real, imag} */,
  {32'hbff66c02, 32'h4048f7fe} /* (15, 30, 15) {real, imag} */,
  {32'h3fc22708, 32'hc08be652} /* (15, 30, 14) {real, imag} */,
  {32'hc0cee376, 32'hc122f9d4} /* (15, 30, 13) {real, imag} */,
  {32'hc0fb40f8, 32'h3eb09e00} /* (15, 30, 12) {real, imag} */,
  {32'h3f6e42e8, 32'h40faeb06} /* (15, 30, 11) {real, imag} */,
  {32'h40de441a, 32'h40c4be1e} /* (15, 30, 10) {real, imag} */,
  {32'hc15177fa, 32'hc171ec78} /* (15, 30, 9) {real, imag} */,
  {32'h41812e38, 32'h4238869f} /* (15, 30, 8) {real, imag} */,
  {32'hc0b6ed96, 32'hc0956dc5} /* (15, 30, 7) {real, imag} */,
  {32'hc1bbffd0, 32'hc20c132a} /* (15, 30, 6) {real, imag} */,
  {32'h4103ec76, 32'h40e96154} /* (15, 30, 5) {real, imag} */,
  {32'hc1a3d818, 32'hc2585694} /* (15, 30, 4) {real, imag} */,
  {32'h4200f102, 32'hc20c7ea2} /* (15, 30, 3) {real, imag} */,
  {32'h433a0394, 32'h4214978c} /* (15, 30, 2) {real, imag} */,
  {32'hc39cc5a7, 32'h429cc922} /* (15, 30, 1) {real, imag} */,
  {32'hc34446ee, 32'hc0618e20} /* (15, 30, 0) {real, imag} */,
  {32'h42687e13, 32'hc0a0f4f0} /* (15, 29, 31) {real, imag} */,
  {32'h4145a74e, 32'h42200cd7} /* (15, 29, 30) {real, imag} */,
  {32'h409d4050, 32'hc1775db8} /* (15, 29, 29) {real, imag} */,
  {32'hc192c4f2, 32'hc1ec8acc} /* (15, 29, 28) {real, imag} */,
  {32'h413b5d54, 32'hc143e139} /* (15, 29, 27) {real, imag} */,
  {32'hc08373ec, 32'hc0cf5ec6} /* (15, 29, 26) {real, imag} */,
  {32'hc1205b99, 32'h4101857c} /* (15, 29, 25) {real, imag} */,
  {32'h40873249, 32'h40d4793f} /* (15, 29, 24) {real, imag} */,
  {32'hc1371e38, 32'hbf70825c} /* (15, 29, 23) {real, imag} */,
  {32'hc0979c0c, 32'hc0999ac6} /* (15, 29, 22) {real, imag} */,
  {32'hc127e2a5, 32'hc11a2dd3} /* (15, 29, 21) {real, imag} */,
  {32'h4091e365, 32'h40b995d2} /* (15, 29, 20) {real, imag} */,
  {32'h4108c562, 32'hc133722d} /* (15, 29, 19) {real, imag} */,
  {32'hbf21b824, 32'hbf8a287a} /* (15, 29, 18) {real, imag} */,
  {32'hc0e17484, 32'h40614d6d} /* (15, 29, 17) {real, imag} */,
  {32'hbf599f38, 32'h408d8b9c} /* (15, 29, 16) {real, imag} */,
  {32'h3fc2587c, 32'hc178e007} /* (15, 29, 15) {real, imag} */,
  {32'h405418f0, 32'h41554048} /* (15, 29, 14) {real, imag} */,
  {32'hbfd85dc6, 32'h4167f592} /* (15, 29, 13) {real, imag} */,
  {32'hc0e0f4ea, 32'hc1b8a196} /* (15, 29, 12) {real, imag} */,
  {32'hc057112c, 32'h4115ea64} /* (15, 29, 11) {real, imag} */,
  {32'h412be82a, 32'h40a6f92a} /* (15, 29, 10) {real, imag} */,
  {32'hc18bfd10, 32'hc0d30932} /* (15, 29, 9) {real, imag} */,
  {32'hc1776c19, 32'h413fae00} /* (15, 29, 8) {real, imag} */,
  {32'hc1afa7cf, 32'hbf6e18a0} /* (15, 29, 7) {real, imag} */,
  {32'hbec9b4c0, 32'hc1b87748} /* (15, 29, 6) {real, imag} */,
  {32'hc0dd8e40, 32'hc12c4008} /* (15, 29, 5) {real, imag} */,
  {32'h41cf13ec, 32'hc17940f6} /* (15, 29, 4) {real, imag} */,
  {32'hc1d71ca0, 32'h410c5562} /* (15, 29, 3) {real, imag} */,
  {32'h4237d485, 32'h419d1ab0} /* (15, 29, 2) {real, imag} */,
  {32'h41835fde, 32'h3d397800} /* (15, 29, 1) {real, imag} */,
  {32'h412d938e, 32'hc1f45722} /* (15, 29, 0) {real, imag} */,
  {32'h42c7996a, 32'hc19f55d5} /* (15, 28, 31) {real, imag} */,
  {32'hc13dcab8, 32'h4236e4eb} /* (15, 28, 30) {real, imag} */,
  {32'hc18ee141, 32'hc1bc9308} /* (15, 28, 29) {real, imag} */,
  {32'hc184f422, 32'hc12c464b} /* (15, 28, 28) {real, imag} */,
  {32'hc1bbe5f9, 32'h415232e4} /* (15, 28, 27) {real, imag} */,
  {32'hc1c13c7e, 32'h41bb5633} /* (15, 28, 26) {real, imag} */,
  {32'h413dc926, 32'hc1e73398} /* (15, 28, 25) {real, imag} */,
  {32'hc1452cb2, 32'h40c349f0} /* (15, 28, 24) {real, imag} */,
  {32'h40b4424c, 32'h40c54cbd} /* (15, 28, 23) {real, imag} */,
  {32'h4170a6e2, 32'h4186eef5} /* (15, 28, 22) {real, imag} */,
  {32'h4140b383, 32'hc0b6149a} /* (15, 28, 21) {real, imag} */,
  {32'h3f8ee8b4, 32'hc02aff94} /* (15, 28, 20) {real, imag} */,
  {32'h414316b5, 32'hbff07f50} /* (15, 28, 19) {real, imag} */,
  {32'hc0e3e2d4, 32'h40bd7ebd} /* (15, 28, 18) {real, imag} */,
  {32'hc082eb07, 32'hc18e0cb9} /* (15, 28, 17) {real, imag} */,
  {32'hc0d91c69, 32'h40b6950c} /* (15, 28, 16) {real, imag} */,
  {32'h4012a4c6, 32'h40aa39e5} /* (15, 28, 15) {real, imag} */,
  {32'h40cb6a14, 32'h40ca8c5e} /* (15, 28, 14) {real, imag} */,
  {32'hc16e9b47, 32'hc0acf6d6} /* (15, 28, 13) {real, imag} */,
  {32'hbe2c5b70, 32'h40cebf23} /* (15, 28, 12) {real, imag} */,
  {32'h3f2b2f62, 32'h40a8e580} /* (15, 28, 11) {real, imag} */,
  {32'hbf874bb6, 32'h40c7aa4c} /* (15, 28, 10) {real, imag} */,
  {32'hc0a34b2e, 32'h3fe84f6e} /* (15, 28, 9) {real, imag} */,
  {32'h40633658, 32'h3e99cdc0} /* (15, 28, 8) {real, imag} */,
  {32'hc10e1cb0, 32'hc214df92} /* (15, 28, 7) {real, imag} */,
  {32'hc1110838, 32'hc18d1f41} /* (15, 28, 6) {real, imag} */,
  {32'hc1a20fc4, 32'hc0a29844} /* (15, 28, 5) {real, imag} */,
  {32'h42006e5c, 32'hc194af2e} /* (15, 28, 4) {real, imag} */,
  {32'h403725e0, 32'h419e83b8} /* (15, 28, 3) {real, imag} */,
  {32'hc19e6d60, 32'h4196f5ba} /* (15, 28, 2) {real, imag} */,
  {32'h421d9fbc, 32'hbfb72c80} /* (15, 28, 1) {real, imag} */,
  {32'hc1dc134a, 32'h4218548b} /* (15, 28, 0) {real, imag} */,
  {32'hc2554f7e, 32'h41374c58} /* (15, 27, 31) {real, imag} */,
  {32'h411b8e68, 32'hc19f5f70} /* (15, 27, 30) {real, imag} */,
  {32'h419041b0, 32'h4195d2e4} /* (15, 27, 29) {real, imag} */,
  {32'h41a29328, 32'h4131d82c} /* (15, 27, 28) {real, imag} */,
  {32'h4114528c, 32'hc0f739e2} /* (15, 27, 27) {real, imag} */,
  {32'h40fec830, 32'h3f707600} /* (15, 27, 26) {real, imag} */,
  {32'hc08fb8ea, 32'h4020ec10} /* (15, 27, 25) {real, imag} */,
  {32'h40a37cce, 32'hc1ca2ad7} /* (15, 27, 24) {real, imag} */,
  {32'hc125f42a, 32'h41596398} /* (15, 27, 23) {real, imag} */,
  {32'hc09a2fca, 32'h4149022a} /* (15, 27, 22) {real, imag} */,
  {32'hc013142e, 32'hc0ee9bb6} /* (15, 27, 21) {real, imag} */,
  {32'hc08d3b8b, 32'h4089d9dc} /* (15, 27, 20) {real, imag} */,
  {32'hc11c9fae, 32'h3fa3f114} /* (15, 27, 19) {real, imag} */,
  {32'hc12a67df, 32'h40a3a5d1} /* (15, 27, 18) {real, imag} */,
  {32'h417cbc4c, 32'hc0021428} /* (15, 27, 17) {real, imag} */,
  {32'hc0feeb64, 32'h400219f4} /* (15, 27, 16) {real, imag} */,
  {32'hc0d9b8a8, 32'h4169f82a} /* (15, 27, 15) {real, imag} */,
  {32'h40c56958, 32'h3f8869b4} /* (15, 27, 14) {real, imag} */,
  {32'hc005f2a7, 32'h4004c9bf} /* (15, 27, 13) {real, imag} */,
  {32'hc030c4dc, 32'h40b5ca5f} /* (15, 27, 12) {real, imag} */,
  {32'h3ea58570, 32'hbfbf9576} /* (15, 27, 11) {real, imag} */,
  {32'h40b86be6, 32'h416881ec} /* (15, 27, 10) {real, imag} */,
  {32'hc121cadc, 32'hc04791d8} /* (15, 27, 9) {real, imag} */,
  {32'hc146b8e2, 32'h3fe5e3b4} /* (15, 27, 8) {real, imag} */,
  {32'hc2248c64, 32'hc0c2bd64} /* (15, 27, 7) {real, imag} */,
  {32'hbf94ffb4, 32'h41286480} /* (15, 27, 6) {real, imag} */,
  {32'h41465102, 32'hc1e2d8af} /* (15, 27, 5) {real, imag} */,
  {32'h404d1a90, 32'hbf779cb8} /* (15, 27, 4) {real, imag} */,
  {32'h3fbfdc1c, 32'hc1a0c403} /* (15, 27, 3) {real, imag} */,
  {32'h4077cc00, 32'h415b8776} /* (15, 27, 2) {real, imag} */,
  {32'hc211640a, 32'hc23dcea6} /* (15, 27, 1) {real, imag} */,
  {32'hc24179e4, 32'h4038dc30} /* (15, 27, 0) {real, imag} */,
  {32'h41a77bff, 32'hc1d5ce2e} /* (15, 26, 31) {real, imag} */,
  {32'h41a767b2, 32'hc1834c19} /* (15, 26, 30) {real, imag} */,
  {32'h41564445, 32'hc0a7c6c5} /* (15, 26, 29) {real, imag} */,
  {32'hc1432d5e, 32'hc08defba} /* (15, 26, 28) {real, imag} */,
  {32'h41472324, 32'h4100d02c} /* (15, 26, 27) {real, imag} */,
  {32'hc0be2efe, 32'hc117208e} /* (15, 26, 26) {real, imag} */,
  {32'hc098c8d2, 32'hbf544c94} /* (15, 26, 25) {real, imag} */,
  {32'hc1813df1, 32'h411cedeb} /* (15, 26, 24) {real, imag} */,
  {32'h411a7126, 32'hc1021f3a} /* (15, 26, 23) {real, imag} */,
  {32'hc10c38f6, 32'hc196ef9e} /* (15, 26, 22) {real, imag} */,
  {32'h40b2ad73, 32'hc0b177f8} /* (15, 26, 21) {real, imag} */,
  {32'h4022c340, 32'hc0efb8be} /* (15, 26, 20) {real, imag} */,
  {32'h3d3a1ce0, 32'hbfd59a68} /* (15, 26, 19) {real, imag} */,
  {32'h40190b4e, 32'hc1386f18} /* (15, 26, 18) {real, imag} */,
  {32'h4100214b, 32'h409a8350} /* (15, 26, 17) {real, imag} */,
  {32'h402fa00a, 32'hc1742f66} /* (15, 26, 16) {real, imag} */,
  {32'h40afda9a, 32'h40bc33da} /* (15, 26, 15) {real, imag} */,
  {32'h412a8d6e, 32'h4089ad78} /* (15, 26, 14) {real, imag} */,
  {32'hc11133e3, 32'h40a15578} /* (15, 26, 13) {real, imag} */,
  {32'hc1ad6aca, 32'hc06cd050} /* (15, 26, 12) {real, imag} */,
  {32'hc085623b, 32'hc116834e} /* (15, 26, 11) {real, imag} */,
  {32'h406b982c, 32'hc0bf6acd} /* (15, 26, 10) {real, imag} */,
  {32'h413916e0, 32'h40b9addc} /* (15, 26, 9) {real, imag} */,
  {32'h3faab5d8, 32'h4152285a} /* (15, 26, 8) {real, imag} */,
  {32'hc1979a1a, 32'hc0b2b79d} /* (15, 26, 7) {real, imag} */,
  {32'hc112b338, 32'h3fe4f512} /* (15, 26, 6) {real, imag} */,
  {32'hc185bbba, 32'hc017e1ae} /* (15, 26, 5) {real, imag} */,
  {32'hc0997bfb, 32'hc07e0b64} /* (15, 26, 4) {real, imag} */,
  {32'hc094832c, 32'hbd9fe200} /* (15, 26, 3) {real, imag} */,
  {32'hc10c4c8c, 32'hc02aa0e2} /* (15, 26, 2) {real, imag} */,
  {32'hc02e55e0, 32'hc0800aec} /* (15, 26, 1) {real, imag} */,
  {32'hc1c276ba, 32'h40ff1662} /* (15, 26, 0) {real, imag} */,
  {32'hc173f4ce, 32'hc23bc676} /* (15, 25, 31) {real, imag} */,
  {32'h40065af0, 32'h40e4b8f3} /* (15, 25, 30) {real, imag} */,
  {32'hc0b8fe40, 32'h419afd12} /* (15, 25, 29) {real, imag} */,
  {32'h40aa9560, 32'h400d7d96} /* (15, 25, 28) {real, imag} */,
  {32'hc10381b0, 32'hbf836770} /* (15, 25, 27) {real, imag} */,
  {32'hc1b76059, 32'hc00575c0} /* (15, 25, 26) {real, imag} */,
  {32'h416723e0, 32'hc172931c} /* (15, 25, 25) {real, imag} */,
  {32'h404734d8, 32'h41c3afac} /* (15, 25, 24) {real, imag} */,
  {32'hc1665b4a, 32'hc09e1e08} /* (15, 25, 23) {real, imag} */,
  {32'hc0d579bb, 32'hc122093c} /* (15, 25, 22) {real, imag} */,
  {32'h40dcd702, 32'hc0eb1839} /* (15, 25, 21) {real, imag} */,
  {32'h3fdb1f98, 32'hc05a05a8} /* (15, 25, 20) {real, imag} */,
  {32'hc05f3f45, 32'h40a71ed0} /* (15, 25, 19) {real, imag} */,
  {32'h40b721ee, 32'hc0e19244} /* (15, 25, 18) {real, imag} */,
  {32'hc1a4a7f4, 32'h40fd1a4a} /* (15, 25, 17) {real, imag} */,
  {32'h40b38f60, 32'h4015410c} /* (15, 25, 16) {real, imag} */,
  {32'h4053c8d6, 32'h406792b3} /* (15, 25, 15) {real, imag} */,
  {32'hc09891b0, 32'h400ecda0} /* (15, 25, 14) {real, imag} */,
  {32'h3f856e3c, 32'h412966a8} /* (15, 25, 13) {real, imag} */,
  {32'h3ef7a16c, 32'h40fd5cd6} /* (15, 25, 12) {real, imag} */,
  {32'hc00b7bd2, 32'hc103f200} /* (15, 25, 11) {real, imag} */,
  {32'h3f86d1ec, 32'hc006a0d2} /* (15, 25, 10) {real, imag} */,
  {32'hc11a118a, 32'hbfe632f0} /* (15, 25, 9) {real, imag} */,
  {32'hc106301e, 32'hbfa71cc0} /* (15, 25, 8) {real, imag} */,
  {32'hbffdae48, 32'h4119eca1} /* (15, 25, 7) {real, imag} */,
  {32'hc0d12498, 32'h3ff655cf} /* (15, 25, 6) {real, imag} */,
  {32'hbfed4d60, 32'h40883c28} /* (15, 25, 5) {real, imag} */,
  {32'hc1574ada, 32'h4139a3a9} /* (15, 25, 4) {real, imag} */,
  {32'hc1215c1a, 32'h40020f95} /* (15, 25, 3) {real, imag} */,
  {32'hc0a4f2e0, 32'h41d2b5d8} /* (15, 25, 2) {real, imag} */,
  {32'h408f8f94, 32'hc1d30667} /* (15, 25, 1) {real, imag} */,
  {32'hc11173b2, 32'h40b3d8de} /* (15, 25, 0) {real, imag} */,
  {32'hc12135f8, 32'hbfa03034} /* (15, 24, 31) {real, imag} */,
  {32'h40d942dc, 32'hc12cadc0} /* (15, 24, 30) {real, imag} */,
  {32'hc123cc91, 32'hc0c32fc6} /* (15, 24, 29) {real, imag} */,
  {32'hc19eede4, 32'h40d5b193} /* (15, 24, 28) {real, imag} */,
  {32'hc161fe98, 32'hbea0e3d0} /* (15, 24, 27) {real, imag} */,
  {32'hc053ecc0, 32'h41ad07a5} /* (15, 24, 26) {real, imag} */,
  {32'hc0bbeffe, 32'h40d624d1} /* (15, 24, 25) {real, imag} */,
  {32'h41b98e6d, 32'h4120452c} /* (15, 24, 24) {real, imag} */,
  {32'hc0c0f554, 32'hc1b17861} /* (15, 24, 23) {real, imag} */,
  {32'h418c8918, 32'hc08277b6} /* (15, 24, 22) {real, imag} */,
  {32'h410946a8, 32'hbffdf039} /* (15, 24, 21) {real, imag} */,
  {32'hc1db646c, 32'hc15cfacc} /* (15, 24, 20) {real, imag} */,
  {32'hc0a8b95b, 32'hc0aac47c} /* (15, 24, 19) {real, imag} */,
  {32'h40c5ee66, 32'h3ec625b0} /* (15, 24, 18) {real, imag} */,
  {32'hbf732558, 32'hbf50199c} /* (15, 24, 17) {real, imag} */,
  {32'h40725459, 32'h4032c0e6} /* (15, 24, 16) {real, imag} */,
  {32'h3de01b00, 32'h418f4e94} /* (15, 24, 15) {real, imag} */,
  {32'hbffa0596, 32'hc0f80001} /* (15, 24, 14) {real, imag} */,
  {32'hc13127b6, 32'h410deb73} /* (15, 24, 13) {real, imag} */,
  {32'h3fe9cbd0, 32'hc1ceaec4} /* (15, 24, 12) {real, imag} */,
  {32'h412f2227, 32'hc089b929} /* (15, 24, 11) {real, imag} */,
  {32'h4199e225, 32'hc005f594} /* (15, 24, 10) {real, imag} */,
  {32'h3dd68e60, 32'hc05a2ef9} /* (15, 24, 9) {real, imag} */,
  {32'h412266ed, 32'h41a9dcbd} /* (15, 24, 8) {real, imag} */,
  {32'hc1288eda, 32'h41943f6a} /* (15, 24, 7) {real, imag} */,
  {32'h415ab47d, 32'hc17b1ad0} /* (15, 24, 6) {real, imag} */,
  {32'h40be9d01, 32'h3e9cc868} /* (15, 24, 5) {real, imag} */,
  {32'h4114b431, 32'hbeea31c8} /* (15, 24, 4) {real, imag} */,
  {32'h4126f42d, 32'hc016e0b0} /* (15, 24, 3) {real, imag} */,
  {32'h41064daf, 32'h40db79ee} /* (15, 24, 2) {real, imag} */,
  {32'hc2429f92, 32'h41e6403c} /* (15, 24, 1) {real, imag} */,
  {32'hc15e19bc, 32'hc178a85e} /* (15, 24, 0) {real, imag} */,
  {32'h408861eb, 32'hc17a34c4} /* (15, 23, 31) {real, imag} */,
  {32'h3fe3c11d, 32'h411d3a9a} /* (15, 23, 30) {real, imag} */,
  {32'h4090f282, 32'hbffb17ec} /* (15, 23, 29) {real, imag} */,
  {32'h40833f1e, 32'hc097cd32} /* (15, 23, 28) {real, imag} */,
  {32'hc13dd375, 32'h3faf994c} /* (15, 23, 27) {real, imag} */,
  {32'h4122def8, 32'h3f65c474} /* (15, 23, 26) {real, imag} */,
  {32'hc18507d4, 32'hc12c7ce9} /* (15, 23, 25) {real, imag} */,
  {32'hc0410ae4, 32'hbeb3cff0} /* (15, 23, 24) {real, imag} */,
  {32'h41f3e339, 32'hc0f880e8} /* (15, 23, 23) {real, imag} */,
  {32'hc13feab6, 32'h417933fa} /* (15, 23, 22) {real, imag} */,
  {32'hc0b6edc6, 32'h40ce0796} /* (15, 23, 21) {real, imag} */,
  {32'h3d8b9040, 32'h4087c416} /* (15, 23, 20) {real, imag} */,
  {32'h418da9e6, 32'hc121560c} /* (15, 23, 19) {real, imag} */,
  {32'hc147de34, 32'hbfe16fb8} /* (15, 23, 18) {real, imag} */,
  {32'h4031e910, 32'h4118f60c} /* (15, 23, 17) {real, imag} */,
  {32'h3f80c388, 32'hc0b1c279} /* (15, 23, 16) {real, imag} */,
  {32'hc0c8a230, 32'h411b818a} /* (15, 23, 15) {real, imag} */,
  {32'hc1ad5a77, 32'h410be229} /* (15, 23, 14) {real, imag} */,
  {32'h412232a6, 32'hc057059e} /* (15, 23, 13) {real, imag} */,
  {32'h409d0e71, 32'hbf8ff480} /* (15, 23, 12) {real, imag} */,
  {32'h41849ac8, 32'hc1220442} /* (15, 23, 11) {real, imag} */,
  {32'hc103ef04, 32'hc10f584f} /* (15, 23, 10) {real, imag} */,
  {32'h3eb7cfc8, 32'hbfadb888} /* (15, 23, 9) {real, imag} */,
  {32'h40660bdc, 32'h41697ce5} /* (15, 23, 8) {real, imag} */,
  {32'h412a85e2, 32'h41158ec2} /* (15, 23, 7) {real, imag} */,
  {32'h412614f0, 32'hc01b0288} /* (15, 23, 6) {real, imag} */,
  {32'h410848ce, 32'h412d4a82} /* (15, 23, 5) {real, imag} */,
  {32'hc06b7816, 32'hc1d003c5} /* (15, 23, 4) {real, imag} */,
  {32'h4146c516, 32'h3f44f5d0} /* (15, 23, 3) {real, imag} */,
  {32'h3f1ffb38, 32'h40405d1c} /* (15, 23, 2) {real, imag} */,
  {32'hc1cbdbc6, 32'h3fe84b0c} /* (15, 23, 1) {real, imag} */,
  {32'h413cd3ad, 32'hc066b44f} /* (15, 23, 0) {real, imag} */,
  {32'h412bde19, 32'h411414fa} /* (15, 22, 31) {real, imag} */,
  {32'hc03a73da, 32'h3e0d84c0} /* (15, 22, 30) {real, imag} */,
  {32'h410a500b, 32'h407b16ae} /* (15, 22, 29) {real, imag} */,
  {32'hc1025d3b, 32'h40bca1ac} /* (15, 22, 28) {real, imag} */,
  {32'hc0f0a26c, 32'h413d3b98} /* (15, 22, 27) {real, imag} */,
  {32'h4108a96e, 32'hc0fd1cd7} /* (15, 22, 26) {real, imag} */,
  {32'h409cabba, 32'hc18ba758} /* (15, 22, 25) {real, imag} */,
  {32'h3fdc6887, 32'hc13171a3} /* (15, 22, 24) {real, imag} */,
  {32'h411f1e9a, 32'h41964328} /* (15, 22, 23) {real, imag} */,
  {32'h406602cf, 32'hc15c5e9a} /* (15, 22, 22) {real, imag} */,
  {32'hc0445f7c, 32'hc1c1c0e9} /* (15, 22, 21) {real, imag} */,
  {32'hc123e690, 32'hc1941c16} /* (15, 22, 20) {real, imag} */,
  {32'h419e5785, 32'h41adbe84} /* (15, 22, 19) {real, imag} */,
  {32'h405cd0fb, 32'h41766fb0} /* (15, 22, 18) {real, imag} */,
  {32'hc1998c8e, 32'h40dd692d} /* (15, 22, 17) {real, imag} */,
  {32'hc068569a, 32'hc17c4d5c} /* (15, 22, 16) {real, imag} */,
  {32'hbfc4aabc, 32'hc0a700cb} /* (15, 22, 15) {real, imag} */,
  {32'h3f690b00, 32'hc114e6cc} /* (15, 22, 14) {real, imag} */,
  {32'h3e32f770, 32'h41cbf15e} /* (15, 22, 13) {real, imag} */,
  {32'hc1035ca8, 32'h412ebba8} /* (15, 22, 12) {real, imag} */,
  {32'hc0e9f173, 32'h419c912c} /* (15, 22, 11) {real, imag} */,
  {32'h40a338dd, 32'hbeacda70} /* (15, 22, 10) {real, imag} */,
  {32'h40ac5b3e, 32'h4031c224} /* (15, 22, 9) {real, imag} */,
  {32'hbf79b418, 32'hc0a84e32} /* (15, 22, 8) {real, imag} */,
  {32'h40aee686, 32'hc11b754f} /* (15, 22, 7) {real, imag} */,
  {32'hc1abaf52, 32'hc0cdf8bc} /* (15, 22, 6) {real, imag} */,
  {32'h404cde35, 32'hc0cb1294} /* (15, 22, 5) {real, imag} */,
  {32'hc0e7dabf, 32'h400ce26c} /* (15, 22, 4) {real, imag} */,
  {32'h3fe2c3ba, 32'h40a0a785} /* (15, 22, 3) {real, imag} */,
  {32'hbec35770, 32'h4185b75f} /* (15, 22, 2) {real, imag} */,
  {32'h40f49bf6, 32'hc1dcd624} /* (15, 22, 1) {real, imag} */,
  {32'hc0c3cad9, 32'hc1c63b8a} /* (15, 22, 0) {real, imag} */,
  {32'hc021a531, 32'h415b11f4} /* (15, 21, 31) {real, imag} */,
  {32'hc082e6dc, 32'h3f8c62d0} /* (15, 21, 30) {real, imag} */,
  {32'hc11f5f3c, 32'h41c38fd4} /* (15, 21, 29) {real, imag} */,
  {32'hc18eb5bc, 32'h3ffad968} /* (15, 21, 28) {real, imag} */,
  {32'h40b388e8, 32'hc148e47d} /* (15, 21, 27) {real, imag} */,
  {32'hc0b0b8c0, 32'h411f6d71} /* (15, 21, 26) {real, imag} */,
  {32'hc11943d2, 32'h3fa04028} /* (15, 21, 25) {real, imag} */,
  {32'hc108699d, 32'hc132c9db} /* (15, 21, 24) {real, imag} */,
  {32'h3fb7a4dc, 32'hbf21c018} /* (15, 21, 23) {real, imag} */,
  {32'h41321d83, 32'h3f8d9cb6} /* (15, 21, 22) {real, imag} */,
  {32'h3fb95fd4, 32'h410c0ef5} /* (15, 21, 21) {real, imag} */,
  {32'hc08184f5, 32'hc10cf2aa} /* (15, 21, 20) {real, imag} */,
  {32'hc10b3301, 32'hc09979b1} /* (15, 21, 19) {real, imag} */,
  {32'h405a1854, 32'h3e9d7444} /* (15, 21, 18) {real, imag} */,
  {32'h411577a3, 32'hc0a44eec} /* (15, 21, 17) {real, imag} */,
  {32'hc05a2314, 32'hc0b9968e} /* (15, 21, 16) {real, imag} */,
  {32'h3e07aae8, 32'hc16ce434} /* (15, 21, 15) {real, imag} */,
  {32'h4187fe86, 32'h40e7af1f} /* (15, 21, 14) {real, imag} */,
  {32'hc127ee3e, 32'h415a8a1c} /* (15, 21, 13) {real, imag} */,
  {32'hc06e7e66, 32'h3fbbe098} /* (15, 21, 12) {real, imag} */,
  {32'h3eb0a4a0, 32'hc180f1b8} /* (15, 21, 11) {real, imag} */,
  {32'h403cbd70, 32'h40896aba} /* (15, 21, 10) {real, imag} */,
  {32'h40159004, 32'h412c0643} /* (15, 21, 9) {real, imag} */,
  {32'h41e039f2, 32'h40f04595} /* (15, 21, 8) {real, imag} */,
  {32'hc12c963e, 32'h416786d5} /* (15, 21, 7) {real, imag} */,
  {32'h41ecd4a3, 32'h3f582c9c} /* (15, 21, 6) {real, imag} */,
  {32'hbe6ba950, 32'h4151fac0} /* (15, 21, 5) {real, imag} */,
  {32'hc1302108, 32'hc0c18964} /* (15, 21, 4) {real, imag} */,
  {32'h400d0332, 32'h406cf89c} /* (15, 21, 3) {real, imag} */,
  {32'hc0d3ba79, 32'hc14f0f14} /* (15, 21, 2) {real, imag} */,
  {32'hc1ca16f4, 32'h412e927c} /* (15, 21, 1) {real, imag} */,
  {32'hc0a5f738, 32'h411b1666} /* (15, 21, 0) {real, imag} */,
  {32'h3f886f98, 32'hc159220e} /* (15, 20, 31) {real, imag} */,
  {32'hc10618a3, 32'h40dab32b} /* (15, 20, 30) {real, imag} */,
  {32'hc11189f4, 32'h418f905a} /* (15, 20, 29) {real, imag} */,
  {32'hc0e3f197, 32'h410f6d50} /* (15, 20, 28) {real, imag} */,
  {32'h4135a953, 32'h40ce7f21} /* (15, 20, 27) {real, imag} */,
  {32'hc00d799f, 32'hc1281c38} /* (15, 20, 26) {real, imag} */,
  {32'h40ec6529, 32'hc052fa2d} /* (15, 20, 25) {real, imag} */,
  {32'h40cb38d4, 32'h410b3488} /* (15, 20, 24) {real, imag} */,
  {32'hc12a70f6, 32'hc1263754} /* (15, 20, 23) {real, imag} */,
  {32'hc127e9e8, 32'hc14ebe68} /* (15, 20, 22) {real, imag} */,
  {32'h41a01eba, 32'h411a93d3} /* (15, 20, 21) {real, imag} */,
  {32'h402d81bf, 32'hbfa657d0} /* (15, 20, 20) {real, imag} */,
  {32'hc0f314ba, 32'h3f7681d0} /* (15, 20, 19) {real, imag} */,
  {32'hc04f24b9, 32'hc12e4e73} /* (15, 20, 18) {real, imag} */,
  {32'h412e5410, 32'h403af877} /* (15, 20, 17) {real, imag} */,
  {32'h40b16a32, 32'h403d4aa8} /* (15, 20, 16) {real, imag} */,
  {32'h413449dc, 32'hbf8e7644} /* (15, 20, 15) {real, imag} */,
  {32'h4087b404, 32'hc147c534} /* (15, 20, 14) {real, imag} */,
  {32'h40e69179, 32'hc139619e} /* (15, 20, 13) {real, imag} */,
  {32'h411687ae, 32'hc035ca75} /* (15, 20, 12) {real, imag} */,
  {32'hc16318b4, 32'hc0e37422} /* (15, 20, 11) {real, imag} */,
  {32'hc056d7dc, 32'h40b4075d} /* (15, 20, 10) {real, imag} */,
  {32'hc0b9ad3b, 32'h407a429a} /* (15, 20, 9) {real, imag} */,
  {32'hc187132c, 32'hc0a6ce30} /* (15, 20, 8) {real, imag} */,
  {32'h411179e0, 32'hc0be7a02} /* (15, 20, 7) {real, imag} */,
  {32'hc0140c78, 32'h41a06f24} /* (15, 20, 6) {real, imag} */,
  {32'h40c89ffa, 32'h412db6fe} /* (15, 20, 5) {real, imag} */,
  {32'h40240939, 32'h412981e3} /* (15, 20, 4) {real, imag} */,
  {32'h412f42f4, 32'h41722d10} /* (15, 20, 3) {real, imag} */,
  {32'h3fc754a7, 32'hc106c7c3} /* (15, 20, 2) {real, imag} */,
  {32'h40ded52e, 32'hc193c004} /* (15, 20, 1) {real, imag} */,
  {32'hc08fafb2, 32'hbf7b80ac} /* (15, 20, 0) {real, imag} */,
  {32'h4144528c, 32'h40955aa4} /* (15, 19, 31) {real, imag} */,
  {32'h4031b308, 32'hc01e3a76} /* (15, 19, 30) {real, imag} */,
  {32'hc0c0a7b6, 32'hc0a4349a} /* (15, 19, 29) {real, imag} */,
  {32'hbf5318f8, 32'hc0c0d10a} /* (15, 19, 28) {real, imag} */,
  {32'hc0e43194, 32'hbe42eae0} /* (15, 19, 27) {real, imag} */,
  {32'h4165323c, 32'h410ad525} /* (15, 19, 26) {real, imag} */,
  {32'hc10b226f, 32'h4045673a} /* (15, 19, 25) {real, imag} */,
  {32'h40cd01c0, 32'h4095d680} /* (15, 19, 24) {real, imag} */,
  {32'hc125cd7f, 32'h41b8d614} /* (15, 19, 23) {real, imag} */,
  {32'hc1a356d8, 32'hbfd235ba} /* (15, 19, 22) {real, imag} */,
  {32'hc07ec47e, 32'hc18bcb15} /* (15, 19, 21) {real, imag} */,
  {32'hc12b972b, 32'h411f006b} /* (15, 19, 20) {real, imag} */,
  {32'hc058563a, 32'hc13a4796} /* (15, 19, 19) {real, imag} */,
  {32'h41524dfb, 32'hc0bb23a0} /* (15, 19, 18) {real, imag} */,
  {32'hbf7a7318, 32'hc0b57bfd} /* (15, 19, 17) {real, imag} */,
  {32'h40690f9c, 32'hc0d999f2} /* (15, 19, 16) {real, imag} */,
  {32'hc04bcfd7, 32'hc0131e2a} /* (15, 19, 15) {real, imag} */,
  {32'hc1227eaa, 32'hc09567e0} /* (15, 19, 14) {real, imag} */,
  {32'h405f08a4, 32'hc13e7b5a} /* (15, 19, 13) {real, imag} */,
  {32'h3fb465ac, 32'h416eab58} /* (15, 19, 12) {real, imag} */,
  {32'hc075d3b7, 32'h413d1e8f} /* (15, 19, 11) {real, imag} */,
  {32'hc093b956, 32'hc09a813b} /* (15, 19, 10) {real, imag} */,
  {32'h40f5b232, 32'h4128ca22} /* (15, 19, 9) {real, imag} */,
  {32'h41762936, 32'hc181c546} /* (15, 19, 8) {real, imag} */,
  {32'hc0a4ad6b, 32'h40e0c0e2} /* (15, 19, 7) {real, imag} */,
  {32'hc180c296, 32'hc0661c9a} /* (15, 19, 6) {real, imag} */,
  {32'h41259ff4, 32'h40703cdc} /* (15, 19, 5) {real, imag} */,
  {32'h410cc830, 32'hbf108a60} /* (15, 19, 4) {real, imag} */,
  {32'hc080e214, 32'h403e024a} /* (15, 19, 3) {real, imag} */,
  {32'hc0cd178f, 32'hc0589e20} /* (15, 19, 2) {real, imag} */,
  {32'h40dd3e34, 32'hc074e2be} /* (15, 19, 1) {real, imag} */,
  {32'h40c2cfda, 32'hc08ba94b} /* (15, 19, 0) {real, imag} */,
  {32'hc003656a, 32'h414faaf2} /* (15, 18, 31) {real, imag} */,
  {32'hc033ae70, 32'hbfaf0228} /* (15, 18, 30) {real, imag} */,
  {32'h3fd53af8, 32'hbed49d80} /* (15, 18, 29) {real, imag} */,
  {32'h4177e942, 32'h412a45b4} /* (15, 18, 28) {real, imag} */,
  {32'hc0db0aa2, 32'hc1b1f232} /* (15, 18, 27) {real, imag} */,
  {32'h3fda10ca, 32'hc0b0575a} /* (15, 18, 26) {real, imag} */,
  {32'h4116a9f6, 32'h41135385} /* (15, 18, 25) {real, imag} */,
  {32'h414f6ace, 32'hc095b549} /* (15, 18, 24) {real, imag} */,
  {32'hbfb3c8a8, 32'hbf6667c0} /* (15, 18, 23) {real, imag} */,
  {32'hc107b5cd, 32'h41a7f712} /* (15, 18, 22) {real, imag} */,
  {32'h4043aa1e, 32'hbf58423c} /* (15, 18, 21) {real, imag} */,
  {32'hbd00b140, 32'h404471b8} /* (15, 18, 20) {real, imag} */,
  {32'hc15dd190, 32'h40ef3170} /* (15, 18, 19) {real, imag} */,
  {32'h401d9f54, 32'h400f7c14} /* (15, 18, 18) {real, imag} */,
  {32'hc131bfd2, 32'h41412d76} /* (15, 18, 17) {real, imag} */,
  {32'hc08acefc, 32'hc09b3a0b} /* (15, 18, 16) {real, imag} */,
  {32'h413e4f8b, 32'h3ffc58d7} /* (15, 18, 15) {real, imag} */,
  {32'hc0a6253c, 32'hc040c25a} /* (15, 18, 14) {real, imag} */,
  {32'h40e86bc9, 32'h40e8fd21} /* (15, 18, 13) {real, imag} */,
  {32'hbeccd440, 32'hc04b3b60} /* (15, 18, 12) {real, imag} */,
  {32'hc0a6f1e6, 32'h41598f3c} /* (15, 18, 11) {real, imag} */,
  {32'h4031f5cf, 32'h409b42ce} /* (15, 18, 10) {real, imag} */,
  {32'h410844a0, 32'hc08f9ec6} /* (15, 18, 9) {real, imag} */,
  {32'hc0281da0, 32'hc095893a} /* (15, 18, 8) {real, imag} */,
  {32'h40f461e5, 32'hc0994466} /* (15, 18, 7) {real, imag} */,
  {32'h41a3e6bf, 32'h412e205e} /* (15, 18, 6) {real, imag} */,
  {32'h4057fe4e, 32'h40f1a578} /* (15, 18, 5) {real, imag} */,
  {32'hc12f7bae, 32'hc033095f} /* (15, 18, 4) {real, imag} */,
  {32'hc053b760, 32'hc08d280e} /* (15, 18, 3) {real, imag} */,
  {32'h40a5dd2c, 32'hc0e6d80c} /* (15, 18, 2) {real, imag} */,
  {32'hc0880169, 32'hc03690b9} /* (15, 18, 1) {real, imag} */,
  {32'h40a8a740, 32'h3f9f55e4} /* (15, 18, 0) {real, imag} */,
  {32'hc026252f, 32'h4000d59b} /* (15, 17, 31) {real, imag} */,
  {32'h41252b5a, 32'h40ad5fb1} /* (15, 17, 30) {real, imag} */,
  {32'hc131fade, 32'h4048657e} /* (15, 17, 29) {real, imag} */,
  {32'h41358e42, 32'hc1311a27} /* (15, 17, 28) {real, imag} */,
  {32'hc091406a, 32'h411507f7} /* (15, 17, 27) {real, imag} */,
  {32'hc0ba2af7, 32'hc11aced4} /* (15, 17, 26) {real, imag} */,
  {32'h3f6ef134, 32'h4175fd4e} /* (15, 17, 25) {real, imag} */,
  {32'h412ad374, 32'h4004b860} /* (15, 17, 24) {real, imag} */,
  {32'hc0d07215, 32'h40bbfc12} /* (15, 17, 23) {real, imag} */,
  {32'h4109bea6, 32'hc11060d2} /* (15, 17, 22) {real, imag} */,
  {32'h40b49f28, 32'hc141f8df} /* (15, 17, 21) {real, imag} */,
  {32'h40b2e04a, 32'hc134f209} /* (15, 17, 20) {real, imag} */,
  {32'hc11f98cf, 32'hc05f9378} /* (15, 17, 19) {real, imag} */,
  {32'h415c3b28, 32'h408131de} /* (15, 17, 18) {real, imag} */,
  {32'h3f9441ba, 32'hc10d8e0b} /* (15, 17, 17) {real, imag} */,
  {32'hc002a65a, 32'h40ac95c4} /* (15, 17, 16) {real, imag} */,
  {32'hc0f99d2d, 32'hc0dd0174} /* (15, 17, 15) {real, imag} */,
  {32'hc1174deb, 32'hc1a5ad7a} /* (15, 17, 14) {real, imag} */,
  {32'h412b3ea4, 32'hc103531c} /* (15, 17, 13) {real, imag} */,
  {32'h410fcba6, 32'hbfc46a22} /* (15, 17, 12) {real, imag} */,
  {32'hbff1460c, 32'hc098ff62} /* (15, 17, 11) {real, imag} */,
  {32'hc11d3b2b, 32'h41494846} /* (15, 17, 10) {real, imag} */,
  {32'h4037f27a, 32'hc01c7d9e} /* (15, 17, 9) {real, imag} */,
  {32'hc17d3c97, 32'h417d9056} /* (15, 17, 8) {real, imag} */,
  {32'hc10466fe, 32'hbfabe760} /* (15, 17, 7) {real, imag} */,
  {32'hc0343282, 32'hc15b0ea9} /* (15, 17, 6) {real, imag} */,
  {32'hc10d420a, 32'hc1423128} /* (15, 17, 5) {real, imag} */,
  {32'h41906119, 32'h4083ec6c} /* (15, 17, 4) {real, imag} */,
  {32'hc0a13ff2, 32'hc03e2f7a} /* (15, 17, 3) {real, imag} */,
  {32'hbf128ba8, 32'h41668018} /* (15, 17, 2) {real, imag} */,
  {32'hc05c69da, 32'h4085c3aa} /* (15, 17, 1) {real, imag} */,
  {32'h406af4fc, 32'hbfc1a4ce} /* (15, 17, 0) {real, imag} */,
  {32'hc103b388, 32'h40da5796} /* (15, 16, 31) {real, imag} */,
  {32'h40705b42, 32'h3f2e0c0e} /* (15, 16, 30) {real, imag} */,
  {32'h40f1de90, 32'h4100c47c} /* (15, 16, 29) {real, imag} */,
  {32'h3ff2695a, 32'h40eb6686} /* (15, 16, 28) {real, imag} */,
  {32'hc03e4145, 32'h4086af9e} /* (15, 16, 27) {real, imag} */,
  {32'h4011fb45, 32'h3ecdb650} /* (15, 16, 26) {real, imag} */,
  {32'h3f1c9398, 32'h3e3d38fc} /* (15, 16, 25) {real, imag} */,
  {32'hc015c203, 32'hc03f1795} /* (15, 16, 24) {real, imag} */,
  {32'hc0eaf1f2, 32'hbff72e90} /* (15, 16, 23) {real, imag} */,
  {32'h40a21f8d, 32'hbf98d14a} /* (15, 16, 22) {real, imag} */,
  {32'h41075eb5, 32'h405a4cce} /* (15, 16, 21) {real, imag} */,
  {32'hc04e479a, 32'hc0ee0dd7} /* (15, 16, 20) {real, imag} */,
  {32'h418a2272, 32'h408c061a} /* (15, 16, 19) {real, imag} */,
  {32'hc085e722, 32'h40b78ef1} /* (15, 16, 18) {real, imag} */,
  {32'h40f79cfc, 32'hc1383e36} /* (15, 16, 17) {real, imag} */,
  {32'h41781d5d, 32'h00000000} /* (15, 16, 16) {real, imag} */,
  {32'h40f79cfc, 32'h41383e36} /* (15, 16, 15) {real, imag} */,
  {32'hc085e722, 32'hc0b78ef1} /* (15, 16, 14) {real, imag} */,
  {32'h418a2272, 32'hc08c061a} /* (15, 16, 13) {real, imag} */,
  {32'hc04e479a, 32'h40ee0dd7} /* (15, 16, 12) {real, imag} */,
  {32'h41075eb5, 32'hc05a4cce} /* (15, 16, 11) {real, imag} */,
  {32'h40a21f8d, 32'h3f98d14a} /* (15, 16, 10) {real, imag} */,
  {32'hc0eaf1f2, 32'h3ff72e90} /* (15, 16, 9) {real, imag} */,
  {32'hc015c203, 32'h403f1795} /* (15, 16, 8) {real, imag} */,
  {32'h3f1c9398, 32'hbe3d38fc} /* (15, 16, 7) {real, imag} */,
  {32'h4011fb45, 32'hbecdb650} /* (15, 16, 6) {real, imag} */,
  {32'hc03e4145, 32'hc086af9e} /* (15, 16, 5) {real, imag} */,
  {32'h3ff2695a, 32'hc0eb6686} /* (15, 16, 4) {real, imag} */,
  {32'h40f1de90, 32'hc100c47c} /* (15, 16, 3) {real, imag} */,
  {32'h40705b42, 32'hbf2e0c0e} /* (15, 16, 2) {real, imag} */,
  {32'hc103b388, 32'hc0da5796} /* (15, 16, 1) {real, imag} */,
  {32'h402f705b, 32'h00000000} /* (15, 16, 0) {real, imag} */,
  {32'hc05c69da, 32'hc085c3aa} /* (15, 15, 31) {real, imag} */,
  {32'hbf128ba8, 32'hc1668018} /* (15, 15, 30) {real, imag} */,
  {32'hc0a13ff2, 32'h403e2f7a} /* (15, 15, 29) {real, imag} */,
  {32'h41906119, 32'hc083ec6c} /* (15, 15, 28) {real, imag} */,
  {32'hc10d420a, 32'h41423128} /* (15, 15, 27) {real, imag} */,
  {32'hc0343282, 32'h415b0ea9} /* (15, 15, 26) {real, imag} */,
  {32'hc10466fe, 32'h3fabe760} /* (15, 15, 25) {real, imag} */,
  {32'hc17d3c97, 32'hc17d9056} /* (15, 15, 24) {real, imag} */,
  {32'h4037f27a, 32'h401c7d9e} /* (15, 15, 23) {real, imag} */,
  {32'hc11d3b2b, 32'hc1494846} /* (15, 15, 22) {real, imag} */,
  {32'hbff1460c, 32'h4098ff62} /* (15, 15, 21) {real, imag} */,
  {32'h410fcba6, 32'h3fc46a22} /* (15, 15, 20) {real, imag} */,
  {32'h412b3ea4, 32'h4103531c} /* (15, 15, 19) {real, imag} */,
  {32'hc1174deb, 32'h41a5ad7a} /* (15, 15, 18) {real, imag} */,
  {32'hc0f99d2d, 32'h40dd0174} /* (15, 15, 17) {real, imag} */,
  {32'hc002a65a, 32'hc0ac95c4} /* (15, 15, 16) {real, imag} */,
  {32'h3f9441ba, 32'h410d8e0b} /* (15, 15, 15) {real, imag} */,
  {32'h415c3b28, 32'hc08131de} /* (15, 15, 14) {real, imag} */,
  {32'hc11f98cf, 32'h405f9378} /* (15, 15, 13) {real, imag} */,
  {32'h40b2e04a, 32'h4134f209} /* (15, 15, 12) {real, imag} */,
  {32'h40b49f28, 32'h4141f8df} /* (15, 15, 11) {real, imag} */,
  {32'h4109bea6, 32'h411060d2} /* (15, 15, 10) {real, imag} */,
  {32'hc0d07215, 32'hc0bbfc12} /* (15, 15, 9) {real, imag} */,
  {32'h412ad374, 32'hc004b860} /* (15, 15, 8) {real, imag} */,
  {32'h3f6ef134, 32'hc175fd4e} /* (15, 15, 7) {real, imag} */,
  {32'hc0ba2af7, 32'h411aced4} /* (15, 15, 6) {real, imag} */,
  {32'hc091406a, 32'hc11507f7} /* (15, 15, 5) {real, imag} */,
  {32'h41358e42, 32'h41311a27} /* (15, 15, 4) {real, imag} */,
  {32'hc131fade, 32'hc048657e} /* (15, 15, 3) {real, imag} */,
  {32'h41252b5a, 32'hc0ad5fb1} /* (15, 15, 2) {real, imag} */,
  {32'hc026252f, 32'hc000d59b} /* (15, 15, 1) {real, imag} */,
  {32'h406af4fc, 32'h3fc1a4ce} /* (15, 15, 0) {real, imag} */,
  {32'hc0880169, 32'h403690b9} /* (15, 14, 31) {real, imag} */,
  {32'h40a5dd2c, 32'h40e6d80c} /* (15, 14, 30) {real, imag} */,
  {32'hc053b760, 32'h408d280e} /* (15, 14, 29) {real, imag} */,
  {32'hc12f7bae, 32'h4033095f} /* (15, 14, 28) {real, imag} */,
  {32'h4057fe4e, 32'hc0f1a578} /* (15, 14, 27) {real, imag} */,
  {32'h41a3e6bf, 32'hc12e205e} /* (15, 14, 26) {real, imag} */,
  {32'h40f461e5, 32'h40994466} /* (15, 14, 25) {real, imag} */,
  {32'hc0281da0, 32'h4095893a} /* (15, 14, 24) {real, imag} */,
  {32'h410844a0, 32'h408f9ec6} /* (15, 14, 23) {real, imag} */,
  {32'h4031f5cf, 32'hc09b42ce} /* (15, 14, 22) {real, imag} */,
  {32'hc0a6f1e6, 32'hc1598f3c} /* (15, 14, 21) {real, imag} */,
  {32'hbeccd440, 32'h404b3b60} /* (15, 14, 20) {real, imag} */,
  {32'h40e86bc9, 32'hc0e8fd21} /* (15, 14, 19) {real, imag} */,
  {32'hc0a6253c, 32'h4040c25a} /* (15, 14, 18) {real, imag} */,
  {32'h413e4f8b, 32'hbffc58d7} /* (15, 14, 17) {real, imag} */,
  {32'hc08acefc, 32'h409b3a0b} /* (15, 14, 16) {real, imag} */,
  {32'hc131bfd2, 32'hc1412d76} /* (15, 14, 15) {real, imag} */,
  {32'h401d9f54, 32'hc00f7c14} /* (15, 14, 14) {real, imag} */,
  {32'hc15dd190, 32'hc0ef3170} /* (15, 14, 13) {real, imag} */,
  {32'hbd00b140, 32'hc04471b8} /* (15, 14, 12) {real, imag} */,
  {32'h4043aa1e, 32'h3f58423c} /* (15, 14, 11) {real, imag} */,
  {32'hc107b5cd, 32'hc1a7f712} /* (15, 14, 10) {real, imag} */,
  {32'hbfb3c8a8, 32'h3f6667c0} /* (15, 14, 9) {real, imag} */,
  {32'h414f6ace, 32'h4095b549} /* (15, 14, 8) {real, imag} */,
  {32'h4116a9f6, 32'hc1135385} /* (15, 14, 7) {real, imag} */,
  {32'h3fda10ca, 32'h40b0575a} /* (15, 14, 6) {real, imag} */,
  {32'hc0db0aa2, 32'h41b1f232} /* (15, 14, 5) {real, imag} */,
  {32'h4177e942, 32'hc12a45b4} /* (15, 14, 4) {real, imag} */,
  {32'h3fd53af8, 32'h3ed49d80} /* (15, 14, 3) {real, imag} */,
  {32'hc033ae70, 32'h3faf0228} /* (15, 14, 2) {real, imag} */,
  {32'hc003656a, 32'hc14faaf2} /* (15, 14, 1) {real, imag} */,
  {32'h40a8a740, 32'hbf9f55e4} /* (15, 14, 0) {real, imag} */,
  {32'h40dd3e34, 32'h4074e2be} /* (15, 13, 31) {real, imag} */,
  {32'hc0cd178f, 32'h40589e20} /* (15, 13, 30) {real, imag} */,
  {32'hc080e214, 32'hc03e024a} /* (15, 13, 29) {real, imag} */,
  {32'h410cc830, 32'h3f108a60} /* (15, 13, 28) {real, imag} */,
  {32'h41259ff4, 32'hc0703cdc} /* (15, 13, 27) {real, imag} */,
  {32'hc180c296, 32'h40661c9a} /* (15, 13, 26) {real, imag} */,
  {32'hc0a4ad6b, 32'hc0e0c0e2} /* (15, 13, 25) {real, imag} */,
  {32'h41762936, 32'h4181c546} /* (15, 13, 24) {real, imag} */,
  {32'h40f5b232, 32'hc128ca22} /* (15, 13, 23) {real, imag} */,
  {32'hc093b956, 32'h409a813b} /* (15, 13, 22) {real, imag} */,
  {32'hc075d3b7, 32'hc13d1e8f} /* (15, 13, 21) {real, imag} */,
  {32'h3fb465ac, 32'hc16eab58} /* (15, 13, 20) {real, imag} */,
  {32'h405f08a4, 32'h413e7b5a} /* (15, 13, 19) {real, imag} */,
  {32'hc1227eaa, 32'h409567e0} /* (15, 13, 18) {real, imag} */,
  {32'hc04bcfd7, 32'h40131e2a} /* (15, 13, 17) {real, imag} */,
  {32'h40690f9c, 32'h40d999f2} /* (15, 13, 16) {real, imag} */,
  {32'hbf7a7318, 32'h40b57bfd} /* (15, 13, 15) {real, imag} */,
  {32'h41524dfb, 32'h40bb23a0} /* (15, 13, 14) {real, imag} */,
  {32'hc058563a, 32'h413a4796} /* (15, 13, 13) {real, imag} */,
  {32'hc12b972b, 32'hc11f006b} /* (15, 13, 12) {real, imag} */,
  {32'hc07ec47e, 32'h418bcb15} /* (15, 13, 11) {real, imag} */,
  {32'hc1a356d8, 32'h3fd235ba} /* (15, 13, 10) {real, imag} */,
  {32'hc125cd7f, 32'hc1b8d614} /* (15, 13, 9) {real, imag} */,
  {32'h40cd01c0, 32'hc095d680} /* (15, 13, 8) {real, imag} */,
  {32'hc10b226f, 32'hc045673a} /* (15, 13, 7) {real, imag} */,
  {32'h4165323c, 32'hc10ad525} /* (15, 13, 6) {real, imag} */,
  {32'hc0e43194, 32'h3e42eae0} /* (15, 13, 5) {real, imag} */,
  {32'hbf5318f8, 32'h40c0d10a} /* (15, 13, 4) {real, imag} */,
  {32'hc0c0a7b6, 32'h40a4349a} /* (15, 13, 3) {real, imag} */,
  {32'h4031b308, 32'h401e3a76} /* (15, 13, 2) {real, imag} */,
  {32'h4144528c, 32'hc0955aa4} /* (15, 13, 1) {real, imag} */,
  {32'h40c2cfda, 32'h408ba94b} /* (15, 13, 0) {real, imag} */,
  {32'h40ded52e, 32'h4193c004} /* (15, 12, 31) {real, imag} */,
  {32'h3fc754a7, 32'h4106c7c3} /* (15, 12, 30) {real, imag} */,
  {32'h412f42f4, 32'hc1722d10} /* (15, 12, 29) {real, imag} */,
  {32'h40240939, 32'hc12981e3} /* (15, 12, 28) {real, imag} */,
  {32'h40c89ffa, 32'hc12db6fe} /* (15, 12, 27) {real, imag} */,
  {32'hc0140c78, 32'hc1a06f24} /* (15, 12, 26) {real, imag} */,
  {32'h411179e0, 32'h40be7a02} /* (15, 12, 25) {real, imag} */,
  {32'hc187132c, 32'h40a6ce30} /* (15, 12, 24) {real, imag} */,
  {32'hc0b9ad3b, 32'hc07a429a} /* (15, 12, 23) {real, imag} */,
  {32'hc056d7dc, 32'hc0b4075d} /* (15, 12, 22) {real, imag} */,
  {32'hc16318b4, 32'h40e37422} /* (15, 12, 21) {real, imag} */,
  {32'h411687ae, 32'h4035ca75} /* (15, 12, 20) {real, imag} */,
  {32'h40e69179, 32'h4139619e} /* (15, 12, 19) {real, imag} */,
  {32'h4087b404, 32'h4147c534} /* (15, 12, 18) {real, imag} */,
  {32'h413449dc, 32'h3f8e7644} /* (15, 12, 17) {real, imag} */,
  {32'h40b16a32, 32'hc03d4aa8} /* (15, 12, 16) {real, imag} */,
  {32'h412e5410, 32'hc03af877} /* (15, 12, 15) {real, imag} */,
  {32'hc04f24b9, 32'h412e4e73} /* (15, 12, 14) {real, imag} */,
  {32'hc0f314ba, 32'hbf7681d0} /* (15, 12, 13) {real, imag} */,
  {32'h402d81bf, 32'h3fa657d0} /* (15, 12, 12) {real, imag} */,
  {32'h41a01eba, 32'hc11a93d3} /* (15, 12, 11) {real, imag} */,
  {32'hc127e9e8, 32'h414ebe68} /* (15, 12, 10) {real, imag} */,
  {32'hc12a70f6, 32'h41263754} /* (15, 12, 9) {real, imag} */,
  {32'h40cb38d4, 32'hc10b3488} /* (15, 12, 8) {real, imag} */,
  {32'h40ec6529, 32'h4052fa2d} /* (15, 12, 7) {real, imag} */,
  {32'hc00d799f, 32'h41281c38} /* (15, 12, 6) {real, imag} */,
  {32'h4135a953, 32'hc0ce7f21} /* (15, 12, 5) {real, imag} */,
  {32'hc0e3f197, 32'hc10f6d50} /* (15, 12, 4) {real, imag} */,
  {32'hc11189f4, 32'hc18f905a} /* (15, 12, 3) {real, imag} */,
  {32'hc10618a3, 32'hc0dab32b} /* (15, 12, 2) {real, imag} */,
  {32'h3f886f98, 32'h4159220e} /* (15, 12, 1) {real, imag} */,
  {32'hc08fafb2, 32'h3f7b80ac} /* (15, 12, 0) {real, imag} */,
  {32'hc1ca16f4, 32'hc12e927c} /* (15, 11, 31) {real, imag} */,
  {32'hc0d3ba79, 32'h414f0f14} /* (15, 11, 30) {real, imag} */,
  {32'h400d0332, 32'hc06cf89c} /* (15, 11, 29) {real, imag} */,
  {32'hc1302108, 32'h40c18964} /* (15, 11, 28) {real, imag} */,
  {32'hbe6ba950, 32'hc151fac0} /* (15, 11, 27) {real, imag} */,
  {32'h41ecd4a3, 32'hbf582c9c} /* (15, 11, 26) {real, imag} */,
  {32'hc12c963e, 32'hc16786d5} /* (15, 11, 25) {real, imag} */,
  {32'h41e039f2, 32'hc0f04595} /* (15, 11, 24) {real, imag} */,
  {32'h40159004, 32'hc12c0643} /* (15, 11, 23) {real, imag} */,
  {32'h403cbd70, 32'hc0896aba} /* (15, 11, 22) {real, imag} */,
  {32'h3eb0a4a0, 32'h4180f1b8} /* (15, 11, 21) {real, imag} */,
  {32'hc06e7e66, 32'hbfbbe098} /* (15, 11, 20) {real, imag} */,
  {32'hc127ee3e, 32'hc15a8a1c} /* (15, 11, 19) {real, imag} */,
  {32'h4187fe86, 32'hc0e7af1f} /* (15, 11, 18) {real, imag} */,
  {32'h3e07aae8, 32'h416ce434} /* (15, 11, 17) {real, imag} */,
  {32'hc05a2314, 32'h40b9968e} /* (15, 11, 16) {real, imag} */,
  {32'h411577a3, 32'h40a44eec} /* (15, 11, 15) {real, imag} */,
  {32'h405a1854, 32'hbe9d7444} /* (15, 11, 14) {real, imag} */,
  {32'hc10b3301, 32'h409979b1} /* (15, 11, 13) {real, imag} */,
  {32'hc08184f5, 32'h410cf2aa} /* (15, 11, 12) {real, imag} */,
  {32'h3fb95fd4, 32'hc10c0ef5} /* (15, 11, 11) {real, imag} */,
  {32'h41321d83, 32'hbf8d9cb6} /* (15, 11, 10) {real, imag} */,
  {32'h3fb7a4dc, 32'h3f21c018} /* (15, 11, 9) {real, imag} */,
  {32'hc108699d, 32'h4132c9db} /* (15, 11, 8) {real, imag} */,
  {32'hc11943d2, 32'hbfa04028} /* (15, 11, 7) {real, imag} */,
  {32'hc0b0b8c0, 32'hc11f6d71} /* (15, 11, 6) {real, imag} */,
  {32'h40b388e8, 32'h4148e47d} /* (15, 11, 5) {real, imag} */,
  {32'hc18eb5bc, 32'hbffad968} /* (15, 11, 4) {real, imag} */,
  {32'hc11f5f3c, 32'hc1c38fd4} /* (15, 11, 3) {real, imag} */,
  {32'hc082e6dc, 32'hbf8c62d0} /* (15, 11, 2) {real, imag} */,
  {32'hc021a531, 32'hc15b11f4} /* (15, 11, 1) {real, imag} */,
  {32'hc0a5f738, 32'hc11b1666} /* (15, 11, 0) {real, imag} */,
  {32'h40f49bf6, 32'h41dcd624} /* (15, 10, 31) {real, imag} */,
  {32'hbec35770, 32'hc185b75f} /* (15, 10, 30) {real, imag} */,
  {32'h3fe2c3ba, 32'hc0a0a785} /* (15, 10, 29) {real, imag} */,
  {32'hc0e7dabf, 32'hc00ce26c} /* (15, 10, 28) {real, imag} */,
  {32'h404cde35, 32'h40cb1294} /* (15, 10, 27) {real, imag} */,
  {32'hc1abaf52, 32'h40cdf8bc} /* (15, 10, 26) {real, imag} */,
  {32'h40aee686, 32'h411b754f} /* (15, 10, 25) {real, imag} */,
  {32'hbf79b418, 32'h40a84e32} /* (15, 10, 24) {real, imag} */,
  {32'h40ac5b3e, 32'hc031c224} /* (15, 10, 23) {real, imag} */,
  {32'h40a338dd, 32'h3eacda70} /* (15, 10, 22) {real, imag} */,
  {32'hc0e9f173, 32'hc19c912c} /* (15, 10, 21) {real, imag} */,
  {32'hc1035ca8, 32'hc12ebba8} /* (15, 10, 20) {real, imag} */,
  {32'h3e32f770, 32'hc1cbf15e} /* (15, 10, 19) {real, imag} */,
  {32'h3f690b00, 32'h4114e6cc} /* (15, 10, 18) {real, imag} */,
  {32'hbfc4aabc, 32'h40a700cb} /* (15, 10, 17) {real, imag} */,
  {32'hc068569a, 32'h417c4d5c} /* (15, 10, 16) {real, imag} */,
  {32'hc1998c8e, 32'hc0dd692d} /* (15, 10, 15) {real, imag} */,
  {32'h405cd0fb, 32'hc1766fb0} /* (15, 10, 14) {real, imag} */,
  {32'h419e5785, 32'hc1adbe84} /* (15, 10, 13) {real, imag} */,
  {32'hc123e690, 32'h41941c16} /* (15, 10, 12) {real, imag} */,
  {32'hc0445f7c, 32'h41c1c0e9} /* (15, 10, 11) {real, imag} */,
  {32'h406602cf, 32'h415c5e9a} /* (15, 10, 10) {real, imag} */,
  {32'h411f1e9a, 32'hc1964328} /* (15, 10, 9) {real, imag} */,
  {32'h3fdc6887, 32'h413171a3} /* (15, 10, 8) {real, imag} */,
  {32'h409cabba, 32'h418ba758} /* (15, 10, 7) {real, imag} */,
  {32'h4108a96e, 32'h40fd1cd7} /* (15, 10, 6) {real, imag} */,
  {32'hc0f0a26c, 32'hc13d3b98} /* (15, 10, 5) {real, imag} */,
  {32'hc1025d3b, 32'hc0bca1ac} /* (15, 10, 4) {real, imag} */,
  {32'h410a500b, 32'hc07b16ae} /* (15, 10, 3) {real, imag} */,
  {32'hc03a73da, 32'hbe0d84c0} /* (15, 10, 2) {real, imag} */,
  {32'h412bde19, 32'hc11414fa} /* (15, 10, 1) {real, imag} */,
  {32'hc0c3cad9, 32'h41c63b8a} /* (15, 10, 0) {real, imag} */,
  {32'hc1cbdbc6, 32'hbfe84b0c} /* (15, 9, 31) {real, imag} */,
  {32'h3f1ffb38, 32'hc0405d1c} /* (15, 9, 30) {real, imag} */,
  {32'h4146c516, 32'hbf44f5d0} /* (15, 9, 29) {real, imag} */,
  {32'hc06b7816, 32'h41d003c5} /* (15, 9, 28) {real, imag} */,
  {32'h410848ce, 32'hc12d4a82} /* (15, 9, 27) {real, imag} */,
  {32'h412614f0, 32'h401b0288} /* (15, 9, 26) {real, imag} */,
  {32'h412a85e2, 32'hc1158ec2} /* (15, 9, 25) {real, imag} */,
  {32'h40660bdc, 32'hc1697ce5} /* (15, 9, 24) {real, imag} */,
  {32'h3eb7cfc8, 32'h3fadb888} /* (15, 9, 23) {real, imag} */,
  {32'hc103ef04, 32'h410f584f} /* (15, 9, 22) {real, imag} */,
  {32'h41849ac8, 32'h41220442} /* (15, 9, 21) {real, imag} */,
  {32'h409d0e71, 32'h3f8ff480} /* (15, 9, 20) {real, imag} */,
  {32'h412232a6, 32'h4057059e} /* (15, 9, 19) {real, imag} */,
  {32'hc1ad5a77, 32'hc10be229} /* (15, 9, 18) {real, imag} */,
  {32'hc0c8a230, 32'hc11b818a} /* (15, 9, 17) {real, imag} */,
  {32'h3f80c388, 32'h40b1c279} /* (15, 9, 16) {real, imag} */,
  {32'h4031e910, 32'hc118f60c} /* (15, 9, 15) {real, imag} */,
  {32'hc147de34, 32'h3fe16fb8} /* (15, 9, 14) {real, imag} */,
  {32'h418da9e6, 32'h4121560c} /* (15, 9, 13) {real, imag} */,
  {32'h3d8b9040, 32'hc087c416} /* (15, 9, 12) {real, imag} */,
  {32'hc0b6edc6, 32'hc0ce0796} /* (15, 9, 11) {real, imag} */,
  {32'hc13feab6, 32'hc17933fa} /* (15, 9, 10) {real, imag} */,
  {32'h41f3e339, 32'h40f880e8} /* (15, 9, 9) {real, imag} */,
  {32'hc0410ae4, 32'h3eb3cff0} /* (15, 9, 8) {real, imag} */,
  {32'hc18507d4, 32'h412c7ce9} /* (15, 9, 7) {real, imag} */,
  {32'h4122def8, 32'hbf65c474} /* (15, 9, 6) {real, imag} */,
  {32'hc13dd375, 32'hbfaf994c} /* (15, 9, 5) {real, imag} */,
  {32'h40833f1e, 32'h4097cd32} /* (15, 9, 4) {real, imag} */,
  {32'h4090f282, 32'h3ffb17ec} /* (15, 9, 3) {real, imag} */,
  {32'h3fe3c11d, 32'hc11d3a9a} /* (15, 9, 2) {real, imag} */,
  {32'h408861eb, 32'h417a34c4} /* (15, 9, 1) {real, imag} */,
  {32'h413cd3ad, 32'h4066b44f} /* (15, 9, 0) {real, imag} */,
  {32'hc2429f92, 32'hc1e6403c} /* (15, 8, 31) {real, imag} */,
  {32'h41064daf, 32'hc0db79ee} /* (15, 8, 30) {real, imag} */,
  {32'h4126f42d, 32'h4016e0b0} /* (15, 8, 29) {real, imag} */,
  {32'h4114b431, 32'h3eea31c8} /* (15, 8, 28) {real, imag} */,
  {32'h40be9d01, 32'hbe9cc868} /* (15, 8, 27) {real, imag} */,
  {32'h415ab47d, 32'h417b1ad0} /* (15, 8, 26) {real, imag} */,
  {32'hc1288eda, 32'hc1943f6a} /* (15, 8, 25) {real, imag} */,
  {32'h412266ed, 32'hc1a9dcbd} /* (15, 8, 24) {real, imag} */,
  {32'h3dd68e60, 32'h405a2ef9} /* (15, 8, 23) {real, imag} */,
  {32'h4199e225, 32'h4005f594} /* (15, 8, 22) {real, imag} */,
  {32'h412f2227, 32'h4089b929} /* (15, 8, 21) {real, imag} */,
  {32'h3fe9cbd0, 32'h41ceaec4} /* (15, 8, 20) {real, imag} */,
  {32'hc13127b6, 32'hc10deb73} /* (15, 8, 19) {real, imag} */,
  {32'hbffa0596, 32'h40f80001} /* (15, 8, 18) {real, imag} */,
  {32'h3de01b00, 32'hc18f4e94} /* (15, 8, 17) {real, imag} */,
  {32'h40725459, 32'hc032c0e6} /* (15, 8, 16) {real, imag} */,
  {32'hbf732558, 32'h3f50199c} /* (15, 8, 15) {real, imag} */,
  {32'h40c5ee66, 32'hbec625b0} /* (15, 8, 14) {real, imag} */,
  {32'hc0a8b95b, 32'h40aac47c} /* (15, 8, 13) {real, imag} */,
  {32'hc1db646c, 32'h415cfacc} /* (15, 8, 12) {real, imag} */,
  {32'h410946a8, 32'h3ffdf039} /* (15, 8, 11) {real, imag} */,
  {32'h418c8918, 32'h408277b6} /* (15, 8, 10) {real, imag} */,
  {32'hc0c0f554, 32'h41b17861} /* (15, 8, 9) {real, imag} */,
  {32'h41b98e6d, 32'hc120452c} /* (15, 8, 8) {real, imag} */,
  {32'hc0bbeffe, 32'hc0d624d1} /* (15, 8, 7) {real, imag} */,
  {32'hc053ecc0, 32'hc1ad07a5} /* (15, 8, 6) {real, imag} */,
  {32'hc161fe98, 32'h3ea0e3d0} /* (15, 8, 5) {real, imag} */,
  {32'hc19eede4, 32'hc0d5b193} /* (15, 8, 4) {real, imag} */,
  {32'hc123cc91, 32'h40c32fc6} /* (15, 8, 3) {real, imag} */,
  {32'h40d942dc, 32'h412cadc0} /* (15, 8, 2) {real, imag} */,
  {32'hc12135f8, 32'h3fa03034} /* (15, 8, 1) {real, imag} */,
  {32'hc15e19bc, 32'h4178a85e} /* (15, 8, 0) {real, imag} */,
  {32'h408f8f94, 32'h41d30667} /* (15, 7, 31) {real, imag} */,
  {32'hc0a4f2e0, 32'hc1d2b5d8} /* (15, 7, 30) {real, imag} */,
  {32'hc1215c1a, 32'hc0020f95} /* (15, 7, 29) {real, imag} */,
  {32'hc1574ada, 32'hc139a3a9} /* (15, 7, 28) {real, imag} */,
  {32'hbfed4d60, 32'hc0883c28} /* (15, 7, 27) {real, imag} */,
  {32'hc0d12498, 32'hbff655cf} /* (15, 7, 26) {real, imag} */,
  {32'hbffdae48, 32'hc119eca1} /* (15, 7, 25) {real, imag} */,
  {32'hc106301e, 32'h3fa71cc0} /* (15, 7, 24) {real, imag} */,
  {32'hc11a118a, 32'h3fe632f0} /* (15, 7, 23) {real, imag} */,
  {32'h3f86d1ec, 32'h4006a0d2} /* (15, 7, 22) {real, imag} */,
  {32'hc00b7bd2, 32'h4103f200} /* (15, 7, 21) {real, imag} */,
  {32'h3ef7a16c, 32'hc0fd5cd6} /* (15, 7, 20) {real, imag} */,
  {32'h3f856e3c, 32'hc12966a8} /* (15, 7, 19) {real, imag} */,
  {32'hc09891b0, 32'hc00ecda0} /* (15, 7, 18) {real, imag} */,
  {32'h4053c8d6, 32'hc06792b3} /* (15, 7, 17) {real, imag} */,
  {32'h40b38f60, 32'hc015410c} /* (15, 7, 16) {real, imag} */,
  {32'hc1a4a7f4, 32'hc0fd1a4a} /* (15, 7, 15) {real, imag} */,
  {32'h40b721ee, 32'h40e19244} /* (15, 7, 14) {real, imag} */,
  {32'hc05f3f45, 32'hc0a71ed0} /* (15, 7, 13) {real, imag} */,
  {32'h3fdb1f98, 32'h405a05a8} /* (15, 7, 12) {real, imag} */,
  {32'h40dcd702, 32'h40eb1839} /* (15, 7, 11) {real, imag} */,
  {32'hc0d579bb, 32'h4122093c} /* (15, 7, 10) {real, imag} */,
  {32'hc1665b4a, 32'h409e1e08} /* (15, 7, 9) {real, imag} */,
  {32'h404734d8, 32'hc1c3afac} /* (15, 7, 8) {real, imag} */,
  {32'h416723e0, 32'h4172931c} /* (15, 7, 7) {real, imag} */,
  {32'hc1b76059, 32'h400575c0} /* (15, 7, 6) {real, imag} */,
  {32'hc10381b0, 32'h3f836770} /* (15, 7, 5) {real, imag} */,
  {32'h40aa9560, 32'hc00d7d96} /* (15, 7, 4) {real, imag} */,
  {32'hc0b8fe40, 32'hc19afd12} /* (15, 7, 3) {real, imag} */,
  {32'h40065af0, 32'hc0e4b8f3} /* (15, 7, 2) {real, imag} */,
  {32'hc173f4ce, 32'h423bc676} /* (15, 7, 1) {real, imag} */,
  {32'hc11173b2, 32'hc0b3d8de} /* (15, 7, 0) {real, imag} */,
  {32'hc02e55e0, 32'h40800aec} /* (15, 6, 31) {real, imag} */,
  {32'hc10c4c8c, 32'h402aa0e2} /* (15, 6, 30) {real, imag} */,
  {32'hc094832c, 32'h3d9fe200} /* (15, 6, 29) {real, imag} */,
  {32'hc0997bfb, 32'h407e0b64} /* (15, 6, 28) {real, imag} */,
  {32'hc185bbba, 32'h4017e1ae} /* (15, 6, 27) {real, imag} */,
  {32'hc112b338, 32'hbfe4f512} /* (15, 6, 26) {real, imag} */,
  {32'hc1979a1a, 32'h40b2b79d} /* (15, 6, 25) {real, imag} */,
  {32'h3faab5d8, 32'hc152285a} /* (15, 6, 24) {real, imag} */,
  {32'h413916e0, 32'hc0b9addc} /* (15, 6, 23) {real, imag} */,
  {32'h406b982c, 32'h40bf6acd} /* (15, 6, 22) {real, imag} */,
  {32'hc085623b, 32'h4116834e} /* (15, 6, 21) {real, imag} */,
  {32'hc1ad6aca, 32'h406cd050} /* (15, 6, 20) {real, imag} */,
  {32'hc11133e3, 32'hc0a15578} /* (15, 6, 19) {real, imag} */,
  {32'h412a8d6e, 32'hc089ad78} /* (15, 6, 18) {real, imag} */,
  {32'h40afda9a, 32'hc0bc33da} /* (15, 6, 17) {real, imag} */,
  {32'h402fa00a, 32'h41742f66} /* (15, 6, 16) {real, imag} */,
  {32'h4100214b, 32'hc09a8350} /* (15, 6, 15) {real, imag} */,
  {32'h40190b4e, 32'h41386f18} /* (15, 6, 14) {real, imag} */,
  {32'h3d3a1ce0, 32'h3fd59a68} /* (15, 6, 13) {real, imag} */,
  {32'h4022c340, 32'h40efb8be} /* (15, 6, 12) {real, imag} */,
  {32'h40b2ad73, 32'h40b177f8} /* (15, 6, 11) {real, imag} */,
  {32'hc10c38f6, 32'h4196ef9e} /* (15, 6, 10) {real, imag} */,
  {32'h411a7126, 32'h41021f3a} /* (15, 6, 9) {real, imag} */,
  {32'hc1813df1, 32'hc11cedeb} /* (15, 6, 8) {real, imag} */,
  {32'hc098c8d2, 32'h3f544c94} /* (15, 6, 7) {real, imag} */,
  {32'hc0be2efe, 32'h4117208e} /* (15, 6, 6) {real, imag} */,
  {32'h41472324, 32'hc100d02c} /* (15, 6, 5) {real, imag} */,
  {32'hc1432d5e, 32'h408defba} /* (15, 6, 4) {real, imag} */,
  {32'h41564445, 32'h40a7c6c5} /* (15, 6, 3) {real, imag} */,
  {32'h41a767b2, 32'h41834c19} /* (15, 6, 2) {real, imag} */,
  {32'h41a77bff, 32'h41d5ce2e} /* (15, 6, 1) {real, imag} */,
  {32'hc1c276ba, 32'hc0ff1662} /* (15, 6, 0) {real, imag} */,
  {32'hc211640a, 32'h423dcea6} /* (15, 5, 31) {real, imag} */,
  {32'h4077cc00, 32'hc15b8776} /* (15, 5, 30) {real, imag} */,
  {32'h3fbfdc1c, 32'h41a0c403} /* (15, 5, 29) {real, imag} */,
  {32'h404d1a90, 32'h3f779cb8} /* (15, 5, 28) {real, imag} */,
  {32'h41465102, 32'h41e2d8af} /* (15, 5, 27) {real, imag} */,
  {32'hbf94ffb4, 32'hc1286480} /* (15, 5, 26) {real, imag} */,
  {32'hc2248c64, 32'h40c2bd64} /* (15, 5, 25) {real, imag} */,
  {32'hc146b8e2, 32'hbfe5e3b4} /* (15, 5, 24) {real, imag} */,
  {32'hc121cadc, 32'h404791d8} /* (15, 5, 23) {real, imag} */,
  {32'h40b86be6, 32'hc16881ec} /* (15, 5, 22) {real, imag} */,
  {32'h3ea58570, 32'h3fbf9576} /* (15, 5, 21) {real, imag} */,
  {32'hc030c4dc, 32'hc0b5ca5f} /* (15, 5, 20) {real, imag} */,
  {32'hc005f2a7, 32'hc004c9bf} /* (15, 5, 19) {real, imag} */,
  {32'h40c56958, 32'hbf8869b4} /* (15, 5, 18) {real, imag} */,
  {32'hc0d9b8a8, 32'hc169f82a} /* (15, 5, 17) {real, imag} */,
  {32'hc0feeb64, 32'hc00219f4} /* (15, 5, 16) {real, imag} */,
  {32'h417cbc4c, 32'h40021428} /* (15, 5, 15) {real, imag} */,
  {32'hc12a67df, 32'hc0a3a5d1} /* (15, 5, 14) {real, imag} */,
  {32'hc11c9fae, 32'hbfa3f114} /* (15, 5, 13) {real, imag} */,
  {32'hc08d3b8b, 32'hc089d9dc} /* (15, 5, 12) {real, imag} */,
  {32'hc013142e, 32'h40ee9bb6} /* (15, 5, 11) {real, imag} */,
  {32'hc09a2fca, 32'hc149022a} /* (15, 5, 10) {real, imag} */,
  {32'hc125f42a, 32'hc1596398} /* (15, 5, 9) {real, imag} */,
  {32'h40a37cce, 32'h41ca2ad7} /* (15, 5, 8) {real, imag} */,
  {32'hc08fb8ea, 32'hc020ec10} /* (15, 5, 7) {real, imag} */,
  {32'h40fec830, 32'hbf707600} /* (15, 5, 6) {real, imag} */,
  {32'h4114528c, 32'h40f739e2} /* (15, 5, 5) {real, imag} */,
  {32'h41a29328, 32'hc131d82c} /* (15, 5, 4) {real, imag} */,
  {32'h419041b0, 32'hc195d2e4} /* (15, 5, 3) {real, imag} */,
  {32'h411b8e68, 32'h419f5f70} /* (15, 5, 2) {real, imag} */,
  {32'hc2554f7e, 32'hc1374c58} /* (15, 5, 1) {real, imag} */,
  {32'hc24179e4, 32'hc038dc30} /* (15, 5, 0) {real, imag} */,
  {32'h421d9fbc, 32'h3fb72c80} /* (15, 4, 31) {real, imag} */,
  {32'hc19e6d60, 32'hc196f5ba} /* (15, 4, 30) {real, imag} */,
  {32'h403725e0, 32'hc19e83b8} /* (15, 4, 29) {real, imag} */,
  {32'h42006e5c, 32'h4194af2e} /* (15, 4, 28) {real, imag} */,
  {32'hc1a20fc4, 32'h40a29844} /* (15, 4, 27) {real, imag} */,
  {32'hc1110838, 32'h418d1f41} /* (15, 4, 26) {real, imag} */,
  {32'hc10e1cb0, 32'h4214df92} /* (15, 4, 25) {real, imag} */,
  {32'h40633658, 32'hbe99cdc0} /* (15, 4, 24) {real, imag} */,
  {32'hc0a34b2e, 32'hbfe84f6e} /* (15, 4, 23) {real, imag} */,
  {32'hbf874bb6, 32'hc0c7aa4c} /* (15, 4, 22) {real, imag} */,
  {32'h3f2b2f62, 32'hc0a8e580} /* (15, 4, 21) {real, imag} */,
  {32'hbe2c5b70, 32'hc0cebf23} /* (15, 4, 20) {real, imag} */,
  {32'hc16e9b47, 32'h40acf6d6} /* (15, 4, 19) {real, imag} */,
  {32'h40cb6a14, 32'hc0ca8c5e} /* (15, 4, 18) {real, imag} */,
  {32'h4012a4c6, 32'hc0aa39e5} /* (15, 4, 17) {real, imag} */,
  {32'hc0d91c69, 32'hc0b6950c} /* (15, 4, 16) {real, imag} */,
  {32'hc082eb07, 32'h418e0cb9} /* (15, 4, 15) {real, imag} */,
  {32'hc0e3e2d4, 32'hc0bd7ebd} /* (15, 4, 14) {real, imag} */,
  {32'h414316b5, 32'h3ff07f50} /* (15, 4, 13) {real, imag} */,
  {32'h3f8ee8b4, 32'h402aff94} /* (15, 4, 12) {real, imag} */,
  {32'h4140b383, 32'h40b6149a} /* (15, 4, 11) {real, imag} */,
  {32'h4170a6e2, 32'hc186eef5} /* (15, 4, 10) {real, imag} */,
  {32'h40b4424c, 32'hc0c54cbd} /* (15, 4, 9) {real, imag} */,
  {32'hc1452cb2, 32'hc0c349f0} /* (15, 4, 8) {real, imag} */,
  {32'h413dc926, 32'h41e73398} /* (15, 4, 7) {real, imag} */,
  {32'hc1c13c7e, 32'hc1bb5633} /* (15, 4, 6) {real, imag} */,
  {32'hc1bbe5f9, 32'hc15232e4} /* (15, 4, 5) {real, imag} */,
  {32'hc184f422, 32'h412c464b} /* (15, 4, 4) {real, imag} */,
  {32'hc18ee141, 32'h41bc9308} /* (15, 4, 3) {real, imag} */,
  {32'hc13dcab8, 32'hc236e4eb} /* (15, 4, 2) {real, imag} */,
  {32'h42c7996a, 32'h419f55d5} /* (15, 4, 1) {real, imag} */,
  {32'hc1dc134a, 32'hc218548b} /* (15, 4, 0) {real, imag} */,
  {32'h41835fde, 32'hbd397800} /* (15, 3, 31) {real, imag} */,
  {32'h4237d485, 32'hc19d1ab0} /* (15, 3, 30) {real, imag} */,
  {32'hc1d71ca0, 32'hc10c5562} /* (15, 3, 29) {real, imag} */,
  {32'h41cf13ec, 32'h417940f6} /* (15, 3, 28) {real, imag} */,
  {32'hc0dd8e40, 32'h412c4008} /* (15, 3, 27) {real, imag} */,
  {32'hbec9b4c0, 32'h41b87748} /* (15, 3, 26) {real, imag} */,
  {32'hc1afa7cf, 32'h3f6e18a0} /* (15, 3, 25) {real, imag} */,
  {32'hc1776c19, 32'hc13fae00} /* (15, 3, 24) {real, imag} */,
  {32'hc18bfd10, 32'h40d30932} /* (15, 3, 23) {real, imag} */,
  {32'h412be82a, 32'hc0a6f92a} /* (15, 3, 22) {real, imag} */,
  {32'hc057112c, 32'hc115ea64} /* (15, 3, 21) {real, imag} */,
  {32'hc0e0f4ea, 32'h41b8a196} /* (15, 3, 20) {real, imag} */,
  {32'hbfd85dc6, 32'hc167f592} /* (15, 3, 19) {real, imag} */,
  {32'h405418f0, 32'hc1554048} /* (15, 3, 18) {real, imag} */,
  {32'h3fc2587c, 32'h4178e007} /* (15, 3, 17) {real, imag} */,
  {32'hbf599f38, 32'hc08d8b9c} /* (15, 3, 16) {real, imag} */,
  {32'hc0e17484, 32'hc0614d6d} /* (15, 3, 15) {real, imag} */,
  {32'hbf21b824, 32'h3f8a287a} /* (15, 3, 14) {real, imag} */,
  {32'h4108c562, 32'h4133722d} /* (15, 3, 13) {real, imag} */,
  {32'h4091e365, 32'hc0b995d2} /* (15, 3, 12) {real, imag} */,
  {32'hc127e2a5, 32'h411a2dd3} /* (15, 3, 11) {real, imag} */,
  {32'hc0979c0c, 32'h40999ac6} /* (15, 3, 10) {real, imag} */,
  {32'hc1371e38, 32'h3f70825c} /* (15, 3, 9) {real, imag} */,
  {32'h40873249, 32'hc0d4793f} /* (15, 3, 8) {real, imag} */,
  {32'hc1205b99, 32'hc101857c} /* (15, 3, 7) {real, imag} */,
  {32'hc08373ec, 32'h40cf5ec6} /* (15, 3, 6) {real, imag} */,
  {32'h413b5d54, 32'h4143e139} /* (15, 3, 5) {real, imag} */,
  {32'hc192c4f2, 32'h41ec8acc} /* (15, 3, 4) {real, imag} */,
  {32'h409d4050, 32'h41775db8} /* (15, 3, 3) {real, imag} */,
  {32'h4145a74e, 32'hc2200cd7} /* (15, 3, 2) {real, imag} */,
  {32'h42687e13, 32'h40a0f4f0} /* (15, 3, 1) {real, imag} */,
  {32'h412d938e, 32'h41f45722} /* (15, 3, 0) {real, imag} */,
  {32'hc39cc5a7, 32'hc29cc922} /* (15, 2, 31) {real, imag} */,
  {32'h433a0394, 32'hc214978c} /* (15, 2, 30) {real, imag} */,
  {32'h4200f102, 32'h420c7ea2} /* (15, 2, 29) {real, imag} */,
  {32'hc1a3d818, 32'h42585694} /* (15, 2, 28) {real, imag} */,
  {32'h4103ec76, 32'hc0e96154} /* (15, 2, 27) {real, imag} */,
  {32'hc1bbffd0, 32'h420c132a} /* (15, 2, 26) {real, imag} */,
  {32'hc0b6ed96, 32'h40956dc5} /* (15, 2, 25) {real, imag} */,
  {32'h41812e38, 32'hc238869f} /* (15, 2, 24) {real, imag} */,
  {32'hc15177fa, 32'h4171ec78} /* (15, 2, 23) {real, imag} */,
  {32'h40de441a, 32'hc0c4be1e} /* (15, 2, 22) {real, imag} */,
  {32'h3f6e42e8, 32'hc0faeb06} /* (15, 2, 21) {real, imag} */,
  {32'hc0fb40f8, 32'hbeb09e00} /* (15, 2, 20) {real, imag} */,
  {32'hc0cee376, 32'h4122f9d4} /* (15, 2, 19) {real, imag} */,
  {32'h3fc22708, 32'h408be652} /* (15, 2, 18) {real, imag} */,
  {32'hbff66c02, 32'hc048f7fe} /* (15, 2, 17) {real, imag} */,
  {32'hc0bb5706, 32'hc0dd9872} /* (15, 2, 16) {real, imag} */,
  {32'h3ee3c278, 32'hc08d37ae} /* (15, 2, 15) {real, imag} */,
  {32'h40bc4161, 32'h41796a64} /* (15, 2, 14) {real, imag} */,
  {32'h40940144, 32'hbfb0bfba} /* (15, 2, 13) {real, imag} */,
  {32'h408e462c, 32'h41486628} /* (15, 2, 12) {real, imag} */,
  {32'hc12d1c62, 32'h4110aedd} /* (15, 2, 11) {real, imag} */,
  {32'hc18bedac, 32'hc1065a68} /* (15, 2, 10) {real, imag} */,
  {32'hc10bf8c0, 32'h41005efe} /* (15, 2, 9) {real, imag} */,
  {32'h41f18c62, 32'h3ff18db0} /* (15, 2, 8) {real, imag} */,
  {32'hbe2ab738, 32'h40d32c30} /* (15, 2, 7) {real, imag} */,
  {32'h4020a6df, 32'h4164eab7} /* (15, 2, 6) {real, imag} */,
  {32'h41bfdd0d, 32'h42279d04} /* (15, 2, 5) {real, imag} */,
  {32'h40e9a620, 32'hc27a85c9} /* (15, 2, 4) {real, imag} */,
  {32'h41ab8b3f, 32'hc10a9278} /* (15, 2, 3) {real, imag} */,
  {32'h42ec5e68, 32'hc1312d1c} /* (15, 2, 2) {real, imag} */,
  {32'hc31dbeae, 32'hc1aa6c18} /* (15, 2, 1) {real, imag} */,
  {32'hc34446ee, 32'h40618e20} /* (15, 2, 0) {real, imag} */,
  {32'h43d60f50, 32'hc3086eb9} /* (15, 1, 31) {real, imag} */,
  {32'hc3104efa, 32'hc218cc8b} /* (15, 1, 30) {real, imag} */,
  {32'hc0c0fadc, 32'h427f0978} /* (15, 1, 29) {real, imag} */,
  {32'h42458192, 32'hc1999196} /* (15, 1, 28) {real, imag} */,
  {32'hc2310238, 32'h41b4d6e6} /* (15, 1, 27) {real, imag} */,
  {32'h41d73571, 32'hc17115ce} /* (15, 1, 26) {real, imag} */,
  {32'hc010a002, 32'h416a7351} /* (15, 1, 25) {real, imag} */,
  {32'hc149a74e, 32'h4135d01a} /* (15, 1, 24) {real, imag} */,
  {32'hc143235a, 32'h4187b618} /* (15, 1, 23) {real, imag} */,
  {32'h4187daa9, 32'hc0a7086c} /* (15, 1, 22) {real, imag} */,
  {32'hc1764074, 32'h4103b3d4} /* (15, 1, 21) {real, imag} */,
  {32'h4160bff3, 32'hbfcbd704} /* (15, 1, 20) {real, imag} */,
  {32'h40c26fe1, 32'h41987dd0} /* (15, 1, 19) {real, imag} */,
  {32'hc0563de8, 32'h410bc191} /* (15, 1, 18) {real, imag} */,
  {32'h412a92c4, 32'hc0562f48} /* (15, 1, 17) {real, imag} */,
  {32'h40aa6adf, 32'hc18bfdf0} /* (15, 1, 16) {real, imag} */,
  {32'hc0fa9b04, 32'h410faaf0} /* (15, 1, 15) {real, imag} */,
  {32'h413ef1c5, 32'hc0ef4662} /* (15, 1, 14) {real, imag} */,
  {32'h4177cc9e, 32'hbf90055a} /* (15, 1, 13) {real, imag} */,
  {32'hc1062490, 32'hc1933f61} /* (15, 1, 12) {real, imag} */,
  {32'hc0f318b2, 32'hbf52feb0} /* (15, 1, 11) {real, imag} */,
  {32'h400bcd7e, 32'hc10aad7a} /* (15, 1, 10) {real, imag} */,
  {32'h3f2a78da, 32'h40b2ed53} /* (15, 1, 9) {real, imag} */,
  {32'hc19c2dfb, 32'hc1a15b96} /* (15, 1, 8) {real, imag} */,
  {32'h41e36749, 32'h4133a78e} /* (15, 1, 7) {real, imag} */,
  {32'h415d400e, 32'hc177816f} /* (15, 1, 6) {real, imag} */,
  {32'hc1470a0a, 32'hc1239f68} /* (15, 1, 5) {real, imag} */,
  {32'hc1c0ee98, 32'h4230abe2} /* (15, 1, 4) {real, imag} */,
  {32'hc27e0c61, 32'h40ef4938} /* (15, 1, 3) {real, imag} */,
  {32'hc3582234, 32'hc3079866} /* (15, 1, 2) {real, imag} */,
  {32'h43deba7e, 32'h43a76652} /* (15, 1, 1) {real, imag} */,
  {32'h43d4b47b, 32'hc2ce2f16} /* (15, 1, 0) {real, imag} */,
  {32'h4313a5c4, 32'hc32feab8} /* (15, 0, 31) {real, imag} */,
  {32'hc2056028, 32'h42de8106} /* (15, 0, 30) {real, imag} */,
  {32'h41dd4a56, 32'hc13a5708} /* (15, 0, 29) {real, imag} */,
  {32'hc245168a, 32'hc1764408} /* (15, 0, 28) {real, imag} */,
  {32'hc2384eee, 32'hc10f2b3e} /* (15, 0, 27) {real, imag} */,
  {32'h40d598be, 32'h408df1cb} /* (15, 0, 26) {real, imag} */,
  {32'h4167edae, 32'hc19d35cb} /* (15, 0, 25) {real, imag} */,
  {32'h3ebcd880, 32'h416e44c6} /* (15, 0, 24) {real, imag} */,
  {32'hc0226794, 32'h3e22be00} /* (15, 0, 23) {real, imag} */,
  {32'hc18e0b00, 32'hc09b5c34} /* (15, 0, 22) {real, imag} */,
  {32'hc10fec97, 32'h40e0fa74} /* (15, 0, 21) {real, imag} */,
  {32'h4163f586, 32'hbf126744} /* (15, 0, 20) {real, imag} */,
  {32'hc1689efa, 32'h4106d76a} /* (15, 0, 19) {real, imag} */,
  {32'h3fe0407c, 32'h41a086e4} /* (15, 0, 18) {real, imag} */,
  {32'h403abbb5, 32'h416647dd} /* (15, 0, 17) {real, imag} */,
  {32'h41751cb0, 32'h00000000} /* (15, 0, 16) {real, imag} */,
  {32'h403abbb5, 32'hc16647dd} /* (15, 0, 15) {real, imag} */,
  {32'h3fe0407c, 32'hc1a086e4} /* (15, 0, 14) {real, imag} */,
  {32'hc1689efa, 32'hc106d76a} /* (15, 0, 13) {real, imag} */,
  {32'h4163f586, 32'h3f126744} /* (15, 0, 12) {real, imag} */,
  {32'hc10fec97, 32'hc0e0fa74} /* (15, 0, 11) {real, imag} */,
  {32'hc18e0b00, 32'h409b5c34} /* (15, 0, 10) {real, imag} */,
  {32'hc0226794, 32'hbe22be00} /* (15, 0, 9) {real, imag} */,
  {32'h3ebcd880, 32'hc16e44c6} /* (15, 0, 8) {real, imag} */,
  {32'h4167edae, 32'h419d35cb} /* (15, 0, 7) {real, imag} */,
  {32'h40d598be, 32'hc08df1cb} /* (15, 0, 6) {real, imag} */,
  {32'hc2384eee, 32'h410f2b3e} /* (15, 0, 5) {real, imag} */,
  {32'hc245168a, 32'h41764408} /* (15, 0, 4) {real, imag} */,
  {32'h41dd4a56, 32'h413a5708} /* (15, 0, 3) {real, imag} */,
  {32'hc2056028, 32'hc2de8106} /* (15, 0, 2) {real, imag} */,
  {32'h4313a5c4, 32'h432feab8} /* (15, 0, 1) {real, imag} */,
  {32'h43e3b4ba, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h449b9faf, 32'hc4442c5e} /* (14, 31, 31) {real, imag} */,
  {32'hc3c4f800, 32'h43ac851c} /* (14, 31, 30) {real, imag} */,
  {32'hc2d292c6, 32'h41346ae2} /* (14, 31, 29) {real, imag} */,
  {32'hc201c90a, 32'hc28b4e7f} /* (14, 31, 28) {real, imag} */,
  {32'hc20e2118, 32'h41fe0fc7} /* (14, 31, 27) {real, imag} */,
  {32'h40462b18, 32'h42428469} /* (14, 31, 26) {real, imag} */,
  {32'h41bba0cb, 32'hc1f5aa6e} /* (14, 31, 25) {real, imag} */,
  {32'hc18d17b2, 32'h414c599e} /* (14, 31, 24) {real, imag} */,
  {32'hbffadf00, 32'hc0f06a1c} /* (14, 31, 23) {real, imag} */,
  {32'hc00ad7d8, 32'h4111c863} /* (14, 31, 22) {real, imag} */,
  {32'h3ec9ea30, 32'h419c8435} /* (14, 31, 21) {real, imag} */,
  {32'h40e6d3df, 32'h40cee9a6} /* (14, 31, 20) {real, imag} */,
  {32'h41a5bc2e, 32'hbda6aab0} /* (14, 31, 19) {real, imag} */,
  {32'hc010b127, 32'h4171a5a8} /* (14, 31, 18) {real, imag} */,
  {32'hc0b7a2e6, 32'hc0969be0} /* (14, 31, 17) {real, imag} */,
  {32'h40cfc513, 32'h4085c5da} /* (14, 31, 16) {real, imag} */,
  {32'hc06a6e9e, 32'hc0eb499e} /* (14, 31, 15) {real, imag} */,
  {32'hbfe14204, 32'hc12444f4} /* (14, 31, 14) {real, imag} */,
  {32'hbfd48f88, 32'h408c41e0} /* (14, 31, 13) {real, imag} */,
  {32'hc08537a0, 32'h408bb386} /* (14, 31, 12) {real, imag} */,
  {32'hc16b1256, 32'hc1fb4b94} /* (14, 31, 11) {real, imag} */,
  {32'h410330a7, 32'h404fd346} /* (14, 31, 10) {real, imag} */,
  {32'hc13d07ec, 32'h405cc148} /* (14, 31, 9) {real, imag} */,
  {32'hc20962fe, 32'hc00a0b3c} /* (14, 31, 8) {real, imag} */,
  {32'h3db42880, 32'hc1e734e8} /* (14, 31, 7) {real, imag} */,
  {32'h41bc57f6, 32'h40b6ba80} /* (14, 31, 6) {real, imag} */,
  {32'hc2a1f3d4, 32'hc1973340} /* (14, 31, 5) {real, imag} */,
  {32'h428bda14, 32'h40b2bcd8} /* (14, 31, 4) {real, imag} */,
  {32'h40625e82, 32'hc2786364} /* (14, 31, 3) {real, imag} */,
  {32'hc38f225e, 32'h418fbbcb} /* (14, 31, 2) {real, imag} */,
  {32'h44754011, 32'h43819160} /* (14, 31, 1) {real, imag} */,
  {32'h448aa966, 32'h417fab80} /* (14, 31, 0) {real, imag} */,
  {32'hc3dce4b0, 32'hc21bfa32} /* (14, 30, 31) {real, imag} */,
  {32'h437ef71b, 32'h41db8362} /* (14, 30, 30) {real, imag} */,
  {32'h40be1bd8, 32'hc0a6f602} /* (14, 30, 29) {real, imag} */,
  {32'hc23a6fd8, 32'h42790b6e} /* (14, 30, 28) {real, imag} */,
  {32'h425387d8, 32'hc29dad09} /* (14, 30, 27) {real, imag} */,
  {32'hc14bac48, 32'hc21a9d6f} /* (14, 30, 26) {real, imag} */,
  {32'hbf366040, 32'hc09e00c3} /* (14, 30, 25) {real, imag} */,
  {32'h4240d158, 32'hc16e1d02} /* (14, 30, 24) {real, imag} */,
  {32'h3f8ca328, 32'hc145aa72} /* (14, 30, 23) {real, imag} */,
  {32'hbf719170, 32'hc078a7ac} /* (14, 30, 22) {real, imag} */,
  {32'h40fab9d2, 32'hc181fa44} /* (14, 30, 21) {real, imag} */,
  {32'hbff1e780, 32'h4115bf64} /* (14, 30, 20) {real, imag} */,
  {32'hc1930e4a, 32'hc128162b} /* (14, 30, 19) {real, imag} */,
  {32'h41bce754, 32'hc0552982} /* (14, 30, 18) {real, imag} */,
  {32'hbf646878, 32'hbfee0fb6} /* (14, 30, 17) {real, imag} */,
  {32'h3fd507f8, 32'h40b23628} /* (14, 30, 16) {real, imag} */,
  {32'h40f98700, 32'hc184d02c} /* (14, 30, 15) {real, imag} */,
  {32'h40c92458, 32'h41903a1c} /* (14, 30, 14) {real, imag} */,
  {32'hc11fbfbf, 32'hc126809e} /* (14, 30, 13) {real, imag} */,
  {32'h40e26fd6, 32'h4138df83} /* (14, 30, 12) {real, imag} */,
  {32'h406be5cd, 32'h408c533c} /* (14, 30, 11) {real, imag} */,
  {32'h40ae2cb8, 32'hc177ca5b} /* (14, 30, 10) {real, imag} */,
  {32'h4032944b, 32'h415eecb2} /* (14, 30, 9) {real, imag} */,
  {32'h409c9cd3, 32'h416373d8} /* (14, 30, 8) {real, imag} */,
  {32'hc1ccc744, 32'hc115f5cf} /* (14, 30, 7) {real, imag} */,
  {32'h405fc6a8, 32'h41b90066} /* (14, 30, 6) {real, imag} */,
  {32'h423befd2, 32'h417e4132} /* (14, 30, 5) {real, imag} */,
  {32'hc24fb7b5, 32'hc2a96ac6} /* (14, 30, 4) {real, imag} */,
  {32'h41384045, 32'hc154297a} /* (14, 30, 3) {real, imag} */,
  {32'h43ca1049, 32'h431496c6} /* (14, 30, 2) {real, imag} */,
  {32'hc4404433, 32'h42800be0} /* (14, 30, 1) {real, imag} */,
  {32'hc3cedef5, 32'h42791f82} /* (14, 30, 0) {real, imag} */,
  {32'h42daa10d, 32'hc28aa287} /* (14, 29, 31) {real, imag} */,
  {32'hc1d7d97b, 32'h427eee7a} /* (14, 29, 30) {real, imag} */,
  {32'h4190bc2d, 32'hc14550dc} /* (14, 29, 29) {real, imag} */,
  {32'hc0f44766, 32'hc1a2b238} /* (14, 29, 28) {real, imag} */,
  {32'h40a551f8, 32'hc20a92a0} /* (14, 29, 27) {real, imag} */,
  {32'h3f1e43c0, 32'h40a74f0c} /* (14, 29, 26) {real, imag} */,
  {32'h41c5b8bc, 32'h40c3492c} /* (14, 29, 25) {real, imag} */,
  {32'h413e50a5, 32'hbf478ec0} /* (14, 29, 24) {real, imag} */,
  {32'hc0df326e, 32'h41eef5bc} /* (14, 29, 23) {real, imag} */,
  {32'hc01a3350, 32'hc09a661c} /* (14, 29, 22) {real, imag} */,
  {32'h413f6950, 32'hc18759ef} /* (14, 29, 21) {real, imag} */,
  {32'h40280470, 32'hc025163c} /* (14, 29, 20) {real, imag} */,
  {32'hbf839296, 32'h3fe41104} /* (14, 29, 19) {real, imag} */,
  {32'h411e6c95, 32'hc0518254} /* (14, 29, 18) {real, imag} */,
  {32'hc0d6e812, 32'hc10848bc} /* (14, 29, 17) {real, imag} */,
  {32'hc0850566, 32'hbfcaaae0} /* (14, 29, 16) {real, imag} */,
  {32'hc0496dfb, 32'hbfa6038c} /* (14, 29, 15) {real, imag} */,
  {32'hbff62d7f, 32'h40aea436} /* (14, 29, 14) {real, imag} */,
  {32'h412c1c13, 32'h409b2ac4} /* (14, 29, 13) {real, imag} */,
  {32'h411a6fe2, 32'hc13a8d5e} /* (14, 29, 12) {real, imag} */,
  {32'hc136a7db, 32'h413b18dc} /* (14, 29, 11) {real, imag} */,
  {32'hc11849e9, 32'hc1bf51fd} /* (14, 29, 10) {real, imag} */,
  {32'hc1a59772, 32'h40e95803} /* (14, 29, 9) {real, imag} */,
  {32'hc13dad1d, 32'h410d8afe} /* (14, 29, 8) {real, imag} */,
  {32'hc0611cb9, 32'h40f19618} /* (14, 29, 7) {real, imag} */,
  {32'hc10bb090, 32'h40529ec8} /* (14, 29, 6) {real, imag} */,
  {32'hc1981f2e, 32'h41048d60} /* (14, 29, 5) {real, imag} */,
  {32'h41cbba10, 32'hc18aeab8} /* (14, 29, 4) {real, imag} */,
  {32'hc11d9938, 32'hc1f94558} /* (14, 29, 3) {real, imag} */,
  {32'h428c3096, 32'h42549870} /* (14, 29, 2) {real, imag} */,
  {32'hc2a04d1c, 32'hc23015a3} /* (14, 29, 1) {real, imag} */,
  {32'h41a3d1be, 32'hc0d22f1e} /* (14, 29, 0) {real, imag} */,
  {32'h4321860a, 32'hc1dfed02} /* (14, 28, 31) {real, imag} */,
  {32'hc27d71c0, 32'h4280cfd4} /* (14, 28, 30) {real, imag} */,
  {32'hc14c4708, 32'hc1b6cea1} /* (14, 28, 29) {real, imag} */,
  {32'h417d4c94, 32'hc1e268e5} /* (14, 28, 28) {real, imag} */,
  {32'hc1a04ab9, 32'h4154b97a} /* (14, 28, 27) {real, imag} */,
  {32'hc1a45d95, 32'hc195fbc3} /* (14, 28, 26) {real, imag} */,
  {32'hc0a2d18d, 32'hc05598ec} /* (14, 28, 25) {real, imag} */,
  {32'hc08b8abd, 32'hc0f6d71a} /* (14, 28, 24) {real, imag} */,
  {32'h4215c679, 32'h40d725db} /* (14, 28, 23) {real, imag} */,
  {32'h411ff1de, 32'hc1acefd6} /* (14, 28, 22) {real, imag} */,
  {32'hc0f23ae4, 32'h40638603} /* (14, 28, 21) {real, imag} */,
  {32'h3f67cb54, 32'h405c865c} /* (14, 28, 20) {real, imag} */,
  {32'hc0c545e5, 32'hc09355fe} /* (14, 28, 19) {real, imag} */,
  {32'hc0aec4c5, 32'h41742284} /* (14, 28, 18) {real, imag} */,
  {32'hbfda3196, 32'h416ed944} /* (14, 28, 17) {real, imag} */,
  {32'h4053392a, 32'h3ea19e58} /* (14, 28, 16) {real, imag} */,
  {32'hc11c6e6b, 32'hc1151f59} /* (14, 28, 15) {real, imag} */,
  {32'hc0cca6f4, 32'hc05820bd} /* (14, 28, 14) {real, imag} */,
  {32'hc15e1de1, 32'h4187f8f1} /* (14, 28, 13) {real, imag} */,
  {32'h3fc17eec, 32'hc066af62} /* (14, 28, 12) {real, imag} */,
  {32'hc0f96f88, 32'hc07a4d25} /* (14, 28, 11) {real, imag} */,
  {32'hc0ba6203, 32'hc0515d70} /* (14, 28, 10) {real, imag} */,
  {32'hc02f57e4, 32'h41142478} /* (14, 28, 9) {real, imag} */,
  {32'hc141fbbe, 32'hc0fe98f2} /* (14, 28, 8) {real, imag} */,
  {32'hc0fe5b74, 32'hc20cc61a} /* (14, 28, 7) {real, imag} */,
  {32'hc04ecff4, 32'hc164c278} /* (14, 28, 6) {real, imag} */,
  {32'hc1944570, 32'hc1bfcf1e} /* (14, 28, 5) {real, imag} */,
  {32'h41d28d42, 32'hc231772c} /* (14, 28, 4) {real, imag} */,
  {32'hc17d9df8, 32'h41127616} /* (14, 28, 3) {real, imag} */,
  {32'hc24f7cae, 32'h429f0bce} /* (14, 28, 2) {real, imag} */,
  {32'h428f529d, 32'hc1d443c0} /* (14, 28, 1) {real, imag} */,
  {32'hc05038b8, 32'h41b63da8} /* (14, 28, 0) {real, imag} */,
  {32'hc2cd3d71, 32'h41a48e40} /* (14, 27, 31) {real, imag} */,
  {32'hbd86c500, 32'hc15e278c} /* (14, 27, 30) {real, imag} */,
  {32'hc05c9e28, 32'hc00d9280} /* (14, 27, 29) {real, imag} */,
  {32'h40f2bc27, 32'h4170e036} /* (14, 27, 28) {real, imag} */,
  {32'h415a6178, 32'hc1ae6b49} /* (14, 27, 27) {real, imag} */,
  {32'h4145672d, 32'h3f115b80} /* (14, 27, 26) {real, imag} */,
  {32'hc0d9279e, 32'hbee41dd8} /* (14, 27, 25) {real, imag} */,
  {32'hc16bae52, 32'hc1467e9e} /* (14, 27, 24) {real, imag} */,
  {32'h4007d2b4, 32'h400eb2d8} /* (14, 27, 23) {real, imag} */,
  {32'h3ff25186, 32'hc17725a7} /* (14, 27, 22) {real, imag} */,
  {32'hbf816d0e, 32'h3f685bc0} /* (14, 27, 21) {real, imag} */,
  {32'hc121158d, 32'hc0837c86} /* (14, 27, 20) {real, imag} */,
  {32'h413f3c45, 32'h4097a45a} /* (14, 27, 19) {real, imag} */,
  {32'h3e356860, 32'hc17cd092} /* (14, 27, 18) {real, imag} */,
  {32'h40db2fab, 32'h3fdb4002} /* (14, 27, 17) {real, imag} */,
  {32'hbfd3ad4e, 32'h4088e3d4} /* (14, 27, 16) {real, imag} */,
  {32'h409313db, 32'hc036a100} /* (14, 27, 15) {real, imag} */,
  {32'h41174fbe, 32'h40e312c4} /* (14, 27, 14) {real, imag} */,
  {32'hbeda2e8a, 32'hc042ad0c} /* (14, 27, 13) {real, imag} */,
  {32'hc0ac88ba, 32'h3fde12dc} /* (14, 27, 12) {real, imag} */,
  {32'h410b0d2c, 32'h3f2a6d28} /* (14, 27, 11) {real, imag} */,
  {32'hbe5edee0, 32'h3ff3fd54} /* (14, 27, 10) {real, imag} */,
  {32'h402f7814, 32'h3fc058d5} /* (14, 27, 9) {real, imag} */,
  {32'h408be2f0, 32'hbf8f8218} /* (14, 27, 8) {real, imag} */,
  {32'hc097b01e, 32'hc103c661} /* (14, 27, 7) {real, imag} */,
  {32'hc105c78e, 32'hc0b95292} /* (14, 27, 6) {real, imag} */,
  {32'h41a12148, 32'h41057d60} /* (14, 27, 5) {real, imag} */,
  {32'hc103166e, 32'h40901be0} /* (14, 27, 4) {real, imag} */,
  {32'hc11bf32b, 32'hc1a13c4d} /* (14, 27, 3) {real, imag} */,
  {32'h40bf196c, 32'hc119df2d} /* (14, 27, 2) {real, imag} */,
  {32'hc28a8fb9, 32'hc2106b62} /* (14, 27, 1) {real, imag} */,
  {32'hc282f9fd, 32'h42203f75} /* (14, 27, 0) {real, imag} */,
  {32'hc1650a4d, 32'h3e1fa320} /* (14, 26, 31) {real, imag} */,
  {32'h41e4a15d, 32'hc107f3d8} /* (14, 26, 30) {real, imag} */,
  {32'h40903f6c, 32'hc19dd5dc} /* (14, 26, 29) {real, imag} */,
  {32'hc124bb72, 32'hc0c1714b} /* (14, 26, 28) {real, imag} */,
  {32'h3f4130a8, 32'h41a68dfc} /* (14, 26, 27) {real, imag} */,
  {32'hc14dae02, 32'hc0870fd2} /* (14, 26, 26) {real, imag} */,
  {32'hbf95af88, 32'h4123e626} /* (14, 26, 25) {real, imag} */,
  {32'h40dc6480, 32'hc11f0860} /* (14, 26, 24) {real, imag} */,
  {32'hc12abd29, 32'hc100f859} /* (14, 26, 23) {real, imag} */,
  {32'h4191b883, 32'hbffffbc2} /* (14, 26, 22) {real, imag} */,
  {32'h4150c398, 32'h410f4176} /* (14, 26, 21) {real, imag} */,
  {32'h40f73050, 32'h40ca2770} /* (14, 26, 20) {real, imag} */,
  {32'h402955b4, 32'h4007b2a4} /* (14, 26, 19) {real, imag} */,
  {32'hc15fa61c, 32'hbeae2298} /* (14, 26, 18) {real, imag} */,
  {32'h4107bd8f, 32'hc02e5980} /* (14, 26, 17) {real, imag} */,
  {32'hbe4b79b8, 32'h3f626804} /* (14, 26, 16) {real, imag} */,
  {32'hc02f6a21, 32'h417e59a8} /* (14, 26, 15) {real, imag} */,
  {32'h401cf1fa, 32'h41198f25} /* (14, 26, 14) {real, imag} */,
  {32'h40d77f42, 32'h41526a7a} /* (14, 26, 13) {real, imag} */,
  {32'hbfd8aac8, 32'hc19249e2} /* (14, 26, 12) {real, imag} */,
  {32'hc088f2e9, 32'hc11cdd25} /* (14, 26, 11) {real, imag} */,
  {32'hc0a93bda, 32'h4189bc72} /* (14, 26, 10) {real, imag} */,
  {32'h40e789e5, 32'hc1903725} /* (14, 26, 9) {real, imag} */,
  {32'hc0077de8, 32'hc10768ad} /* (14, 26, 8) {real, imag} */,
  {32'hc1a93a68, 32'h41fe66ad} /* (14, 26, 7) {real, imag} */,
  {32'h40dabdea, 32'hc1b663df} /* (14, 26, 6) {real, imag} */,
  {32'hc114de72, 32'hc0de7216} /* (14, 26, 5) {real, imag} */,
  {32'hc14cac08, 32'h4103f7fe} /* (14, 26, 4) {real, imag} */,
  {32'hc20a773c, 32'h41870b6e} /* (14, 26, 3) {real, imag} */,
  {32'h41c93076, 32'hc0a54934} /* (14, 26, 2) {real, imag} */,
  {32'h412c37d9, 32'hc113cbb8} /* (14, 26, 1) {real, imag} */,
  {32'hc1324388, 32'hc070aaa4} /* (14, 26, 0) {real, imag} */,
  {32'hc0f51c4e, 32'hc1e36c2e} /* (14, 25, 31) {real, imag} */,
  {32'h40956b2c, 32'h419833ce} /* (14, 25, 30) {real, imag} */,
  {32'hc088a118, 32'h40ff7a2c} /* (14, 25, 29) {real, imag} */,
  {32'hc1ee6cac, 32'hc184a701} /* (14, 25, 28) {real, imag} */,
  {32'hc109f044, 32'h4096c99a} /* (14, 25, 27) {real, imag} */,
  {32'h412bf63a, 32'h412c81a8} /* (14, 25, 26) {real, imag} */,
  {32'hc0edb2b6, 32'h415a94f4} /* (14, 25, 25) {real, imag} */,
  {32'h4115c152, 32'h41b0954c} /* (14, 25, 24) {real, imag} */,
  {32'hc129c79b, 32'h419a7a14} /* (14, 25, 23) {real, imag} */,
  {32'hbfb37cac, 32'hc1b3a45c} /* (14, 25, 22) {real, imag} */,
  {32'hc09670a6, 32'hc085bc8b} /* (14, 25, 21) {real, imag} */,
  {32'hc18a9490, 32'hc17f0658} /* (14, 25, 20) {real, imag} */,
  {32'h3fcd5a2c, 32'hc1c32e6d} /* (14, 25, 19) {real, imag} */,
  {32'hc0a6c378, 32'hbe95b040} /* (14, 25, 18) {real, imag} */,
  {32'h4103890f, 32'hc0a5e198} /* (14, 25, 17) {real, imag} */,
  {32'h4129d26c, 32'hc1668c96} /* (14, 25, 16) {real, imag} */,
  {32'h41204da6, 32'h3fa0e598} /* (14, 25, 15) {real, imag} */,
  {32'hc08fd3ed, 32'h3ff1fa00} /* (14, 25, 14) {real, imag} */,
  {32'h412b7bc6, 32'hc118d94d} /* (14, 25, 13) {real, imag} */,
  {32'h41b69b24, 32'h41db02b9} /* (14, 25, 12) {real, imag} */,
  {32'h412cba39, 32'h40bc2ff9} /* (14, 25, 11) {real, imag} */,
  {32'h41084198, 32'hc0470696} /* (14, 25, 10) {real, imag} */,
  {32'hc10ee0e5, 32'hc1059fef} /* (14, 25, 9) {real, imag} */,
  {32'hbf5ffd68, 32'h3fdb750a} /* (14, 25, 8) {real, imag} */,
  {32'hc11c5816, 32'hc080fda0} /* (14, 25, 7) {real, imag} */,
  {32'hc1a8b55b, 32'h3fff4468} /* (14, 25, 6) {real, imag} */,
  {32'hc187d4d8, 32'hc1ebc854} /* (14, 25, 5) {real, imag} */,
  {32'hc10eef98, 32'h41259c4d} /* (14, 25, 4) {real, imag} */,
  {32'h40765ea0, 32'h4080ace5} /* (14, 25, 3) {real, imag} */,
  {32'hc0a10d46, 32'h41ea0730} /* (14, 25, 2) {real, imag} */,
  {32'h41e64b91, 32'h41a8ec68} /* (14, 25, 1) {real, imag} */,
  {32'hbff1350c, 32'hc21d80aa} /* (14, 25, 0) {real, imag} */,
  {32'hc1aea470, 32'h420a9226} /* (14, 24, 31) {real, imag} */,
  {32'h41b65f51, 32'hc06e5a60} /* (14, 24, 30) {real, imag} */,
  {32'hc0b0765f, 32'hc0c1c104} /* (14, 24, 29) {real, imag} */,
  {32'hc1cc9cd6, 32'hc0087159} /* (14, 24, 28) {real, imag} */,
  {32'hbfff0ef6, 32'hc1c88ef6} /* (14, 24, 27) {real, imag} */,
  {32'h401923af, 32'hbfb254ec} /* (14, 24, 26) {real, imag} */,
  {32'h4108f3c7, 32'hc0c6f734} /* (14, 24, 25) {real, imag} */,
  {32'hbf2db8c0, 32'hbe0b3bc0} /* (14, 24, 24) {real, imag} */,
  {32'hc0cf55fd, 32'hc044726f} /* (14, 24, 23) {real, imag} */,
  {32'hc1e3d422, 32'hc0c6dfd0} /* (14, 24, 22) {real, imag} */,
  {32'h4190ff78, 32'h40ec41ea} /* (14, 24, 21) {real, imag} */,
  {32'hc13784c2, 32'h41350657} /* (14, 24, 20) {real, imag} */,
  {32'hbf2c4510, 32'h40bc17f3} /* (14, 24, 19) {real, imag} */,
  {32'h4099a760, 32'hc09b7eae} /* (14, 24, 18) {real, imag} */,
  {32'hc1194266, 32'h417160dd} /* (14, 24, 17) {real, imag} */,
  {32'hc0db26aa, 32'hc0d3c248} /* (14, 24, 16) {real, imag} */,
  {32'hc086c192, 32'hc12a9510} /* (14, 24, 15) {real, imag} */,
  {32'h3f31ff88, 32'h3fa6cf1c} /* (14, 24, 14) {real, imag} */,
  {32'h405579c4, 32'hc1286238} /* (14, 24, 13) {real, imag} */,
  {32'hc14012a8, 32'hc0b3907d} /* (14, 24, 12) {real, imag} */,
  {32'h4150918c, 32'h3f44b998} /* (14, 24, 11) {real, imag} */,
  {32'h40b0e129, 32'h4191a2dc} /* (14, 24, 10) {real, imag} */,
  {32'hc03e9ce8, 32'h41526e8f} /* (14, 24, 9) {real, imag} */,
  {32'h3e0a84e8, 32'h40cb9b90} /* (14, 24, 8) {real, imag} */,
  {32'h414d44c3, 32'hc08da6a8} /* (14, 24, 7) {real, imag} */,
  {32'h4161e62d, 32'hbfa7a084} /* (14, 24, 6) {real, imag} */,
  {32'h41c04486, 32'h3f86343a} /* (14, 24, 5) {real, imag} */,
  {32'hc1393fa0, 32'hc11ca426} /* (14, 24, 4) {real, imag} */,
  {32'h413f9e15, 32'h40ef409a} /* (14, 24, 3) {real, imag} */,
  {32'h41aeaa56, 32'hc1998e3b} /* (14, 24, 2) {real, imag} */,
  {32'hc28b4cde, 32'h421379d5} /* (14, 24, 1) {real, imag} */,
  {32'hc1ba0d4e, 32'h40e4e9e6} /* (14, 24, 0) {real, imag} */,
  {32'h3f9144c0, 32'h3ff2ffb8} /* (14, 23, 31) {real, imag} */,
  {32'h4096cdaf, 32'h40d7fdf8} /* (14, 23, 30) {real, imag} */,
  {32'hc0f27797, 32'hc11d50a5} /* (14, 23, 29) {real, imag} */,
  {32'hc0bb1f17, 32'hc1499d1d} /* (14, 23, 28) {real, imag} */,
  {32'h413dc41b, 32'h413ab2c3} /* (14, 23, 27) {real, imag} */,
  {32'hc0a1a11a, 32'h419afbba} /* (14, 23, 26) {real, imag} */,
  {32'hc1b582ae, 32'hc111940a} /* (14, 23, 25) {real, imag} */,
  {32'hc158d8f3, 32'hc147ad17} /* (14, 23, 24) {real, imag} */,
  {32'h40da1cc1, 32'h400b4bec} /* (14, 23, 23) {real, imag} */,
  {32'hc080633b, 32'hc16fc54c} /* (14, 23, 22) {real, imag} */,
  {32'hc111e473, 32'hc14988be} /* (14, 23, 21) {real, imag} */,
  {32'hc1141b13, 32'h40c1febe} /* (14, 23, 20) {real, imag} */,
  {32'h40cd795c, 32'h41180da8} /* (14, 23, 19) {real, imag} */,
  {32'hc1231163, 32'hbf7c4b64} /* (14, 23, 18) {real, imag} */,
  {32'hbf800f72, 32'h4186e588} /* (14, 23, 17) {real, imag} */,
  {32'hc09735ab, 32'hc02e30ec} /* (14, 23, 16) {real, imag} */,
  {32'hc127d911, 32'h40ea68e0} /* (14, 23, 15) {real, imag} */,
  {32'h41aa6e97, 32'h41972b7f} /* (14, 23, 14) {real, imag} */,
  {32'h41915c1c, 32'h415e164f} /* (14, 23, 13) {real, imag} */,
  {32'hc04f694a, 32'hbedb8520} /* (14, 23, 12) {real, imag} */,
  {32'hc1b61464, 32'hc126f738} /* (14, 23, 11) {real, imag} */,
  {32'hc1391550, 32'hc0fa17ce} /* (14, 23, 10) {real, imag} */,
  {32'hc103d0fb, 32'h4038e3e4} /* (14, 23, 9) {real, imag} */,
  {32'h40c9773a, 32'h411ecf6c} /* (14, 23, 8) {real, imag} */,
  {32'h41cc817f, 32'hc1163ba8} /* (14, 23, 7) {real, imag} */,
  {32'h41033108, 32'h40445c80} /* (14, 23, 6) {real, imag} */,
  {32'hc1a61ebf, 32'h4138b3c8} /* (14, 23, 5) {real, imag} */,
  {32'h414414a9, 32'hc0dfa954} /* (14, 23, 4) {real, imag} */,
  {32'h41009193, 32'hc06a286f} /* (14, 23, 3) {real, imag} */,
  {32'hc017aa20, 32'h416eec56} /* (14, 23, 2) {real, imag} */,
  {32'hc0a59db5, 32'hc185d1b4} /* (14, 23, 1) {real, imag} */,
  {32'h40ef8717, 32'hc0b4ceba} /* (14, 23, 0) {real, imag} */,
  {32'h41e70a46, 32'hc08f2d3b} /* (14, 22, 31) {real, imag} */,
  {32'hc0b89566, 32'h3f88d198} /* (14, 22, 30) {real, imag} */,
  {32'hc0894436, 32'hc0997633} /* (14, 22, 29) {real, imag} */,
  {32'hbf94d510, 32'h419810cc} /* (14, 22, 28) {real, imag} */,
  {32'h4178faf0, 32'h3da17f00} /* (14, 22, 27) {real, imag} */,
  {32'h410955ea, 32'hbff669ec} /* (14, 22, 26) {real, imag} */,
  {32'h41236ee6, 32'hc033e555} /* (14, 22, 25) {real, imag} */,
  {32'hbffb5fc8, 32'h3fbef619} /* (14, 22, 24) {real, imag} */,
  {32'h4082e1b3, 32'h4184af94} /* (14, 22, 23) {real, imag} */,
  {32'h40270212, 32'h41686cb2} /* (14, 22, 22) {real, imag} */,
  {32'h41948a6d, 32'h401fa698} /* (14, 22, 21) {real, imag} */,
  {32'h3eea5ca0, 32'hc1339646} /* (14, 22, 20) {real, imag} */,
  {32'hc0625868, 32'h41645687} /* (14, 22, 19) {real, imag} */,
  {32'h3fe63f28, 32'hc0b8e038} /* (14, 22, 18) {real, imag} */,
  {32'hc18e4ea6, 32'hc151fe88} /* (14, 22, 17) {real, imag} */,
  {32'hc102234b, 32'h41190e8d} /* (14, 22, 16) {real, imag} */,
  {32'h40a48a77, 32'h41a5e7c5} /* (14, 22, 15) {real, imag} */,
  {32'h4081dda2, 32'h4001bd8e} /* (14, 22, 14) {real, imag} */,
  {32'hc0e0b663, 32'hc0256ee2} /* (14, 22, 13) {real, imag} */,
  {32'hbdd116e0, 32'h4122dc9c} /* (14, 22, 12) {real, imag} */,
  {32'h408b2ac3, 32'h41669055} /* (14, 22, 11) {real, imag} */,
  {32'h3f76f910, 32'hc07cdb92} /* (14, 22, 10) {real, imag} */,
  {32'h41155a53, 32'hc1bc4af6} /* (14, 22, 9) {real, imag} */,
  {32'hc12a9ed4, 32'hc11acb56} /* (14, 22, 8) {real, imag} */,
  {32'h41aea7ae, 32'hc1c2a69e} /* (14, 22, 7) {real, imag} */,
  {32'h41b985d9, 32'hc09a9b70} /* (14, 22, 6) {real, imag} */,
  {32'hc101bdd8, 32'h40dd8994} /* (14, 22, 5) {real, imag} */,
  {32'hc1aa1715, 32'hc09f50f4} /* (14, 22, 4) {real, imag} */,
  {32'hc02e4d7a, 32'hbf360260} /* (14, 22, 3) {real, imag} */,
  {32'h40579e20, 32'h41b0250c} /* (14, 22, 2) {real, imag} */,
  {32'hc092e34a, 32'hc10f28c3} /* (14, 22, 1) {real, imag} */,
  {32'h41229090, 32'hc1cefe2b} /* (14, 22, 0) {real, imag} */,
  {32'h3f2b12da, 32'h41fbaf2a} /* (14, 21, 31) {real, imag} */,
  {32'hc0145138, 32'hc155eb35} /* (14, 21, 30) {real, imag} */,
  {32'hc09daa61, 32'hc10076b6} /* (14, 21, 29) {real, imag} */,
  {32'h3ffbaf97, 32'h41104fba} /* (14, 21, 28) {real, imag} */,
  {32'hc09754a3, 32'hc0e42ca6} /* (14, 21, 27) {real, imag} */,
  {32'h4182d79c, 32'hc15c5786} /* (14, 21, 26) {real, imag} */,
  {32'h415775a8, 32'hc17afa1b} /* (14, 21, 25) {real, imag} */,
  {32'h4045fc20, 32'hc09d54b8} /* (14, 21, 24) {real, imag} */,
  {32'hc0aaeb46, 32'h3f600658} /* (14, 21, 23) {real, imag} */,
  {32'h4079b8a2, 32'h41b622c2} /* (14, 21, 22) {real, imag} */,
  {32'hc0daef2a, 32'h416d6f43} /* (14, 21, 21) {real, imag} */,
  {32'h40f03928, 32'h405ddc29} /* (14, 21, 20) {real, imag} */,
  {32'h416a0856, 32'h400f1dea} /* (14, 21, 19) {real, imag} */,
  {32'h41790ef0, 32'hc162ec17} /* (14, 21, 18) {real, imag} */,
  {32'h4104cf07, 32'hbfe8e494} /* (14, 21, 17) {real, imag} */,
  {32'hc17ab361, 32'h3fc0e98a} /* (14, 21, 16) {real, imag} */,
  {32'hc0bf3d1a, 32'hc00ee391} /* (14, 21, 15) {real, imag} */,
  {32'h40586fe5, 32'h3f10166e} /* (14, 21, 14) {real, imag} */,
  {32'hc1818b8d, 32'hc109ce17} /* (14, 21, 13) {real, imag} */,
  {32'hc0b52ea2, 32'hc0971131} /* (14, 21, 12) {real, imag} */,
  {32'h41330e8a, 32'hc1b9a82d} /* (14, 21, 11) {real, imag} */,
  {32'hbeffe100, 32'h40a2f092} /* (14, 21, 10) {real, imag} */,
  {32'h416d133e, 32'h4165aad3} /* (14, 21, 9) {real, imag} */,
  {32'h41544e2f, 32'h418e26d8} /* (14, 21, 8) {real, imag} */,
  {32'h411027f2, 32'h4161efce} /* (14, 21, 7) {real, imag} */,
  {32'hc011eb64, 32'h40b10b6b} /* (14, 21, 6) {real, imag} */,
  {32'h41c4d613, 32'hc18eda24} /* (14, 21, 5) {real, imag} */,
  {32'hbf7deb44, 32'hc10658b2} /* (14, 21, 4) {real, imag} */,
  {32'hc18ca28e, 32'hbf78ba58} /* (14, 21, 3) {real, imag} */,
  {32'hc030a0e4, 32'hc198fa90} /* (14, 21, 2) {real, imag} */,
  {32'hc1c43bc0, 32'h406ad3be} /* (14, 21, 1) {real, imag} */,
  {32'hc1906db5, 32'h41f66e78} /* (14, 21, 0) {real, imag} */,
  {32'h4180fceb, 32'hc04c4d48} /* (14, 20, 31) {real, imag} */,
  {32'h4085882c, 32'hbf5641f0} /* (14, 20, 30) {real, imag} */,
  {32'hc068c3eb, 32'hc125ac4a} /* (14, 20, 29) {real, imag} */,
  {32'h4146ac00, 32'h40b3d437} /* (14, 20, 28) {real, imag} */,
  {32'hc0919b36, 32'hbf91d10d} /* (14, 20, 27) {real, imag} */,
  {32'h4071a94f, 32'h413914c1} /* (14, 20, 26) {real, imag} */,
  {32'h41509ac1, 32'hbfcc4e50} /* (14, 20, 25) {real, imag} */,
  {32'hc12bab96, 32'h411a2f5c} /* (14, 20, 24) {real, imag} */,
  {32'hc10fed94, 32'hc19568eb} /* (14, 20, 23) {real, imag} */,
  {32'hc0a2390f, 32'hc0b94af9} /* (14, 20, 22) {real, imag} */,
  {32'hc1177a16, 32'hc06ecae2} /* (14, 20, 21) {real, imag} */,
  {32'hc13c2880, 32'h40fdaffe} /* (14, 20, 20) {real, imag} */,
  {32'hbe450088, 32'h40d84515} /* (14, 20, 19) {real, imag} */,
  {32'hc0ad15f8, 32'h4023df9a} /* (14, 20, 18) {real, imag} */,
  {32'hc1424eaf, 32'h4015fac4} /* (14, 20, 17) {real, imag} */,
  {32'hbfc3a4ec, 32'h403d1d18} /* (14, 20, 16) {real, imag} */,
  {32'hc11fa2d2, 32'h3f41ef8e} /* (14, 20, 15) {real, imag} */,
  {32'hc06ef3c0, 32'h410befa5} /* (14, 20, 14) {real, imag} */,
  {32'h411e32d6, 32'hc17d7a7e} /* (14, 20, 13) {real, imag} */,
  {32'hc16ac9f4, 32'hc02d35da} /* (14, 20, 12) {real, imag} */,
  {32'h40eb8024, 32'h40d726a7} /* (14, 20, 11) {real, imag} */,
  {32'h4102973a, 32'h3fd213bc} /* (14, 20, 10) {real, imag} */,
  {32'hc0fbe71f, 32'hc08b31d6} /* (14, 20, 9) {real, imag} */,
  {32'h414091b1, 32'hc0ebd58c} /* (14, 20, 8) {real, imag} */,
  {32'h3f9cfaae, 32'h411ec116} /* (14, 20, 7) {real, imag} */,
  {32'hc114b019, 32'hc0816204} /* (14, 20, 6) {real, imag} */,
  {32'h3fec36fe, 32'h4147e1b3} /* (14, 20, 5) {real, imag} */,
  {32'h4034dfe9, 32'h410d1f42} /* (14, 20, 4) {real, imag} */,
  {32'h3f6dff10, 32'h4057e6ee} /* (14, 20, 3) {real, imag} */,
  {32'h4091835f, 32'hc194468e} /* (14, 20, 2) {real, imag} */,
  {32'hc0e4bf90, 32'hbfb0e358} /* (14, 20, 1) {real, imag} */,
  {32'h4150862e, 32'h40a4bb46} /* (14, 20, 0) {real, imag} */,
  {32'h41050d3c, 32'hc14bedda} /* (14, 19, 31) {real, imag} */,
  {32'h40b1d12c, 32'hc0ea931b} /* (14, 19, 30) {real, imag} */,
  {32'h3d55cbe0, 32'hc0ec8c86} /* (14, 19, 29) {real, imag} */,
  {32'hc0cff28f, 32'hbfdb15a0} /* (14, 19, 28) {real, imag} */,
  {32'hc04bd2c4, 32'hc11a3d0f} /* (14, 19, 27) {real, imag} */,
  {32'h40d64742, 32'h40ea1520} /* (14, 19, 26) {real, imag} */,
  {32'hbfc4980c, 32'h3fe5c6ac} /* (14, 19, 25) {real, imag} */,
  {32'hc09f361f, 32'hc0bad620} /* (14, 19, 24) {real, imag} */,
  {32'hc0c296f8, 32'hc09212bc} /* (14, 19, 23) {real, imag} */,
  {32'h40dd079c, 32'h4080f852} /* (14, 19, 22) {real, imag} */,
  {32'hbfb345d0, 32'h412ad11c} /* (14, 19, 21) {real, imag} */,
  {32'hbf6edd6c, 32'hc1861bb1} /* (14, 19, 20) {real, imag} */,
  {32'h3efd4a70, 32'hc0a59fc9} /* (14, 19, 19) {real, imag} */,
  {32'h417e3368, 32'h41025e56} /* (14, 19, 18) {real, imag} */,
  {32'hc1c5d546, 32'hc08c5787} /* (14, 19, 17) {real, imag} */,
  {32'h4058d8ac, 32'hc09ae742} /* (14, 19, 16) {real, imag} */,
  {32'h40187ce6, 32'hc0ec2d28} /* (14, 19, 15) {real, imag} */,
  {32'hc1863cd1, 32'h4127723e} /* (14, 19, 14) {real, imag} */,
  {32'hc169dcd9, 32'h40ec664a} /* (14, 19, 13) {real, imag} */,
  {32'h415fb897, 32'h417ab5b4} /* (14, 19, 12) {real, imag} */,
  {32'h406dafc9, 32'hc06580c8} /* (14, 19, 11) {real, imag} */,
  {32'hc0813e79, 32'hc0dce3de} /* (14, 19, 10) {real, imag} */,
  {32'hc0e248c9, 32'hc1094285} /* (14, 19, 9) {real, imag} */,
  {32'hc010cd97, 32'hbe1dace0} /* (14, 19, 8) {real, imag} */,
  {32'h414c208f, 32'hbf2edd70} /* (14, 19, 7) {real, imag} */,
  {32'hc1675cca, 32'h4198c5a4} /* (14, 19, 6) {real, imag} */,
  {32'hc1892253, 32'h40896ad0} /* (14, 19, 5) {real, imag} */,
  {32'h4053c1f5, 32'h40b7be22} /* (14, 19, 4) {real, imag} */,
  {32'h3ff4d69e, 32'h40bbfe9a} /* (14, 19, 3) {real, imag} */,
  {32'hbff3304a, 32'hc0e9b071} /* (14, 19, 2) {real, imag} */,
  {32'h3c52d700, 32'h412e2e74} /* (14, 19, 1) {real, imag} */,
  {32'hc1846821, 32'hc0f289fa} /* (14, 19, 0) {real, imag} */,
  {32'hbf408828, 32'h413d712e} /* (14, 18, 31) {real, imag} */,
  {32'hc12e7ff9, 32'hc19a24c6} /* (14, 18, 30) {real, imag} */,
  {32'h41296f4a, 32'h403f4790} /* (14, 18, 29) {real, imag} */,
  {32'hc0870ba9, 32'h404f86c6} /* (14, 18, 28) {real, imag} */,
  {32'hc043c230, 32'h40d2649e} /* (14, 18, 27) {real, imag} */,
  {32'h41261c82, 32'hc146b524} /* (14, 18, 26) {real, imag} */,
  {32'hc139afc6, 32'h3f53f450} /* (14, 18, 25) {real, imag} */,
  {32'hc0c81cf9, 32'h41258db0} /* (14, 18, 24) {real, imag} */,
  {32'hc10e67cd, 32'h401d5d0c} /* (14, 18, 23) {real, imag} */,
  {32'h41b8424a, 32'h4109969e} /* (14, 18, 22) {real, imag} */,
  {32'h412dd80a, 32'h4119cafa} /* (14, 18, 21) {real, imag} */,
  {32'h411af5d1, 32'h401286ac} /* (14, 18, 20) {real, imag} */,
  {32'h409ef2a2, 32'h4188ca88} /* (14, 18, 19) {real, imag} */,
  {32'h417f1194, 32'h3fbd0df8} /* (14, 18, 18) {real, imag} */,
  {32'h4115d91b, 32'hbf2b82e0} /* (14, 18, 17) {real, imag} */,
  {32'h3fddbe32, 32'hc015ec8c} /* (14, 18, 16) {real, imag} */,
  {32'h41d50c56, 32'hc0a1e6bc} /* (14, 18, 15) {real, imag} */,
  {32'h419a3c40, 32'hc1072e9e} /* (14, 18, 14) {real, imag} */,
  {32'hc00bcdf0, 32'hc13705a2} /* (14, 18, 13) {real, imag} */,
  {32'h4077ff15, 32'hc0e6a297} /* (14, 18, 12) {real, imag} */,
  {32'h404d408e, 32'h41029b12} /* (14, 18, 11) {real, imag} */,
  {32'hc17181a8, 32'h407bab6e} /* (14, 18, 10) {real, imag} */,
  {32'hc062104e, 32'h4150b406} /* (14, 18, 9) {real, imag} */,
  {32'hc1552756, 32'h40cd9b58} /* (14, 18, 8) {real, imag} */,
  {32'hc0d6ff30, 32'h412b995e} /* (14, 18, 7) {real, imag} */,
  {32'h41b8f986, 32'hbfe978b1} /* (14, 18, 6) {real, imag} */,
  {32'hc00f7a2e, 32'h413b15d4} /* (14, 18, 5) {real, imag} */,
  {32'h40b1745c, 32'hc10f3ab9} /* (14, 18, 4) {real, imag} */,
  {32'hbfed6c8a, 32'hc0585e70} /* (14, 18, 3) {real, imag} */,
  {32'hc0c16bf7, 32'h3ea9f5f8} /* (14, 18, 2) {real, imag} */,
  {32'hc0f3e3a1, 32'h41297002} /* (14, 18, 1) {real, imag} */,
  {32'hbfb20d0c, 32'h40566b82} /* (14, 18, 0) {real, imag} */,
  {32'h40a25ee0, 32'hc0e5b531} /* (14, 17, 31) {real, imag} */,
  {32'hbfc8ffee, 32'h3fecc0c0} /* (14, 17, 30) {real, imag} */,
  {32'h4155405b, 32'hc08b2d48} /* (14, 17, 29) {real, imag} */,
  {32'hbfd3dc0a, 32'h4081c56d} /* (14, 17, 28) {real, imag} */,
  {32'hc0ec9e2c, 32'h411cbcd4} /* (14, 17, 27) {real, imag} */,
  {32'hc0893268, 32'hc0d566c8} /* (14, 17, 26) {real, imag} */,
  {32'hbf14fe98, 32'hc0af02a1} /* (14, 17, 25) {real, imag} */,
  {32'h415c1589, 32'hc070f942} /* (14, 17, 24) {real, imag} */,
  {32'h4136a390, 32'hc0fd3f63} /* (14, 17, 23) {real, imag} */,
  {32'h409f2fe8, 32'h40129914} /* (14, 17, 22) {real, imag} */,
  {32'hbdbf4ec0, 32'hc0604242} /* (14, 17, 21) {real, imag} */,
  {32'h3f632658, 32'h412dbed0} /* (14, 17, 20) {real, imag} */,
  {32'h3ef26280, 32'h3fcdb3d0} /* (14, 17, 19) {real, imag} */,
  {32'hc04719b6, 32'h411d8547} /* (14, 17, 18) {real, imag} */,
  {32'hc053e797, 32'h3f821152} /* (14, 17, 17) {real, imag} */,
  {32'h3e863834, 32'h411e5da7} /* (14, 17, 16) {real, imag} */,
  {32'h3ea32620, 32'h41324c42} /* (14, 17, 15) {real, imag} */,
  {32'hc0f88386, 32'h3fe6e62c} /* (14, 17, 14) {real, imag} */,
  {32'hc1727710, 32'h4080cd18} /* (14, 17, 13) {real, imag} */,
  {32'hc0beaf50, 32'hbff90bd0} /* (14, 17, 12) {real, imag} */,
  {32'h40b38b8a, 32'hc1455026} /* (14, 17, 11) {real, imag} */,
  {32'h41037e0b, 32'hc05314e5} /* (14, 17, 10) {real, imag} */,
  {32'hc041941c, 32'hbf2176b0} /* (14, 17, 9) {real, imag} */,
  {32'hbf533504, 32'h413a0931} /* (14, 17, 8) {real, imag} */,
  {32'hc0bbf4e1, 32'h40381332} /* (14, 17, 7) {real, imag} */,
  {32'hc10fadc1, 32'h41599cc6} /* (14, 17, 6) {real, imag} */,
  {32'hc05ce9c6, 32'hc037ac25} /* (14, 17, 5) {real, imag} */,
  {32'hbfef5589, 32'hc138e043} /* (14, 17, 4) {real, imag} */,
  {32'h4105718e, 32'hc10b85cb} /* (14, 17, 3) {real, imag} */,
  {32'hc0554486, 32'hbfdef4d0} /* (14, 17, 2) {real, imag} */,
  {32'h405d73f4, 32'hc0a3013e} /* (14, 17, 1) {real, imag} */,
  {32'hc1265459, 32'hc0c861aa} /* (14, 17, 0) {real, imag} */,
  {32'h401825b8, 32'h405e34c7} /* (14, 16, 31) {real, imag} */,
  {32'hc1157375, 32'hc0568c54} /* (14, 16, 30) {real, imag} */,
  {32'hc0d670b2, 32'hbfc1e020} /* (14, 16, 29) {real, imag} */,
  {32'h40db552e, 32'h40dd02f8} /* (14, 16, 28) {real, imag} */,
  {32'h3f94c8e1, 32'h4054dc5a} /* (14, 16, 27) {real, imag} */,
  {32'hc001aa3d, 32'h4082d6d8} /* (14, 16, 26) {real, imag} */,
  {32'h4035329d, 32'hbfc867c0} /* (14, 16, 25) {real, imag} */,
  {32'hc04f12f6, 32'hbfc91dfc} /* (14, 16, 24) {real, imag} */,
  {32'h3faa85ad, 32'hbfa68b9c} /* (14, 16, 23) {real, imag} */,
  {32'h40ff0d25, 32'h416018b0} /* (14, 16, 22) {real, imag} */,
  {32'h40b54561, 32'hc147adcf} /* (14, 16, 21) {real, imag} */,
  {32'hc09039f0, 32'hc02fbb12} /* (14, 16, 20) {real, imag} */,
  {32'hc10a03c6, 32'h41058d41} /* (14, 16, 19) {real, imag} */,
  {32'h3f196eec, 32'hc086b67c} /* (14, 16, 18) {real, imag} */,
  {32'hc09f3ff2, 32'hc1214de1} /* (14, 16, 17) {real, imag} */,
  {32'hc0f68552, 32'h00000000} /* (14, 16, 16) {real, imag} */,
  {32'hc09f3ff2, 32'h41214de1} /* (14, 16, 15) {real, imag} */,
  {32'h3f196eec, 32'h4086b67c} /* (14, 16, 14) {real, imag} */,
  {32'hc10a03c6, 32'hc1058d41} /* (14, 16, 13) {real, imag} */,
  {32'hc09039f0, 32'h402fbb12} /* (14, 16, 12) {real, imag} */,
  {32'h40b54561, 32'h4147adcf} /* (14, 16, 11) {real, imag} */,
  {32'h40ff0d25, 32'hc16018b0} /* (14, 16, 10) {real, imag} */,
  {32'h3faa85ad, 32'h3fa68b9c} /* (14, 16, 9) {real, imag} */,
  {32'hc04f12f6, 32'h3fc91dfc} /* (14, 16, 8) {real, imag} */,
  {32'h4035329d, 32'h3fc867c0} /* (14, 16, 7) {real, imag} */,
  {32'hc001aa3d, 32'hc082d6d8} /* (14, 16, 6) {real, imag} */,
  {32'h3f94c8e1, 32'hc054dc5a} /* (14, 16, 5) {real, imag} */,
  {32'h40db552e, 32'hc0dd02f8} /* (14, 16, 4) {real, imag} */,
  {32'hc0d670b2, 32'h3fc1e020} /* (14, 16, 3) {real, imag} */,
  {32'hc1157375, 32'h40568c54} /* (14, 16, 2) {real, imag} */,
  {32'h401825b8, 32'hc05e34c7} /* (14, 16, 1) {real, imag} */,
  {32'h40e99a4c, 32'h00000000} /* (14, 16, 0) {real, imag} */,
  {32'h405d73f4, 32'h40a3013e} /* (14, 15, 31) {real, imag} */,
  {32'hc0554486, 32'h3fdef4d0} /* (14, 15, 30) {real, imag} */,
  {32'h4105718e, 32'h410b85cb} /* (14, 15, 29) {real, imag} */,
  {32'hbfef5589, 32'h4138e043} /* (14, 15, 28) {real, imag} */,
  {32'hc05ce9c6, 32'h4037ac25} /* (14, 15, 27) {real, imag} */,
  {32'hc10fadc1, 32'hc1599cc6} /* (14, 15, 26) {real, imag} */,
  {32'hc0bbf4e1, 32'hc0381332} /* (14, 15, 25) {real, imag} */,
  {32'hbf533504, 32'hc13a0931} /* (14, 15, 24) {real, imag} */,
  {32'hc041941c, 32'h3f2176b0} /* (14, 15, 23) {real, imag} */,
  {32'h41037e0b, 32'h405314e5} /* (14, 15, 22) {real, imag} */,
  {32'h40b38b8a, 32'h41455026} /* (14, 15, 21) {real, imag} */,
  {32'hc0beaf50, 32'h3ff90bd0} /* (14, 15, 20) {real, imag} */,
  {32'hc1727710, 32'hc080cd18} /* (14, 15, 19) {real, imag} */,
  {32'hc0f88386, 32'hbfe6e62c} /* (14, 15, 18) {real, imag} */,
  {32'h3ea32620, 32'hc1324c42} /* (14, 15, 17) {real, imag} */,
  {32'h3e863834, 32'hc11e5da7} /* (14, 15, 16) {real, imag} */,
  {32'hc053e797, 32'hbf821152} /* (14, 15, 15) {real, imag} */,
  {32'hc04719b6, 32'hc11d8547} /* (14, 15, 14) {real, imag} */,
  {32'h3ef26280, 32'hbfcdb3d0} /* (14, 15, 13) {real, imag} */,
  {32'h3f632658, 32'hc12dbed0} /* (14, 15, 12) {real, imag} */,
  {32'hbdbf4ec0, 32'h40604242} /* (14, 15, 11) {real, imag} */,
  {32'h409f2fe8, 32'hc0129914} /* (14, 15, 10) {real, imag} */,
  {32'h4136a390, 32'h40fd3f63} /* (14, 15, 9) {real, imag} */,
  {32'h415c1589, 32'h4070f942} /* (14, 15, 8) {real, imag} */,
  {32'hbf14fe98, 32'h40af02a1} /* (14, 15, 7) {real, imag} */,
  {32'hc0893268, 32'h40d566c8} /* (14, 15, 6) {real, imag} */,
  {32'hc0ec9e2c, 32'hc11cbcd4} /* (14, 15, 5) {real, imag} */,
  {32'hbfd3dc0a, 32'hc081c56d} /* (14, 15, 4) {real, imag} */,
  {32'h4155405b, 32'h408b2d48} /* (14, 15, 3) {real, imag} */,
  {32'hbfc8ffee, 32'hbfecc0c0} /* (14, 15, 2) {real, imag} */,
  {32'h40a25ee0, 32'h40e5b531} /* (14, 15, 1) {real, imag} */,
  {32'hc1265459, 32'h40c861aa} /* (14, 15, 0) {real, imag} */,
  {32'hc0f3e3a1, 32'hc1297002} /* (14, 14, 31) {real, imag} */,
  {32'hc0c16bf7, 32'hbea9f5f8} /* (14, 14, 30) {real, imag} */,
  {32'hbfed6c8a, 32'h40585e70} /* (14, 14, 29) {real, imag} */,
  {32'h40b1745c, 32'h410f3ab9} /* (14, 14, 28) {real, imag} */,
  {32'hc00f7a2e, 32'hc13b15d4} /* (14, 14, 27) {real, imag} */,
  {32'h41b8f986, 32'h3fe978b1} /* (14, 14, 26) {real, imag} */,
  {32'hc0d6ff30, 32'hc12b995e} /* (14, 14, 25) {real, imag} */,
  {32'hc1552756, 32'hc0cd9b58} /* (14, 14, 24) {real, imag} */,
  {32'hc062104e, 32'hc150b406} /* (14, 14, 23) {real, imag} */,
  {32'hc17181a8, 32'hc07bab6e} /* (14, 14, 22) {real, imag} */,
  {32'h404d408e, 32'hc1029b12} /* (14, 14, 21) {real, imag} */,
  {32'h4077ff15, 32'h40e6a297} /* (14, 14, 20) {real, imag} */,
  {32'hc00bcdf0, 32'h413705a2} /* (14, 14, 19) {real, imag} */,
  {32'h419a3c40, 32'h41072e9e} /* (14, 14, 18) {real, imag} */,
  {32'h41d50c56, 32'h40a1e6bc} /* (14, 14, 17) {real, imag} */,
  {32'h3fddbe32, 32'h4015ec8c} /* (14, 14, 16) {real, imag} */,
  {32'h4115d91b, 32'h3f2b82e0} /* (14, 14, 15) {real, imag} */,
  {32'h417f1194, 32'hbfbd0df8} /* (14, 14, 14) {real, imag} */,
  {32'h409ef2a2, 32'hc188ca88} /* (14, 14, 13) {real, imag} */,
  {32'h411af5d1, 32'hc01286ac} /* (14, 14, 12) {real, imag} */,
  {32'h412dd80a, 32'hc119cafa} /* (14, 14, 11) {real, imag} */,
  {32'h41b8424a, 32'hc109969e} /* (14, 14, 10) {real, imag} */,
  {32'hc10e67cd, 32'hc01d5d0c} /* (14, 14, 9) {real, imag} */,
  {32'hc0c81cf9, 32'hc1258db0} /* (14, 14, 8) {real, imag} */,
  {32'hc139afc6, 32'hbf53f450} /* (14, 14, 7) {real, imag} */,
  {32'h41261c82, 32'h4146b524} /* (14, 14, 6) {real, imag} */,
  {32'hc043c230, 32'hc0d2649e} /* (14, 14, 5) {real, imag} */,
  {32'hc0870ba9, 32'hc04f86c6} /* (14, 14, 4) {real, imag} */,
  {32'h41296f4a, 32'hc03f4790} /* (14, 14, 3) {real, imag} */,
  {32'hc12e7ff9, 32'h419a24c6} /* (14, 14, 2) {real, imag} */,
  {32'hbf408828, 32'hc13d712e} /* (14, 14, 1) {real, imag} */,
  {32'hbfb20d0c, 32'hc0566b82} /* (14, 14, 0) {real, imag} */,
  {32'h3c52d700, 32'hc12e2e74} /* (14, 13, 31) {real, imag} */,
  {32'hbff3304a, 32'h40e9b071} /* (14, 13, 30) {real, imag} */,
  {32'h3ff4d69e, 32'hc0bbfe9a} /* (14, 13, 29) {real, imag} */,
  {32'h4053c1f5, 32'hc0b7be22} /* (14, 13, 28) {real, imag} */,
  {32'hc1892253, 32'hc0896ad0} /* (14, 13, 27) {real, imag} */,
  {32'hc1675cca, 32'hc198c5a4} /* (14, 13, 26) {real, imag} */,
  {32'h414c208f, 32'h3f2edd70} /* (14, 13, 25) {real, imag} */,
  {32'hc010cd97, 32'h3e1dace0} /* (14, 13, 24) {real, imag} */,
  {32'hc0e248c9, 32'h41094285} /* (14, 13, 23) {real, imag} */,
  {32'hc0813e79, 32'h40dce3de} /* (14, 13, 22) {real, imag} */,
  {32'h406dafc9, 32'h406580c8} /* (14, 13, 21) {real, imag} */,
  {32'h415fb897, 32'hc17ab5b4} /* (14, 13, 20) {real, imag} */,
  {32'hc169dcd9, 32'hc0ec664a} /* (14, 13, 19) {real, imag} */,
  {32'hc1863cd1, 32'hc127723e} /* (14, 13, 18) {real, imag} */,
  {32'h40187ce6, 32'h40ec2d28} /* (14, 13, 17) {real, imag} */,
  {32'h4058d8ac, 32'h409ae742} /* (14, 13, 16) {real, imag} */,
  {32'hc1c5d546, 32'h408c5787} /* (14, 13, 15) {real, imag} */,
  {32'h417e3368, 32'hc1025e56} /* (14, 13, 14) {real, imag} */,
  {32'h3efd4a70, 32'h40a59fc9} /* (14, 13, 13) {real, imag} */,
  {32'hbf6edd6c, 32'h41861bb1} /* (14, 13, 12) {real, imag} */,
  {32'hbfb345d0, 32'hc12ad11c} /* (14, 13, 11) {real, imag} */,
  {32'h40dd079c, 32'hc080f852} /* (14, 13, 10) {real, imag} */,
  {32'hc0c296f8, 32'h409212bc} /* (14, 13, 9) {real, imag} */,
  {32'hc09f361f, 32'h40bad620} /* (14, 13, 8) {real, imag} */,
  {32'hbfc4980c, 32'hbfe5c6ac} /* (14, 13, 7) {real, imag} */,
  {32'h40d64742, 32'hc0ea1520} /* (14, 13, 6) {real, imag} */,
  {32'hc04bd2c4, 32'h411a3d0f} /* (14, 13, 5) {real, imag} */,
  {32'hc0cff28f, 32'h3fdb15a0} /* (14, 13, 4) {real, imag} */,
  {32'h3d55cbe0, 32'h40ec8c86} /* (14, 13, 3) {real, imag} */,
  {32'h40b1d12c, 32'h40ea931b} /* (14, 13, 2) {real, imag} */,
  {32'h41050d3c, 32'h414bedda} /* (14, 13, 1) {real, imag} */,
  {32'hc1846821, 32'h40f289fa} /* (14, 13, 0) {real, imag} */,
  {32'hc0e4bf90, 32'h3fb0e358} /* (14, 12, 31) {real, imag} */,
  {32'h4091835f, 32'h4194468e} /* (14, 12, 30) {real, imag} */,
  {32'h3f6dff10, 32'hc057e6ee} /* (14, 12, 29) {real, imag} */,
  {32'h4034dfe9, 32'hc10d1f42} /* (14, 12, 28) {real, imag} */,
  {32'h3fec36fe, 32'hc147e1b3} /* (14, 12, 27) {real, imag} */,
  {32'hc114b019, 32'h40816204} /* (14, 12, 26) {real, imag} */,
  {32'h3f9cfaae, 32'hc11ec116} /* (14, 12, 25) {real, imag} */,
  {32'h414091b1, 32'h40ebd58c} /* (14, 12, 24) {real, imag} */,
  {32'hc0fbe71f, 32'h408b31d6} /* (14, 12, 23) {real, imag} */,
  {32'h4102973a, 32'hbfd213bc} /* (14, 12, 22) {real, imag} */,
  {32'h40eb8024, 32'hc0d726a7} /* (14, 12, 21) {real, imag} */,
  {32'hc16ac9f4, 32'h402d35da} /* (14, 12, 20) {real, imag} */,
  {32'h411e32d6, 32'h417d7a7e} /* (14, 12, 19) {real, imag} */,
  {32'hc06ef3c0, 32'hc10befa5} /* (14, 12, 18) {real, imag} */,
  {32'hc11fa2d2, 32'hbf41ef8e} /* (14, 12, 17) {real, imag} */,
  {32'hbfc3a4ec, 32'hc03d1d18} /* (14, 12, 16) {real, imag} */,
  {32'hc1424eaf, 32'hc015fac4} /* (14, 12, 15) {real, imag} */,
  {32'hc0ad15f8, 32'hc023df9a} /* (14, 12, 14) {real, imag} */,
  {32'hbe450088, 32'hc0d84515} /* (14, 12, 13) {real, imag} */,
  {32'hc13c2880, 32'hc0fdaffe} /* (14, 12, 12) {real, imag} */,
  {32'hc1177a16, 32'h406ecae2} /* (14, 12, 11) {real, imag} */,
  {32'hc0a2390f, 32'h40b94af9} /* (14, 12, 10) {real, imag} */,
  {32'hc10fed94, 32'h419568eb} /* (14, 12, 9) {real, imag} */,
  {32'hc12bab96, 32'hc11a2f5c} /* (14, 12, 8) {real, imag} */,
  {32'h41509ac1, 32'h3fcc4e50} /* (14, 12, 7) {real, imag} */,
  {32'h4071a94f, 32'hc13914c1} /* (14, 12, 6) {real, imag} */,
  {32'hc0919b36, 32'h3f91d10d} /* (14, 12, 5) {real, imag} */,
  {32'h4146ac00, 32'hc0b3d437} /* (14, 12, 4) {real, imag} */,
  {32'hc068c3eb, 32'h4125ac4a} /* (14, 12, 3) {real, imag} */,
  {32'h4085882c, 32'h3f5641f0} /* (14, 12, 2) {real, imag} */,
  {32'h4180fceb, 32'h404c4d48} /* (14, 12, 1) {real, imag} */,
  {32'h4150862e, 32'hc0a4bb46} /* (14, 12, 0) {real, imag} */,
  {32'hc1c43bc0, 32'hc06ad3be} /* (14, 11, 31) {real, imag} */,
  {32'hc030a0e4, 32'h4198fa90} /* (14, 11, 30) {real, imag} */,
  {32'hc18ca28e, 32'h3f78ba58} /* (14, 11, 29) {real, imag} */,
  {32'hbf7deb44, 32'h410658b2} /* (14, 11, 28) {real, imag} */,
  {32'h41c4d613, 32'h418eda24} /* (14, 11, 27) {real, imag} */,
  {32'hc011eb64, 32'hc0b10b6b} /* (14, 11, 26) {real, imag} */,
  {32'h411027f2, 32'hc161efce} /* (14, 11, 25) {real, imag} */,
  {32'h41544e2f, 32'hc18e26d8} /* (14, 11, 24) {real, imag} */,
  {32'h416d133e, 32'hc165aad3} /* (14, 11, 23) {real, imag} */,
  {32'hbeffe100, 32'hc0a2f092} /* (14, 11, 22) {real, imag} */,
  {32'h41330e8a, 32'h41b9a82d} /* (14, 11, 21) {real, imag} */,
  {32'hc0b52ea2, 32'h40971131} /* (14, 11, 20) {real, imag} */,
  {32'hc1818b8d, 32'h4109ce17} /* (14, 11, 19) {real, imag} */,
  {32'h40586fe5, 32'hbf10166e} /* (14, 11, 18) {real, imag} */,
  {32'hc0bf3d1a, 32'h400ee391} /* (14, 11, 17) {real, imag} */,
  {32'hc17ab361, 32'hbfc0e98a} /* (14, 11, 16) {real, imag} */,
  {32'h4104cf07, 32'h3fe8e494} /* (14, 11, 15) {real, imag} */,
  {32'h41790ef0, 32'h4162ec17} /* (14, 11, 14) {real, imag} */,
  {32'h416a0856, 32'hc00f1dea} /* (14, 11, 13) {real, imag} */,
  {32'h40f03928, 32'hc05ddc29} /* (14, 11, 12) {real, imag} */,
  {32'hc0daef2a, 32'hc16d6f43} /* (14, 11, 11) {real, imag} */,
  {32'h4079b8a2, 32'hc1b622c2} /* (14, 11, 10) {real, imag} */,
  {32'hc0aaeb46, 32'hbf600658} /* (14, 11, 9) {real, imag} */,
  {32'h4045fc20, 32'h409d54b8} /* (14, 11, 8) {real, imag} */,
  {32'h415775a8, 32'h417afa1b} /* (14, 11, 7) {real, imag} */,
  {32'h4182d79c, 32'h415c5786} /* (14, 11, 6) {real, imag} */,
  {32'hc09754a3, 32'h40e42ca6} /* (14, 11, 5) {real, imag} */,
  {32'h3ffbaf97, 32'hc1104fba} /* (14, 11, 4) {real, imag} */,
  {32'hc09daa61, 32'h410076b6} /* (14, 11, 3) {real, imag} */,
  {32'hc0145138, 32'h4155eb35} /* (14, 11, 2) {real, imag} */,
  {32'h3f2b12da, 32'hc1fbaf2a} /* (14, 11, 1) {real, imag} */,
  {32'hc1906db5, 32'hc1f66e78} /* (14, 11, 0) {real, imag} */,
  {32'hc092e34a, 32'h410f28c3} /* (14, 10, 31) {real, imag} */,
  {32'h40579e20, 32'hc1b0250c} /* (14, 10, 30) {real, imag} */,
  {32'hc02e4d7a, 32'h3f360260} /* (14, 10, 29) {real, imag} */,
  {32'hc1aa1715, 32'h409f50f4} /* (14, 10, 28) {real, imag} */,
  {32'hc101bdd8, 32'hc0dd8994} /* (14, 10, 27) {real, imag} */,
  {32'h41b985d9, 32'h409a9b70} /* (14, 10, 26) {real, imag} */,
  {32'h41aea7ae, 32'h41c2a69e} /* (14, 10, 25) {real, imag} */,
  {32'hc12a9ed4, 32'h411acb56} /* (14, 10, 24) {real, imag} */,
  {32'h41155a53, 32'h41bc4af6} /* (14, 10, 23) {real, imag} */,
  {32'h3f76f910, 32'h407cdb92} /* (14, 10, 22) {real, imag} */,
  {32'h408b2ac3, 32'hc1669055} /* (14, 10, 21) {real, imag} */,
  {32'hbdd116e0, 32'hc122dc9c} /* (14, 10, 20) {real, imag} */,
  {32'hc0e0b663, 32'h40256ee2} /* (14, 10, 19) {real, imag} */,
  {32'h4081dda2, 32'hc001bd8e} /* (14, 10, 18) {real, imag} */,
  {32'h40a48a77, 32'hc1a5e7c5} /* (14, 10, 17) {real, imag} */,
  {32'hc102234b, 32'hc1190e8d} /* (14, 10, 16) {real, imag} */,
  {32'hc18e4ea6, 32'h4151fe88} /* (14, 10, 15) {real, imag} */,
  {32'h3fe63f28, 32'h40b8e038} /* (14, 10, 14) {real, imag} */,
  {32'hc0625868, 32'hc1645687} /* (14, 10, 13) {real, imag} */,
  {32'h3eea5ca0, 32'h41339646} /* (14, 10, 12) {real, imag} */,
  {32'h41948a6d, 32'hc01fa698} /* (14, 10, 11) {real, imag} */,
  {32'h40270212, 32'hc1686cb2} /* (14, 10, 10) {real, imag} */,
  {32'h4082e1b3, 32'hc184af94} /* (14, 10, 9) {real, imag} */,
  {32'hbffb5fc8, 32'hbfbef619} /* (14, 10, 8) {real, imag} */,
  {32'h41236ee6, 32'h4033e555} /* (14, 10, 7) {real, imag} */,
  {32'h410955ea, 32'h3ff669ec} /* (14, 10, 6) {real, imag} */,
  {32'h4178faf0, 32'hbda17f00} /* (14, 10, 5) {real, imag} */,
  {32'hbf94d510, 32'hc19810cc} /* (14, 10, 4) {real, imag} */,
  {32'hc0894436, 32'h40997633} /* (14, 10, 3) {real, imag} */,
  {32'hc0b89566, 32'hbf88d198} /* (14, 10, 2) {real, imag} */,
  {32'h41e70a46, 32'h408f2d3b} /* (14, 10, 1) {real, imag} */,
  {32'h41229090, 32'h41cefe2b} /* (14, 10, 0) {real, imag} */,
  {32'hc0a59db5, 32'h4185d1b4} /* (14, 9, 31) {real, imag} */,
  {32'hc017aa20, 32'hc16eec56} /* (14, 9, 30) {real, imag} */,
  {32'h41009193, 32'h406a286f} /* (14, 9, 29) {real, imag} */,
  {32'h414414a9, 32'h40dfa954} /* (14, 9, 28) {real, imag} */,
  {32'hc1a61ebf, 32'hc138b3c8} /* (14, 9, 27) {real, imag} */,
  {32'h41033108, 32'hc0445c80} /* (14, 9, 26) {real, imag} */,
  {32'h41cc817f, 32'h41163ba8} /* (14, 9, 25) {real, imag} */,
  {32'h40c9773a, 32'hc11ecf6c} /* (14, 9, 24) {real, imag} */,
  {32'hc103d0fb, 32'hc038e3e4} /* (14, 9, 23) {real, imag} */,
  {32'hc1391550, 32'h40fa17ce} /* (14, 9, 22) {real, imag} */,
  {32'hc1b61464, 32'h4126f738} /* (14, 9, 21) {real, imag} */,
  {32'hc04f694a, 32'h3edb8520} /* (14, 9, 20) {real, imag} */,
  {32'h41915c1c, 32'hc15e164f} /* (14, 9, 19) {real, imag} */,
  {32'h41aa6e97, 32'hc1972b7f} /* (14, 9, 18) {real, imag} */,
  {32'hc127d911, 32'hc0ea68e0} /* (14, 9, 17) {real, imag} */,
  {32'hc09735ab, 32'h402e30ec} /* (14, 9, 16) {real, imag} */,
  {32'hbf800f72, 32'hc186e588} /* (14, 9, 15) {real, imag} */,
  {32'hc1231163, 32'h3f7c4b64} /* (14, 9, 14) {real, imag} */,
  {32'h40cd795c, 32'hc1180da8} /* (14, 9, 13) {real, imag} */,
  {32'hc1141b13, 32'hc0c1febe} /* (14, 9, 12) {real, imag} */,
  {32'hc111e473, 32'h414988be} /* (14, 9, 11) {real, imag} */,
  {32'hc080633b, 32'h416fc54c} /* (14, 9, 10) {real, imag} */,
  {32'h40da1cc1, 32'hc00b4bec} /* (14, 9, 9) {real, imag} */,
  {32'hc158d8f3, 32'h4147ad17} /* (14, 9, 8) {real, imag} */,
  {32'hc1b582ae, 32'h4111940a} /* (14, 9, 7) {real, imag} */,
  {32'hc0a1a11a, 32'hc19afbba} /* (14, 9, 6) {real, imag} */,
  {32'h413dc41b, 32'hc13ab2c3} /* (14, 9, 5) {real, imag} */,
  {32'hc0bb1f17, 32'h41499d1d} /* (14, 9, 4) {real, imag} */,
  {32'hc0f27797, 32'h411d50a5} /* (14, 9, 3) {real, imag} */,
  {32'h4096cdaf, 32'hc0d7fdf8} /* (14, 9, 2) {real, imag} */,
  {32'h3f9144c0, 32'hbff2ffb8} /* (14, 9, 1) {real, imag} */,
  {32'h40ef8717, 32'h40b4ceba} /* (14, 9, 0) {real, imag} */,
  {32'hc28b4cde, 32'hc21379d5} /* (14, 8, 31) {real, imag} */,
  {32'h41aeaa56, 32'h41998e3b} /* (14, 8, 30) {real, imag} */,
  {32'h413f9e15, 32'hc0ef409a} /* (14, 8, 29) {real, imag} */,
  {32'hc1393fa0, 32'h411ca426} /* (14, 8, 28) {real, imag} */,
  {32'h41c04486, 32'hbf86343a} /* (14, 8, 27) {real, imag} */,
  {32'h4161e62d, 32'h3fa7a084} /* (14, 8, 26) {real, imag} */,
  {32'h414d44c3, 32'h408da6a8} /* (14, 8, 25) {real, imag} */,
  {32'h3e0a84e8, 32'hc0cb9b90} /* (14, 8, 24) {real, imag} */,
  {32'hc03e9ce8, 32'hc1526e8f} /* (14, 8, 23) {real, imag} */,
  {32'h40b0e129, 32'hc191a2dc} /* (14, 8, 22) {real, imag} */,
  {32'h4150918c, 32'hbf44b998} /* (14, 8, 21) {real, imag} */,
  {32'hc14012a8, 32'h40b3907d} /* (14, 8, 20) {real, imag} */,
  {32'h405579c4, 32'h41286238} /* (14, 8, 19) {real, imag} */,
  {32'h3f31ff88, 32'hbfa6cf1c} /* (14, 8, 18) {real, imag} */,
  {32'hc086c192, 32'h412a9510} /* (14, 8, 17) {real, imag} */,
  {32'hc0db26aa, 32'h40d3c248} /* (14, 8, 16) {real, imag} */,
  {32'hc1194266, 32'hc17160dd} /* (14, 8, 15) {real, imag} */,
  {32'h4099a760, 32'h409b7eae} /* (14, 8, 14) {real, imag} */,
  {32'hbf2c4510, 32'hc0bc17f3} /* (14, 8, 13) {real, imag} */,
  {32'hc13784c2, 32'hc1350657} /* (14, 8, 12) {real, imag} */,
  {32'h4190ff78, 32'hc0ec41ea} /* (14, 8, 11) {real, imag} */,
  {32'hc1e3d422, 32'h40c6dfd0} /* (14, 8, 10) {real, imag} */,
  {32'hc0cf55fd, 32'h4044726f} /* (14, 8, 9) {real, imag} */,
  {32'hbf2db8c0, 32'h3e0b3bc0} /* (14, 8, 8) {real, imag} */,
  {32'h4108f3c7, 32'h40c6f734} /* (14, 8, 7) {real, imag} */,
  {32'h401923af, 32'h3fb254ec} /* (14, 8, 6) {real, imag} */,
  {32'hbfff0ef6, 32'h41c88ef6} /* (14, 8, 5) {real, imag} */,
  {32'hc1cc9cd6, 32'h40087159} /* (14, 8, 4) {real, imag} */,
  {32'hc0b0765f, 32'h40c1c104} /* (14, 8, 3) {real, imag} */,
  {32'h41b65f51, 32'h406e5a60} /* (14, 8, 2) {real, imag} */,
  {32'hc1aea470, 32'hc20a9226} /* (14, 8, 1) {real, imag} */,
  {32'hc1ba0d4e, 32'hc0e4e9e6} /* (14, 8, 0) {real, imag} */,
  {32'h41e64b91, 32'hc1a8ec68} /* (14, 7, 31) {real, imag} */,
  {32'hc0a10d46, 32'hc1ea0730} /* (14, 7, 30) {real, imag} */,
  {32'h40765ea0, 32'hc080ace5} /* (14, 7, 29) {real, imag} */,
  {32'hc10eef98, 32'hc1259c4d} /* (14, 7, 28) {real, imag} */,
  {32'hc187d4d8, 32'h41ebc854} /* (14, 7, 27) {real, imag} */,
  {32'hc1a8b55b, 32'hbfff4468} /* (14, 7, 26) {real, imag} */,
  {32'hc11c5816, 32'h4080fda0} /* (14, 7, 25) {real, imag} */,
  {32'hbf5ffd68, 32'hbfdb750a} /* (14, 7, 24) {real, imag} */,
  {32'hc10ee0e5, 32'h41059fef} /* (14, 7, 23) {real, imag} */,
  {32'h41084198, 32'h40470696} /* (14, 7, 22) {real, imag} */,
  {32'h412cba39, 32'hc0bc2ff9} /* (14, 7, 21) {real, imag} */,
  {32'h41b69b24, 32'hc1db02b9} /* (14, 7, 20) {real, imag} */,
  {32'h412b7bc6, 32'h4118d94d} /* (14, 7, 19) {real, imag} */,
  {32'hc08fd3ed, 32'hbff1fa00} /* (14, 7, 18) {real, imag} */,
  {32'h41204da6, 32'hbfa0e598} /* (14, 7, 17) {real, imag} */,
  {32'h4129d26c, 32'h41668c96} /* (14, 7, 16) {real, imag} */,
  {32'h4103890f, 32'h40a5e198} /* (14, 7, 15) {real, imag} */,
  {32'hc0a6c378, 32'h3e95b040} /* (14, 7, 14) {real, imag} */,
  {32'h3fcd5a2c, 32'h41c32e6d} /* (14, 7, 13) {real, imag} */,
  {32'hc18a9490, 32'h417f0658} /* (14, 7, 12) {real, imag} */,
  {32'hc09670a6, 32'h4085bc8b} /* (14, 7, 11) {real, imag} */,
  {32'hbfb37cac, 32'h41b3a45c} /* (14, 7, 10) {real, imag} */,
  {32'hc129c79b, 32'hc19a7a14} /* (14, 7, 9) {real, imag} */,
  {32'h4115c152, 32'hc1b0954c} /* (14, 7, 8) {real, imag} */,
  {32'hc0edb2b6, 32'hc15a94f4} /* (14, 7, 7) {real, imag} */,
  {32'h412bf63a, 32'hc12c81a8} /* (14, 7, 6) {real, imag} */,
  {32'hc109f044, 32'hc096c99a} /* (14, 7, 5) {real, imag} */,
  {32'hc1ee6cac, 32'h4184a701} /* (14, 7, 4) {real, imag} */,
  {32'hc088a118, 32'hc0ff7a2c} /* (14, 7, 3) {real, imag} */,
  {32'h40956b2c, 32'hc19833ce} /* (14, 7, 2) {real, imag} */,
  {32'hc0f51c4e, 32'h41e36c2e} /* (14, 7, 1) {real, imag} */,
  {32'hbff1350c, 32'h421d80aa} /* (14, 7, 0) {real, imag} */,
  {32'h412c37d9, 32'h4113cbb8} /* (14, 6, 31) {real, imag} */,
  {32'h41c93076, 32'h40a54934} /* (14, 6, 30) {real, imag} */,
  {32'hc20a773c, 32'hc1870b6e} /* (14, 6, 29) {real, imag} */,
  {32'hc14cac08, 32'hc103f7fe} /* (14, 6, 28) {real, imag} */,
  {32'hc114de72, 32'h40de7216} /* (14, 6, 27) {real, imag} */,
  {32'h40dabdea, 32'h41b663df} /* (14, 6, 26) {real, imag} */,
  {32'hc1a93a68, 32'hc1fe66ad} /* (14, 6, 25) {real, imag} */,
  {32'hc0077de8, 32'h410768ad} /* (14, 6, 24) {real, imag} */,
  {32'h40e789e5, 32'h41903725} /* (14, 6, 23) {real, imag} */,
  {32'hc0a93bda, 32'hc189bc72} /* (14, 6, 22) {real, imag} */,
  {32'hc088f2e9, 32'h411cdd25} /* (14, 6, 21) {real, imag} */,
  {32'hbfd8aac8, 32'h419249e2} /* (14, 6, 20) {real, imag} */,
  {32'h40d77f42, 32'hc1526a7a} /* (14, 6, 19) {real, imag} */,
  {32'h401cf1fa, 32'hc1198f25} /* (14, 6, 18) {real, imag} */,
  {32'hc02f6a21, 32'hc17e59a8} /* (14, 6, 17) {real, imag} */,
  {32'hbe4b79b8, 32'hbf626804} /* (14, 6, 16) {real, imag} */,
  {32'h4107bd8f, 32'h402e5980} /* (14, 6, 15) {real, imag} */,
  {32'hc15fa61c, 32'h3eae2298} /* (14, 6, 14) {real, imag} */,
  {32'h402955b4, 32'hc007b2a4} /* (14, 6, 13) {real, imag} */,
  {32'h40f73050, 32'hc0ca2770} /* (14, 6, 12) {real, imag} */,
  {32'h4150c398, 32'hc10f4176} /* (14, 6, 11) {real, imag} */,
  {32'h4191b883, 32'h3ffffbc2} /* (14, 6, 10) {real, imag} */,
  {32'hc12abd29, 32'h4100f859} /* (14, 6, 9) {real, imag} */,
  {32'h40dc6480, 32'h411f0860} /* (14, 6, 8) {real, imag} */,
  {32'hbf95af88, 32'hc123e626} /* (14, 6, 7) {real, imag} */,
  {32'hc14dae02, 32'h40870fd2} /* (14, 6, 6) {real, imag} */,
  {32'h3f4130a8, 32'hc1a68dfc} /* (14, 6, 5) {real, imag} */,
  {32'hc124bb72, 32'h40c1714b} /* (14, 6, 4) {real, imag} */,
  {32'h40903f6c, 32'h419dd5dc} /* (14, 6, 3) {real, imag} */,
  {32'h41e4a15d, 32'h4107f3d8} /* (14, 6, 2) {real, imag} */,
  {32'hc1650a4d, 32'hbe1fa320} /* (14, 6, 1) {real, imag} */,
  {32'hc1324388, 32'h4070aaa4} /* (14, 6, 0) {real, imag} */,
  {32'hc28a8fb9, 32'h42106b62} /* (14, 5, 31) {real, imag} */,
  {32'h40bf196c, 32'h4119df2d} /* (14, 5, 30) {real, imag} */,
  {32'hc11bf32b, 32'h41a13c4d} /* (14, 5, 29) {real, imag} */,
  {32'hc103166e, 32'hc0901be0} /* (14, 5, 28) {real, imag} */,
  {32'h41a12148, 32'hc1057d60} /* (14, 5, 27) {real, imag} */,
  {32'hc105c78e, 32'h40b95292} /* (14, 5, 26) {real, imag} */,
  {32'hc097b01e, 32'h4103c661} /* (14, 5, 25) {real, imag} */,
  {32'h408be2f0, 32'h3f8f8218} /* (14, 5, 24) {real, imag} */,
  {32'h402f7814, 32'hbfc058d5} /* (14, 5, 23) {real, imag} */,
  {32'hbe5edee0, 32'hbff3fd54} /* (14, 5, 22) {real, imag} */,
  {32'h410b0d2c, 32'hbf2a6d28} /* (14, 5, 21) {real, imag} */,
  {32'hc0ac88ba, 32'hbfde12dc} /* (14, 5, 20) {real, imag} */,
  {32'hbeda2e8a, 32'h4042ad0c} /* (14, 5, 19) {real, imag} */,
  {32'h41174fbe, 32'hc0e312c4} /* (14, 5, 18) {real, imag} */,
  {32'h409313db, 32'h4036a100} /* (14, 5, 17) {real, imag} */,
  {32'hbfd3ad4e, 32'hc088e3d4} /* (14, 5, 16) {real, imag} */,
  {32'h40db2fab, 32'hbfdb4002} /* (14, 5, 15) {real, imag} */,
  {32'h3e356860, 32'h417cd092} /* (14, 5, 14) {real, imag} */,
  {32'h413f3c45, 32'hc097a45a} /* (14, 5, 13) {real, imag} */,
  {32'hc121158d, 32'h40837c86} /* (14, 5, 12) {real, imag} */,
  {32'hbf816d0e, 32'hbf685bc0} /* (14, 5, 11) {real, imag} */,
  {32'h3ff25186, 32'h417725a7} /* (14, 5, 10) {real, imag} */,
  {32'h4007d2b4, 32'hc00eb2d8} /* (14, 5, 9) {real, imag} */,
  {32'hc16bae52, 32'h41467e9e} /* (14, 5, 8) {real, imag} */,
  {32'hc0d9279e, 32'h3ee41dd8} /* (14, 5, 7) {real, imag} */,
  {32'h4145672d, 32'hbf115b80} /* (14, 5, 6) {real, imag} */,
  {32'h415a6178, 32'h41ae6b49} /* (14, 5, 5) {real, imag} */,
  {32'h40f2bc27, 32'hc170e036} /* (14, 5, 4) {real, imag} */,
  {32'hc05c9e28, 32'h400d9280} /* (14, 5, 3) {real, imag} */,
  {32'hbd86c500, 32'h415e278c} /* (14, 5, 2) {real, imag} */,
  {32'hc2cd3d71, 32'hc1a48e40} /* (14, 5, 1) {real, imag} */,
  {32'hc282f9fd, 32'hc2203f75} /* (14, 5, 0) {real, imag} */,
  {32'h428f529d, 32'h41d443c0} /* (14, 4, 31) {real, imag} */,
  {32'hc24f7cae, 32'hc29f0bce} /* (14, 4, 30) {real, imag} */,
  {32'hc17d9df8, 32'hc1127616} /* (14, 4, 29) {real, imag} */,
  {32'h41d28d42, 32'h4231772c} /* (14, 4, 28) {real, imag} */,
  {32'hc1944570, 32'h41bfcf1e} /* (14, 4, 27) {real, imag} */,
  {32'hc04ecff4, 32'h4164c278} /* (14, 4, 26) {real, imag} */,
  {32'hc0fe5b74, 32'h420cc61a} /* (14, 4, 25) {real, imag} */,
  {32'hc141fbbe, 32'h40fe98f2} /* (14, 4, 24) {real, imag} */,
  {32'hc02f57e4, 32'hc1142478} /* (14, 4, 23) {real, imag} */,
  {32'hc0ba6203, 32'h40515d70} /* (14, 4, 22) {real, imag} */,
  {32'hc0f96f88, 32'h407a4d25} /* (14, 4, 21) {real, imag} */,
  {32'h3fc17eec, 32'h4066af62} /* (14, 4, 20) {real, imag} */,
  {32'hc15e1de1, 32'hc187f8f1} /* (14, 4, 19) {real, imag} */,
  {32'hc0cca6f4, 32'h405820bd} /* (14, 4, 18) {real, imag} */,
  {32'hc11c6e6b, 32'h41151f59} /* (14, 4, 17) {real, imag} */,
  {32'h4053392a, 32'hbea19e58} /* (14, 4, 16) {real, imag} */,
  {32'hbfda3196, 32'hc16ed944} /* (14, 4, 15) {real, imag} */,
  {32'hc0aec4c5, 32'hc1742284} /* (14, 4, 14) {real, imag} */,
  {32'hc0c545e5, 32'h409355fe} /* (14, 4, 13) {real, imag} */,
  {32'h3f67cb54, 32'hc05c865c} /* (14, 4, 12) {real, imag} */,
  {32'hc0f23ae4, 32'hc0638603} /* (14, 4, 11) {real, imag} */,
  {32'h411ff1de, 32'h41acefd6} /* (14, 4, 10) {real, imag} */,
  {32'h4215c679, 32'hc0d725db} /* (14, 4, 9) {real, imag} */,
  {32'hc08b8abd, 32'h40f6d71a} /* (14, 4, 8) {real, imag} */,
  {32'hc0a2d18d, 32'h405598ec} /* (14, 4, 7) {real, imag} */,
  {32'hc1a45d95, 32'h4195fbc3} /* (14, 4, 6) {real, imag} */,
  {32'hc1a04ab9, 32'hc154b97a} /* (14, 4, 5) {real, imag} */,
  {32'h417d4c94, 32'h41e268e5} /* (14, 4, 4) {real, imag} */,
  {32'hc14c4708, 32'h41b6cea1} /* (14, 4, 3) {real, imag} */,
  {32'hc27d71c0, 32'hc280cfd4} /* (14, 4, 2) {real, imag} */,
  {32'h4321860a, 32'h41dfed02} /* (14, 4, 1) {real, imag} */,
  {32'hc05038b8, 32'hc1b63da8} /* (14, 4, 0) {real, imag} */,
  {32'hc2a04d1c, 32'h423015a3} /* (14, 3, 31) {real, imag} */,
  {32'h428c3096, 32'hc2549870} /* (14, 3, 30) {real, imag} */,
  {32'hc11d9938, 32'h41f94558} /* (14, 3, 29) {real, imag} */,
  {32'h41cbba10, 32'h418aeab8} /* (14, 3, 28) {real, imag} */,
  {32'hc1981f2e, 32'hc1048d60} /* (14, 3, 27) {real, imag} */,
  {32'hc10bb090, 32'hc0529ec8} /* (14, 3, 26) {real, imag} */,
  {32'hc0611cb9, 32'hc0f19618} /* (14, 3, 25) {real, imag} */,
  {32'hc13dad1d, 32'hc10d8afe} /* (14, 3, 24) {real, imag} */,
  {32'hc1a59772, 32'hc0e95803} /* (14, 3, 23) {real, imag} */,
  {32'hc11849e9, 32'h41bf51fd} /* (14, 3, 22) {real, imag} */,
  {32'hc136a7db, 32'hc13b18dc} /* (14, 3, 21) {real, imag} */,
  {32'h411a6fe2, 32'h413a8d5e} /* (14, 3, 20) {real, imag} */,
  {32'h412c1c13, 32'hc09b2ac4} /* (14, 3, 19) {real, imag} */,
  {32'hbff62d7f, 32'hc0aea436} /* (14, 3, 18) {real, imag} */,
  {32'hc0496dfb, 32'h3fa6038c} /* (14, 3, 17) {real, imag} */,
  {32'hc0850566, 32'h3fcaaae0} /* (14, 3, 16) {real, imag} */,
  {32'hc0d6e812, 32'h410848bc} /* (14, 3, 15) {real, imag} */,
  {32'h411e6c95, 32'h40518254} /* (14, 3, 14) {real, imag} */,
  {32'hbf839296, 32'hbfe41104} /* (14, 3, 13) {real, imag} */,
  {32'h40280470, 32'h4025163c} /* (14, 3, 12) {real, imag} */,
  {32'h413f6950, 32'h418759ef} /* (14, 3, 11) {real, imag} */,
  {32'hc01a3350, 32'h409a661c} /* (14, 3, 10) {real, imag} */,
  {32'hc0df326e, 32'hc1eef5bc} /* (14, 3, 9) {real, imag} */,
  {32'h413e50a5, 32'h3f478ec0} /* (14, 3, 8) {real, imag} */,
  {32'h41c5b8bc, 32'hc0c3492c} /* (14, 3, 7) {real, imag} */,
  {32'h3f1e43c0, 32'hc0a74f0c} /* (14, 3, 6) {real, imag} */,
  {32'h40a551f8, 32'h420a92a0} /* (14, 3, 5) {real, imag} */,
  {32'hc0f44766, 32'h41a2b238} /* (14, 3, 4) {real, imag} */,
  {32'h4190bc2d, 32'h414550dc} /* (14, 3, 3) {real, imag} */,
  {32'hc1d7d97b, 32'hc27eee7a} /* (14, 3, 2) {real, imag} */,
  {32'h42daa10d, 32'h428aa287} /* (14, 3, 1) {real, imag} */,
  {32'h41a3d1be, 32'h40d22f1e} /* (14, 3, 0) {real, imag} */,
  {32'hc4404433, 32'hc2800be0} /* (14, 2, 31) {real, imag} */,
  {32'h43ca1049, 32'hc31496c6} /* (14, 2, 30) {real, imag} */,
  {32'h41384045, 32'h4154297a} /* (14, 2, 29) {real, imag} */,
  {32'hc24fb7b5, 32'h42a96ac6} /* (14, 2, 28) {real, imag} */,
  {32'h423befd2, 32'hc17e4132} /* (14, 2, 27) {real, imag} */,
  {32'h405fc6a8, 32'hc1b90066} /* (14, 2, 26) {real, imag} */,
  {32'hc1ccc744, 32'h4115f5cf} /* (14, 2, 25) {real, imag} */,
  {32'h409c9cd3, 32'hc16373d8} /* (14, 2, 24) {real, imag} */,
  {32'h4032944b, 32'hc15eecb2} /* (14, 2, 23) {real, imag} */,
  {32'h40ae2cb8, 32'h4177ca5b} /* (14, 2, 22) {real, imag} */,
  {32'h406be5cd, 32'hc08c533c} /* (14, 2, 21) {real, imag} */,
  {32'h40e26fd6, 32'hc138df83} /* (14, 2, 20) {real, imag} */,
  {32'hc11fbfbf, 32'h4126809e} /* (14, 2, 19) {real, imag} */,
  {32'h40c92458, 32'hc1903a1c} /* (14, 2, 18) {real, imag} */,
  {32'h40f98700, 32'h4184d02c} /* (14, 2, 17) {real, imag} */,
  {32'h3fd507f8, 32'hc0b23628} /* (14, 2, 16) {real, imag} */,
  {32'hbf646878, 32'h3fee0fb6} /* (14, 2, 15) {real, imag} */,
  {32'h41bce754, 32'h40552982} /* (14, 2, 14) {real, imag} */,
  {32'hc1930e4a, 32'h4128162b} /* (14, 2, 13) {real, imag} */,
  {32'hbff1e780, 32'hc115bf64} /* (14, 2, 12) {real, imag} */,
  {32'h40fab9d2, 32'h4181fa44} /* (14, 2, 11) {real, imag} */,
  {32'hbf719170, 32'h4078a7ac} /* (14, 2, 10) {real, imag} */,
  {32'h3f8ca328, 32'h4145aa72} /* (14, 2, 9) {real, imag} */,
  {32'h4240d158, 32'h416e1d02} /* (14, 2, 8) {real, imag} */,
  {32'hbf366040, 32'h409e00c3} /* (14, 2, 7) {real, imag} */,
  {32'hc14bac48, 32'h421a9d6f} /* (14, 2, 6) {real, imag} */,
  {32'h425387d8, 32'h429dad09} /* (14, 2, 5) {real, imag} */,
  {32'hc23a6fd8, 32'hc2790b6e} /* (14, 2, 4) {real, imag} */,
  {32'h40be1bd8, 32'h40a6f602} /* (14, 2, 3) {real, imag} */,
  {32'h437ef71b, 32'hc1db8362} /* (14, 2, 2) {real, imag} */,
  {32'hc3dce4b0, 32'h421bfa32} /* (14, 2, 1) {real, imag} */,
  {32'hc3cedef5, 32'hc2791f82} /* (14, 2, 0) {real, imag} */,
  {32'h44754011, 32'hc3819160} /* (14, 1, 31) {real, imag} */,
  {32'hc38f225e, 32'hc18fbbcb} /* (14, 1, 30) {real, imag} */,
  {32'h40625e82, 32'h42786364} /* (14, 1, 29) {real, imag} */,
  {32'h428bda14, 32'hc0b2bcd8} /* (14, 1, 28) {real, imag} */,
  {32'hc2a1f3d4, 32'h41973340} /* (14, 1, 27) {real, imag} */,
  {32'h41bc57f6, 32'hc0b6ba80} /* (14, 1, 26) {real, imag} */,
  {32'h3db42880, 32'h41e734e8} /* (14, 1, 25) {real, imag} */,
  {32'hc20962fe, 32'h400a0b3c} /* (14, 1, 24) {real, imag} */,
  {32'hc13d07ec, 32'hc05cc148} /* (14, 1, 23) {real, imag} */,
  {32'h410330a7, 32'hc04fd346} /* (14, 1, 22) {real, imag} */,
  {32'hc16b1256, 32'h41fb4b94} /* (14, 1, 21) {real, imag} */,
  {32'hc08537a0, 32'hc08bb386} /* (14, 1, 20) {real, imag} */,
  {32'hbfd48f88, 32'hc08c41e0} /* (14, 1, 19) {real, imag} */,
  {32'hbfe14204, 32'h412444f4} /* (14, 1, 18) {real, imag} */,
  {32'hc06a6e9e, 32'h40eb499e} /* (14, 1, 17) {real, imag} */,
  {32'h40cfc513, 32'hc085c5da} /* (14, 1, 16) {real, imag} */,
  {32'hc0b7a2e6, 32'h40969be0} /* (14, 1, 15) {real, imag} */,
  {32'hc010b127, 32'hc171a5a8} /* (14, 1, 14) {real, imag} */,
  {32'h41a5bc2e, 32'h3da6aab0} /* (14, 1, 13) {real, imag} */,
  {32'h40e6d3df, 32'hc0cee9a6} /* (14, 1, 12) {real, imag} */,
  {32'h3ec9ea30, 32'hc19c8435} /* (14, 1, 11) {real, imag} */,
  {32'hc00ad7d8, 32'hc111c863} /* (14, 1, 10) {real, imag} */,
  {32'hbffadf00, 32'h40f06a1c} /* (14, 1, 9) {real, imag} */,
  {32'hc18d17b2, 32'hc14c599e} /* (14, 1, 8) {real, imag} */,
  {32'h41bba0cb, 32'h41f5aa6e} /* (14, 1, 7) {real, imag} */,
  {32'h40462b18, 32'hc2428469} /* (14, 1, 6) {real, imag} */,
  {32'hc20e2118, 32'hc1fe0fc7} /* (14, 1, 5) {real, imag} */,
  {32'hc201c90a, 32'h428b4e7f} /* (14, 1, 4) {real, imag} */,
  {32'hc2d292c6, 32'hc1346ae2} /* (14, 1, 3) {real, imag} */,
  {32'hc3c4f800, 32'hc3ac851c} /* (14, 1, 2) {real, imag} */,
  {32'h449b9faf, 32'h44442c5e} /* (14, 1, 1) {real, imag} */,
  {32'h448aa966, 32'hc17fab80} /* (14, 1, 0) {real, imag} */,
  {32'h4421fa34, 32'hc40d8503} /* (14, 0, 31) {real, imag} */,
  {32'hc2f3e1ad, 32'h434e8f90} /* (14, 0, 30) {real, imag} */,
  {32'h4128c798, 32'h408f08a0} /* (14, 0, 29) {real, imag} */,
  {32'hc18721a9, 32'h415d747f} /* (14, 0, 28) {real, imag} */,
  {32'hc2736b84, 32'h4141dbec} /* (14, 0, 27) {real, imag} */,
  {32'h3ee20210, 32'hc0fc444c} /* (14, 0, 26) {real, imag} */,
  {32'hc115e2c2, 32'hc0f52606} /* (14, 0, 25) {real, imag} */,
  {32'h41a89dfb, 32'h418819f4} /* (14, 0, 24) {real, imag} */,
  {32'hc166cc03, 32'h40d88449} /* (14, 0, 23) {real, imag} */,
  {32'hc1744116, 32'hc1cf10b5} /* (14, 0, 22) {real, imag} */,
  {32'hc161921f, 32'h3ec09550} /* (14, 0, 21) {real, imag} */,
  {32'h418c5a07, 32'h412bcc18} /* (14, 0, 20) {real, imag} */,
  {32'h3f12ab38, 32'hc0b7d640} /* (14, 0, 19) {real, imag} */,
  {32'hc1608057, 32'h4122d0d7} /* (14, 0, 18) {real, imag} */,
  {32'hc0681d9e, 32'h411bcf86} /* (14, 0, 17) {real, imag} */,
  {32'h4076c459, 32'h00000000} /* (14, 0, 16) {real, imag} */,
  {32'hc0681d9e, 32'hc11bcf86} /* (14, 0, 15) {real, imag} */,
  {32'hc1608057, 32'hc122d0d7} /* (14, 0, 14) {real, imag} */,
  {32'h3f12ab38, 32'h40b7d640} /* (14, 0, 13) {real, imag} */,
  {32'h418c5a07, 32'hc12bcc18} /* (14, 0, 12) {real, imag} */,
  {32'hc161921f, 32'hbec09550} /* (14, 0, 11) {real, imag} */,
  {32'hc1744116, 32'h41cf10b5} /* (14, 0, 10) {real, imag} */,
  {32'hc166cc03, 32'hc0d88449} /* (14, 0, 9) {real, imag} */,
  {32'h41a89dfb, 32'hc18819f4} /* (14, 0, 8) {real, imag} */,
  {32'hc115e2c2, 32'h40f52606} /* (14, 0, 7) {real, imag} */,
  {32'h3ee20210, 32'h40fc444c} /* (14, 0, 6) {real, imag} */,
  {32'hc2736b84, 32'hc141dbec} /* (14, 0, 5) {real, imag} */,
  {32'hc18721a9, 32'hc15d747f} /* (14, 0, 4) {real, imag} */,
  {32'h4128c798, 32'hc08f08a0} /* (14, 0, 3) {real, imag} */,
  {32'hc2f3e1ad, 32'hc34e8f90} /* (14, 0, 2) {real, imag} */,
  {32'h4421fa34, 32'h440d8503} /* (14, 0, 1) {real, imag} */,
  {32'h448f1b02, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h44e1b185, 32'hc4886478} /* (13, 31, 31) {real, imag} */,
  {32'hc402e8c4, 32'h43ec369e} /* (13, 31, 30) {real, imag} */,
  {32'hc2b4c27d, 32'h40dada78} /* (13, 31, 29) {real, imag} */,
  {32'hc1ae13db, 32'hc2a3767e} /* (13, 31, 28) {real, imag} */,
  {32'hc25abc92, 32'h41a7d83a} /* (13, 31, 27) {real, imag} */,
  {32'hc126abd0, 32'h423c441e} /* (13, 31, 26) {real, imag} */,
  {32'h4204747f, 32'hc0e777a5} /* (13, 31, 25) {real, imag} */,
  {32'hc0f87749, 32'h423a3654} /* (13, 31, 24) {real, imag} */,
  {32'h402cbf30, 32'hc0a3a6f9} /* (13, 31, 23) {real, imag} */,
  {32'h40d5f99e, 32'h40d461a2} /* (13, 31, 22) {real, imag} */,
  {32'hc1684b84, 32'hc0d87810} /* (13, 31, 21) {real, imag} */,
  {32'h41832e1e, 32'h40209c45} /* (13, 31, 20) {real, imag} */,
  {32'hc0091a82, 32'h40927560} /* (13, 31, 19) {real, imag} */,
  {32'h40daa498, 32'hc142f752} /* (13, 31, 18) {real, imag} */,
  {32'hc095677c, 32'h40d04219} /* (13, 31, 17) {real, imag} */,
  {32'h3f9e4d7a, 32'hc06b9c43} /* (13, 31, 16) {real, imag} */,
  {32'hc0eb603b, 32'h413797e4} /* (13, 31, 15) {real, imag} */,
  {32'hbf76c148, 32'hc11373e6} /* (13, 31, 14) {real, imag} */,
  {32'h403a2386, 32'h41080944} /* (13, 31, 13) {real, imag} */,
  {32'hc0c962ea, 32'h4096c8ee} /* (13, 31, 12) {real, imag} */,
  {32'h40f7833e, 32'hc1d130c4} /* (13, 31, 11) {real, imag} */,
  {32'h4156a2ef, 32'hc167e2aa} /* (13, 31, 10) {real, imag} */,
  {32'hc1e65271, 32'hc11d0d82} /* (13, 31, 9) {real, imag} */,
  {32'hc1c5ff5d, 32'hc1e73836} /* (13, 31, 8) {real, imag} */,
  {32'h40cf47b6, 32'hc08a0662} /* (13, 31, 7) {real, imag} */,
  {32'h41f15cf4, 32'hbf731240} /* (13, 31, 6) {real, imag} */,
  {32'hc2d0536d, 32'hc1939335} /* (13, 31, 5) {real, imag} */,
  {32'h428aae68, 32'hc18e8612} /* (13, 31, 4) {real, imag} */,
  {32'h407b94b8, 32'hc2490d33} /* (13, 31, 3) {real, imag} */,
  {32'hc3b454ff, 32'h3ddbd280} /* (13, 31, 2) {real, imag} */,
  {32'h44aa3b02, 32'h439bc8b7} /* (13, 31, 1) {real, imag} */,
  {32'h44d0d69a, 32'hc289118f} /* (13, 31, 0) {real, imag} */,
  {32'hc41114de, 32'hc2828f76} /* (13, 30, 31) {real, imag} */,
  {32'h439f13b5, 32'h42b25670} /* (13, 30, 30) {real, imag} */,
  {32'h4130d0ee, 32'hc1176950} /* (13, 30, 29) {real, imag} */,
  {32'hc2a94460, 32'h4280e95a} /* (13, 30, 28) {real, imag} */,
  {32'h422d1202, 32'hc292c31d} /* (13, 30, 27) {real, imag} */,
  {32'h40c2dbcf, 32'hc1a0b9a9} /* (13, 30, 26) {real, imag} */,
  {32'hc184c831, 32'h4148bc52} /* (13, 30, 25) {real, imag} */,
  {32'h41b20941, 32'h40c89240} /* (13, 30, 24) {real, imag} */,
  {32'hc129a519, 32'h411a11d5} /* (13, 30, 23) {real, imag} */,
  {32'hc073e737, 32'hc02ed053} /* (13, 30, 22) {real, imag} */,
  {32'h400a8dfa, 32'hc10e0133} /* (13, 30, 21) {real, imag} */,
  {32'h4144da32, 32'h3f99dd4a} /* (13, 30, 20) {real, imag} */,
  {32'hc0441c38, 32'h3ff27df8} /* (13, 30, 19) {real, imag} */,
  {32'h4086d73e, 32'h3f477020} /* (13, 30, 18) {real, imag} */,
  {32'hc07a6fe6, 32'hc000c659} /* (13, 30, 17) {real, imag} */,
  {32'h404048ba, 32'h4109ff00} /* (13, 30, 16) {real, imag} */,
  {32'h40a71e94, 32'h4071e27c} /* (13, 30, 15) {real, imag} */,
  {32'h40d2eaa6, 32'h40b9d64a} /* (13, 30, 14) {real, imag} */,
  {32'hc13d2edf, 32'hc13dddff} /* (13, 30, 13) {real, imag} */,
  {32'hc108a3c5, 32'h3f823a6c} /* (13, 30, 12) {real, imag} */,
  {32'h41c5c5b7, 32'h41965722} /* (13, 30, 11) {real, imag} */,
  {32'h3ffbe8a6, 32'hc0c51894} /* (13, 30, 10) {real, imag} */,
  {32'hc1aa734e, 32'hc01195c8} /* (13, 30, 9) {real, imag} */,
  {32'h418a2f20, 32'h421cc432} /* (13, 30, 8) {real, imag} */,
  {32'hc1bf6962, 32'hc1268bfe} /* (13, 30, 7) {real, imag} */,
  {32'h41f1b084, 32'h41964333} /* (13, 30, 6) {real, imag} */,
  {32'h4252dfd8, 32'h422eb7d0} /* (13, 30, 5) {real, imag} */,
  {32'hc27c727d, 32'hc29aa5a0} /* (13, 30, 4) {real, imag} */,
  {32'h418ee477, 32'hc236c940} /* (13, 30, 3) {real, imag} */,
  {32'h4400fd8c, 32'h433c423d} /* (13, 30, 2) {real, imag} */,
  {32'hc4815e68, 32'h42018fb5} /* (13, 30, 1) {real, imag} */,
  {32'hc400e086, 32'h4281dfa2} /* (13, 30, 0) {real, imag} */,
  {32'h431fb372, 32'hc2be16a3} /* (13, 29, 31) {real, imag} */,
  {32'hc1fe4c2e, 32'h428f0f16} /* (13, 29, 30) {real, imag} */,
  {32'h40081768, 32'hc16725fc} /* (13, 29, 29) {real, imag} */,
  {32'hc0f1406c, 32'hc11adfc1} /* (13, 29, 28) {real, imag} */,
  {32'h4092de62, 32'hc2015ec2} /* (13, 29, 27) {real, imag} */,
  {32'h409ada3e, 32'h40d748a0} /* (13, 29, 26) {real, imag} */,
  {32'h41873f7e, 32'hc0d45d4e} /* (13, 29, 25) {real, imag} */,
  {32'h41544653, 32'h40e32b28} /* (13, 29, 24) {real, imag} */,
  {32'hc1a665ad, 32'h41c5a785} /* (13, 29, 23) {real, imag} */,
  {32'hc1355213, 32'hc0c8641c} /* (13, 29, 22) {real, imag} */,
  {32'h419c4002, 32'h40aebbca} /* (13, 29, 21) {real, imag} */,
  {32'h410734c1, 32'h413ae193} /* (13, 29, 20) {real, imag} */,
  {32'hbfe28a90, 32'hc0d394ce} /* (13, 29, 19) {real, imag} */,
  {32'hc1140fbd, 32'hc0dfb95f} /* (13, 29, 18) {real, imag} */,
  {32'h41062dcb, 32'h41759eb1} /* (13, 29, 17) {real, imag} */,
  {32'h408c217f, 32'h4017d838} /* (13, 29, 16) {real, imag} */,
  {32'hc09b4100, 32'hc1306c75} /* (13, 29, 15) {real, imag} */,
  {32'hc0519008, 32'hc0f9caa6} /* (13, 29, 14) {real, imag} */,
  {32'hc0976c15, 32'h4122b43e} /* (13, 29, 13) {real, imag} */,
  {32'hc10bb8bf, 32'h4144d7fd} /* (13, 29, 12) {real, imag} */,
  {32'hc0aea28d, 32'h40b53435} /* (13, 29, 11) {real, imag} */,
  {32'h4054200c, 32'hc19f8cf4} /* (13, 29, 10) {real, imag} */,
  {32'h3d640c80, 32'hc0e8fc8d} /* (13, 29, 9) {real, imag} */,
  {32'h4112f958, 32'h419f822c} /* (13, 29, 8) {real, imag} */,
  {32'h417954ec, 32'hc1045988} /* (13, 29, 7) {real, imag} */,
  {32'hc1def5ef, 32'hbf0bc6b0} /* (13, 29, 6) {real, imag} */,
  {32'hc1166041, 32'hc10d634d} /* (13, 29, 5) {real, imag} */,
  {32'h42019c62, 32'hc1e10618} /* (13, 29, 4) {real, imag} */,
  {32'hc1442026, 32'hc1ae3352} /* (13, 29, 3) {real, imag} */,
  {32'h42b1e709, 32'h429ad8bc} /* (13, 29, 2) {real, imag} */,
  {32'hc323e835, 32'hc2361e82} /* (13, 29, 1) {real, imag} */,
  {32'h3fa660e0, 32'h416acc22} /* (13, 29, 0) {real, imag} */,
  {32'h434134bb, 32'hc1a3fbe6} /* (13, 28, 31) {real, imag} */,
  {32'hc2738a88, 32'h4294fddf} /* (13, 28, 30) {real, imag} */,
  {32'hc13d5dd2, 32'hc1c66230} /* (13, 28, 29) {real, imag} */,
  {32'hc115f132, 32'hc1950263} /* (13, 28, 28) {real, imag} */,
  {32'hc115d4a8, 32'h4212b3a1} /* (13, 28, 27) {real, imag} */,
  {32'hc134e8dc, 32'hc115d063} /* (13, 28, 26) {real, imag} */,
  {32'hc138111a, 32'h40ef40a5} /* (13, 28, 25) {real, imag} */,
  {32'h3e88b118, 32'h41a796ce} /* (13, 28, 24) {real, imag} */,
  {32'h412bf314, 32'hbe9fd3e0} /* (13, 28, 23) {real, imag} */,
  {32'hc172e426, 32'hbfd37064} /* (13, 28, 22) {real, imag} */,
  {32'h41672d82, 32'hc05c4be5} /* (13, 28, 21) {real, imag} */,
  {32'hc03c8419, 32'hc135cf08} /* (13, 28, 20) {real, imag} */,
  {32'h410f1810, 32'h41182688} /* (13, 28, 19) {real, imag} */,
  {32'hbff32c70, 32'h414bbd1f} /* (13, 28, 18) {real, imag} */,
  {32'h40de528c, 32'h40061a46} /* (13, 28, 17) {real, imag} */,
  {32'h3fdec480, 32'hc0bf1d7d} /* (13, 28, 16) {real, imag} */,
  {32'h4117c6a2, 32'h3f210444} /* (13, 28, 15) {real, imag} */,
  {32'h40ab6e14, 32'hc16ace81} /* (13, 28, 14) {real, imag} */,
  {32'h413c092b, 32'h414bc68e} /* (13, 28, 13) {real, imag} */,
  {32'hc15910d7, 32'h41522389} /* (13, 28, 12) {real, imag} */,
  {32'hc162338a, 32'hc1164ae7} /* (13, 28, 11) {real, imag} */,
  {32'h40a75a64, 32'h3e133c00} /* (13, 28, 10) {real, imag} */,
  {32'h408589ea, 32'h418d8598} /* (13, 28, 9) {real, imag} */,
  {32'h3fdd60bc, 32'h41bf91f0} /* (13, 28, 8) {real, imag} */,
  {32'h40b60ff3, 32'hc0feea37} /* (13, 28, 7) {real, imag} */,
  {32'hc0d001d2, 32'h40c8ca52} /* (13, 28, 6) {real, imag} */,
  {32'hc19a2cce, 32'h4101cccb} /* (13, 28, 5) {real, imag} */,
  {32'h4258e3ca, 32'hc1ffa87d} /* (13, 28, 4) {real, imag} */,
  {32'hc1ae96af, 32'h41408be4} /* (13, 28, 3) {real, imag} */,
  {32'hc2ae7a55, 32'h42a671e1} /* (13, 28, 2) {real, imag} */,
  {32'h42763424, 32'hc27eb9e1} /* (13, 28, 1) {real, imag} */,
  {32'h41380e20, 32'h412ec639} /* (13, 28, 0) {real, imag} */,
  {32'hc2c6f1cc, 32'h422f97c2} /* (13, 27, 31) {real, imag} */,
  {32'h40e5bdfc, 32'hc2162bd2} /* (13, 27, 30) {real, imag} */,
  {32'hc0144124, 32'hc1524846} /* (13, 27, 29) {real, imag} */,
  {32'h41173b86, 32'h414777c2} /* (13, 27, 28) {real, imag} */,
  {32'h412eb203, 32'h3e5f9100} /* (13, 27, 27) {real, imag} */,
  {32'hc0b6526f, 32'hc2047398} /* (13, 27, 26) {real, imag} */,
  {32'h411c90d6, 32'h415b972a} /* (13, 27, 25) {real, imag} */,
  {32'hc0dc47e2, 32'hc0cb32e7} /* (13, 27, 24) {real, imag} */,
  {32'h4175407a, 32'h3f0607c0} /* (13, 27, 23) {real, imag} */,
  {32'hbff75528, 32'hc001d2b2} /* (13, 27, 22) {real, imag} */,
  {32'h40acc1d8, 32'hc180485e} /* (13, 27, 21) {real, imag} */,
  {32'h41a9452e, 32'h41dbfb07} /* (13, 27, 20) {real, imag} */,
  {32'hc1167bc6, 32'h412c0b6e} /* (13, 27, 19) {real, imag} */,
  {32'h3fd29ed2, 32'hc09929b3} /* (13, 27, 18) {real, imag} */,
  {32'hc1b9ec88, 32'hc09ed446} /* (13, 27, 17) {real, imag} */,
  {32'hc08e8f1e, 32'h4121450c} /* (13, 27, 16) {real, imag} */,
  {32'h40cbab56, 32'hbf157c20} /* (13, 27, 15) {real, imag} */,
  {32'h40adddfe, 32'h40e8ec86} /* (13, 27, 14) {real, imag} */,
  {32'hc13ad052, 32'h40d59138} /* (13, 27, 13) {real, imag} */,
  {32'hc16795e5, 32'hc0f08931} /* (13, 27, 12) {real, imag} */,
  {32'h41878da4, 32'h40f0f856} /* (13, 27, 11) {real, imag} */,
  {32'h4111f752, 32'hc042755a} /* (13, 27, 10) {real, imag} */,
  {32'h3ec89760, 32'hc20c54eb} /* (13, 27, 9) {real, imag} */,
  {32'hbff696ac, 32'h41a39c88} /* (13, 27, 8) {real, imag} */,
  {32'h40e1e970, 32'h412f145e} /* (13, 27, 7) {real, imag} */,
  {32'h412384c4, 32'hc101ae72} /* (13, 27, 6) {real, imag} */,
  {32'h4203f2be, 32'hc11c3dfb} /* (13, 27, 5) {real, imag} */,
  {32'hc1972e40, 32'hc106de6e} /* (13, 27, 4) {real, imag} */,
  {32'h40dc56b6, 32'hc1ad358a} /* (13, 27, 3) {real, imag} */,
  {32'h41813790, 32'hc138a0b9} /* (13, 27, 2) {real, imag} */,
  {32'hc2b63146, 32'h4081a5b4} /* (13, 27, 1) {real, imag} */,
  {32'hc26f3a4c, 32'h4212d780} /* (13, 27, 0) {real, imag} */,
  {32'hc1c455c4, 32'h41b2da9a} /* (13, 26, 31) {real, imag} */,
  {32'h41f7b36e, 32'hc149b3ee} /* (13, 26, 30) {real, imag} */,
  {32'hbff39ad0, 32'hc0f469ec} /* (13, 26, 29) {real, imag} */,
  {32'hc1af4012, 32'hc085c350} /* (13, 26, 28) {real, imag} */,
  {32'hc1ac545c, 32'h41a2170a} /* (13, 26, 27) {real, imag} */,
  {32'hc1543b88, 32'h41af63c4} /* (13, 26, 26) {real, imag} */,
  {32'hc16fb5fe, 32'hc0c11700} /* (13, 26, 25) {real, imag} */,
  {32'h41baa759, 32'hbf9bdf78} /* (13, 26, 24) {real, imag} */,
  {32'hc1316944, 32'hc15c55bc} /* (13, 26, 23) {real, imag} */,
  {32'hc011fb8b, 32'h41a2e4eb} /* (13, 26, 22) {real, imag} */,
  {32'hbf4e3ed0, 32'hc1da7a4e} /* (13, 26, 21) {real, imag} */,
  {32'h40764150, 32'h40159ac3} /* (13, 26, 20) {real, imag} */,
  {32'h41835f85, 32'hc05c0136} /* (13, 26, 19) {real, imag} */,
  {32'h4103e04a, 32'h41280c0f} /* (13, 26, 18) {real, imag} */,
  {32'h40b8ad38, 32'h410f9a67} /* (13, 26, 17) {real, imag} */,
  {32'hc133c81d, 32'h3fa4bdec} /* (13, 26, 16) {real, imag} */,
  {32'hc09c5098, 32'hbf83a1c8} /* (13, 26, 15) {real, imag} */,
  {32'h411bf044, 32'h4137df40} /* (13, 26, 14) {real, imag} */,
  {32'h41095335, 32'hc13ec5c2} /* (13, 26, 13) {real, imag} */,
  {32'hc09db331, 32'hc0119c30} /* (13, 26, 12) {real, imag} */,
  {32'hbf048af8, 32'h402a0f5e} /* (13, 26, 11) {real, imag} */,
  {32'h4055be40, 32'hc198c41e} /* (13, 26, 10) {real, imag} */,
  {32'h400229a9, 32'h40ce1962} /* (13, 26, 9) {real, imag} */,
  {32'h3f849590, 32'hbf4f6850} /* (13, 26, 8) {real, imag} */,
  {32'h3ff944b4, 32'h415b0ebc} /* (13, 26, 7) {real, imag} */,
  {32'h415bfc44, 32'hc0c79ad8} /* (13, 26, 6) {real, imag} */,
  {32'h41ac914a, 32'hbfe336be} /* (13, 26, 5) {real, imag} */,
  {32'hc0ee3792, 32'h41157319} /* (13, 26, 4) {real, imag} */,
  {32'h40757450, 32'h419817bb} /* (13, 26, 3) {real, imag} */,
  {32'h4229db9c, 32'h41c76efd} /* (13, 26, 2) {real, imag} */,
  {32'hc1664e1a, 32'h408adba3} /* (13, 26, 1) {real, imag} */,
  {32'h40f6795a, 32'hc1b60a7b} /* (13, 26, 0) {real, imag} */,
  {32'h4169c74d, 32'hc23f104b} /* (13, 25, 31) {real, imag} */,
  {32'h4167deae, 32'h4166f549} /* (13, 25, 30) {real, imag} */,
  {32'hc0446cfc, 32'hc1543637} /* (13, 25, 29) {real, imag} */,
  {32'hc1a86111, 32'hc08cb928} /* (13, 25, 28) {real, imag} */,
  {32'h4161087c, 32'h401e804a} /* (13, 25, 27) {real, imag} */,
  {32'h41450506, 32'h3fadf2d8} /* (13, 25, 26) {real, imag} */,
  {32'h3ff833a8, 32'h40234031} /* (13, 25, 25) {real, imag} */,
  {32'hc17e0184, 32'h40b5bd42} /* (13, 25, 24) {real, imag} */,
  {32'hc09566b0, 32'hc10e7455} /* (13, 25, 23) {real, imag} */,
  {32'hc0a5bddc, 32'hc12ae05d} /* (13, 25, 22) {real, imag} */,
  {32'hc09a5f72, 32'hbf846b2e} /* (13, 25, 21) {real, imag} */,
  {32'h40e93226, 32'h4122d604} /* (13, 25, 20) {real, imag} */,
  {32'h3fd1b3c8, 32'h41687e1b} /* (13, 25, 19) {real, imag} */,
  {32'h40295782, 32'h3f396acc} /* (13, 25, 18) {real, imag} */,
  {32'h40ca45a5, 32'hc00b3fe8} /* (13, 25, 17) {real, imag} */,
  {32'hc14d3524, 32'hc091d20c} /* (13, 25, 16) {real, imag} */,
  {32'h40b01ccf, 32'hc14a9326} /* (13, 25, 15) {real, imag} */,
  {32'hc030bc38, 32'hc187df6a} /* (13, 25, 14) {real, imag} */,
  {32'hc01e3db2, 32'hc0f5a208} /* (13, 25, 13) {real, imag} */,
  {32'h415c767b, 32'hbead32a0} /* (13, 25, 12) {real, imag} */,
  {32'hc12d4107, 32'h4164d3b6} /* (13, 25, 11) {real, imag} */,
  {32'h3fe5382a, 32'hc122babc} /* (13, 25, 10) {real, imag} */,
  {32'h40e3b5a9, 32'h415238b5} /* (13, 25, 9) {real, imag} */,
  {32'h40bf1851, 32'h400a33e2} /* (13, 25, 8) {real, imag} */,
  {32'h410b5e9b, 32'hbf0895f8} /* (13, 25, 7) {real, imag} */,
  {32'hc0ce8e8b, 32'hbd210700} /* (13, 25, 6) {real, imag} */,
  {32'hc0feb5ac, 32'hc1734fdc} /* (13, 25, 5) {real, imag} */,
  {32'hc108dfd9, 32'h3e9577b0} /* (13, 25, 4) {real, imag} */,
  {32'hc0412d74, 32'h418d8e94} /* (13, 25, 3) {real, imag} */,
  {32'h4123de80, 32'h413004e8} /* (13, 25, 2) {real, imag} */,
  {32'h414d5d92, 32'h40b6d18f} /* (13, 25, 1) {real, imag} */,
  {32'hc0c1bbab, 32'hc19745c3} /* (13, 25, 0) {real, imag} */,
  {32'hc22f2eba, 32'h41c285bf} /* (13, 24, 31) {real, imag} */,
  {32'h41ee168a, 32'h41c566d0} /* (13, 24, 30) {real, imag} */,
  {32'h41ab6674, 32'h4085acd5} /* (13, 24, 29) {real, imag} */,
  {32'hc17f26c8, 32'h41b75150} /* (13, 24, 28) {real, imag} */,
  {32'hbfe24394, 32'hc10d3d73} /* (13, 24, 27) {real, imag} */,
  {32'h417df968, 32'h3ff33aa4} /* (13, 24, 26) {real, imag} */,
  {32'hc0e27e16, 32'h3f743fe4} /* (13, 24, 25) {real, imag} */,
  {32'h40bc68aa, 32'hc05ec6c6} /* (13, 24, 24) {real, imag} */,
  {32'hc1033544, 32'hc0a7c22e} /* (13, 24, 23) {real, imag} */,
  {32'hc15c900a, 32'h40c3f10e} /* (13, 24, 22) {real, imag} */,
  {32'h421db97e, 32'h41737893} /* (13, 24, 21) {real, imag} */,
  {32'h4137d65b, 32'hc11b9e99} /* (13, 24, 20) {real, imag} */,
  {32'h4105eec9, 32'h4115ed24} /* (13, 24, 19) {real, imag} */,
  {32'h4085cd18, 32'h41014a58} /* (13, 24, 18) {real, imag} */,
  {32'h3ff288a8, 32'hc06b9f65} /* (13, 24, 17) {real, imag} */,
  {32'h4006819b, 32'hc1d56a2c} /* (13, 24, 16) {real, imag} */,
  {32'hc097df1d, 32'h40252309} /* (13, 24, 15) {real, imag} */,
  {32'h40671316, 32'hbfcfbf30} /* (13, 24, 14) {real, imag} */,
  {32'h4134266c, 32'hc08cd034} /* (13, 24, 13) {real, imag} */,
  {32'hc11b07d9, 32'h4083730e} /* (13, 24, 12) {real, imag} */,
  {32'h416bbe2a, 32'hbfa54296} /* (13, 24, 11) {real, imag} */,
  {32'hc1ce4388, 32'hc1811a72} /* (13, 24, 10) {real, imag} */,
  {32'h40bc2698, 32'hc1160ba1} /* (13, 24, 9) {real, imag} */,
  {32'h4208647e, 32'h410d5614} /* (13, 24, 8) {real, imag} */,
  {32'h413a8a2f, 32'h3e140f88} /* (13, 24, 7) {real, imag} */,
  {32'hc026b85a, 32'h411b6cd0} /* (13, 24, 6) {real, imag} */,
  {32'h41fc592c, 32'hc0d03528} /* (13, 24, 5) {real, imag} */,
  {32'h3d88a380, 32'hc1c8c3f1} /* (13, 24, 4) {real, imag} */,
  {32'h41aeb311, 32'h41a33ae5} /* (13, 24, 3) {real, imag} */,
  {32'h419b81c7, 32'hc1c1a334} /* (13, 24, 2) {real, imag} */,
  {32'hc24f58c9, 32'h41d8d77e} /* (13, 24, 1) {real, imag} */,
  {32'hc1af2008, 32'h4184792d} /* (13, 24, 0) {real, imag} */,
  {32'hc1080924, 32'hc1b4aedd} /* (13, 23, 31) {real, imag} */,
  {32'hbf84cb04, 32'h418cea07} /* (13, 23, 30) {real, imag} */,
  {32'hbf87f916, 32'h4122b074} /* (13, 23, 29) {real, imag} */,
  {32'hc1098ff6, 32'hc16895be} /* (13, 23, 28) {real, imag} */,
  {32'h41163c95, 32'h413d15b0} /* (13, 23, 27) {real, imag} */,
  {32'hc15ca715, 32'h41356770} /* (13, 23, 26) {real, imag} */,
  {32'h40c58030, 32'hc1df3370} /* (13, 23, 25) {real, imag} */,
  {32'hc0570b94, 32'hc082e662} /* (13, 23, 24) {real, imag} */,
  {32'hc14e9714, 32'hc17b700d} /* (13, 23, 23) {real, imag} */,
  {32'hc12fb682, 32'h411ac6fa} /* (13, 23, 22) {real, imag} */,
  {32'h41424fe6, 32'hbe7b2660} /* (13, 23, 21) {real, imag} */,
  {32'hc0a97dab, 32'hc106ea06} /* (13, 23, 20) {real, imag} */,
  {32'hc01e5efa, 32'hc138f85d} /* (13, 23, 19) {real, imag} */,
  {32'h41b1bf8d, 32'h3f83d4b8} /* (13, 23, 18) {real, imag} */,
  {32'hc12a80fb, 32'h4101612c} /* (13, 23, 17) {real, imag} */,
  {32'hc0eabf9a, 32'hc127d7c8} /* (13, 23, 16) {real, imag} */,
  {32'hc14002a4, 32'hc1877b3f} /* (13, 23, 15) {real, imag} */,
  {32'hc0a1cd9e, 32'h410dddbe} /* (13, 23, 14) {real, imag} */,
  {32'h4103ac4e, 32'hbed32780} /* (13, 23, 13) {real, imag} */,
  {32'h40744b37, 32'h4141a116} /* (13, 23, 12) {real, imag} */,
  {32'hc19c89b2, 32'h40241e4d} /* (13, 23, 11) {real, imag} */,
  {32'hc02645ae, 32'hc0c5fc3f} /* (13, 23, 10) {real, imag} */,
  {32'h418e1bf5, 32'hc15be339} /* (13, 23, 9) {real, imag} */,
  {32'hc037ded2, 32'hc186331b} /* (13, 23, 8) {real, imag} */,
  {32'hc1024eaf, 32'h4092e09c} /* (13, 23, 7) {real, imag} */,
  {32'hbf0a5f70, 32'hc034fcf9} /* (13, 23, 6) {real, imag} */,
  {32'hc18fadd6, 32'hc0ff303e} /* (13, 23, 5) {real, imag} */,
  {32'h41c802d2, 32'h40b72d2a} /* (13, 23, 4) {real, imag} */,
  {32'h4159941a, 32'hbeba3180} /* (13, 23, 3) {real, imag} */,
  {32'h41a18c14, 32'h4166f0fe} /* (13, 23, 2) {real, imag} */,
  {32'h3ef59ad0, 32'hc15f00bd} /* (13, 23, 1) {real, imag} */,
  {32'hc053332f, 32'h415469e4} /* (13, 23, 0) {real, imag} */,
  {32'h41adc711, 32'hc0455a7c} /* (13, 22, 31) {real, imag} */,
  {32'hbf8666a0, 32'h41aeea29} /* (13, 22, 30) {real, imag} */,
  {32'hc0c2680c, 32'h41582738} /* (13, 22, 29) {real, imag} */,
  {32'h41946580, 32'hbfa180c8} /* (13, 22, 28) {real, imag} */,
  {32'h40354b56, 32'hc10bc7c1} /* (13, 22, 27) {real, imag} */,
  {32'hc18819c7, 32'hc08e4ff8} /* (13, 22, 26) {real, imag} */,
  {32'h41bcdc03, 32'hc0cb21b2} /* (13, 22, 25) {real, imag} */,
  {32'hc1b72f7e, 32'hc1913b78} /* (13, 22, 24) {real, imag} */,
  {32'h4180c720, 32'h40ce1d96} /* (13, 22, 23) {real, imag} */,
  {32'hbf95e1b8, 32'h410abcfb} /* (13, 22, 22) {real, imag} */,
  {32'h41a6130f, 32'hc10f9e3a} /* (13, 22, 21) {real, imag} */,
  {32'hc1d2cade, 32'hc0323997} /* (13, 22, 20) {real, imag} */,
  {32'hc140b2da, 32'h3f677738} /* (13, 22, 19) {real, imag} */,
  {32'hc11572b4, 32'h419b9d76} /* (13, 22, 18) {real, imag} */,
  {32'h40997282, 32'hc1847c52} /* (13, 22, 17) {real, imag} */,
  {32'h410cbc64, 32'hc10898c4} /* (13, 22, 16) {real, imag} */,
  {32'h412a81dc, 32'hbfa96c30} /* (13, 22, 15) {real, imag} */,
  {32'hc11fe6e2, 32'hbe65d1d0} /* (13, 22, 14) {real, imag} */,
  {32'h3f820a7c, 32'hc1b469d6} /* (13, 22, 13) {real, imag} */,
  {32'hc16f42cc, 32'hc0490442} /* (13, 22, 12) {real, imag} */,
  {32'hc127cfd8, 32'hc00d4ed0} /* (13, 22, 11) {real, imag} */,
  {32'h40d484eb, 32'h410c8177} /* (13, 22, 10) {real, imag} */,
  {32'h40cf7b84, 32'h3dbacf40} /* (13, 22, 9) {real, imag} */,
  {32'hc107b5ba, 32'hc0be29d8} /* (13, 22, 8) {real, imag} */,
  {32'hc135893a, 32'hc01277a2} /* (13, 22, 7) {real, imag} */,
  {32'h40c4d813, 32'hc1711c7e} /* (13, 22, 6) {real, imag} */,
  {32'h40df293c, 32'hc1321a0b} /* (13, 22, 5) {real, imag} */,
  {32'h40294be6, 32'h419b0f5b} /* (13, 22, 4) {real, imag} */,
  {32'hc0a7593d, 32'h4005be93} /* (13, 22, 3) {real, imag} */,
  {32'h412494da, 32'h413e2712} /* (13, 22, 2) {real, imag} */,
  {32'hbff30f36, 32'hc1a14af6} /* (13, 22, 1) {real, imag} */,
  {32'h413196e6, 32'hc15bb700} /* (13, 22, 0) {real, imag} */,
  {32'hc1339b49, 32'h41265f06} /* (13, 21, 31) {real, imag} */,
  {32'hc1cb90c4, 32'hc0c25e86} /* (13, 21, 30) {real, imag} */,
  {32'h4124024d, 32'h413c1d6d} /* (13, 21, 29) {real, imag} */,
  {32'h3f9bb8ea, 32'h4189e496} /* (13, 21, 28) {real, imag} */,
  {32'h40cd29f8, 32'hc0407806} /* (13, 21, 27) {real, imag} */,
  {32'hc0c105f6, 32'hc1177122} /* (13, 21, 26) {real, imag} */,
  {32'hc0a5dc36, 32'h411a48fa} /* (13, 21, 25) {real, imag} */,
  {32'h418ec45d, 32'h40503761} /* (13, 21, 24) {real, imag} */,
  {32'h4181cddc, 32'h4108e343} /* (13, 21, 23) {real, imag} */,
  {32'h4001ff48, 32'h41b62de9} /* (13, 21, 22) {real, imag} */,
  {32'hc0ce0f58, 32'h4024e4db} /* (13, 21, 21) {real, imag} */,
  {32'hc153cf73, 32'h408dac17} /* (13, 21, 20) {real, imag} */,
  {32'h41023aed, 32'h40b2ac36} /* (13, 21, 19) {real, imag} */,
  {32'h40c3b4ba, 32'hc100818e} /* (13, 21, 18) {real, imag} */,
  {32'hbfa69eec, 32'hc0bc3a6c} /* (13, 21, 17) {real, imag} */,
  {32'hc02b358d, 32'h411f04ac} /* (13, 21, 16) {real, imag} */,
  {32'h408754f7, 32'hc049a734} /* (13, 21, 15) {real, imag} */,
  {32'hc0c3e76e, 32'hc099ed15} /* (13, 21, 14) {real, imag} */,
  {32'h3f8a85a6, 32'h4096c683} /* (13, 21, 13) {real, imag} */,
  {32'h419794b1, 32'hc10f9875} /* (13, 21, 12) {real, imag} */,
  {32'hc03fdb08, 32'hc0d1e87f} /* (13, 21, 11) {real, imag} */,
  {32'hc0498028, 32'h4126a11d} /* (13, 21, 10) {real, imag} */,
  {32'h40c30698, 32'h412324b2} /* (13, 21, 9) {real, imag} */,
  {32'hc11680e4, 32'h4198614e} /* (13, 21, 8) {real, imag} */,
  {32'h411f9d51, 32'h41acde1a} /* (13, 21, 7) {real, imag} */,
  {32'hc01f3a3c, 32'h3f727d84} /* (13, 21, 6) {real, imag} */,
  {32'h4204d9dc, 32'hc184f27a} /* (13, 21, 5) {real, imag} */,
  {32'hc0579494, 32'hc0d9dc14} /* (13, 21, 4) {real, imag} */,
  {32'h4126345a, 32'h40f9e231} /* (13, 21, 3) {real, imag} */,
  {32'hc0841063, 32'hc1951ef5} /* (13, 21, 2) {real, imag} */,
  {32'hc18dfeed, 32'h40a2fd42} /* (13, 21, 1) {real, imag} */,
  {32'hc1a3ae54, 32'h415b33d4} /* (13, 21, 0) {real, imag} */,
  {32'h417dd74f, 32'hc0ffc88c} /* (13, 20, 31) {real, imag} */,
  {32'hc08a0feb, 32'hc1160ccd} /* (13, 20, 30) {real, imag} */,
  {32'h40da1ee7, 32'hc069a56a} /* (13, 20, 29) {real, imag} */,
  {32'h40992131, 32'h411b2403} /* (13, 20, 28) {real, imag} */,
  {32'hc0bd8fc8, 32'h41172f61} /* (13, 20, 27) {real, imag} */,
  {32'hbf57901c, 32'h410c0bc6} /* (13, 20, 26) {real, imag} */,
  {32'h3fc36848, 32'hc10e1f20} /* (13, 20, 25) {real, imag} */,
  {32'h41371681, 32'h41be037c} /* (13, 20, 24) {real, imag} */,
  {32'h412217ba, 32'hc0291fee} /* (13, 20, 23) {real, imag} */,
  {32'h4193741a, 32'hc1134163} /* (13, 20, 22) {real, imag} */,
  {32'h3f92aac6, 32'hbfa2a7d8} /* (13, 20, 21) {real, imag} */,
  {32'hc19831b2, 32'h40dcea3e} /* (13, 20, 20) {real, imag} */,
  {32'h40c512d5, 32'h4025ad64} /* (13, 20, 19) {real, imag} */,
  {32'hc12abd7b, 32'hbeacac80} /* (13, 20, 18) {real, imag} */,
  {32'h40fd51f2, 32'hc115e1fa} /* (13, 20, 17) {real, imag} */,
  {32'h414256c7, 32'hbdfa4e60} /* (13, 20, 16) {real, imag} */,
  {32'hc187c8cd, 32'hbfb3ed4e} /* (13, 20, 15) {real, imag} */,
  {32'hc04b03c4, 32'h41819fd7} /* (13, 20, 14) {real, imag} */,
  {32'h40046a60, 32'h40f352dc} /* (13, 20, 13) {real, imag} */,
  {32'hc07c01e5, 32'hc0e1b8c2} /* (13, 20, 12) {real, imag} */,
  {32'h4189a971, 32'hc09101f4} /* (13, 20, 11) {real, imag} */,
  {32'hc15799aa, 32'hc1225968} /* (13, 20, 10) {real, imag} */,
  {32'h41018a04, 32'h4199007c} /* (13, 20, 9) {real, imag} */,
  {32'h3f7e79e0, 32'h40a2e54e} /* (13, 20, 8) {real, imag} */,
  {32'h40ad3606, 32'h410e89d7} /* (13, 20, 7) {real, imag} */,
  {32'hc1200f58, 32'h4125303a} /* (13, 20, 6) {real, imag} */,
  {32'h4016ccbf, 32'hc1629c9c} /* (13, 20, 5) {real, imag} */,
  {32'h404cd2bc, 32'h40202eae} /* (13, 20, 4) {real, imag} */,
  {32'h409acb6b, 32'h40a7677b} /* (13, 20, 3) {real, imag} */,
  {32'h4118bb7a, 32'hc10f194c} /* (13, 20, 2) {real, imag} */,
  {32'hc0f714dd, 32'hc1420c3a} /* (13, 20, 1) {real, imag} */,
  {32'h411577c5, 32'hc0be5094} /* (13, 20, 0) {real, imag} */,
  {32'hbf577128, 32'hc10e54f4} /* (13, 19, 31) {real, imag} */,
  {32'h414d7fca, 32'h40227610} /* (13, 19, 30) {real, imag} */,
  {32'hc0c0ccfa, 32'hc0d00e12} /* (13, 19, 29) {real, imag} */,
  {32'h40ed2ce4, 32'h413f26f6} /* (13, 19, 28) {real, imag} */,
  {32'h408bdb40, 32'hc09f1380} /* (13, 19, 27) {real, imag} */,
  {32'hc169dc64, 32'hbf7449ff} /* (13, 19, 26) {real, imag} */,
  {32'h418b46ce, 32'h3f8d89be} /* (13, 19, 25) {real, imag} */,
  {32'hc1096f89, 32'hbe0a9530} /* (13, 19, 24) {real, imag} */,
  {32'h419370d2, 32'hc1403763} /* (13, 19, 23) {real, imag} */,
  {32'h3ff72da0, 32'hc18ac702} /* (13, 19, 22) {real, imag} */,
  {32'h418f5569, 32'h4199e6de} /* (13, 19, 21) {real, imag} */,
  {32'hc14e3f00, 32'h4151db15} /* (13, 19, 20) {real, imag} */,
  {32'hc0df2ce5, 32'h40a79e87} /* (13, 19, 19) {real, imag} */,
  {32'hc1196368, 32'h40c79c64} /* (13, 19, 18) {real, imag} */,
  {32'h410bdef0, 32'hbfdbdf38} /* (13, 19, 17) {real, imag} */,
  {32'h4009ee53, 32'hc004d1d2} /* (13, 19, 16) {real, imag} */,
  {32'hc0e88e7a, 32'hc0c9c748} /* (13, 19, 15) {real, imag} */,
  {32'hc088c2fc, 32'hc1092e43} /* (13, 19, 14) {real, imag} */,
  {32'h408cf60d, 32'h414de788} /* (13, 19, 13) {real, imag} */,
  {32'h41140bfc, 32'hc19850d8} /* (13, 19, 12) {real, imag} */,
  {32'hc0e44154, 32'h3d8bc040} /* (13, 19, 11) {real, imag} */,
  {32'h411d8683, 32'h40802bf2} /* (13, 19, 10) {real, imag} */,
  {32'hc159ff89, 32'h41b57e97} /* (13, 19, 9) {real, imag} */,
  {32'h3e02ff60, 32'h40df9bc2} /* (13, 19, 8) {real, imag} */,
  {32'hbba1f800, 32'h414d6056} /* (13, 19, 7) {real, imag} */,
  {32'h407ef437, 32'hc0f68747} /* (13, 19, 6) {real, imag} */,
  {32'h3e5fc4e0, 32'h4071bf63} /* (13, 19, 5) {real, imag} */,
  {32'h3e360550, 32'hbff866a0} /* (13, 19, 4) {real, imag} */,
  {32'hc0a8e77a, 32'hc0ac6b89} /* (13, 19, 3) {real, imag} */,
  {32'h4025c2fe, 32'h4105f5b2} /* (13, 19, 2) {real, imag} */,
  {32'h410d8ba8, 32'h3ff57bee} /* (13, 19, 1) {real, imag} */,
  {32'hc0be72e7, 32'hc1201e94} /* (13, 19, 0) {real, imag} */,
  {32'hc0cc06da, 32'h40de18c0} /* (13, 18, 31) {real, imag} */,
  {32'hc1342df6, 32'h40266c61} /* (13, 18, 30) {real, imag} */,
  {32'h405ad5c6, 32'hc1381d8f} /* (13, 18, 29) {real, imag} */,
  {32'h3fd4ab8a, 32'h40a0e2de} /* (13, 18, 28) {real, imag} */,
  {32'hbfb01364, 32'h41186912} /* (13, 18, 27) {real, imag} */,
  {32'h40f724b4, 32'h4145a8c8} /* (13, 18, 26) {real, imag} */,
  {32'h4067134b, 32'hc0464a78} /* (13, 18, 25) {real, imag} */,
  {32'h4198e5ce, 32'h40fedd0b} /* (13, 18, 24) {real, imag} */,
  {32'h4107939f, 32'hc0bedeaa} /* (13, 18, 23) {real, imag} */,
  {32'h40c9e630, 32'hc0d5e684} /* (13, 18, 22) {real, imag} */,
  {32'hc038c0e2, 32'h415754be} /* (13, 18, 21) {real, imag} */,
  {32'h4153fc98, 32'hc094a579} /* (13, 18, 20) {real, imag} */,
  {32'hbf4a35ec, 32'h40675ae9} /* (13, 18, 19) {real, imag} */,
  {32'hc197d4bb, 32'hc14a884e} /* (13, 18, 18) {real, imag} */,
  {32'h3f2ec848, 32'h41001454} /* (13, 18, 17) {real, imag} */,
  {32'hc0f242fe, 32'h4112f976} /* (13, 18, 16) {real, imag} */,
  {32'hc07678ef, 32'h41602056} /* (13, 18, 15) {real, imag} */,
  {32'h405cf84b, 32'hc092d94d} /* (13, 18, 14) {real, imag} */,
  {32'h4029df13, 32'h40d6e8c6} /* (13, 18, 13) {real, imag} */,
  {32'h41638884, 32'hc0588530} /* (13, 18, 12) {real, imag} */,
  {32'h40ac6de1, 32'hc17d9373} /* (13, 18, 11) {real, imag} */,
  {32'h40f8ddf3, 32'hc07feecf} /* (13, 18, 10) {real, imag} */,
  {32'hc0becf51, 32'hc138e88d} /* (13, 18, 9) {real, imag} */,
  {32'h40b8dec9, 32'h40a961fe} /* (13, 18, 8) {real, imag} */,
  {32'hbff591dd, 32'h41524851} /* (13, 18, 7) {real, imag} */,
  {32'hc1073512, 32'hc12f93c2} /* (13, 18, 6) {real, imag} */,
  {32'h407e47ed, 32'h40f5d1b9} /* (13, 18, 5) {real, imag} */,
  {32'hc0099b6d, 32'h4068024c} /* (13, 18, 4) {real, imag} */,
  {32'hbf03d60e, 32'hc0f6715a} /* (13, 18, 3) {real, imag} */,
  {32'h4013633c, 32'hc0fe5396} /* (13, 18, 2) {real, imag} */,
  {32'hbf869910, 32'h41213749} /* (13, 18, 1) {real, imag} */,
  {32'h414368f6, 32'hc021809a} /* (13, 18, 0) {real, imag} */,
  {32'hc002e4c3, 32'hc0b4d510} /* (13, 17, 31) {real, imag} */,
  {32'hbf20749a, 32'h3ffb6ff4} /* (13, 17, 30) {real, imag} */,
  {32'hc0ae56c0, 32'h3f689162} /* (13, 17, 29) {real, imag} */,
  {32'hbf336080, 32'h4103cfdb} /* (13, 17, 28) {real, imag} */,
  {32'h40d9ea56, 32'hc08d647c} /* (13, 17, 27) {real, imag} */,
  {32'hc03dd78c, 32'h40933e4c} /* (13, 17, 26) {real, imag} */,
  {32'hbe44fa00, 32'h3fb3b460} /* (13, 17, 25) {real, imag} */,
  {32'h400c08e7, 32'hc02c70a5} /* (13, 17, 24) {real, imag} */,
  {32'hbf3a45e0, 32'h40f16a8c} /* (13, 17, 23) {real, imag} */,
  {32'hc14cbf40, 32'hc0a29c18} /* (13, 17, 22) {real, imag} */,
  {32'h40623768, 32'hc132a45c} /* (13, 17, 21) {real, imag} */,
  {32'h41284c1f, 32'hc0e2201f} /* (13, 17, 20) {real, imag} */,
  {32'h4173e296, 32'h41234b35} /* (13, 17, 19) {real, imag} */,
  {32'hc000bb80, 32'hc0e31441} /* (13, 17, 18) {real, imag} */,
  {32'h408e47a4, 32'h40fdc46f} /* (13, 17, 17) {real, imag} */,
  {32'h40498102, 32'hc165651c} /* (13, 17, 16) {real, imag} */,
  {32'h4177f109, 32'h3c0cfd00} /* (13, 17, 15) {real, imag} */,
  {32'h407ed566, 32'hbf801847} /* (13, 17, 14) {real, imag} */,
  {32'h3f3526e8, 32'h40e99656} /* (13, 17, 13) {real, imag} */,
  {32'hc0906268, 32'h3e2540c0} /* (13, 17, 12) {real, imag} */,
  {32'hbb5f6600, 32'h40f65f3e} /* (13, 17, 11) {real, imag} */,
  {32'hc0418bcd, 32'h415fef96} /* (13, 17, 10) {real, imag} */,
  {32'h40cabc93, 32'h40a4dd00} /* (13, 17, 9) {real, imag} */,
  {32'h40ce3534, 32'hc115c48a} /* (13, 17, 8) {real, imag} */,
  {32'h40c084a6, 32'h40111c80} /* (13, 17, 7) {real, imag} */,
  {32'h3ed06588, 32'hc00b80b8} /* (13, 17, 6) {real, imag} */,
  {32'hbed064e0, 32'h40318b88} /* (13, 17, 5) {real, imag} */,
  {32'hc02dd383, 32'hc08732db} /* (13, 17, 4) {real, imag} */,
  {32'h407f7780, 32'hc17e5476} /* (13, 17, 3) {real, imag} */,
  {32'hc0c29cbb, 32'hc10d56aa} /* (13, 17, 2) {real, imag} */,
  {32'hc0e2ec0d, 32'hbfb5c15d} /* (13, 17, 1) {real, imag} */,
  {32'hc01ffe99, 32'hc1917b54} /* (13, 17, 0) {real, imag} */,
  {32'hc0a90dca, 32'hc089a814} /* (13, 16, 31) {real, imag} */,
  {32'hc034709d, 32'hc09296ad} /* (13, 16, 30) {real, imag} */,
  {32'hc0ad5425, 32'hc13c1497} /* (13, 16, 29) {real, imag} */,
  {32'h3e0f268c, 32'hc1098ede} /* (13, 16, 28) {real, imag} */,
  {32'h411624b4, 32'h4090476c} /* (13, 16, 27) {real, imag} */,
  {32'hc05105e4, 32'h40a57725} /* (13, 16, 26) {real, imag} */,
  {32'hc13975ce, 32'h3fb0b5f2} /* (13, 16, 25) {real, imag} */,
  {32'h3e2ddba0, 32'hc0bed29e} /* (13, 16, 24) {real, imag} */,
  {32'h4000c653, 32'hc1827f50} /* (13, 16, 23) {real, imag} */,
  {32'h40e430da, 32'hc0b2d6a3} /* (13, 16, 22) {real, imag} */,
  {32'h40a9cb18, 32'hc10bf90a} /* (13, 16, 21) {real, imag} */,
  {32'hc0e90af8, 32'h40d948a0} /* (13, 16, 20) {real, imag} */,
  {32'hc18eb076, 32'hc0d4038b} /* (13, 16, 19) {real, imag} */,
  {32'hc019ef09, 32'hc159b9cf} /* (13, 16, 18) {real, imag} */,
  {32'h40fbc62e, 32'h40812948} /* (13, 16, 17) {real, imag} */,
  {32'hc0cf80e2, 32'h00000000} /* (13, 16, 16) {real, imag} */,
  {32'h40fbc62e, 32'hc0812948} /* (13, 16, 15) {real, imag} */,
  {32'hc019ef09, 32'h4159b9cf} /* (13, 16, 14) {real, imag} */,
  {32'hc18eb076, 32'h40d4038b} /* (13, 16, 13) {real, imag} */,
  {32'hc0e90af8, 32'hc0d948a0} /* (13, 16, 12) {real, imag} */,
  {32'h40a9cb18, 32'h410bf90a} /* (13, 16, 11) {real, imag} */,
  {32'h40e430da, 32'h40b2d6a3} /* (13, 16, 10) {real, imag} */,
  {32'h4000c653, 32'h41827f50} /* (13, 16, 9) {real, imag} */,
  {32'h3e2ddba0, 32'h40bed29e} /* (13, 16, 8) {real, imag} */,
  {32'hc13975ce, 32'hbfb0b5f2} /* (13, 16, 7) {real, imag} */,
  {32'hc05105e4, 32'hc0a57725} /* (13, 16, 6) {real, imag} */,
  {32'h411624b4, 32'hc090476c} /* (13, 16, 5) {real, imag} */,
  {32'h3e0f268c, 32'h41098ede} /* (13, 16, 4) {real, imag} */,
  {32'hc0ad5425, 32'h413c1497} /* (13, 16, 3) {real, imag} */,
  {32'hc034709d, 32'h409296ad} /* (13, 16, 2) {real, imag} */,
  {32'hc0a90dca, 32'h4089a814} /* (13, 16, 1) {real, imag} */,
  {32'h410812b7, 32'h00000000} /* (13, 16, 0) {real, imag} */,
  {32'hc0e2ec0d, 32'h3fb5c15d} /* (13, 15, 31) {real, imag} */,
  {32'hc0c29cbb, 32'h410d56aa} /* (13, 15, 30) {real, imag} */,
  {32'h407f7780, 32'h417e5476} /* (13, 15, 29) {real, imag} */,
  {32'hc02dd383, 32'h408732db} /* (13, 15, 28) {real, imag} */,
  {32'hbed064e0, 32'hc0318b88} /* (13, 15, 27) {real, imag} */,
  {32'h3ed06588, 32'h400b80b8} /* (13, 15, 26) {real, imag} */,
  {32'h40c084a6, 32'hc0111c80} /* (13, 15, 25) {real, imag} */,
  {32'h40ce3534, 32'h4115c48a} /* (13, 15, 24) {real, imag} */,
  {32'h40cabc93, 32'hc0a4dd00} /* (13, 15, 23) {real, imag} */,
  {32'hc0418bcd, 32'hc15fef96} /* (13, 15, 22) {real, imag} */,
  {32'hbb5f6600, 32'hc0f65f3e} /* (13, 15, 21) {real, imag} */,
  {32'hc0906268, 32'hbe2540c0} /* (13, 15, 20) {real, imag} */,
  {32'h3f3526e8, 32'hc0e99656} /* (13, 15, 19) {real, imag} */,
  {32'h407ed566, 32'h3f801847} /* (13, 15, 18) {real, imag} */,
  {32'h4177f109, 32'hbc0cfd00} /* (13, 15, 17) {real, imag} */,
  {32'h40498102, 32'h4165651c} /* (13, 15, 16) {real, imag} */,
  {32'h408e47a4, 32'hc0fdc46f} /* (13, 15, 15) {real, imag} */,
  {32'hc000bb80, 32'h40e31441} /* (13, 15, 14) {real, imag} */,
  {32'h4173e296, 32'hc1234b35} /* (13, 15, 13) {real, imag} */,
  {32'h41284c1f, 32'h40e2201f} /* (13, 15, 12) {real, imag} */,
  {32'h40623768, 32'h4132a45c} /* (13, 15, 11) {real, imag} */,
  {32'hc14cbf40, 32'h40a29c18} /* (13, 15, 10) {real, imag} */,
  {32'hbf3a45e0, 32'hc0f16a8c} /* (13, 15, 9) {real, imag} */,
  {32'h400c08e7, 32'h402c70a5} /* (13, 15, 8) {real, imag} */,
  {32'hbe44fa00, 32'hbfb3b460} /* (13, 15, 7) {real, imag} */,
  {32'hc03dd78c, 32'hc0933e4c} /* (13, 15, 6) {real, imag} */,
  {32'h40d9ea56, 32'h408d647c} /* (13, 15, 5) {real, imag} */,
  {32'hbf336080, 32'hc103cfdb} /* (13, 15, 4) {real, imag} */,
  {32'hc0ae56c0, 32'hbf689162} /* (13, 15, 3) {real, imag} */,
  {32'hbf20749a, 32'hbffb6ff4} /* (13, 15, 2) {real, imag} */,
  {32'hc002e4c3, 32'h40b4d510} /* (13, 15, 1) {real, imag} */,
  {32'hc01ffe99, 32'h41917b54} /* (13, 15, 0) {real, imag} */,
  {32'hbf869910, 32'hc1213749} /* (13, 14, 31) {real, imag} */,
  {32'h4013633c, 32'h40fe5396} /* (13, 14, 30) {real, imag} */,
  {32'hbf03d60e, 32'h40f6715a} /* (13, 14, 29) {real, imag} */,
  {32'hc0099b6d, 32'hc068024c} /* (13, 14, 28) {real, imag} */,
  {32'h407e47ed, 32'hc0f5d1b9} /* (13, 14, 27) {real, imag} */,
  {32'hc1073512, 32'h412f93c2} /* (13, 14, 26) {real, imag} */,
  {32'hbff591dd, 32'hc1524851} /* (13, 14, 25) {real, imag} */,
  {32'h40b8dec9, 32'hc0a961fe} /* (13, 14, 24) {real, imag} */,
  {32'hc0becf51, 32'h4138e88d} /* (13, 14, 23) {real, imag} */,
  {32'h40f8ddf3, 32'h407feecf} /* (13, 14, 22) {real, imag} */,
  {32'h40ac6de1, 32'h417d9373} /* (13, 14, 21) {real, imag} */,
  {32'h41638884, 32'h40588530} /* (13, 14, 20) {real, imag} */,
  {32'h4029df13, 32'hc0d6e8c6} /* (13, 14, 19) {real, imag} */,
  {32'h405cf84b, 32'h4092d94d} /* (13, 14, 18) {real, imag} */,
  {32'hc07678ef, 32'hc1602056} /* (13, 14, 17) {real, imag} */,
  {32'hc0f242fe, 32'hc112f976} /* (13, 14, 16) {real, imag} */,
  {32'h3f2ec848, 32'hc1001454} /* (13, 14, 15) {real, imag} */,
  {32'hc197d4bb, 32'h414a884e} /* (13, 14, 14) {real, imag} */,
  {32'hbf4a35ec, 32'hc0675ae9} /* (13, 14, 13) {real, imag} */,
  {32'h4153fc98, 32'h4094a579} /* (13, 14, 12) {real, imag} */,
  {32'hc038c0e2, 32'hc15754be} /* (13, 14, 11) {real, imag} */,
  {32'h40c9e630, 32'h40d5e684} /* (13, 14, 10) {real, imag} */,
  {32'h4107939f, 32'h40bedeaa} /* (13, 14, 9) {real, imag} */,
  {32'h4198e5ce, 32'hc0fedd0b} /* (13, 14, 8) {real, imag} */,
  {32'h4067134b, 32'h40464a78} /* (13, 14, 7) {real, imag} */,
  {32'h40f724b4, 32'hc145a8c8} /* (13, 14, 6) {real, imag} */,
  {32'hbfb01364, 32'hc1186912} /* (13, 14, 5) {real, imag} */,
  {32'h3fd4ab8a, 32'hc0a0e2de} /* (13, 14, 4) {real, imag} */,
  {32'h405ad5c6, 32'h41381d8f} /* (13, 14, 3) {real, imag} */,
  {32'hc1342df6, 32'hc0266c61} /* (13, 14, 2) {real, imag} */,
  {32'hc0cc06da, 32'hc0de18c0} /* (13, 14, 1) {real, imag} */,
  {32'h414368f6, 32'h4021809a} /* (13, 14, 0) {real, imag} */,
  {32'h410d8ba8, 32'hbff57bee} /* (13, 13, 31) {real, imag} */,
  {32'h4025c2fe, 32'hc105f5b2} /* (13, 13, 30) {real, imag} */,
  {32'hc0a8e77a, 32'h40ac6b89} /* (13, 13, 29) {real, imag} */,
  {32'h3e360550, 32'h3ff866a0} /* (13, 13, 28) {real, imag} */,
  {32'h3e5fc4e0, 32'hc071bf63} /* (13, 13, 27) {real, imag} */,
  {32'h407ef437, 32'h40f68747} /* (13, 13, 26) {real, imag} */,
  {32'hbba1f800, 32'hc14d6056} /* (13, 13, 25) {real, imag} */,
  {32'h3e02ff60, 32'hc0df9bc2} /* (13, 13, 24) {real, imag} */,
  {32'hc159ff89, 32'hc1b57e97} /* (13, 13, 23) {real, imag} */,
  {32'h411d8683, 32'hc0802bf2} /* (13, 13, 22) {real, imag} */,
  {32'hc0e44154, 32'hbd8bc040} /* (13, 13, 21) {real, imag} */,
  {32'h41140bfc, 32'h419850d8} /* (13, 13, 20) {real, imag} */,
  {32'h408cf60d, 32'hc14de788} /* (13, 13, 19) {real, imag} */,
  {32'hc088c2fc, 32'h41092e43} /* (13, 13, 18) {real, imag} */,
  {32'hc0e88e7a, 32'h40c9c748} /* (13, 13, 17) {real, imag} */,
  {32'h4009ee53, 32'h4004d1d2} /* (13, 13, 16) {real, imag} */,
  {32'h410bdef0, 32'h3fdbdf38} /* (13, 13, 15) {real, imag} */,
  {32'hc1196368, 32'hc0c79c64} /* (13, 13, 14) {real, imag} */,
  {32'hc0df2ce5, 32'hc0a79e87} /* (13, 13, 13) {real, imag} */,
  {32'hc14e3f00, 32'hc151db15} /* (13, 13, 12) {real, imag} */,
  {32'h418f5569, 32'hc199e6de} /* (13, 13, 11) {real, imag} */,
  {32'h3ff72da0, 32'h418ac702} /* (13, 13, 10) {real, imag} */,
  {32'h419370d2, 32'h41403763} /* (13, 13, 9) {real, imag} */,
  {32'hc1096f89, 32'h3e0a9530} /* (13, 13, 8) {real, imag} */,
  {32'h418b46ce, 32'hbf8d89be} /* (13, 13, 7) {real, imag} */,
  {32'hc169dc64, 32'h3f7449ff} /* (13, 13, 6) {real, imag} */,
  {32'h408bdb40, 32'h409f1380} /* (13, 13, 5) {real, imag} */,
  {32'h40ed2ce4, 32'hc13f26f6} /* (13, 13, 4) {real, imag} */,
  {32'hc0c0ccfa, 32'h40d00e12} /* (13, 13, 3) {real, imag} */,
  {32'h414d7fca, 32'hc0227610} /* (13, 13, 2) {real, imag} */,
  {32'hbf577128, 32'h410e54f4} /* (13, 13, 1) {real, imag} */,
  {32'hc0be72e7, 32'h41201e94} /* (13, 13, 0) {real, imag} */,
  {32'hc0f714dd, 32'h41420c3a} /* (13, 12, 31) {real, imag} */,
  {32'h4118bb7a, 32'h410f194c} /* (13, 12, 30) {real, imag} */,
  {32'h409acb6b, 32'hc0a7677b} /* (13, 12, 29) {real, imag} */,
  {32'h404cd2bc, 32'hc0202eae} /* (13, 12, 28) {real, imag} */,
  {32'h4016ccbf, 32'h41629c9c} /* (13, 12, 27) {real, imag} */,
  {32'hc1200f58, 32'hc125303a} /* (13, 12, 26) {real, imag} */,
  {32'h40ad3606, 32'hc10e89d7} /* (13, 12, 25) {real, imag} */,
  {32'h3f7e79e0, 32'hc0a2e54e} /* (13, 12, 24) {real, imag} */,
  {32'h41018a04, 32'hc199007c} /* (13, 12, 23) {real, imag} */,
  {32'hc15799aa, 32'h41225968} /* (13, 12, 22) {real, imag} */,
  {32'h4189a971, 32'h409101f4} /* (13, 12, 21) {real, imag} */,
  {32'hc07c01e5, 32'h40e1b8c2} /* (13, 12, 20) {real, imag} */,
  {32'h40046a60, 32'hc0f352dc} /* (13, 12, 19) {real, imag} */,
  {32'hc04b03c4, 32'hc1819fd7} /* (13, 12, 18) {real, imag} */,
  {32'hc187c8cd, 32'h3fb3ed4e} /* (13, 12, 17) {real, imag} */,
  {32'h414256c7, 32'h3dfa4e60} /* (13, 12, 16) {real, imag} */,
  {32'h40fd51f2, 32'h4115e1fa} /* (13, 12, 15) {real, imag} */,
  {32'hc12abd7b, 32'h3eacac80} /* (13, 12, 14) {real, imag} */,
  {32'h40c512d5, 32'hc025ad64} /* (13, 12, 13) {real, imag} */,
  {32'hc19831b2, 32'hc0dcea3e} /* (13, 12, 12) {real, imag} */,
  {32'h3f92aac6, 32'h3fa2a7d8} /* (13, 12, 11) {real, imag} */,
  {32'h4193741a, 32'h41134163} /* (13, 12, 10) {real, imag} */,
  {32'h412217ba, 32'h40291fee} /* (13, 12, 9) {real, imag} */,
  {32'h41371681, 32'hc1be037c} /* (13, 12, 8) {real, imag} */,
  {32'h3fc36848, 32'h410e1f20} /* (13, 12, 7) {real, imag} */,
  {32'hbf57901c, 32'hc10c0bc6} /* (13, 12, 6) {real, imag} */,
  {32'hc0bd8fc8, 32'hc1172f61} /* (13, 12, 5) {real, imag} */,
  {32'h40992131, 32'hc11b2403} /* (13, 12, 4) {real, imag} */,
  {32'h40da1ee7, 32'h4069a56a} /* (13, 12, 3) {real, imag} */,
  {32'hc08a0feb, 32'h41160ccd} /* (13, 12, 2) {real, imag} */,
  {32'h417dd74f, 32'h40ffc88c} /* (13, 12, 1) {real, imag} */,
  {32'h411577c5, 32'h40be5094} /* (13, 12, 0) {real, imag} */,
  {32'hc18dfeed, 32'hc0a2fd42} /* (13, 11, 31) {real, imag} */,
  {32'hc0841063, 32'h41951ef5} /* (13, 11, 30) {real, imag} */,
  {32'h4126345a, 32'hc0f9e231} /* (13, 11, 29) {real, imag} */,
  {32'hc0579494, 32'h40d9dc14} /* (13, 11, 28) {real, imag} */,
  {32'h4204d9dc, 32'h4184f27a} /* (13, 11, 27) {real, imag} */,
  {32'hc01f3a3c, 32'hbf727d84} /* (13, 11, 26) {real, imag} */,
  {32'h411f9d51, 32'hc1acde1a} /* (13, 11, 25) {real, imag} */,
  {32'hc11680e4, 32'hc198614e} /* (13, 11, 24) {real, imag} */,
  {32'h40c30698, 32'hc12324b2} /* (13, 11, 23) {real, imag} */,
  {32'hc0498028, 32'hc126a11d} /* (13, 11, 22) {real, imag} */,
  {32'hc03fdb08, 32'h40d1e87f} /* (13, 11, 21) {real, imag} */,
  {32'h419794b1, 32'h410f9875} /* (13, 11, 20) {real, imag} */,
  {32'h3f8a85a6, 32'hc096c683} /* (13, 11, 19) {real, imag} */,
  {32'hc0c3e76e, 32'h4099ed15} /* (13, 11, 18) {real, imag} */,
  {32'h408754f7, 32'h4049a734} /* (13, 11, 17) {real, imag} */,
  {32'hc02b358d, 32'hc11f04ac} /* (13, 11, 16) {real, imag} */,
  {32'hbfa69eec, 32'h40bc3a6c} /* (13, 11, 15) {real, imag} */,
  {32'h40c3b4ba, 32'h4100818e} /* (13, 11, 14) {real, imag} */,
  {32'h41023aed, 32'hc0b2ac36} /* (13, 11, 13) {real, imag} */,
  {32'hc153cf73, 32'hc08dac17} /* (13, 11, 12) {real, imag} */,
  {32'hc0ce0f58, 32'hc024e4db} /* (13, 11, 11) {real, imag} */,
  {32'h4001ff48, 32'hc1b62de9} /* (13, 11, 10) {real, imag} */,
  {32'h4181cddc, 32'hc108e343} /* (13, 11, 9) {real, imag} */,
  {32'h418ec45d, 32'hc0503761} /* (13, 11, 8) {real, imag} */,
  {32'hc0a5dc36, 32'hc11a48fa} /* (13, 11, 7) {real, imag} */,
  {32'hc0c105f6, 32'h41177122} /* (13, 11, 6) {real, imag} */,
  {32'h40cd29f8, 32'h40407806} /* (13, 11, 5) {real, imag} */,
  {32'h3f9bb8ea, 32'hc189e496} /* (13, 11, 4) {real, imag} */,
  {32'h4124024d, 32'hc13c1d6d} /* (13, 11, 3) {real, imag} */,
  {32'hc1cb90c4, 32'h40c25e86} /* (13, 11, 2) {real, imag} */,
  {32'hc1339b49, 32'hc1265f06} /* (13, 11, 1) {real, imag} */,
  {32'hc1a3ae54, 32'hc15b33d4} /* (13, 11, 0) {real, imag} */,
  {32'hbff30f36, 32'h41a14af6} /* (13, 10, 31) {real, imag} */,
  {32'h412494da, 32'hc13e2712} /* (13, 10, 30) {real, imag} */,
  {32'hc0a7593d, 32'hc005be93} /* (13, 10, 29) {real, imag} */,
  {32'h40294be6, 32'hc19b0f5b} /* (13, 10, 28) {real, imag} */,
  {32'h40df293c, 32'h41321a0b} /* (13, 10, 27) {real, imag} */,
  {32'h40c4d813, 32'h41711c7e} /* (13, 10, 26) {real, imag} */,
  {32'hc135893a, 32'h401277a2} /* (13, 10, 25) {real, imag} */,
  {32'hc107b5ba, 32'h40be29d8} /* (13, 10, 24) {real, imag} */,
  {32'h40cf7b84, 32'hbdbacf40} /* (13, 10, 23) {real, imag} */,
  {32'h40d484eb, 32'hc10c8177} /* (13, 10, 22) {real, imag} */,
  {32'hc127cfd8, 32'h400d4ed0} /* (13, 10, 21) {real, imag} */,
  {32'hc16f42cc, 32'h40490442} /* (13, 10, 20) {real, imag} */,
  {32'h3f820a7c, 32'h41b469d6} /* (13, 10, 19) {real, imag} */,
  {32'hc11fe6e2, 32'h3e65d1d0} /* (13, 10, 18) {real, imag} */,
  {32'h412a81dc, 32'h3fa96c30} /* (13, 10, 17) {real, imag} */,
  {32'h410cbc64, 32'h410898c4} /* (13, 10, 16) {real, imag} */,
  {32'h40997282, 32'h41847c52} /* (13, 10, 15) {real, imag} */,
  {32'hc11572b4, 32'hc19b9d76} /* (13, 10, 14) {real, imag} */,
  {32'hc140b2da, 32'hbf677738} /* (13, 10, 13) {real, imag} */,
  {32'hc1d2cade, 32'h40323997} /* (13, 10, 12) {real, imag} */,
  {32'h41a6130f, 32'h410f9e3a} /* (13, 10, 11) {real, imag} */,
  {32'hbf95e1b8, 32'hc10abcfb} /* (13, 10, 10) {real, imag} */,
  {32'h4180c720, 32'hc0ce1d96} /* (13, 10, 9) {real, imag} */,
  {32'hc1b72f7e, 32'h41913b78} /* (13, 10, 8) {real, imag} */,
  {32'h41bcdc03, 32'h40cb21b2} /* (13, 10, 7) {real, imag} */,
  {32'hc18819c7, 32'h408e4ff8} /* (13, 10, 6) {real, imag} */,
  {32'h40354b56, 32'h410bc7c1} /* (13, 10, 5) {real, imag} */,
  {32'h41946580, 32'h3fa180c8} /* (13, 10, 4) {real, imag} */,
  {32'hc0c2680c, 32'hc1582738} /* (13, 10, 3) {real, imag} */,
  {32'hbf8666a0, 32'hc1aeea29} /* (13, 10, 2) {real, imag} */,
  {32'h41adc711, 32'h40455a7c} /* (13, 10, 1) {real, imag} */,
  {32'h413196e6, 32'h415bb700} /* (13, 10, 0) {real, imag} */,
  {32'h3ef59ad0, 32'h415f00bd} /* (13, 9, 31) {real, imag} */,
  {32'h41a18c14, 32'hc166f0fe} /* (13, 9, 30) {real, imag} */,
  {32'h4159941a, 32'h3eba3180} /* (13, 9, 29) {real, imag} */,
  {32'h41c802d2, 32'hc0b72d2a} /* (13, 9, 28) {real, imag} */,
  {32'hc18fadd6, 32'h40ff303e} /* (13, 9, 27) {real, imag} */,
  {32'hbf0a5f70, 32'h4034fcf9} /* (13, 9, 26) {real, imag} */,
  {32'hc1024eaf, 32'hc092e09c} /* (13, 9, 25) {real, imag} */,
  {32'hc037ded2, 32'h4186331b} /* (13, 9, 24) {real, imag} */,
  {32'h418e1bf5, 32'h415be339} /* (13, 9, 23) {real, imag} */,
  {32'hc02645ae, 32'h40c5fc3f} /* (13, 9, 22) {real, imag} */,
  {32'hc19c89b2, 32'hc0241e4d} /* (13, 9, 21) {real, imag} */,
  {32'h40744b37, 32'hc141a116} /* (13, 9, 20) {real, imag} */,
  {32'h4103ac4e, 32'h3ed32780} /* (13, 9, 19) {real, imag} */,
  {32'hc0a1cd9e, 32'hc10dddbe} /* (13, 9, 18) {real, imag} */,
  {32'hc14002a4, 32'h41877b3f} /* (13, 9, 17) {real, imag} */,
  {32'hc0eabf9a, 32'h4127d7c8} /* (13, 9, 16) {real, imag} */,
  {32'hc12a80fb, 32'hc101612c} /* (13, 9, 15) {real, imag} */,
  {32'h41b1bf8d, 32'hbf83d4b8} /* (13, 9, 14) {real, imag} */,
  {32'hc01e5efa, 32'h4138f85d} /* (13, 9, 13) {real, imag} */,
  {32'hc0a97dab, 32'h4106ea06} /* (13, 9, 12) {real, imag} */,
  {32'h41424fe6, 32'h3e7b2660} /* (13, 9, 11) {real, imag} */,
  {32'hc12fb682, 32'hc11ac6fa} /* (13, 9, 10) {real, imag} */,
  {32'hc14e9714, 32'h417b700d} /* (13, 9, 9) {real, imag} */,
  {32'hc0570b94, 32'h4082e662} /* (13, 9, 8) {real, imag} */,
  {32'h40c58030, 32'h41df3370} /* (13, 9, 7) {real, imag} */,
  {32'hc15ca715, 32'hc1356770} /* (13, 9, 6) {real, imag} */,
  {32'h41163c95, 32'hc13d15b0} /* (13, 9, 5) {real, imag} */,
  {32'hc1098ff6, 32'h416895be} /* (13, 9, 4) {real, imag} */,
  {32'hbf87f916, 32'hc122b074} /* (13, 9, 3) {real, imag} */,
  {32'hbf84cb04, 32'hc18cea07} /* (13, 9, 2) {real, imag} */,
  {32'hc1080924, 32'h41b4aedd} /* (13, 9, 1) {real, imag} */,
  {32'hc053332f, 32'hc15469e4} /* (13, 9, 0) {real, imag} */,
  {32'hc24f58c9, 32'hc1d8d77e} /* (13, 8, 31) {real, imag} */,
  {32'h419b81c7, 32'h41c1a334} /* (13, 8, 30) {real, imag} */,
  {32'h41aeb311, 32'hc1a33ae5} /* (13, 8, 29) {real, imag} */,
  {32'h3d88a380, 32'h41c8c3f1} /* (13, 8, 28) {real, imag} */,
  {32'h41fc592c, 32'h40d03528} /* (13, 8, 27) {real, imag} */,
  {32'hc026b85a, 32'hc11b6cd0} /* (13, 8, 26) {real, imag} */,
  {32'h413a8a2f, 32'hbe140f88} /* (13, 8, 25) {real, imag} */,
  {32'h4208647e, 32'hc10d5614} /* (13, 8, 24) {real, imag} */,
  {32'h40bc2698, 32'h41160ba1} /* (13, 8, 23) {real, imag} */,
  {32'hc1ce4388, 32'h41811a72} /* (13, 8, 22) {real, imag} */,
  {32'h416bbe2a, 32'h3fa54296} /* (13, 8, 21) {real, imag} */,
  {32'hc11b07d9, 32'hc083730e} /* (13, 8, 20) {real, imag} */,
  {32'h4134266c, 32'h408cd034} /* (13, 8, 19) {real, imag} */,
  {32'h40671316, 32'h3fcfbf30} /* (13, 8, 18) {real, imag} */,
  {32'hc097df1d, 32'hc0252309} /* (13, 8, 17) {real, imag} */,
  {32'h4006819b, 32'h41d56a2c} /* (13, 8, 16) {real, imag} */,
  {32'h3ff288a8, 32'h406b9f65} /* (13, 8, 15) {real, imag} */,
  {32'h4085cd18, 32'hc1014a58} /* (13, 8, 14) {real, imag} */,
  {32'h4105eec9, 32'hc115ed24} /* (13, 8, 13) {real, imag} */,
  {32'h4137d65b, 32'h411b9e99} /* (13, 8, 12) {real, imag} */,
  {32'h421db97e, 32'hc1737893} /* (13, 8, 11) {real, imag} */,
  {32'hc15c900a, 32'hc0c3f10e} /* (13, 8, 10) {real, imag} */,
  {32'hc1033544, 32'h40a7c22e} /* (13, 8, 9) {real, imag} */,
  {32'h40bc68aa, 32'h405ec6c6} /* (13, 8, 8) {real, imag} */,
  {32'hc0e27e16, 32'hbf743fe4} /* (13, 8, 7) {real, imag} */,
  {32'h417df968, 32'hbff33aa4} /* (13, 8, 6) {real, imag} */,
  {32'hbfe24394, 32'h410d3d73} /* (13, 8, 5) {real, imag} */,
  {32'hc17f26c8, 32'hc1b75150} /* (13, 8, 4) {real, imag} */,
  {32'h41ab6674, 32'hc085acd5} /* (13, 8, 3) {real, imag} */,
  {32'h41ee168a, 32'hc1c566d0} /* (13, 8, 2) {real, imag} */,
  {32'hc22f2eba, 32'hc1c285bf} /* (13, 8, 1) {real, imag} */,
  {32'hc1af2008, 32'hc184792d} /* (13, 8, 0) {real, imag} */,
  {32'h414d5d92, 32'hc0b6d18f} /* (13, 7, 31) {real, imag} */,
  {32'h4123de80, 32'hc13004e8} /* (13, 7, 30) {real, imag} */,
  {32'hc0412d74, 32'hc18d8e94} /* (13, 7, 29) {real, imag} */,
  {32'hc108dfd9, 32'hbe9577b0} /* (13, 7, 28) {real, imag} */,
  {32'hc0feb5ac, 32'h41734fdc} /* (13, 7, 27) {real, imag} */,
  {32'hc0ce8e8b, 32'h3d210700} /* (13, 7, 26) {real, imag} */,
  {32'h410b5e9b, 32'h3f0895f8} /* (13, 7, 25) {real, imag} */,
  {32'h40bf1851, 32'hc00a33e2} /* (13, 7, 24) {real, imag} */,
  {32'h40e3b5a9, 32'hc15238b5} /* (13, 7, 23) {real, imag} */,
  {32'h3fe5382a, 32'h4122babc} /* (13, 7, 22) {real, imag} */,
  {32'hc12d4107, 32'hc164d3b6} /* (13, 7, 21) {real, imag} */,
  {32'h415c767b, 32'h3ead32a0} /* (13, 7, 20) {real, imag} */,
  {32'hc01e3db2, 32'h40f5a208} /* (13, 7, 19) {real, imag} */,
  {32'hc030bc38, 32'h4187df6a} /* (13, 7, 18) {real, imag} */,
  {32'h40b01ccf, 32'h414a9326} /* (13, 7, 17) {real, imag} */,
  {32'hc14d3524, 32'h4091d20c} /* (13, 7, 16) {real, imag} */,
  {32'h40ca45a5, 32'h400b3fe8} /* (13, 7, 15) {real, imag} */,
  {32'h40295782, 32'hbf396acc} /* (13, 7, 14) {real, imag} */,
  {32'h3fd1b3c8, 32'hc1687e1b} /* (13, 7, 13) {real, imag} */,
  {32'h40e93226, 32'hc122d604} /* (13, 7, 12) {real, imag} */,
  {32'hc09a5f72, 32'h3f846b2e} /* (13, 7, 11) {real, imag} */,
  {32'hc0a5bddc, 32'h412ae05d} /* (13, 7, 10) {real, imag} */,
  {32'hc09566b0, 32'h410e7455} /* (13, 7, 9) {real, imag} */,
  {32'hc17e0184, 32'hc0b5bd42} /* (13, 7, 8) {real, imag} */,
  {32'h3ff833a8, 32'hc0234031} /* (13, 7, 7) {real, imag} */,
  {32'h41450506, 32'hbfadf2d8} /* (13, 7, 6) {real, imag} */,
  {32'h4161087c, 32'hc01e804a} /* (13, 7, 5) {real, imag} */,
  {32'hc1a86111, 32'h408cb928} /* (13, 7, 4) {real, imag} */,
  {32'hc0446cfc, 32'h41543637} /* (13, 7, 3) {real, imag} */,
  {32'h4167deae, 32'hc166f549} /* (13, 7, 2) {real, imag} */,
  {32'h4169c74d, 32'h423f104b} /* (13, 7, 1) {real, imag} */,
  {32'hc0c1bbab, 32'h419745c3} /* (13, 7, 0) {real, imag} */,
  {32'hc1664e1a, 32'hc08adba3} /* (13, 6, 31) {real, imag} */,
  {32'h4229db9c, 32'hc1c76efd} /* (13, 6, 30) {real, imag} */,
  {32'h40757450, 32'hc19817bb} /* (13, 6, 29) {real, imag} */,
  {32'hc0ee3792, 32'hc1157319} /* (13, 6, 28) {real, imag} */,
  {32'h41ac914a, 32'h3fe336be} /* (13, 6, 27) {real, imag} */,
  {32'h415bfc44, 32'h40c79ad8} /* (13, 6, 26) {real, imag} */,
  {32'h3ff944b4, 32'hc15b0ebc} /* (13, 6, 25) {real, imag} */,
  {32'h3f849590, 32'h3f4f6850} /* (13, 6, 24) {real, imag} */,
  {32'h400229a9, 32'hc0ce1962} /* (13, 6, 23) {real, imag} */,
  {32'h4055be40, 32'h4198c41e} /* (13, 6, 22) {real, imag} */,
  {32'hbf048af8, 32'hc02a0f5e} /* (13, 6, 21) {real, imag} */,
  {32'hc09db331, 32'h40119c30} /* (13, 6, 20) {real, imag} */,
  {32'h41095335, 32'h413ec5c2} /* (13, 6, 19) {real, imag} */,
  {32'h411bf044, 32'hc137df40} /* (13, 6, 18) {real, imag} */,
  {32'hc09c5098, 32'h3f83a1c8} /* (13, 6, 17) {real, imag} */,
  {32'hc133c81d, 32'hbfa4bdec} /* (13, 6, 16) {real, imag} */,
  {32'h40b8ad38, 32'hc10f9a67} /* (13, 6, 15) {real, imag} */,
  {32'h4103e04a, 32'hc1280c0f} /* (13, 6, 14) {real, imag} */,
  {32'h41835f85, 32'h405c0136} /* (13, 6, 13) {real, imag} */,
  {32'h40764150, 32'hc0159ac3} /* (13, 6, 12) {real, imag} */,
  {32'hbf4e3ed0, 32'h41da7a4e} /* (13, 6, 11) {real, imag} */,
  {32'hc011fb8b, 32'hc1a2e4eb} /* (13, 6, 10) {real, imag} */,
  {32'hc1316944, 32'h415c55bc} /* (13, 6, 9) {real, imag} */,
  {32'h41baa759, 32'h3f9bdf78} /* (13, 6, 8) {real, imag} */,
  {32'hc16fb5fe, 32'h40c11700} /* (13, 6, 7) {real, imag} */,
  {32'hc1543b88, 32'hc1af63c4} /* (13, 6, 6) {real, imag} */,
  {32'hc1ac545c, 32'hc1a2170a} /* (13, 6, 5) {real, imag} */,
  {32'hc1af4012, 32'h4085c350} /* (13, 6, 4) {real, imag} */,
  {32'hbff39ad0, 32'h40f469ec} /* (13, 6, 3) {real, imag} */,
  {32'h41f7b36e, 32'h4149b3ee} /* (13, 6, 2) {real, imag} */,
  {32'hc1c455c4, 32'hc1b2da9a} /* (13, 6, 1) {real, imag} */,
  {32'h40f6795a, 32'h41b60a7b} /* (13, 6, 0) {real, imag} */,
  {32'hc2b63146, 32'hc081a5b4} /* (13, 5, 31) {real, imag} */,
  {32'h41813790, 32'h4138a0b9} /* (13, 5, 30) {real, imag} */,
  {32'h40dc56b6, 32'h41ad358a} /* (13, 5, 29) {real, imag} */,
  {32'hc1972e40, 32'h4106de6e} /* (13, 5, 28) {real, imag} */,
  {32'h4203f2be, 32'h411c3dfb} /* (13, 5, 27) {real, imag} */,
  {32'h412384c4, 32'h4101ae72} /* (13, 5, 26) {real, imag} */,
  {32'h40e1e970, 32'hc12f145e} /* (13, 5, 25) {real, imag} */,
  {32'hbff696ac, 32'hc1a39c88} /* (13, 5, 24) {real, imag} */,
  {32'h3ec89760, 32'h420c54eb} /* (13, 5, 23) {real, imag} */,
  {32'h4111f752, 32'h4042755a} /* (13, 5, 22) {real, imag} */,
  {32'h41878da4, 32'hc0f0f856} /* (13, 5, 21) {real, imag} */,
  {32'hc16795e5, 32'h40f08931} /* (13, 5, 20) {real, imag} */,
  {32'hc13ad052, 32'hc0d59138} /* (13, 5, 19) {real, imag} */,
  {32'h40adddfe, 32'hc0e8ec86} /* (13, 5, 18) {real, imag} */,
  {32'h40cbab56, 32'h3f157c20} /* (13, 5, 17) {real, imag} */,
  {32'hc08e8f1e, 32'hc121450c} /* (13, 5, 16) {real, imag} */,
  {32'hc1b9ec88, 32'h409ed446} /* (13, 5, 15) {real, imag} */,
  {32'h3fd29ed2, 32'h409929b3} /* (13, 5, 14) {real, imag} */,
  {32'hc1167bc6, 32'hc12c0b6e} /* (13, 5, 13) {real, imag} */,
  {32'h41a9452e, 32'hc1dbfb07} /* (13, 5, 12) {real, imag} */,
  {32'h40acc1d8, 32'h4180485e} /* (13, 5, 11) {real, imag} */,
  {32'hbff75528, 32'h4001d2b2} /* (13, 5, 10) {real, imag} */,
  {32'h4175407a, 32'hbf0607c0} /* (13, 5, 9) {real, imag} */,
  {32'hc0dc47e2, 32'h40cb32e7} /* (13, 5, 8) {real, imag} */,
  {32'h411c90d6, 32'hc15b972a} /* (13, 5, 7) {real, imag} */,
  {32'hc0b6526f, 32'h42047398} /* (13, 5, 6) {real, imag} */,
  {32'h412eb203, 32'hbe5f9100} /* (13, 5, 5) {real, imag} */,
  {32'h41173b86, 32'hc14777c2} /* (13, 5, 4) {real, imag} */,
  {32'hc0144124, 32'h41524846} /* (13, 5, 3) {real, imag} */,
  {32'h40e5bdfc, 32'h42162bd2} /* (13, 5, 2) {real, imag} */,
  {32'hc2c6f1cc, 32'hc22f97c2} /* (13, 5, 1) {real, imag} */,
  {32'hc26f3a4c, 32'hc212d780} /* (13, 5, 0) {real, imag} */,
  {32'h42763424, 32'h427eb9e1} /* (13, 4, 31) {real, imag} */,
  {32'hc2ae7a55, 32'hc2a671e1} /* (13, 4, 30) {real, imag} */,
  {32'hc1ae96af, 32'hc1408be4} /* (13, 4, 29) {real, imag} */,
  {32'h4258e3ca, 32'h41ffa87d} /* (13, 4, 28) {real, imag} */,
  {32'hc19a2cce, 32'hc101cccb} /* (13, 4, 27) {real, imag} */,
  {32'hc0d001d2, 32'hc0c8ca52} /* (13, 4, 26) {real, imag} */,
  {32'h40b60ff3, 32'h40feea37} /* (13, 4, 25) {real, imag} */,
  {32'h3fdd60bc, 32'hc1bf91f0} /* (13, 4, 24) {real, imag} */,
  {32'h408589ea, 32'hc18d8598} /* (13, 4, 23) {real, imag} */,
  {32'h40a75a64, 32'hbe133c00} /* (13, 4, 22) {real, imag} */,
  {32'hc162338a, 32'h41164ae7} /* (13, 4, 21) {real, imag} */,
  {32'hc15910d7, 32'hc1522389} /* (13, 4, 20) {real, imag} */,
  {32'h413c092b, 32'hc14bc68e} /* (13, 4, 19) {real, imag} */,
  {32'h40ab6e14, 32'h416ace81} /* (13, 4, 18) {real, imag} */,
  {32'h4117c6a2, 32'hbf210444} /* (13, 4, 17) {real, imag} */,
  {32'h3fdec480, 32'h40bf1d7d} /* (13, 4, 16) {real, imag} */,
  {32'h40de528c, 32'hc0061a46} /* (13, 4, 15) {real, imag} */,
  {32'hbff32c70, 32'hc14bbd1f} /* (13, 4, 14) {real, imag} */,
  {32'h410f1810, 32'hc1182688} /* (13, 4, 13) {real, imag} */,
  {32'hc03c8419, 32'h4135cf08} /* (13, 4, 12) {real, imag} */,
  {32'h41672d82, 32'h405c4be5} /* (13, 4, 11) {real, imag} */,
  {32'hc172e426, 32'h3fd37064} /* (13, 4, 10) {real, imag} */,
  {32'h412bf314, 32'h3e9fd3e0} /* (13, 4, 9) {real, imag} */,
  {32'h3e88b118, 32'hc1a796ce} /* (13, 4, 8) {real, imag} */,
  {32'hc138111a, 32'hc0ef40a5} /* (13, 4, 7) {real, imag} */,
  {32'hc134e8dc, 32'h4115d063} /* (13, 4, 6) {real, imag} */,
  {32'hc115d4a8, 32'hc212b3a1} /* (13, 4, 5) {real, imag} */,
  {32'hc115f132, 32'h41950263} /* (13, 4, 4) {real, imag} */,
  {32'hc13d5dd2, 32'h41c66230} /* (13, 4, 3) {real, imag} */,
  {32'hc2738a88, 32'hc294fddf} /* (13, 4, 2) {real, imag} */,
  {32'h434134bb, 32'h41a3fbe6} /* (13, 4, 1) {real, imag} */,
  {32'h41380e20, 32'hc12ec639} /* (13, 4, 0) {real, imag} */,
  {32'hc323e835, 32'h42361e82} /* (13, 3, 31) {real, imag} */,
  {32'h42b1e709, 32'hc29ad8bc} /* (13, 3, 30) {real, imag} */,
  {32'hc1442026, 32'h41ae3352} /* (13, 3, 29) {real, imag} */,
  {32'h42019c62, 32'h41e10618} /* (13, 3, 28) {real, imag} */,
  {32'hc1166041, 32'h410d634d} /* (13, 3, 27) {real, imag} */,
  {32'hc1def5ef, 32'h3f0bc6b0} /* (13, 3, 26) {real, imag} */,
  {32'h417954ec, 32'h41045988} /* (13, 3, 25) {real, imag} */,
  {32'h4112f958, 32'hc19f822c} /* (13, 3, 24) {real, imag} */,
  {32'h3d640c80, 32'h40e8fc8d} /* (13, 3, 23) {real, imag} */,
  {32'h4054200c, 32'h419f8cf4} /* (13, 3, 22) {real, imag} */,
  {32'hc0aea28d, 32'hc0b53435} /* (13, 3, 21) {real, imag} */,
  {32'hc10bb8bf, 32'hc144d7fd} /* (13, 3, 20) {real, imag} */,
  {32'hc0976c15, 32'hc122b43e} /* (13, 3, 19) {real, imag} */,
  {32'hc0519008, 32'h40f9caa6} /* (13, 3, 18) {real, imag} */,
  {32'hc09b4100, 32'h41306c75} /* (13, 3, 17) {real, imag} */,
  {32'h408c217f, 32'hc017d838} /* (13, 3, 16) {real, imag} */,
  {32'h41062dcb, 32'hc1759eb1} /* (13, 3, 15) {real, imag} */,
  {32'hc1140fbd, 32'h40dfb95f} /* (13, 3, 14) {real, imag} */,
  {32'hbfe28a90, 32'h40d394ce} /* (13, 3, 13) {real, imag} */,
  {32'h410734c1, 32'hc13ae193} /* (13, 3, 12) {real, imag} */,
  {32'h419c4002, 32'hc0aebbca} /* (13, 3, 11) {real, imag} */,
  {32'hc1355213, 32'h40c8641c} /* (13, 3, 10) {real, imag} */,
  {32'hc1a665ad, 32'hc1c5a785} /* (13, 3, 9) {real, imag} */,
  {32'h41544653, 32'hc0e32b28} /* (13, 3, 8) {real, imag} */,
  {32'h41873f7e, 32'h40d45d4e} /* (13, 3, 7) {real, imag} */,
  {32'h409ada3e, 32'hc0d748a0} /* (13, 3, 6) {real, imag} */,
  {32'h4092de62, 32'h42015ec2} /* (13, 3, 5) {real, imag} */,
  {32'hc0f1406c, 32'h411adfc1} /* (13, 3, 4) {real, imag} */,
  {32'h40081768, 32'h416725fc} /* (13, 3, 3) {real, imag} */,
  {32'hc1fe4c2e, 32'hc28f0f16} /* (13, 3, 2) {real, imag} */,
  {32'h431fb372, 32'h42be16a3} /* (13, 3, 1) {real, imag} */,
  {32'h3fa660e0, 32'hc16acc22} /* (13, 3, 0) {real, imag} */,
  {32'hc4815e68, 32'hc2018fb5} /* (13, 2, 31) {real, imag} */,
  {32'h4400fd8c, 32'hc33c423d} /* (13, 2, 30) {real, imag} */,
  {32'h418ee477, 32'h4236c940} /* (13, 2, 29) {real, imag} */,
  {32'hc27c727d, 32'h429aa5a0} /* (13, 2, 28) {real, imag} */,
  {32'h4252dfd8, 32'hc22eb7d0} /* (13, 2, 27) {real, imag} */,
  {32'h41f1b084, 32'hc1964333} /* (13, 2, 26) {real, imag} */,
  {32'hc1bf6962, 32'h41268bfe} /* (13, 2, 25) {real, imag} */,
  {32'h418a2f20, 32'hc21cc432} /* (13, 2, 24) {real, imag} */,
  {32'hc1aa734e, 32'h401195c8} /* (13, 2, 23) {real, imag} */,
  {32'h3ffbe8a6, 32'h40c51894} /* (13, 2, 22) {real, imag} */,
  {32'h41c5c5b7, 32'hc1965722} /* (13, 2, 21) {real, imag} */,
  {32'hc108a3c5, 32'hbf823a6c} /* (13, 2, 20) {real, imag} */,
  {32'hc13d2edf, 32'h413dddff} /* (13, 2, 19) {real, imag} */,
  {32'h40d2eaa6, 32'hc0b9d64a} /* (13, 2, 18) {real, imag} */,
  {32'h40a71e94, 32'hc071e27c} /* (13, 2, 17) {real, imag} */,
  {32'h404048ba, 32'hc109ff00} /* (13, 2, 16) {real, imag} */,
  {32'hc07a6fe6, 32'h4000c659} /* (13, 2, 15) {real, imag} */,
  {32'h4086d73e, 32'hbf477020} /* (13, 2, 14) {real, imag} */,
  {32'hc0441c38, 32'hbff27df8} /* (13, 2, 13) {real, imag} */,
  {32'h4144da32, 32'hbf99dd4a} /* (13, 2, 12) {real, imag} */,
  {32'h400a8dfa, 32'h410e0133} /* (13, 2, 11) {real, imag} */,
  {32'hc073e737, 32'h402ed053} /* (13, 2, 10) {real, imag} */,
  {32'hc129a519, 32'hc11a11d5} /* (13, 2, 9) {real, imag} */,
  {32'h41b20941, 32'hc0c89240} /* (13, 2, 8) {real, imag} */,
  {32'hc184c831, 32'hc148bc52} /* (13, 2, 7) {real, imag} */,
  {32'h40c2dbcf, 32'h41a0b9a9} /* (13, 2, 6) {real, imag} */,
  {32'h422d1202, 32'h4292c31d} /* (13, 2, 5) {real, imag} */,
  {32'hc2a94460, 32'hc280e95a} /* (13, 2, 4) {real, imag} */,
  {32'h4130d0ee, 32'h41176950} /* (13, 2, 3) {real, imag} */,
  {32'h439f13b5, 32'hc2b25670} /* (13, 2, 2) {real, imag} */,
  {32'hc41114de, 32'h42828f76} /* (13, 2, 1) {real, imag} */,
  {32'hc400e086, 32'hc281dfa2} /* (13, 2, 0) {real, imag} */,
  {32'h44aa3b02, 32'hc39bc8b7} /* (13, 1, 31) {real, imag} */,
  {32'hc3b454ff, 32'hbddbd280} /* (13, 1, 30) {real, imag} */,
  {32'h407b94b8, 32'h42490d33} /* (13, 1, 29) {real, imag} */,
  {32'h428aae68, 32'h418e8612} /* (13, 1, 28) {real, imag} */,
  {32'hc2d0536d, 32'h41939335} /* (13, 1, 27) {real, imag} */,
  {32'h41f15cf4, 32'h3f731240} /* (13, 1, 26) {real, imag} */,
  {32'h40cf47b6, 32'h408a0662} /* (13, 1, 25) {real, imag} */,
  {32'hc1c5ff5d, 32'h41e73836} /* (13, 1, 24) {real, imag} */,
  {32'hc1e65271, 32'h411d0d82} /* (13, 1, 23) {real, imag} */,
  {32'h4156a2ef, 32'h4167e2aa} /* (13, 1, 22) {real, imag} */,
  {32'h40f7833e, 32'h41d130c4} /* (13, 1, 21) {real, imag} */,
  {32'hc0c962ea, 32'hc096c8ee} /* (13, 1, 20) {real, imag} */,
  {32'h403a2386, 32'hc1080944} /* (13, 1, 19) {real, imag} */,
  {32'hbf76c148, 32'h411373e6} /* (13, 1, 18) {real, imag} */,
  {32'hc0eb603b, 32'hc13797e4} /* (13, 1, 17) {real, imag} */,
  {32'h3f9e4d7a, 32'h406b9c43} /* (13, 1, 16) {real, imag} */,
  {32'hc095677c, 32'hc0d04219} /* (13, 1, 15) {real, imag} */,
  {32'h40daa498, 32'h4142f752} /* (13, 1, 14) {real, imag} */,
  {32'hc0091a82, 32'hc0927560} /* (13, 1, 13) {real, imag} */,
  {32'h41832e1e, 32'hc0209c45} /* (13, 1, 12) {real, imag} */,
  {32'hc1684b84, 32'h40d87810} /* (13, 1, 11) {real, imag} */,
  {32'h40d5f99e, 32'hc0d461a2} /* (13, 1, 10) {real, imag} */,
  {32'h402cbf30, 32'h40a3a6f9} /* (13, 1, 9) {real, imag} */,
  {32'hc0f87749, 32'hc23a3654} /* (13, 1, 8) {real, imag} */,
  {32'h4204747f, 32'h40e777a5} /* (13, 1, 7) {real, imag} */,
  {32'hc126abd0, 32'hc23c441e} /* (13, 1, 6) {real, imag} */,
  {32'hc25abc92, 32'hc1a7d83a} /* (13, 1, 5) {real, imag} */,
  {32'hc1ae13db, 32'h42a3767e} /* (13, 1, 4) {real, imag} */,
  {32'hc2b4c27d, 32'hc0dada78} /* (13, 1, 3) {real, imag} */,
  {32'hc402e8c4, 32'hc3ec369e} /* (13, 1, 2) {real, imag} */,
  {32'h44e1b185, 32'h44886478} /* (13, 1, 1) {real, imag} */,
  {32'h44d0d69a, 32'h4289118f} /* (13, 1, 0) {real, imag} */,
  {32'h447a1af5, 32'hc4598278} /* (13, 0, 31) {real, imag} */,
  {32'hc332fb1d, 32'h4384ef35} /* (13, 0, 30) {real, imag} */,
  {32'hc1f68721, 32'hbe620200} /* (13, 0, 29) {real, imag} */,
  {32'h409d109e, 32'h41ac3145} /* (13, 0, 28) {real, imag} */,
  {32'hc256f2b6, 32'hc1715a62} /* (13, 0, 27) {real, imag} */,
  {32'h40255f1a, 32'hc1df5d9e} /* (13, 0, 26) {real, imag} */,
  {32'hc051d744, 32'hc1eaa92c} /* (13, 0, 25) {real, imag} */,
  {32'h414054a7, 32'h41c57d3e} /* (13, 0, 24) {real, imag} */,
  {32'hc1322841, 32'h4189bb5e} /* (13, 0, 23) {real, imag} */,
  {32'hc1a6f5f7, 32'hc0d839a9} /* (13, 0, 22) {real, imag} */,
  {32'hc1876cb2, 32'hbfdb4c0c} /* (13, 0, 21) {real, imag} */,
  {32'h40012962, 32'h400b0f61} /* (13, 0, 20) {real, imag} */,
  {32'h40c141ed, 32'hc1dab894} /* (13, 0, 19) {real, imag} */,
  {32'hbfa46338, 32'h41781e04} /* (13, 0, 18) {real, imag} */,
  {32'h40e22d90, 32'h4134fbaf} /* (13, 0, 17) {real, imag} */,
  {32'hc122e0fd, 32'h00000000} /* (13, 0, 16) {real, imag} */,
  {32'h40e22d90, 32'hc134fbaf} /* (13, 0, 15) {real, imag} */,
  {32'hbfa46338, 32'hc1781e04} /* (13, 0, 14) {real, imag} */,
  {32'h40c141ed, 32'h41dab894} /* (13, 0, 13) {real, imag} */,
  {32'h40012962, 32'hc00b0f61} /* (13, 0, 12) {real, imag} */,
  {32'hc1876cb2, 32'h3fdb4c0c} /* (13, 0, 11) {real, imag} */,
  {32'hc1a6f5f7, 32'h40d839a9} /* (13, 0, 10) {real, imag} */,
  {32'hc1322841, 32'hc189bb5e} /* (13, 0, 9) {real, imag} */,
  {32'h414054a7, 32'hc1c57d3e} /* (13, 0, 8) {real, imag} */,
  {32'hc051d744, 32'h41eaa92c} /* (13, 0, 7) {real, imag} */,
  {32'h40255f1a, 32'h41df5d9e} /* (13, 0, 6) {real, imag} */,
  {32'hc256f2b6, 32'h41715a62} /* (13, 0, 5) {real, imag} */,
  {32'h409d109e, 32'hc1ac3145} /* (13, 0, 4) {real, imag} */,
  {32'hc1f68721, 32'h3e620200} /* (13, 0, 3) {real, imag} */,
  {32'hc332fb1d, 32'hc384ef35} /* (13, 0, 2) {real, imag} */,
  {32'h447a1af5, 32'h44598278} /* (13, 0, 1) {real, imag} */,
  {32'h44cde24c, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h450a1a57, 32'hc4a42047} /* (12, 31, 31) {real, imag} */,
  {32'hc4178599, 32'h44040624} /* (12, 31, 30) {real, imag} */,
  {32'hc17c7a62, 32'h3eb1b2c0} /* (12, 31, 29) {real, imag} */,
  {32'hc1d5e5f8, 32'hc28a5466} /* (12, 31, 28) {real, imag} */,
  {32'hc297b820, 32'h41330fcc} /* (12, 31, 27) {real, imag} */,
  {32'hbfbdca10, 32'h41f86efc} /* (12, 31, 26) {real, imag} */,
  {32'h419c62ee, 32'hc0fe0faa} /* (12, 31, 25) {real, imag} */,
  {32'hc118265b, 32'h422d55c8} /* (12, 31, 24) {real, imag} */,
  {32'hc0818bd4, 32'h40b55bcb} /* (12, 31, 23) {real, imag} */,
  {32'hc110a74c, 32'h40627cf8} /* (12, 31, 22) {real, imag} */,
  {32'hbf86ff92, 32'h41aca6b3} /* (12, 31, 21) {real, imag} */,
  {32'h41091fa2, 32'h416dba92} /* (12, 31, 20) {real, imag} */,
  {32'hc023e17f, 32'h4035f07d} /* (12, 31, 19) {real, imag} */,
  {32'h40ca4ffc, 32'h4051755e} /* (12, 31, 18) {real, imag} */,
  {32'h410515ae, 32'hc0d3341d} /* (12, 31, 17) {real, imag} */,
  {32'h3f1d3b54, 32'hc0045edd} /* (12, 31, 16) {real, imag} */,
  {32'h4124ae14, 32'hc11f5256} /* (12, 31, 15) {real, imag} */,
  {32'h418bc016, 32'hc09f11d7} /* (12, 31, 14) {real, imag} */,
  {32'hc0bb366d, 32'hc13b3332} /* (12, 31, 13) {real, imag} */,
  {32'hc1b4d5fa, 32'hc0148662} /* (12, 31, 12) {real, imag} */,
  {32'hc1ba5049, 32'hc1d08e26} /* (12, 31, 11) {real, imag} */,
  {32'h41d95c2a, 32'hc1d1dde3} /* (12, 31, 10) {real, imag} */,
  {32'hc1870fa2, 32'h40eff2d8} /* (12, 31, 9) {real, imag} */,
  {32'hc163a5e7, 32'h3fc53760} /* (12, 31, 8) {real, imag} */,
  {32'h3ef52830, 32'h40c3bb92} /* (12, 31, 7) {real, imag} */,
  {32'h4137bf7e, 32'h3fc3a2e8} /* (12, 31, 6) {real, imag} */,
  {32'hc302d0df, 32'h4192267f} /* (12, 31, 5) {real, imag} */,
  {32'h42a8dd31, 32'hc243f438} /* (12, 31, 4) {real, imag} */,
  {32'h3ecc7e60, 32'hc1d14ad1} /* (12, 31, 3) {real, imag} */,
  {32'hc3c996dd, 32'hc19d7d75} /* (12, 31, 2) {real, imag} */,
  {32'h44c82ad4, 32'h439e442a} /* (12, 31, 1) {real, imag} */,
  {32'h45027137, 32'hc2fc5dd8} /* (12, 31, 0) {real, imag} */,
  {32'hc4277074, 32'hc29ec049} /* (12, 30, 31) {real, imag} */,
  {32'h43b3884d, 32'h430b266a} /* (12, 30, 30) {real, imag} */,
  {32'h416ad44f, 32'hc04dec46} /* (12, 30, 29) {real, imag} */,
  {32'hc2bf031d, 32'h42613fe7} /* (12, 30, 28) {real, imag} */,
  {32'h421fe174, 32'hc294b361} /* (12, 30, 27) {real, imag} */,
  {32'h40d54688, 32'hc1edd322} /* (12, 30, 26) {real, imag} */,
  {32'hc1baad82, 32'h40af3b90} /* (12, 30, 25) {real, imag} */,
  {32'h41923302, 32'hc16edf45} /* (12, 30, 24) {real, imag} */,
  {32'hc15da304, 32'h3fd6421c} /* (12, 30, 23) {real, imag} */,
  {32'hc09c5747, 32'h4003ad38} /* (12, 30, 22) {real, imag} */,
  {32'h40035d5e, 32'hc1d94946} /* (12, 30, 21) {real, imag} */,
  {32'h40c9d1cf, 32'hc17f73f2} /* (12, 30, 20) {real, imag} */,
  {32'h3f580674, 32'h40876737} /* (12, 30, 19) {real, imag} */,
  {32'h419fb44e, 32'hc1b52066} /* (12, 30, 18) {real, imag} */,
  {32'hc1370633, 32'h409610f8} /* (12, 30, 17) {real, imag} */,
  {32'h402fd85c, 32'hc05e13b1} /* (12, 30, 16) {real, imag} */,
  {32'hc1223768, 32'hc11c3d1c} /* (12, 30, 15) {real, imag} */,
  {32'h3f07fa99, 32'h41956b41} /* (12, 30, 14) {real, imag} */,
  {32'h3e64a3a0, 32'hc0c07170} /* (12, 30, 13) {real, imag} */,
  {32'hc18883d2, 32'hc024e536} /* (12, 30, 12) {real, imag} */,
  {32'h41982ee2, 32'h40e80d46} /* (12, 30, 11) {real, imag} */,
  {32'hbf2616c0, 32'hc11de8c6} /* (12, 30, 10) {real, imag} */,
  {32'hc155106e, 32'hc062f3b2} /* (12, 30, 9) {real, imag} */,
  {32'h409fef56, 32'h422d5feb} /* (12, 30, 8) {real, imag} */,
  {32'hc1a564aa, 32'hc01e9024} /* (12, 30, 7) {real, imag} */,
  {32'h41c01a4f, 32'h40038ca4} /* (12, 30, 6) {real, imag} */,
  {32'h420a77f5, 32'h427ff0ed} /* (12, 30, 5) {real, imag} */,
  {32'hc1ddc005, 32'hc264f300} /* (12, 30, 4) {real, imag} */,
  {32'h414652fa, 32'hc1d9fe6a} /* (12, 30, 3) {real, imag} */,
  {32'h4410d81c, 32'h431eaae8} /* (12, 30, 2) {real, imag} */,
  {32'hc497a83c, 32'h4178cf0d} /* (12, 30, 1) {real, imag} */,
  {32'hc4170c5e, 32'h42ae9758} /* (12, 30, 0) {real, imag} */,
  {32'h4312a3e9, 32'hc2ea5577} /* (12, 29, 31) {real, imag} */,
  {32'hc128edd3, 32'h42cfd050} /* (12, 29, 30) {real, imag} */,
  {32'hc1a2e696, 32'h403b32f8} /* (12, 29, 29) {real, imag} */,
  {32'hc1a7b10e, 32'hc04836a2} /* (12, 29, 28) {real, imag} */,
  {32'h3f6fd260, 32'hc20c5d78} /* (12, 29, 27) {real, imag} */,
  {32'h41e0d454, 32'hc1a74a15} /* (12, 29, 26) {real, imag} */,
  {32'h41421172, 32'h41840ec2} /* (12, 29, 25) {real, imag} */,
  {32'hc11f6a52, 32'hc191faf9} /* (12, 29, 24) {real, imag} */,
  {32'hc0f32a41, 32'hbfa1388e} /* (12, 29, 23) {real, imag} */,
  {32'h415aeefa, 32'h40d73c36} /* (12, 29, 22) {real, imag} */,
  {32'h3e1b77f8, 32'hbff0360a} /* (12, 29, 21) {real, imag} */,
  {32'hbf777728, 32'hc1002321} /* (12, 29, 20) {real, imag} */,
  {32'h40e0bfcd, 32'hbf411428} /* (12, 29, 19) {real, imag} */,
  {32'h4140d174, 32'h41b66366} /* (12, 29, 18) {real, imag} */,
  {32'h3d26f400, 32'h402872c3} /* (12, 29, 17) {real, imag} */,
  {32'h3fab2892, 32'hc103207f} /* (12, 29, 16) {real, imag} */,
  {32'hbefd6064, 32'hc130ecf8} /* (12, 29, 15) {real, imag} */,
  {32'hc131414e, 32'h414da552} /* (12, 29, 14) {real, imag} */,
  {32'hc0b8b918, 32'h40cad76c} /* (12, 29, 13) {real, imag} */,
  {32'hc09c74ba, 32'hbf7e70c4} /* (12, 29, 12) {real, imag} */,
  {32'hc10648f9, 32'hc0093eac} /* (12, 29, 11) {real, imag} */,
  {32'h400f9476, 32'h40f131d8} /* (12, 29, 10) {real, imag} */,
  {32'h41c0d3d6, 32'hc089f5b6} /* (12, 29, 9) {real, imag} */,
  {32'h41b30560, 32'h41ccfaf7} /* (12, 29, 8) {real, imag} */,
  {32'h40e79dbc, 32'hc02aa85f} /* (12, 29, 7) {real, imag} */,
  {32'hc0af6f4c, 32'hc17ea88b} /* (12, 29, 6) {real, imag} */,
  {32'hc1a6ba80, 32'hc083b5f0} /* (12, 29, 5) {real, imag} */,
  {32'h4245e4f9, 32'hc223d5ea} /* (12, 29, 4) {real, imag} */,
  {32'hc1c2fd55, 32'hc171830f} /* (12, 29, 3) {real, imag} */,
  {32'h428bdc71, 32'h42f6a746} /* (12, 29, 2) {real, imag} */,
  {32'hc32f9341, 32'hc286f384} /* (12, 29, 1) {real, imag} */,
  {32'hc10d2149, 32'hc0c7578c} /* (12, 29, 0) {real, imag} */,
  {32'h4337d9a4, 32'hc2032bea} /* (12, 28, 31) {real, imag} */,
  {32'hc28a8819, 32'h42a57cce} /* (12, 28, 30) {real, imag} */,
  {32'h41a63a80, 32'hc10b4e3e} /* (12, 28, 29) {real, imag} */,
  {32'h3fcab608, 32'hc15d0d77} /* (12, 28, 28) {real, imag} */,
  {32'h418753c1, 32'h42469815} /* (12, 28, 27) {real, imag} */,
  {32'hc164fdca, 32'hc153d029} /* (12, 28, 26) {real, imag} */,
  {32'hbff00cdf, 32'h3ffd57e8} /* (12, 28, 25) {real, imag} */,
  {32'h3fa5d519, 32'h421f6337} /* (12, 28, 24) {real, imag} */,
  {32'hc1868d64, 32'hbf9128a8} /* (12, 28, 23) {real, imag} */,
  {32'hbf8847ca, 32'hc1b29544} /* (12, 28, 22) {real, imag} */,
  {32'hc162df5e, 32'h40d92f7f} /* (12, 28, 21) {real, imag} */,
  {32'hc16678b6, 32'h3f8de550} /* (12, 28, 20) {real, imag} */,
  {32'hc08fada2, 32'hc11db3ae} /* (12, 28, 19) {real, imag} */,
  {32'h40dd89da, 32'h40fea952} /* (12, 28, 18) {real, imag} */,
  {32'hc04c54b7, 32'hc05d78bf} /* (12, 28, 17) {real, imag} */,
  {32'h3fb7afbe, 32'h3fbb251e} /* (12, 28, 16) {real, imag} */,
  {32'h4082338f, 32'hc1835316} /* (12, 28, 15) {real, imag} */,
  {32'hc13ff452, 32'hc047fd40} /* (12, 28, 14) {real, imag} */,
  {32'hbefd0cf0, 32'h40dcf40a} /* (12, 28, 13) {real, imag} */,
  {32'h412cc460, 32'h40c9beae} /* (12, 28, 12) {real, imag} */,
  {32'hc1311b24, 32'hc1be53de} /* (12, 28, 11) {real, imag} */,
  {32'hc046726b, 32'h40eb4496} /* (12, 28, 10) {real, imag} */,
  {32'hc10eedca, 32'h4156346c} /* (12, 28, 9) {real, imag} */,
  {32'h4123a800, 32'h41637b8e} /* (12, 28, 8) {real, imag} */,
  {32'h41c1bb7c, 32'hbf87b904} /* (12, 28, 7) {real, imag} */,
  {32'hbfb09fd0, 32'h40e1f966} /* (12, 28, 6) {real, imag} */,
  {32'hc1a1bf81, 32'h4209961c} /* (12, 28, 5) {real, imag} */,
  {32'h420d7230, 32'hc0d87f00} /* (12, 28, 4) {real, imag} */,
  {32'h4115a513, 32'h411e767e} /* (12, 28, 3) {real, imag} */,
  {32'hc2dcea31, 32'h429ef263} /* (12, 28, 2) {real, imag} */,
  {32'h41f27b0d, 32'hc286c60a} /* (12, 28, 1) {real, imag} */,
  {32'h4223de4b, 32'h40ad0483} /* (12, 28, 0) {real, imag} */,
  {32'hc28f1aa0, 32'h429778cd} /* (12, 27, 31) {real, imag} */,
  {32'h4196b9ec, 32'hc23e9b2e} /* (12, 27, 30) {real, imag} */,
  {32'h3f969efc, 32'h41247fc8} /* (12, 27, 29) {real, imag} */,
  {32'hc0518a98, 32'h420fa1ff} /* (12, 27, 28) {real, imag} */,
  {32'h4222f932, 32'hc1ca88df} /* (12, 27, 27) {real, imag} */,
  {32'h410ef28b, 32'hc0b88fac} /* (12, 27, 26) {real, imag} */,
  {32'hc156146b, 32'h40549664} /* (12, 27, 25) {real, imag} */,
  {32'h413e32db, 32'h3fbd766c} /* (12, 27, 24) {real, imag} */,
  {32'h41ca58fd, 32'hc1a897eb} /* (12, 27, 23) {real, imag} */,
  {32'hc11a86c0, 32'hc14bbc92} /* (12, 27, 22) {real, imag} */,
  {32'h40ef5cb0, 32'hc13b6d1c} /* (12, 27, 21) {real, imag} */,
  {32'h41646224, 32'h3faa26f8} /* (12, 27, 20) {real, imag} */,
  {32'hc0e751e9, 32'hc0e34ba0} /* (12, 27, 19) {real, imag} */,
  {32'hc1a7de4e, 32'hc0d2b6f0} /* (12, 27, 18) {real, imag} */,
  {32'h40096b4e, 32'hbfb23a2e} /* (12, 27, 17) {real, imag} */,
  {32'h40faf88e, 32'hbe299bc0} /* (12, 27, 16) {real, imag} */,
  {32'h403a5002, 32'h40ff7cd6} /* (12, 27, 15) {real, imag} */,
  {32'hc10e6636, 32'h404b7434} /* (12, 27, 14) {real, imag} */,
  {32'hc04710e5, 32'hc1bbc358} /* (12, 27, 13) {real, imag} */,
  {32'h40a19a58, 32'h406bb680} /* (12, 27, 12) {real, imag} */,
  {32'h4195e960, 32'h3fe3c09e} /* (12, 27, 11) {real, imag} */,
  {32'h4136a4df, 32'h40ce5ece} /* (12, 27, 10) {real, imag} */,
  {32'h413bef24, 32'h402990b2} /* (12, 27, 9) {real, imag} */,
  {32'h41646d1a, 32'h41a14e6a} /* (12, 27, 8) {real, imag} */,
  {32'h4111643e, 32'h417be684} /* (12, 27, 7) {real, imag} */,
  {32'hc08a0898, 32'h404530d6} /* (12, 27, 6) {real, imag} */,
  {32'h413d4f8e, 32'hc1db9038} /* (12, 27, 5) {real, imag} */,
  {32'hc15d801a, 32'hc21fcc3e} /* (12, 27, 4) {real, imag} */,
  {32'hc0546108, 32'hbe714600} /* (12, 27, 3) {real, imag} */,
  {32'h41a0296b, 32'hc1439b3d} /* (12, 27, 2) {real, imag} */,
  {32'hc2d779ce, 32'h4181bdaa} /* (12, 27, 1) {real, imag} */,
  {32'hc2b36c5a, 32'h41d1c64b} /* (12, 27, 0) {real, imag} */,
  {32'h41c0688c, 32'h41256c48} /* (12, 26, 31) {real, imag} */,
  {32'h40e21dd1, 32'h40a82dc7} /* (12, 26, 30) {real, imag} */,
  {32'hbfda4105, 32'hc15058cc} /* (12, 26, 29) {real, imag} */,
  {32'h41276cbc, 32'h4186d6ae} /* (12, 26, 28) {real, imag} */,
  {32'h416c1961, 32'h41eb224e} /* (12, 26, 27) {real, imag} */,
  {32'h3f8748fe, 32'h418dff78} /* (12, 26, 26) {real, imag} */,
  {32'hc1209ccd, 32'hc0c3c6fc} /* (12, 26, 25) {real, imag} */,
  {32'h40f6e78d, 32'h411d95cf} /* (12, 26, 24) {real, imag} */,
  {32'hc1f1ccb5, 32'h4020763e} /* (12, 26, 23) {real, imag} */,
  {32'hc194698a, 32'h41435a5e} /* (12, 26, 22) {real, imag} */,
  {32'hc022c197, 32'hbf15855c} /* (12, 26, 21) {real, imag} */,
  {32'hbfd79764, 32'hc0ab156b} /* (12, 26, 20) {real, imag} */,
  {32'hc0b7ac2e, 32'hc0cb43c5} /* (12, 26, 19) {real, imag} */,
  {32'h4115d21d, 32'h414410c2} /* (12, 26, 18) {real, imag} */,
  {32'h40293c3f, 32'h3f4e4a20} /* (12, 26, 17) {real, imag} */,
  {32'hc0f8fa08, 32'hc07247e3} /* (12, 26, 16) {real, imag} */,
  {32'h40f80efa, 32'h41106fff} /* (12, 26, 15) {real, imag} */,
  {32'hc1277344, 32'h40178d2d} /* (12, 26, 14) {real, imag} */,
  {32'h4145368a, 32'hc16748ca} /* (12, 26, 13) {real, imag} */,
  {32'h41025b10, 32'h3fdda844} /* (12, 26, 12) {real, imag} */,
  {32'h3ff59cd4, 32'h40498209} /* (12, 26, 11) {real, imag} */,
  {32'h41d6f712, 32'h4130ef90} /* (12, 26, 10) {real, imag} */,
  {32'hbf2dade8, 32'h4091acab} /* (12, 26, 9) {real, imag} */,
  {32'hc12c8ba4, 32'hc0ae2e86} /* (12, 26, 8) {real, imag} */,
  {32'h3f95db3c, 32'h40fa869f} /* (12, 26, 7) {real, imag} */,
  {32'hbf527f58, 32'hc10adc55} /* (12, 26, 6) {real, imag} */,
  {32'hc04d6dd6, 32'hc177188a} /* (12, 26, 5) {real, imag} */,
  {32'hc0a373d8, 32'h418ec897} /* (12, 26, 4) {real, imag} */,
  {32'h4170c5af, 32'h418cd5b2} /* (12, 26, 3) {real, imag} */,
  {32'h42070773, 32'h402dedc6} /* (12, 26, 2) {real, imag} */,
  {32'h4148d60a, 32'h4189383b} /* (12, 26, 1) {real, imag} */,
  {32'h40d79f30, 32'hc1892917} /* (12, 26, 0) {real, imag} */,
  {32'h41b2866c, 32'hc19a62ae} /* (12, 25, 31) {real, imag} */,
  {32'hc12ad936, 32'h410de49f} /* (12, 25, 30) {real, imag} */,
  {32'hc1abaeea, 32'hc1a19736} /* (12, 25, 29) {real, imag} */,
  {32'hc109305b, 32'hc1c35708} /* (12, 25, 28) {real, imag} */,
  {32'hbe104e60, 32'hc0edab12} /* (12, 25, 27) {real, imag} */,
  {32'h410e4e3f, 32'h3ed027e0} /* (12, 25, 26) {real, imag} */,
  {32'hc0ee6d63, 32'hbffc670f} /* (12, 25, 25) {real, imag} */,
  {32'h41373284, 32'h40492c72} /* (12, 25, 24) {real, imag} */,
  {32'hc129ec26, 32'h41102867} /* (12, 25, 23) {real, imag} */,
  {32'h4137f084, 32'hc0ceae74} /* (12, 25, 22) {real, imag} */,
  {32'h41c6678c, 32'h4109de8a} /* (12, 25, 21) {real, imag} */,
  {32'h4076e958, 32'h3fea1e50} /* (12, 25, 20) {real, imag} */,
  {32'hbfcee135, 32'h41a09ca0} /* (12, 25, 19) {real, imag} */,
  {32'hc0bfcbee, 32'h3f8a4222} /* (12, 25, 18) {real, imag} */,
  {32'h41195c5a, 32'h405a43c5} /* (12, 25, 17) {real, imag} */,
  {32'hc13a4e07, 32'hc11ec426} /* (12, 25, 16) {real, imag} */,
  {32'hc0baef45, 32'hc107c313} /* (12, 25, 15) {real, imag} */,
  {32'h3f39c740, 32'hc0d03f0a} /* (12, 25, 14) {real, imag} */,
  {32'hc0db93a7, 32'hc0d40646} /* (12, 25, 13) {real, imag} */,
  {32'h40cba3a8, 32'hc10a611a} /* (12, 25, 12) {real, imag} */,
  {32'h41b1bf63, 32'h4130db68} /* (12, 25, 11) {real, imag} */,
  {32'hc0494967, 32'hc19576f0} /* (12, 25, 10) {real, imag} */,
  {32'hc168ce72, 32'h40ecdbfa} /* (12, 25, 9) {real, imag} */,
  {32'hc0c69ca6, 32'h416da232} /* (12, 25, 8) {real, imag} */,
  {32'h418e6da7, 32'hc180ff3c} /* (12, 25, 7) {real, imag} */,
  {32'h3fd8d4d9, 32'hc114ef5a} /* (12, 25, 6) {real, imag} */,
  {32'hc00de3ca, 32'h4159da9e} /* (12, 25, 5) {real, imag} */,
  {32'hbe771ae0, 32'hc100fbe1} /* (12, 25, 4) {real, imag} */,
  {32'hc0a66d90, 32'hc01902ab} /* (12, 25, 3) {real, imag} */,
  {32'h400ba543, 32'h41a83cd6} /* (12, 25, 2) {real, imag} */,
  {32'h418864b8, 32'h4186813c} /* (12, 25, 1) {real, imag} */,
  {32'h3f8a5948, 32'hc11dbf1c} /* (12, 25, 0) {real, imag} */,
  {32'hc2271c54, 32'hc0336e38} /* (12, 24, 31) {real, imag} */,
  {32'h411f72d3, 32'hc19c418b} /* (12, 24, 30) {real, imag} */,
  {32'hc0cc5146, 32'hc0d2beb6} /* (12, 24, 29) {real, imag} */,
  {32'hc1fe4fbb, 32'h4201c3e9} /* (12, 24, 28) {real, imag} */,
  {32'h41b8f709, 32'h41125a6d} /* (12, 24, 27) {real, imag} */,
  {32'h413bce2b, 32'h416fa4ac} /* (12, 24, 26) {real, imag} */,
  {32'hc1902ce7, 32'h3fa94934} /* (12, 24, 25) {real, imag} */,
  {32'h41296b24, 32'h402807c6} /* (12, 24, 24) {real, imag} */,
  {32'h4077b3d4, 32'hbf832c72} /* (12, 24, 23) {real, imag} */,
  {32'h4198462c, 32'hc0575580} /* (12, 24, 22) {real, imag} */,
  {32'h408d3d5d, 32'h4191cd84} /* (12, 24, 21) {real, imag} */,
  {32'h41214265, 32'hc1f0923e} /* (12, 24, 20) {real, imag} */,
  {32'hc1dfd550, 32'hc182e46c} /* (12, 24, 19) {real, imag} */,
  {32'hc1090ca4, 32'h413d1332} /* (12, 24, 18) {real, imag} */,
  {32'h4072397a, 32'hc150a0ba} /* (12, 24, 17) {real, imag} */,
  {32'h408bee82, 32'h40832daf} /* (12, 24, 16) {real, imag} */,
  {32'h40f55ed6, 32'h40845e9e} /* (12, 24, 15) {real, imag} */,
  {32'h4185b8f0, 32'hbfa29cb2} /* (12, 24, 14) {real, imag} */,
  {32'hc1602cc6, 32'h410ace42} /* (12, 24, 13) {real, imag} */,
  {32'h41843314, 32'h40c0ca62} /* (12, 24, 12) {real, imag} */,
  {32'h418af3dd, 32'h3e0b2610} /* (12, 24, 11) {real, imag} */,
  {32'hc14c24f9, 32'hc18b88c2} /* (12, 24, 10) {real, imag} */,
  {32'h3fcaf790, 32'h411e647d} /* (12, 24, 9) {real, imag} */,
  {32'h40265bd6, 32'hc114c569} /* (12, 24, 8) {real, imag} */,
  {32'h3fbb2a06, 32'h412a99d8} /* (12, 24, 7) {real, imag} */,
  {32'h4057b212, 32'hc1189799} /* (12, 24, 6) {real, imag} */,
  {32'h41ac1f4b, 32'h411a1a5d} /* (12, 24, 5) {real, imag} */,
  {32'h4109fe48, 32'h4180a829} /* (12, 24, 4) {real, imag} */,
  {32'h403e2a16, 32'h417d3084} /* (12, 24, 3) {real, imag} */,
  {32'h41e7b91d, 32'hc14f02ca} /* (12, 24, 2) {real, imag} */,
  {32'hc2368768, 32'h41c3492a} /* (12, 24, 1) {real, imag} */,
  {32'hc1a18586, 32'h41e59562} /* (12, 24, 0) {real, imag} */,
  {32'h420c88e0, 32'hc17ba136} /* (12, 23, 31) {real, imag} */,
  {32'hc132cf29, 32'h41450dc2} /* (12, 23, 30) {real, imag} */,
  {32'h4194694d, 32'h41a73b66} /* (12, 23, 29) {real, imag} */,
  {32'hc123440a, 32'hc10694be} /* (12, 23, 28) {real, imag} */,
  {32'hc10e991e, 32'hc16c5cd1} /* (12, 23, 27) {real, imag} */,
  {32'hc18d0231, 32'hc156ed2e} /* (12, 23, 26) {real, imag} */,
  {32'h41347e58, 32'hc1010b1f} /* (12, 23, 25) {real, imag} */,
  {32'hbfc8f9b8, 32'h408550f6} /* (12, 23, 24) {real, imag} */,
  {32'h41a8d9da, 32'h4081fdc0} /* (12, 23, 23) {real, imag} */,
  {32'hc144eb94, 32'h41104fb8} /* (12, 23, 22) {real, imag} */,
  {32'hc17ee0a2, 32'h3fe47501} /* (12, 23, 21) {real, imag} */,
  {32'hc105bdbf, 32'h40c26312} /* (12, 23, 20) {real, imag} */,
  {32'hc14508e0, 32'hc10603a0} /* (12, 23, 19) {real, imag} */,
  {32'h40afeba0, 32'h4081e7d2} /* (12, 23, 18) {real, imag} */,
  {32'h404f1389, 32'hbdf37140} /* (12, 23, 17) {real, imag} */,
  {32'hbf159970, 32'hc0c8ca82} /* (12, 23, 16) {real, imag} */,
  {32'h4062ee80, 32'hc0d6a21a} /* (12, 23, 15) {real, imag} */,
  {32'h402be536, 32'h4096da72} /* (12, 23, 14) {real, imag} */,
  {32'h416b7e76, 32'hc050ba5d} /* (12, 23, 13) {real, imag} */,
  {32'h40acd43c, 32'hbf088848} /* (12, 23, 12) {real, imag} */,
  {32'hc0d4d71b, 32'hc05e34ba} /* (12, 23, 11) {real, imag} */,
  {32'h404731f8, 32'h40c52e51} /* (12, 23, 10) {real, imag} */,
  {32'h4067e15b, 32'hc144c022} /* (12, 23, 9) {real, imag} */,
  {32'hc1e9029f, 32'h4073fe1a} /* (12, 23, 8) {real, imag} */,
  {32'hc10bfbea, 32'h40b09ac7} /* (12, 23, 7) {real, imag} */,
  {32'hc011b4d8, 32'hc0176184} /* (12, 23, 6) {real, imag} */,
  {32'hc15fdec0, 32'hc09180ca} /* (12, 23, 5) {real, imag} */,
  {32'h40930aa4, 32'h411f0be6} /* (12, 23, 4) {real, imag} */,
  {32'h406fb2a9, 32'h40f5a3de} /* (12, 23, 3) {real, imag} */,
  {32'h40f139b0, 32'h408ba34c} /* (12, 23, 2) {real, imag} */,
  {32'hc1ac26a2, 32'hc1581372} /* (12, 23, 1) {real, imag} */,
  {32'hc0d846d4, 32'h41362a85} /* (12, 23, 0) {real, imag} */,
  {32'h407e1902, 32'hc0dc5910} /* (12, 22, 31) {real, imag} */,
  {32'hc0ab7df5, 32'h41d16798} /* (12, 22, 30) {real, imag} */,
  {32'h4055a988, 32'h3fa4b378} /* (12, 22, 29) {real, imag} */,
  {32'hc12b3b36, 32'hc1be0441} /* (12, 22, 28) {real, imag} */,
  {32'h4192f1d9, 32'h418ec082} /* (12, 22, 27) {real, imag} */,
  {32'h40265c2a, 32'h41802e80} /* (12, 22, 26) {real, imag} */,
  {32'h4106ba6c, 32'hc178915e} /* (12, 22, 25) {real, imag} */,
  {32'hbfd82168, 32'h40815e4e} /* (12, 22, 24) {real, imag} */,
  {32'h4093d84c, 32'h40148162} /* (12, 22, 23) {real, imag} */,
  {32'hc163e382, 32'hc10fcf0f} /* (12, 22, 22) {real, imag} */,
  {32'h3ff092a0, 32'h40f888d9} /* (12, 22, 21) {real, imag} */,
  {32'hc0ad19d0, 32'h41655c6c} /* (12, 22, 20) {real, imag} */,
  {32'h4066aef2, 32'h412f487a} /* (12, 22, 19) {real, imag} */,
  {32'h3f227404, 32'h3fad560c} /* (12, 22, 18) {real, imag} */,
  {32'h41051009, 32'hc13a4702} /* (12, 22, 17) {real, imag} */,
  {32'hc16c8e7e, 32'hc07c09dd} /* (12, 22, 16) {real, imag} */,
  {32'hc044ab12, 32'h408a335e} /* (12, 22, 15) {real, imag} */,
  {32'hbf4ae3b0, 32'hc10ad5ee} /* (12, 22, 14) {real, imag} */,
  {32'h413b9b44, 32'h40b4e42a} /* (12, 22, 13) {real, imag} */,
  {32'h3fa06ae4, 32'h401c2027} /* (12, 22, 12) {real, imag} */,
  {32'h414faca5, 32'h41587aac} /* (12, 22, 11) {real, imag} */,
  {32'h411a7328, 32'hbf5635a8} /* (12, 22, 10) {real, imag} */,
  {32'hc1a078e2, 32'hc16f731e} /* (12, 22, 9) {real, imag} */,
  {32'h417c55c3, 32'h417c540c} /* (12, 22, 8) {real, imag} */,
  {32'hc1839a38, 32'hc07ccb74} /* (12, 22, 7) {real, imag} */,
  {32'h4041c780, 32'h415dd260} /* (12, 22, 6) {real, imag} */,
  {32'hc15de302, 32'hc1206066} /* (12, 22, 5) {real, imag} */,
  {32'h4087cbfa, 32'hc08c8678} /* (12, 22, 4) {real, imag} */,
  {32'hc0e26c69, 32'h40f32102} /* (12, 22, 3) {real, imag} */,
  {32'hc088eda4, 32'hbbf3f800} /* (12, 22, 2) {real, imag} */,
  {32'h404abc3a, 32'hc17acf8d} /* (12, 22, 1) {real, imag} */,
  {32'hbfcdcbf4, 32'h4017835a} /* (12, 22, 0) {real, imag} */,
  {32'hc2034f73, 32'h4183b45a} /* (12, 21, 31) {real, imag} */,
  {32'hc15f6022, 32'hc08e3276} /* (12, 21, 30) {real, imag} */,
  {32'h41cc6d1a, 32'h40afa69c} /* (12, 21, 29) {real, imag} */,
  {32'h3f826e04, 32'hbf3ce460} /* (12, 21, 28) {real, imag} */,
  {32'hc0decbde, 32'hc13b6016} /* (12, 21, 27) {real, imag} */,
  {32'hc07d1fda, 32'h41852fba} /* (12, 21, 26) {real, imag} */,
  {32'h40a28a16, 32'hc0d698ec} /* (12, 21, 25) {real, imag} */,
  {32'hbf8f15a0, 32'hbf821db8} /* (12, 21, 24) {real, imag} */,
  {32'hbf2f3f30, 32'h4184f9f2} /* (12, 21, 23) {real, imag} */,
  {32'h3e8c34a0, 32'hc0d3f7b6} /* (12, 21, 22) {real, imag} */,
  {32'hbf5c20a8, 32'hc1669013} /* (12, 21, 21) {real, imag} */,
  {32'hc13219e8, 32'h4012b9ce} /* (12, 21, 20) {real, imag} */,
  {32'h405eaaac, 32'h40933988} /* (12, 21, 19) {real, imag} */,
  {32'hc07aa75d, 32'h413de7ae} /* (12, 21, 18) {real, imag} */,
  {32'hc0df6904, 32'h408f6480} /* (12, 21, 17) {real, imag} */,
  {32'hc155b970, 32'h40cbf572} /* (12, 21, 16) {real, imag} */,
  {32'h40f092f5, 32'hc1109226} /* (12, 21, 15) {real, imag} */,
  {32'hc1486a28, 32'h3fc17662} /* (12, 21, 14) {real, imag} */,
  {32'h41c734fa, 32'hbf4d33dc} /* (12, 21, 13) {real, imag} */,
  {32'hc0a6ae40, 32'h415eb3c2} /* (12, 21, 12) {real, imag} */,
  {32'h414bbf9e, 32'hc167477e} /* (12, 21, 11) {real, imag} */,
  {32'h40e54954, 32'hbfe7e868} /* (12, 21, 10) {real, imag} */,
  {32'h40ca8dd2, 32'hc12e6fc1} /* (12, 21, 9) {real, imag} */,
  {32'h41539253, 32'hc10fdd7c} /* (12, 21, 8) {real, imag} */,
  {32'hc1eb4003, 32'h419f3120} /* (12, 21, 7) {real, imag} */,
  {32'h412ba9e8, 32'hbffbf840} /* (12, 21, 6) {real, imag} */,
  {32'h40ed1526, 32'h416b689e} /* (12, 21, 5) {real, imag} */,
  {32'hbf5a4168, 32'hbf3040c0} /* (12, 21, 4) {real, imag} */,
  {32'h3fe45410, 32'h404cb406} /* (12, 21, 3) {real, imag} */,
  {32'h40d363fc, 32'hc12be2e8} /* (12, 21, 2) {real, imag} */,
  {32'hc13fcec4, 32'h41967562} /* (12, 21, 1) {real, imag} */,
  {32'hc18a8386, 32'h40be7d22} /* (12, 21, 0) {real, imag} */,
  {32'h40f337c8, 32'h3f1418a0} /* (12, 20, 31) {real, imag} */,
  {32'hc1266d18, 32'hc024d354} /* (12, 20, 30) {real, imag} */,
  {32'hc023b7c8, 32'h41661765} /* (12, 20, 29) {real, imag} */,
  {32'hc06a3c6c, 32'hc15f0697} /* (12, 20, 28) {real, imag} */,
  {32'hc11436e9, 32'hc09e677e} /* (12, 20, 27) {real, imag} */,
  {32'hc0867068, 32'h405b58c5} /* (12, 20, 26) {real, imag} */,
  {32'h3f405360, 32'hc1049ec0} /* (12, 20, 25) {real, imag} */,
  {32'h40cd632e, 32'h3eb02380} /* (12, 20, 24) {real, imag} */,
  {32'h3de10580, 32'hc1afb08a} /* (12, 20, 23) {real, imag} */,
  {32'h41a5f23c, 32'hc18e306e} /* (12, 20, 22) {real, imag} */,
  {32'hbfa70f42, 32'hc1786d17} /* (12, 20, 21) {real, imag} */,
  {32'h4194f2aa, 32'h40b4e7f0} /* (12, 20, 20) {real, imag} */,
  {32'h3ffd2d48, 32'h410ac66a} /* (12, 20, 19) {real, imag} */,
  {32'h4101f0a9, 32'hbffdb680} /* (12, 20, 18) {real, imag} */,
  {32'hc1487338, 32'h41b45976} /* (12, 20, 17) {real, imag} */,
  {32'hbf8dc800, 32'hc11a3c52} /* (12, 20, 16) {real, imag} */,
  {32'h3f17fe48, 32'hc02c5759} /* (12, 20, 15) {real, imag} */,
  {32'hc0eeb2ab, 32'hc19872ae} /* (12, 20, 14) {real, imag} */,
  {32'hc02d76ca, 32'hc087159a} /* (12, 20, 13) {real, imag} */,
  {32'h4143922c, 32'h416bcc95} /* (12, 20, 12) {real, imag} */,
  {32'hc1080318, 32'h40fef1de} /* (12, 20, 11) {real, imag} */,
  {32'hc01d0888, 32'h4192ca60} /* (12, 20, 10) {real, imag} */,
  {32'h40d78f7f, 32'h411e9134} /* (12, 20, 9) {real, imag} */,
  {32'h406170ae, 32'hc0457417} /* (12, 20, 8) {real, imag} */,
  {32'h413f21a0, 32'hc12eb222} /* (12, 20, 7) {real, imag} */,
  {32'hc1c00daa, 32'hc11d8693} /* (12, 20, 6) {real, imag} */,
  {32'h411a6eef, 32'hc10e1ac0} /* (12, 20, 5) {real, imag} */,
  {32'hc1a18d62, 32'h41185a0e} /* (12, 20, 4) {real, imag} */,
  {32'h4091ea00, 32'h41a198bc} /* (12, 20, 3) {real, imag} */,
  {32'hc141bcf4, 32'h40d708b8} /* (12, 20, 2) {real, imag} */,
  {32'hc0be874d, 32'hc01329a6} /* (12, 20, 1) {real, imag} */,
  {32'h4172f83e, 32'hc0ad0092} /* (12, 20, 0) {real, imag} */,
  {32'h4003ccea, 32'hc04277a7} /* (12, 19, 31) {real, imag} */,
  {32'h410f0c9d, 32'h3f7f1520} /* (12, 19, 30) {real, imag} */,
  {32'hc0a39940, 32'h40d401b2} /* (12, 19, 29) {real, imag} */,
  {32'h4086036e, 32'hc1c010a4} /* (12, 19, 28) {real, imag} */,
  {32'h4137ee46, 32'h40c70ab4} /* (12, 19, 27) {real, imag} */,
  {32'hc0ddb408, 32'h409b1316} /* (12, 19, 26) {real, imag} */,
  {32'h418cfb45, 32'h40851d0a} /* (12, 19, 25) {real, imag} */,
  {32'hbe9b0ff0, 32'h40f9c87e} /* (12, 19, 24) {real, imag} */,
  {32'hc0e3249d, 32'hbdfebee0} /* (12, 19, 23) {real, imag} */,
  {32'hc1180126, 32'h41029b13} /* (12, 19, 22) {real, imag} */,
  {32'hc0b3bc6a, 32'h408834a9} /* (12, 19, 21) {real, imag} */,
  {32'h41344d4f, 32'h413251eb} /* (12, 19, 20) {real, imag} */,
  {32'h4161cc70, 32'hc0ff0e7c} /* (12, 19, 19) {real, imag} */,
  {32'hc03db11c, 32'h411f5429} /* (12, 19, 18) {real, imag} */,
  {32'h411492f8, 32'h4034e552} /* (12, 19, 17) {real, imag} */,
  {32'hc10062f2, 32'hbf093d2c} /* (12, 19, 16) {real, imag} */,
  {32'h3fa1a1d2, 32'h4039fbc8} /* (12, 19, 15) {real, imag} */,
  {32'h411ab7a6, 32'hc0c7ad18} /* (12, 19, 14) {real, imag} */,
  {32'h3f5bcea4, 32'h4071e649} /* (12, 19, 13) {real, imag} */,
  {32'hbf2ec320, 32'hbee3d140} /* (12, 19, 12) {real, imag} */,
  {32'hc0bf0222, 32'hbfe7d49c} /* (12, 19, 11) {real, imag} */,
  {32'h41a25326, 32'hc1ad1844} /* (12, 19, 10) {real, imag} */,
  {32'hc13814f6, 32'h3f89dc84} /* (12, 19, 9) {real, imag} */,
  {32'h400cd287, 32'hc0b8f510} /* (12, 19, 8) {real, imag} */,
  {32'h412f3170, 32'h407731c8} /* (12, 19, 7) {real, imag} */,
  {32'h40cea723, 32'hbfbb1a57} /* (12, 19, 6) {real, imag} */,
  {32'hc1644dd6, 32'h4183020a} /* (12, 19, 5) {real, imag} */,
  {32'h40caeecc, 32'hc04f1528} /* (12, 19, 4) {real, imag} */,
  {32'h3eedc580, 32'hbfa54666} /* (12, 19, 3) {real, imag} */,
  {32'hc09b5811, 32'hc0b4f2dd} /* (12, 19, 2) {real, imag} */,
  {32'h40d8c7cf, 32'hc10a5177} /* (12, 19, 1) {real, imag} */,
  {32'h4013f162, 32'hc0a09a76} /* (12, 19, 0) {real, imag} */,
  {32'hc0817e78, 32'h3fdd81ce} /* (12, 18, 31) {real, imag} */,
  {32'h4090307c, 32'hc07d2cdc} /* (12, 18, 30) {real, imag} */,
  {32'hc0b4a66b, 32'h40af07a3} /* (12, 18, 29) {real, imag} */,
  {32'hc13b83d0, 32'h3f8bf2ec} /* (12, 18, 28) {real, imag} */,
  {32'hc0d3b863, 32'hc1b32638} /* (12, 18, 27) {real, imag} */,
  {32'hc0b6f300, 32'hc003f87c} /* (12, 18, 26) {real, imag} */,
  {32'h4031cd35, 32'h410b6377} /* (12, 18, 25) {real, imag} */,
  {32'hc0034c0c, 32'h4087dcc4} /* (12, 18, 24) {real, imag} */,
  {32'hbd93c0c0, 32'hc162cb74} /* (12, 18, 23) {real, imag} */,
  {32'hc0a56c3d, 32'h415d488a} /* (12, 18, 22) {real, imag} */,
  {32'hc1595416, 32'hc19ad53a} /* (12, 18, 21) {real, imag} */,
  {32'h40b93705, 32'h410d30c8} /* (12, 18, 20) {real, imag} */,
  {32'h411b8c15, 32'h4183ba70} /* (12, 18, 19) {real, imag} */,
  {32'h40d3911a, 32'hbff3eff0} /* (12, 18, 18) {real, imag} */,
  {32'h400f7ed8, 32'hc14dac09} /* (12, 18, 17) {real, imag} */,
  {32'h418acf87, 32'h4145cea3} /* (12, 18, 16) {real, imag} */,
  {32'hbe11f8e0, 32'h40e10868} /* (12, 18, 15) {real, imag} */,
  {32'hbf4920b4, 32'h4040929f} /* (12, 18, 14) {real, imag} */,
  {32'hc0c16301, 32'hc1753cf4} /* (12, 18, 13) {real, imag} */,
  {32'hc0a9b85a, 32'hc0b146cd} /* (12, 18, 12) {real, imag} */,
  {32'hc0ffcd52, 32'h40a1c17b} /* (12, 18, 11) {real, imag} */,
  {32'hbf9c6788, 32'hbfa5a96a} /* (12, 18, 10) {real, imag} */,
  {32'h411e4a18, 32'h40ca374c} /* (12, 18, 9) {real, imag} */,
  {32'h4137ecc2, 32'h411c6160} /* (12, 18, 8) {real, imag} */,
  {32'hbe740fc0, 32'h40544ca6} /* (12, 18, 7) {real, imag} */,
  {32'hc0bc2b9c, 32'h3f59e61c} /* (12, 18, 6) {real, imag} */,
  {32'hc172c10e, 32'hc1ab7596} /* (12, 18, 5) {real, imag} */,
  {32'hc16664b1, 32'h40fd9d26} /* (12, 18, 4) {real, imag} */,
  {32'h3fb908a6, 32'h4004b85e} /* (12, 18, 3) {real, imag} */,
  {32'h401b15e6, 32'h4048a5b4} /* (12, 18, 2) {real, imag} */,
  {32'hc0e79179, 32'hbfd78598} /* (12, 18, 1) {real, imag} */,
  {32'h3fac0611, 32'h411af71e} /* (12, 18, 0) {real, imag} */,
  {32'hc06dbe28, 32'hc0af7bf5} /* (12, 17, 31) {real, imag} */,
  {32'hc14b0194, 32'h40b97bf6} /* (12, 17, 30) {real, imag} */,
  {32'h409c4aaa, 32'hbeee4ce8} /* (12, 17, 29) {real, imag} */,
  {32'hc0046534, 32'hc056f5f3} /* (12, 17, 28) {real, imag} */,
  {32'h3f41e67c, 32'h40db53d2} /* (12, 17, 27) {real, imag} */,
  {32'h409853fd, 32'hc18a42a2} /* (12, 17, 26) {real, imag} */,
  {32'h406c32e3, 32'h40c5d243} /* (12, 17, 25) {real, imag} */,
  {32'hc1662a82, 32'hc163aed8} /* (12, 17, 24) {real, imag} */,
  {32'hbfdf34dc, 32'h41428782} /* (12, 17, 23) {real, imag} */,
  {32'hc07399a7, 32'h3fda526e} /* (12, 17, 22) {real, imag} */,
  {32'h41548c87, 32'h408daf24} /* (12, 17, 21) {real, imag} */,
  {32'h4061c8b7, 32'hc0042c9c} /* (12, 17, 20) {real, imag} */,
  {32'hc0a7082e, 32'hc1088e34} /* (12, 17, 19) {real, imag} */,
  {32'h4083ada6, 32'hc094c1c4} /* (12, 17, 18) {real, imag} */,
  {32'hc060e474, 32'hc018584e} /* (12, 17, 17) {real, imag} */,
  {32'hc0cf8362, 32'hc0e54ba5} /* (12, 17, 16) {real, imag} */,
  {32'hc0f61406, 32'hbff0824c} /* (12, 17, 15) {real, imag} */,
  {32'hc13b465c, 32'h408719aa} /* (12, 17, 14) {real, imag} */,
  {32'hc08d21eb, 32'hbfda4218} /* (12, 17, 13) {real, imag} */,
  {32'hc1053d36, 32'h3f1759dc} /* (12, 17, 12) {real, imag} */,
  {32'h4042cd1e, 32'hc070813e} /* (12, 17, 11) {real, imag} */,
  {32'h41447398, 32'h414e63bd} /* (12, 17, 10) {real, imag} */,
  {32'hbf8f6096, 32'hc0115f1c} /* (12, 17, 9) {real, imag} */,
  {32'hbf826fa4, 32'h40a6ae6a} /* (12, 17, 8) {real, imag} */,
  {32'hc1577d76, 32'h40d90872} /* (12, 17, 7) {real, imag} */,
  {32'hc118b0dd, 32'h40e26087} /* (12, 17, 6) {real, imag} */,
  {32'h4021a312, 32'hc0667816} /* (12, 17, 5) {real, imag} */,
  {32'h41371132, 32'h40d2f912} /* (12, 17, 4) {real, imag} */,
  {32'hc08b4282, 32'hbea561e0} /* (12, 17, 3) {real, imag} */,
  {32'hc0a5fdf8, 32'h3fa41f1e} /* (12, 17, 2) {real, imag} */,
  {32'h409982a7, 32'hc01742f6} /* (12, 17, 1) {real, imag} */,
  {32'h4101092f, 32'hc0fbc172} /* (12, 17, 0) {real, imag} */,
  {32'hc0b7ab8a, 32'h402e1d4e} /* (12, 16, 31) {real, imag} */,
  {32'hc0a8b886, 32'h40b4cb12} /* (12, 16, 30) {real, imag} */,
  {32'hc07f2b97, 32'h4041d87e} /* (12, 16, 29) {real, imag} */,
  {32'h408aa74e, 32'h4147d54a} /* (12, 16, 28) {real, imag} */,
  {32'h40469758, 32'h408a1e37} /* (12, 16, 27) {real, imag} */,
  {32'hc07a28e6, 32'hc08b5b4e} /* (12, 16, 26) {real, imag} */,
  {32'h416167c4, 32'hbe7dfec0} /* (12, 16, 25) {real, imag} */,
  {32'h411e6992, 32'hc03047ef} /* (12, 16, 24) {real, imag} */,
  {32'h40a1e68a, 32'h41568856} /* (12, 16, 23) {real, imag} */,
  {32'hbfb24c68, 32'h40acc2cf} /* (12, 16, 22) {real, imag} */,
  {32'hc1027a9f, 32'h4031efa0} /* (12, 16, 21) {real, imag} */,
  {32'hc0695eae, 32'hc03df524} /* (12, 16, 20) {real, imag} */,
  {32'h3f4c5ba0, 32'hc01d366b} /* (12, 16, 19) {real, imag} */,
  {32'h41418d42, 32'h3f8e0240} /* (12, 16, 18) {real, imag} */,
  {32'h4172caaa, 32'h40492da0} /* (12, 16, 17) {real, imag} */,
  {32'h40896b48, 32'h00000000} /* (12, 16, 16) {real, imag} */,
  {32'h4172caaa, 32'hc0492da0} /* (12, 16, 15) {real, imag} */,
  {32'h41418d42, 32'hbf8e0240} /* (12, 16, 14) {real, imag} */,
  {32'h3f4c5ba0, 32'h401d366b} /* (12, 16, 13) {real, imag} */,
  {32'hc0695eae, 32'h403df524} /* (12, 16, 12) {real, imag} */,
  {32'hc1027a9f, 32'hc031efa0} /* (12, 16, 11) {real, imag} */,
  {32'hbfb24c68, 32'hc0acc2cf} /* (12, 16, 10) {real, imag} */,
  {32'h40a1e68a, 32'hc1568856} /* (12, 16, 9) {real, imag} */,
  {32'h411e6992, 32'h403047ef} /* (12, 16, 8) {real, imag} */,
  {32'h416167c4, 32'h3e7dfec0} /* (12, 16, 7) {real, imag} */,
  {32'hc07a28e6, 32'h408b5b4e} /* (12, 16, 6) {real, imag} */,
  {32'h40469758, 32'hc08a1e37} /* (12, 16, 5) {real, imag} */,
  {32'h408aa74e, 32'hc147d54a} /* (12, 16, 4) {real, imag} */,
  {32'hc07f2b97, 32'hc041d87e} /* (12, 16, 3) {real, imag} */,
  {32'hc0a8b886, 32'hc0b4cb12} /* (12, 16, 2) {real, imag} */,
  {32'hc0b7ab8a, 32'hc02e1d4e} /* (12, 16, 1) {real, imag} */,
  {32'h40d392c0, 32'h00000000} /* (12, 16, 0) {real, imag} */,
  {32'h409982a7, 32'h401742f6} /* (12, 15, 31) {real, imag} */,
  {32'hc0a5fdf8, 32'hbfa41f1e} /* (12, 15, 30) {real, imag} */,
  {32'hc08b4282, 32'h3ea561e0} /* (12, 15, 29) {real, imag} */,
  {32'h41371132, 32'hc0d2f912} /* (12, 15, 28) {real, imag} */,
  {32'h4021a312, 32'h40667816} /* (12, 15, 27) {real, imag} */,
  {32'hc118b0dd, 32'hc0e26087} /* (12, 15, 26) {real, imag} */,
  {32'hc1577d76, 32'hc0d90872} /* (12, 15, 25) {real, imag} */,
  {32'hbf826fa4, 32'hc0a6ae6a} /* (12, 15, 24) {real, imag} */,
  {32'hbf8f6096, 32'h40115f1c} /* (12, 15, 23) {real, imag} */,
  {32'h41447398, 32'hc14e63bd} /* (12, 15, 22) {real, imag} */,
  {32'h4042cd1e, 32'h4070813e} /* (12, 15, 21) {real, imag} */,
  {32'hc1053d36, 32'hbf1759dc} /* (12, 15, 20) {real, imag} */,
  {32'hc08d21eb, 32'h3fda4218} /* (12, 15, 19) {real, imag} */,
  {32'hc13b465c, 32'hc08719aa} /* (12, 15, 18) {real, imag} */,
  {32'hc0f61406, 32'h3ff0824c} /* (12, 15, 17) {real, imag} */,
  {32'hc0cf8362, 32'h40e54ba5} /* (12, 15, 16) {real, imag} */,
  {32'hc060e474, 32'h4018584e} /* (12, 15, 15) {real, imag} */,
  {32'h4083ada6, 32'h4094c1c4} /* (12, 15, 14) {real, imag} */,
  {32'hc0a7082e, 32'h41088e34} /* (12, 15, 13) {real, imag} */,
  {32'h4061c8b7, 32'h40042c9c} /* (12, 15, 12) {real, imag} */,
  {32'h41548c87, 32'hc08daf24} /* (12, 15, 11) {real, imag} */,
  {32'hc07399a7, 32'hbfda526e} /* (12, 15, 10) {real, imag} */,
  {32'hbfdf34dc, 32'hc1428782} /* (12, 15, 9) {real, imag} */,
  {32'hc1662a82, 32'h4163aed8} /* (12, 15, 8) {real, imag} */,
  {32'h406c32e3, 32'hc0c5d243} /* (12, 15, 7) {real, imag} */,
  {32'h409853fd, 32'h418a42a2} /* (12, 15, 6) {real, imag} */,
  {32'h3f41e67c, 32'hc0db53d2} /* (12, 15, 5) {real, imag} */,
  {32'hc0046534, 32'h4056f5f3} /* (12, 15, 4) {real, imag} */,
  {32'h409c4aaa, 32'h3eee4ce8} /* (12, 15, 3) {real, imag} */,
  {32'hc14b0194, 32'hc0b97bf6} /* (12, 15, 2) {real, imag} */,
  {32'hc06dbe28, 32'h40af7bf5} /* (12, 15, 1) {real, imag} */,
  {32'h4101092f, 32'h40fbc172} /* (12, 15, 0) {real, imag} */,
  {32'hc0e79179, 32'h3fd78598} /* (12, 14, 31) {real, imag} */,
  {32'h401b15e6, 32'hc048a5b4} /* (12, 14, 30) {real, imag} */,
  {32'h3fb908a6, 32'hc004b85e} /* (12, 14, 29) {real, imag} */,
  {32'hc16664b1, 32'hc0fd9d26} /* (12, 14, 28) {real, imag} */,
  {32'hc172c10e, 32'h41ab7596} /* (12, 14, 27) {real, imag} */,
  {32'hc0bc2b9c, 32'hbf59e61c} /* (12, 14, 26) {real, imag} */,
  {32'hbe740fc0, 32'hc0544ca6} /* (12, 14, 25) {real, imag} */,
  {32'h4137ecc2, 32'hc11c6160} /* (12, 14, 24) {real, imag} */,
  {32'h411e4a18, 32'hc0ca374c} /* (12, 14, 23) {real, imag} */,
  {32'hbf9c6788, 32'h3fa5a96a} /* (12, 14, 22) {real, imag} */,
  {32'hc0ffcd52, 32'hc0a1c17b} /* (12, 14, 21) {real, imag} */,
  {32'hc0a9b85a, 32'h40b146cd} /* (12, 14, 20) {real, imag} */,
  {32'hc0c16301, 32'h41753cf4} /* (12, 14, 19) {real, imag} */,
  {32'hbf4920b4, 32'hc040929f} /* (12, 14, 18) {real, imag} */,
  {32'hbe11f8e0, 32'hc0e10868} /* (12, 14, 17) {real, imag} */,
  {32'h418acf87, 32'hc145cea3} /* (12, 14, 16) {real, imag} */,
  {32'h400f7ed8, 32'h414dac09} /* (12, 14, 15) {real, imag} */,
  {32'h40d3911a, 32'h3ff3eff0} /* (12, 14, 14) {real, imag} */,
  {32'h411b8c15, 32'hc183ba70} /* (12, 14, 13) {real, imag} */,
  {32'h40b93705, 32'hc10d30c8} /* (12, 14, 12) {real, imag} */,
  {32'hc1595416, 32'h419ad53a} /* (12, 14, 11) {real, imag} */,
  {32'hc0a56c3d, 32'hc15d488a} /* (12, 14, 10) {real, imag} */,
  {32'hbd93c0c0, 32'h4162cb74} /* (12, 14, 9) {real, imag} */,
  {32'hc0034c0c, 32'hc087dcc4} /* (12, 14, 8) {real, imag} */,
  {32'h4031cd35, 32'hc10b6377} /* (12, 14, 7) {real, imag} */,
  {32'hc0b6f300, 32'h4003f87c} /* (12, 14, 6) {real, imag} */,
  {32'hc0d3b863, 32'h41b32638} /* (12, 14, 5) {real, imag} */,
  {32'hc13b83d0, 32'hbf8bf2ec} /* (12, 14, 4) {real, imag} */,
  {32'hc0b4a66b, 32'hc0af07a3} /* (12, 14, 3) {real, imag} */,
  {32'h4090307c, 32'h407d2cdc} /* (12, 14, 2) {real, imag} */,
  {32'hc0817e78, 32'hbfdd81ce} /* (12, 14, 1) {real, imag} */,
  {32'h3fac0611, 32'hc11af71e} /* (12, 14, 0) {real, imag} */,
  {32'h40d8c7cf, 32'h410a5177} /* (12, 13, 31) {real, imag} */,
  {32'hc09b5811, 32'h40b4f2dd} /* (12, 13, 30) {real, imag} */,
  {32'h3eedc580, 32'h3fa54666} /* (12, 13, 29) {real, imag} */,
  {32'h40caeecc, 32'h404f1528} /* (12, 13, 28) {real, imag} */,
  {32'hc1644dd6, 32'hc183020a} /* (12, 13, 27) {real, imag} */,
  {32'h40cea723, 32'h3fbb1a57} /* (12, 13, 26) {real, imag} */,
  {32'h412f3170, 32'hc07731c8} /* (12, 13, 25) {real, imag} */,
  {32'h400cd287, 32'h40b8f510} /* (12, 13, 24) {real, imag} */,
  {32'hc13814f6, 32'hbf89dc84} /* (12, 13, 23) {real, imag} */,
  {32'h41a25326, 32'h41ad1844} /* (12, 13, 22) {real, imag} */,
  {32'hc0bf0222, 32'h3fe7d49c} /* (12, 13, 21) {real, imag} */,
  {32'hbf2ec320, 32'h3ee3d140} /* (12, 13, 20) {real, imag} */,
  {32'h3f5bcea4, 32'hc071e649} /* (12, 13, 19) {real, imag} */,
  {32'h411ab7a6, 32'h40c7ad18} /* (12, 13, 18) {real, imag} */,
  {32'h3fa1a1d2, 32'hc039fbc8} /* (12, 13, 17) {real, imag} */,
  {32'hc10062f2, 32'h3f093d2c} /* (12, 13, 16) {real, imag} */,
  {32'h411492f8, 32'hc034e552} /* (12, 13, 15) {real, imag} */,
  {32'hc03db11c, 32'hc11f5429} /* (12, 13, 14) {real, imag} */,
  {32'h4161cc70, 32'h40ff0e7c} /* (12, 13, 13) {real, imag} */,
  {32'h41344d4f, 32'hc13251eb} /* (12, 13, 12) {real, imag} */,
  {32'hc0b3bc6a, 32'hc08834a9} /* (12, 13, 11) {real, imag} */,
  {32'hc1180126, 32'hc1029b13} /* (12, 13, 10) {real, imag} */,
  {32'hc0e3249d, 32'h3dfebee0} /* (12, 13, 9) {real, imag} */,
  {32'hbe9b0ff0, 32'hc0f9c87e} /* (12, 13, 8) {real, imag} */,
  {32'h418cfb45, 32'hc0851d0a} /* (12, 13, 7) {real, imag} */,
  {32'hc0ddb408, 32'hc09b1316} /* (12, 13, 6) {real, imag} */,
  {32'h4137ee46, 32'hc0c70ab4} /* (12, 13, 5) {real, imag} */,
  {32'h4086036e, 32'h41c010a4} /* (12, 13, 4) {real, imag} */,
  {32'hc0a39940, 32'hc0d401b2} /* (12, 13, 3) {real, imag} */,
  {32'h410f0c9d, 32'hbf7f1520} /* (12, 13, 2) {real, imag} */,
  {32'h4003ccea, 32'h404277a7} /* (12, 13, 1) {real, imag} */,
  {32'h4013f162, 32'h40a09a76} /* (12, 13, 0) {real, imag} */,
  {32'hc0be874d, 32'h401329a6} /* (12, 12, 31) {real, imag} */,
  {32'hc141bcf4, 32'hc0d708b8} /* (12, 12, 30) {real, imag} */,
  {32'h4091ea00, 32'hc1a198bc} /* (12, 12, 29) {real, imag} */,
  {32'hc1a18d62, 32'hc1185a0e} /* (12, 12, 28) {real, imag} */,
  {32'h411a6eef, 32'h410e1ac0} /* (12, 12, 27) {real, imag} */,
  {32'hc1c00daa, 32'h411d8693} /* (12, 12, 26) {real, imag} */,
  {32'h413f21a0, 32'h412eb222} /* (12, 12, 25) {real, imag} */,
  {32'h406170ae, 32'h40457417} /* (12, 12, 24) {real, imag} */,
  {32'h40d78f7f, 32'hc11e9134} /* (12, 12, 23) {real, imag} */,
  {32'hc01d0888, 32'hc192ca60} /* (12, 12, 22) {real, imag} */,
  {32'hc1080318, 32'hc0fef1de} /* (12, 12, 21) {real, imag} */,
  {32'h4143922c, 32'hc16bcc95} /* (12, 12, 20) {real, imag} */,
  {32'hc02d76ca, 32'h4087159a} /* (12, 12, 19) {real, imag} */,
  {32'hc0eeb2ab, 32'h419872ae} /* (12, 12, 18) {real, imag} */,
  {32'h3f17fe48, 32'h402c5759} /* (12, 12, 17) {real, imag} */,
  {32'hbf8dc800, 32'h411a3c52} /* (12, 12, 16) {real, imag} */,
  {32'hc1487338, 32'hc1b45976} /* (12, 12, 15) {real, imag} */,
  {32'h4101f0a9, 32'h3ffdb680} /* (12, 12, 14) {real, imag} */,
  {32'h3ffd2d48, 32'hc10ac66a} /* (12, 12, 13) {real, imag} */,
  {32'h4194f2aa, 32'hc0b4e7f0} /* (12, 12, 12) {real, imag} */,
  {32'hbfa70f42, 32'h41786d17} /* (12, 12, 11) {real, imag} */,
  {32'h41a5f23c, 32'h418e306e} /* (12, 12, 10) {real, imag} */,
  {32'h3de10580, 32'h41afb08a} /* (12, 12, 9) {real, imag} */,
  {32'h40cd632e, 32'hbeb02380} /* (12, 12, 8) {real, imag} */,
  {32'h3f405360, 32'h41049ec0} /* (12, 12, 7) {real, imag} */,
  {32'hc0867068, 32'hc05b58c5} /* (12, 12, 6) {real, imag} */,
  {32'hc11436e9, 32'h409e677e} /* (12, 12, 5) {real, imag} */,
  {32'hc06a3c6c, 32'h415f0697} /* (12, 12, 4) {real, imag} */,
  {32'hc023b7c8, 32'hc1661765} /* (12, 12, 3) {real, imag} */,
  {32'hc1266d18, 32'h4024d354} /* (12, 12, 2) {real, imag} */,
  {32'h40f337c8, 32'hbf1418a0} /* (12, 12, 1) {real, imag} */,
  {32'h4172f83e, 32'h40ad0092} /* (12, 12, 0) {real, imag} */,
  {32'hc13fcec4, 32'hc1967562} /* (12, 11, 31) {real, imag} */,
  {32'h40d363fc, 32'h412be2e8} /* (12, 11, 30) {real, imag} */,
  {32'h3fe45410, 32'hc04cb406} /* (12, 11, 29) {real, imag} */,
  {32'hbf5a4168, 32'h3f3040c0} /* (12, 11, 28) {real, imag} */,
  {32'h40ed1526, 32'hc16b689e} /* (12, 11, 27) {real, imag} */,
  {32'h412ba9e8, 32'h3ffbf840} /* (12, 11, 26) {real, imag} */,
  {32'hc1eb4003, 32'hc19f3120} /* (12, 11, 25) {real, imag} */,
  {32'h41539253, 32'h410fdd7c} /* (12, 11, 24) {real, imag} */,
  {32'h40ca8dd2, 32'h412e6fc1} /* (12, 11, 23) {real, imag} */,
  {32'h40e54954, 32'h3fe7e868} /* (12, 11, 22) {real, imag} */,
  {32'h414bbf9e, 32'h4167477e} /* (12, 11, 21) {real, imag} */,
  {32'hc0a6ae40, 32'hc15eb3c2} /* (12, 11, 20) {real, imag} */,
  {32'h41c734fa, 32'h3f4d33dc} /* (12, 11, 19) {real, imag} */,
  {32'hc1486a28, 32'hbfc17662} /* (12, 11, 18) {real, imag} */,
  {32'h40f092f5, 32'h41109226} /* (12, 11, 17) {real, imag} */,
  {32'hc155b970, 32'hc0cbf572} /* (12, 11, 16) {real, imag} */,
  {32'hc0df6904, 32'hc08f6480} /* (12, 11, 15) {real, imag} */,
  {32'hc07aa75d, 32'hc13de7ae} /* (12, 11, 14) {real, imag} */,
  {32'h405eaaac, 32'hc0933988} /* (12, 11, 13) {real, imag} */,
  {32'hc13219e8, 32'hc012b9ce} /* (12, 11, 12) {real, imag} */,
  {32'hbf5c20a8, 32'h41669013} /* (12, 11, 11) {real, imag} */,
  {32'h3e8c34a0, 32'h40d3f7b6} /* (12, 11, 10) {real, imag} */,
  {32'hbf2f3f30, 32'hc184f9f2} /* (12, 11, 9) {real, imag} */,
  {32'hbf8f15a0, 32'h3f821db8} /* (12, 11, 8) {real, imag} */,
  {32'h40a28a16, 32'h40d698ec} /* (12, 11, 7) {real, imag} */,
  {32'hc07d1fda, 32'hc1852fba} /* (12, 11, 6) {real, imag} */,
  {32'hc0decbde, 32'h413b6016} /* (12, 11, 5) {real, imag} */,
  {32'h3f826e04, 32'h3f3ce460} /* (12, 11, 4) {real, imag} */,
  {32'h41cc6d1a, 32'hc0afa69c} /* (12, 11, 3) {real, imag} */,
  {32'hc15f6022, 32'h408e3276} /* (12, 11, 2) {real, imag} */,
  {32'hc2034f73, 32'hc183b45a} /* (12, 11, 1) {real, imag} */,
  {32'hc18a8386, 32'hc0be7d22} /* (12, 11, 0) {real, imag} */,
  {32'h404abc3a, 32'h417acf8d} /* (12, 10, 31) {real, imag} */,
  {32'hc088eda4, 32'h3bf3f800} /* (12, 10, 30) {real, imag} */,
  {32'hc0e26c69, 32'hc0f32102} /* (12, 10, 29) {real, imag} */,
  {32'h4087cbfa, 32'h408c8678} /* (12, 10, 28) {real, imag} */,
  {32'hc15de302, 32'h41206066} /* (12, 10, 27) {real, imag} */,
  {32'h4041c780, 32'hc15dd260} /* (12, 10, 26) {real, imag} */,
  {32'hc1839a38, 32'h407ccb74} /* (12, 10, 25) {real, imag} */,
  {32'h417c55c3, 32'hc17c540c} /* (12, 10, 24) {real, imag} */,
  {32'hc1a078e2, 32'h416f731e} /* (12, 10, 23) {real, imag} */,
  {32'h411a7328, 32'h3f5635a8} /* (12, 10, 22) {real, imag} */,
  {32'h414faca5, 32'hc1587aac} /* (12, 10, 21) {real, imag} */,
  {32'h3fa06ae4, 32'hc01c2027} /* (12, 10, 20) {real, imag} */,
  {32'h413b9b44, 32'hc0b4e42a} /* (12, 10, 19) {real, imag} */,
  {32'hbf4ae3b0, 32'h410ad5ee} /* (12, 10, 18) {real, imag} */,
  {32'hc044ab12, 32'hc08a335e} /* (12, 10, 17) {real, imag} */,
  {32'hc16c8e7e, 32'h407c09dd} /* (12, 10, 16) {real, imag} */,
  {32'h41051009, 32'h413a4702} /* (12, 10, 15) {real, imag} */,
  {32'h3f227404, 32'hbfad560c} /* (12, 10, 14) {real, imag} */,
  {32'h4066aef2, 32'hc12f487a} /* (12, 10, 13) {real, imag} */,
  {32'hc0ad19d0, 32'hc1655c6c} /* (12, 10, 12) {real, imag} */,
  {32'h3ff092a0, 32'hc0f888d9} /* (12, 10, 11) {real, imag} */,
  {32'hc163e382, 32'h410fcf0f} /* (12, 10, 10) {real, imag} */,
  {32'h4093d84c, 32'hc0148162} /* (12, 10, 9) {real, imag} */,
  {32'hbfd82168, 32'hc0815e4e} /* (12, 10, 8) {real, imag} */,
  {32'h4106ba6c, 32'h4178915e} /* (12, 10, 7) {real, imag} */,
  {32'h40265c2a, 32'hc1802e80} /* (12, 10, 6) {real, imag} */,
  {32'h4192f1d9, 32'hc18ec082} /* (12, 10, 5) {real, imag} */,
  {32'hc12b3b36, 32'h41be0441} /* (12, 10, 4) {real, imag} */,
  {32'h4055a988, 32'hbfa4b378} /* (12, 10, 3) {real, imag} */,
  {32'hc0ab7df5, 32'hc1d16798} /* (12, 10, 2) {real, imag} */,
  {32'h407e1902, 32'h40dc5910} /* (12, 10, 1) {real, imag} */,
  {32'hbfcdcbf4, 32'hc017835a} /* (12, 10, 0) {real, imag} */,
  {32'hc1ac26a2, 32'h41581372} /* (12, 9, 31) {real, imag} */,
  {32'h40f139b0, 32'hc08ba34c} /* (12, 9, 30) {real, imag} */,
  {32'h406fb2a9, 32'hc0f5a3de} /* (12, 9, 29) {real, imag} */,
  {32'h40930aa4, 32'hc11f0be6} /* (12, 9, 28) {real, imag} */,
  {32'hc15fdec0, 32'h409180ca} /* (12, 9, 27) {real, imag} */,
  {32'hc011b4d8, 32'h40176184} /* (12, 9, 26) {real, imag} */,
  {32'hc10bfbea, 32'hc0b09ac7} /* (12, 9, 25) {real, imag} */,
  {32'hc1e9029f, 32'hc073fe1a} /* (12, 9, 24) {real, imag} */,
  {32'h4067e15b, 32'h4144c022} /* (12, 9, 23) {real, imag} */,
  {32'h404731f8, 32'hc0c52e51} /* (12, 9, 22) {real, imag} */,
  {32'hc0d4d71b, 32'h405e34ba} /* (12, 9, 21) {real, imag} */,
  {32'h40acd43c, 32'h3f088848} /* (12, 9, 20) {real, imag} */,
  {32'h416b7e76, 32'h4050ba5d} /* (12, 9, 19) {real, imag} */,
  {32'h402be536, 32'hc096da72} /* (12, 9, 18) {real, imag} */,
  {32'h4062ee80, 32'h40d6a21a} /* (12, 9, 17) {real, imag} */,
  {32'hbf159970, 32'h40c8ca82} /* (12, 9, 16) {real, imag} */,
  {32'h404f1389, 32'h3df37140} /* (12, 9, 15) {real, imag} */,
  {32'h40afeba0, 32'hc081e7d2} /* (12, 9, 14) {real, imag} */,
  {32'hc14508e0, 32'h410603a0} /* (12, 9, 13) {real, imag} */,
  {32'hc105bdbf, 32'hc0c26312} /* (12, 9, 12) {real, imag} */,
  {32'hc17ee0a2, 32'hbfe47501} /* (12, 9, 11) {real, imag} */,
  {32'hc144eb94, 32'hc1104fb8} /* (12, 9, 10) {real, imag} */,
  {32'h41a8d9da, 32'hc081fdc0} /* (12, 9, 9) {real, imag} */,
  {32'hbfc8f9b8, 32'hc08550f6} /* (12, 9, 8) {real, imag} */,
  {32'h41347e58, 32'h41010b1f} /* (12, 9, 7) {real, imag} */,
  {32'hc18d0231, 32'h4156ed2e} /* (12, 9, 6) {real, imag} */,
  {32'hc10e991e, 32'h416c5cd1} /* (12, 9, 5) {real, imag} */,
  {32'hc123440a, 32'h410694be} /* (12, 9, 4) {real, imag} */,
  {32'h4194694d, 32'hc1a73b66} /* (12, 9, 3) {real, imag} */,
  {32'hc132cf29, 32'hc1450dc2} /* (12, 9, 2) {real, imag} */,
  {32'h420c88e0, 32'h417ba136} /* (12, 9, 1) {real, imag} */,
  {32'hc0d846d4, 32'hc1362a85} /* (12, 9, 0) {real, imag} */,
  {32'hc2368768, 32'hc1c3492a} /* (12, 8, 31) {real, imag} */,
  {32'h41e7b91d, 32'h414f02ca} /* (12, 8, 30) {real, imag} */,
  {32'h403e2a16, 32'hc17d3084} /* (12, 8, 29) {real, imag} */,
  {32'h4109fe48, 32'hc180a829} /* (12, 8, 28) {real, imag} */,
  {32'h41ac1f4b, 32'hc11a1a5d} /* (12, 8, 27) {real, imag} */,
  {32'h4057b212, 32'h41189799} /* (12, 8, 26) {real, imag} */,
  {32'h3fbb2a06, 32'hc12a99d8} /* (12, 8, 25) {real, imag} */,
  {32'h40265bd6, 32'h4114c569} /* (12, 8, 24) {real, imag} */,
  {32'h3fcaf790, 32'hc11e647d} /* (12, 8, 23) {real, imag} */,
  {32'hc14c24f9, 32'h418b88c2} /* (12, 8, 22) {real, imag} */,
  {32'h418af3dd, 32'hbe0b2610} /* (12, 8, 21) {real, imag} */,
  {32'h41843314, 32'hc0c0ca62} /* (12, 8, 20) {real, imag} */,
  {32'hc1602cc6, 32'hc10ace42} /* (12, 8, 19) {real, imag} */,
  {32'h4185b8f0, 32'h3fa29cb2} /* (12, 8, 18) {real, imag} */,
  {32'h40f55ed6, 32'hc0845e9e} /* (12, 8, 17) {real, imag} */,
  {32'h408bee82, 32'hc0832daf} /* (12, 8, 16) {real, imag} */,
  {32'h4072397a, 32'h4150a0ba} /* (12, 8, 15) {real, imag} */,
  {32'hc1090ca4, 32'hc13d1332} /* (12, 8, 14) {real, imag} */,
  {32'hc1dfd550, 32'h4182e46c} /* (12, 8, 13) {real, imag} */,
  {32'h41214265, 32'h41f0923e} /* (12, 8, 12) {real, imag} */,
  {32'h408d3d5d, 32'hc191cd84} /* (12, 8, 11) {real, imag} */,
  {32'h4198462c, 32'h40575580} /* (12, 8, 10) {real, imag} */,
  {32'h4077b3d4, 32'h3f832c72} /* (12, 8, 9) {real, imag} */,
  {32'h41296b24, 32'hc02807c6} /* (12, 8, 8) {real, imag} */,
  {32'hc1902ce7, 32'hbfa94934} /* (12, 8, 7) {real, imag} */,
  {32'h413bce2b, 32'hc16fa4ac} /* (12, 8, 6) {real, imag} */,
  {32'h41b8f709, 32'hc1125a6d} /* (12, 8, 5) {real, imag} */,
  {32'hc1fe4fbb, 32'hc201c3e9} /* (12, 8, 4) {real, imag} */,
  {32'hc0cc5146, 32'h40d2beb6} /* (12, 8, 3) {real, imag} */,
  {32'h411f72d3, 32'h419c418b} /* (12, 8, 2) {real, imag} */,
  {32'hc2271c54, 32'h40336e38} /* (12, 8, 1) {real, imag} */,
  {32'hc1a18586, 32'hc1e59562} /* (12, 8, 0) {real, imag} */,
  {32'h418864b8, 32'hc186813c} /* (12, 7, 31) {real, imag} */,
  {32'h400ba543, 32'hc1a83cd6} /* (12, 7, 30) {real, imag} */,
  {32'hc0a66d90, 32'h401902ab} /* (12, 7, 29) {real, imag} */,
  {32'hbe771ae0, 32'h4100fbe1} /* (12, 7, 28) {real, imag} */,
  {32'hc00de3ca, 32'hc159da9e} /* (12, 7, 27) {real, imag} */,
  {32'h3fd8d4d9, 32'h4114ef5a} /* (12, 7, 26) {real, imag} */,
  {32'h418e6da7, 32'h4180ff3c} /* (12, 7, 25) {real, imag} */,
  {32'hc0c69ca6, 32'hc16da232} /* (12, 7, 24) {real, imag} */,
  {32'hc168ce72, 32'hc0ecdbfa} /* (12, 7, 23) {real, imag} */,
  {32'hc0494967, 32'h419576f0} /* (12, 7, 22) {real, imag} */,
  {32'h41b1bf63, 32'hc130db68} /* (12, 7, 21) {real, imag} */,
  {32'h40cba3a8, 32'h410a611a} /* (12, 7, 20) {real, imag} */,
  {32'hc0db93a7, 32'h40d40646} /* (12, 7, 19) {real, imag} */,
  {32'h3f39c740, 32'h40d03f0a} /* (12, 7, 18) {real, imag} */,
  {32'hc0baef45, 32'h4107c313} /* (12, 7, 17) {real, imag} */,
  {32'hc13a4e07, 32'h411ec426} /* (12, 7, 16) {real, imag} */,
  {32'h41195c5a, 32'hc05a43c5} /* (12, 7, 15) {real, imag} */,
  {32'hc0bfcbee, 32'hbf8a4222} /* (12, 7, 14) {real, imag} */,
  {32'hbfcee135, 32'hc1a09ca0} /* (12, 7, 13) {real, imag} */,
  {32'h4076e958, 32'hbfea1e50} /* (12, 7, 12) {real, imag} */,
  {32'h41c6678c, 32'hc109de8a} /* (12, 7, 11) {real, imag} */,
  {32'h4137f084, 32'h40ceae74} /* (12, 7, 10) {real, imag} */,
  {32'hc129ec26, 32'hc1102867} /* (12, 7, 9) {real, imag} */,
  {32'h41373284, 32'hc0492c72} /* (12, 7, 8) {real, imag} */,
  {32'hc0ee6d63, 32'h3ffc670f} /* (12, 7, 7) {real, imag} */,
  {32'h410e4e3f, 32'hbed027e0} /* (12, 7, 6) {real, imag} */,
  {32'hbe104e60, 32'h40edab12} /* (12, 7, 5) {real, imag} */,
  {32'hc109305b, 32'h41c35708} /* (12, 7, 4) {real, imag} */,
  {32'hc1abaeea, 32'h41a19736} /* (12, 7, 3) {real, imag} */,
  {32'hc12ad936, 32'hc10de49f} /* (12, 7, 2) {real, imag} */,
  {32'h41b2866c, 32'h419a62ae} /* (12, 7, 1) {real, imag} */,
  {32'h3f8a5948, 32'h411dbf1c} /* (12, 7, 0) {real, imag} */,
  {32'h4148d60a, 32'hc189383b} /* (12, 6, 31) {real, imag} */,
  {32'h42070773, 32'hc02dedc6} /* (12, 6, 30) {real, imag} */,
  {32'h4170c5af, 32'hc18cd5b2} /* (12, 6, 29) {real, imag} */,
  {32'hc0a373d8, 32'hc18ec897} /* (12, 6, 28) {real, imag} */,
  {32'hc04d6dd6, 32'h4177188a} /* (12, 6, 27) {real, imag} */,
  {32'hbf527f58, 32'h410adc55} /* (12, 6, 26) {real, imag} */,
  {32'h3f95db3c, 32'hc0fa869f} /* (12, 6, 25) {real, imag} */,
  {32'hc12c8ba4, 32'h40ae2e86} /* (12, 6, 24) {real, imag} */,
  {32'hbf2dade8, 32'hc091acab} /* (12, 6, 23) {real, imag} */,
  {32'h41d6f712, 32'hc130ef90} /* (12, 6, 22) {real, imag} */,
  {32'h3ff59cd4, 32'hc0498209} /* (12, 6, 21) {real, imag} */,
  {32'h41025b10, 32'hbfdda844} /* (12, 6, 20) {real, imag} */,
  {32'h4145368a, 32'h416748ca} /* (12, 6, 19) {real, imag} */,
  {32'hc1277344, 32'hc0178d2d} /* (12, 6, 18) {real, imag} */,
  {32'h40f80efa, 32'hc1106fff} /* (12, 6, 17) {real, imag} */,
  {32'hc0f8fa08, 32'h407247e3} /* (12, 6, 16) {real, imag} */,
  {32'h40293c3f, 32'hbf4e4a20} /* (12, 6, 15) {real, imag} */,
  {32'h4115d21d, 32'hc14410c2} /* (12, 6, 14) {real, imag} */,
  {32'hc0b7ac2e, 32'h40cb43c5} /* (12, 6, 13) {real, imag} */,
  {32'hbfd79764, 32'h40ab156b} /* (12, 6, 12) {real, imag} */,
  {32'hc022c197, 32'h3f15855c} /* (12, 6, 11) {real, imag} */,
  {32'hc194698a, 32'hc1435a5e} /* (12, 6, 10) {real, imag} */,
  {32'hc1f1ccb5, 32'hc020763e} /* (12, 6, 9) {real, imag} */,
  {32'h40f6e78d, 32'hc11d95cf} /* (12, 6, 8) {real, imag} */,
  {32'hc1209ccd, 32'h40c3c6fc} /* (12, 6, 7) {real, imag} */,
  {32'h3f8748fe, 32'hc18dff78} /* (12, 6, 6) {real, imag} */,
  {32'h416c1961, 32'hc1eb224e} /* (12, 6, 5) {real, imag} */,
  {32'h41276cbc, 32'hc186d6ae} /* (12, 6, 4) {real, imag} */,
  {32'hbfda4105, 32'h415058cc} /* (12, 6, 3) {real, imag} */,
  {32'h40e21dd1, 32'hc0a82dc7} /* (12, 6, 2) {real, imag} */,
  {32'h41c0688c, 32'hc1256c48} /* (12, 6, 1) {real, imag} */,
  {32'h40d79f30, 32'h41892917} /* (12, 6, 0) {real, imag} */,
  {32'hc2d779ce, 32'hc181bdaa} /* (12, 5, 31) {real, imag} */,
  {32'h41a0296b, 32'h41439b3d} /* (12, 5, 30) {real, imag} */,
  {32'hc0546108, 32'h3e714600} /* (12, 5, 29) {real, imag} */,
  {32'hc15d801a, 32'h421fcc3e} /* (12, 5, 28) {real, imag} */,
  {32'h413d4f8e, 32'h41db9038} /* (12, 5, 27) {real, imag} */,
  {32'hc08a0898, 32'hc04530d6} /* (12, 5, 26) {real, imag} */,
  {32'h4111643e, 32'hc17be684} /* (12, 5, 25) {real, imag} */,
  {32'h41646d1a, 32'hc1a14e6a} /* (12, 5, 24) {real, imag} */,
  {32'h413bef24, 32'hc02990b2} /* (12, 5, 23) {real, imag} */,
  {32'h4136a4df, 32'hc0ce5ece} /* (12, 5, 22) {real, imag} */,
  {32'h4195e960, 32'hbfe3c09e} /* (12, 5, 21) {real, imag} */,
  {32'h40a19a58, 32'hc06bb680} /* (12, 5, 20) {real, imag} */,
  {32'hc04710e5, 32'h41bbc358} /* (12, 5, 19) {real, imag} */,
  {32'hc10e6636, 32'hc04b7434} /* (12, 5, 18) {real, imag} */,
  {32'h403a5002, 32'hc0ff7cd6} /* (12, 5, 17) {real, imag} */,
  {32'h40faf88e, 32'h3e299bc0} /* (12, 5, 16) {real, imag} */,
  {32'h40096b4e, 32'h3fb23a2e} /* (12, 5, 15) {real, imag} */,
  {32'hc1a7de4e, 32'h40d2b6f0} /* (12, 5, 14) {real, imag} */,
  {32'hc0e751e9, 32'h40e34ba0} /* (12, 5, 13) {real, imag} */,
  {32'h41646224, 32'hbfaa26f8} /* (12, 5, 12) {real, imag} */,
  {32'h40ef5cb0, 32'h413b6d1c} /* (12, 5, 11) {real, imag} */,
  {32'hc11a86c0, 32'h414bbc92} /* (12, 5, 10) {real, imag} */,
  {32'h41ca58fd, 32'h41a897eb} /* (12, 5, 9) {real, imag} */,
  {32'h413e32db, 32'hbfbd766c} /* (12, 5, 8) {real, imag} */,
  {32'hc156146b, 32'hc0549664} /* (12, 5, 7) {real, imag} */,
  {32'h410ef28b, 32'h40b88fac} /* (12, 5, 6) {real, imag} */,
  {32'h4222f932, 32'h41ca88df} /* (12, 5, 5) {real, imag} */,
  {32'hc0518a98, 32'hc20fa1ff} /* (12, 5, 4) {real, imag} */,
  {32'h3f969efc, 32'hc1247fc8} /* (12, 5, 3) {real, imag} */,
  {32'h4196b9ec, 32'h423e9b2e} /* (12, 5, 2) {real, imag} */,
  {32'hc28f1aa0, 32'hc29778cd} /* (12, 5, 1) {real, imag} */,
  {32'hc2b36c5a, 32'hc1d1c64b} /* (12, 5, 0) {real, imag} */,
  {32'h41f27b0d, 32'h4286c60a} /* (12, 4, 31) {real, imag} */,
  {32'hc2dcea31, 32'hc29ef263} /* (12, 4, 30) {real, imag} */,
  {32'h4115a513, 32'hc11e767e} /* (12, 4, 29) {real, imag} */,
  {32'h420d7230, 32'h40d87f00} /* (12, 4, 28) {real, imag} */,
  {32'hc1a1bf81, 32'hc209961c} /* (12, 4, 27) {real, imag} */,
  {32'hbfb09fd0, 32'hc0e1f966} /* (12, 4, 26) {real, imag} */,
  {32'h41c1bb7c, 32'h3f87b904} /* (12, 4, 25) {real, imag} */,
  {32'h4123a800, 32'hc1637b8e} /* (12, 4, 24) {real, imag} */,
  {32'hc10eedca, 32'hc156346c} /* (12, 4, 23) {real, imag} */,
  {32'hc046726b, 32'hc0eb4496} /* (12, 4, 22) {real, imag} */,
  {32'hc1311b24, 32'h41be53de} /* (12, 4, 21) {real, imag} */,
  {32'h412cc460, 32'hc0c9beae} /* (12, 4, 20) {real, imag} */,
  {32'hbefd0cf0, 32'hc0dcf40a} /* (12, 4, 19) {real, imag} */,
  {32'hc13ff452, 32'h4047fd40} /* (12, 4, 18) {real, imag} */,
  {32'h4082338f, 32'h41835316} /* (12, 4, 17) {real, imag} */,
  {32'h3fb7afbe, 32'hbfbb251e} /* (12, 4, 16) {real, imag} */,
  {32'hc04c54b7, 32'h405d78bf} /* (12, 4, 15) {real, imag} */,
  {32'h40dd89da, 32'hc0fea952} /* (12, 4, 14) {real, imag} */,
  {32'hc08fada2, 32'h411db3ae} /* (12, 4, 13) {real, imag} */,
  {32'hc16678b6, 32'hbf8de550} /* (12, 4, 12) {real, imag} */,
  {32'hc162df5e, 32'hc0d92f7f} /* (12, 4, 11) {real, imag} */,
  {32'hbf8847ca, 32'h41b29544} /* (12, 4, 10) {real, imag} */,
  {32'hc1868d64, 32'h3f9128a8} /* (12, 4, 9) {real, imag} */,
  {32'h3fa5d519, 32'hc21f6337} /* (12, 4, 8) {real, imag} */,
  {32'hbff00cdf, 32'hbffd57e8} /* (12, 4, 7) {real, imag} */,
  {32'hc164fdca, 32'h4153d029} /* (12, 4, 6) {real, imag} */,
  {32'h418753c1, 32'hc2469815} /* (12, 4, 5) {real, imag} */,
  {32'h3fcab608, 32'h415d0d77} /* (12, 4, 4) {real, imag} */,
  {32'h41a63a80, 32'h410b4e3e} /* (12, 4, 3) {real, imag} */,
  {32'hc28a8819, 32'hc2a57cce} /* (12, 4, 2) {real, imag} */,
  {32'h4337d9a4, 32'h42032bea} /* (12, 4, 1) {real, imag} */,
  {32'h4223de4b, 32'hc0ad0483} /* (12, 4, 0) {real, imag} */,
  {32'hc32f9341, 32'h4286f384} /* (12, 3, 31) {real, imag} */,
  {32'h428bdc71, 32'hc2f6a746} /* (12, 3, 30) {real, imag} */,
  {32'hc1c2fd55, 32'h4171830f} /* (12, 3, 29) {real, imag} */,
  {32'h4245e4f9, 32'h4223d5ea} /* (12, 3, 28) {real, imag} */,
  {32'hc1a6ba80, 32'h4083b5f0} /* (12, 3, 27) {real, imag} */,
  {32'hc0af6f4c, 32'h417ea88b} /* (12, 3, 26) {real, imag} */,
  {32'h40e79dbc, 32'h402aa85f} /* (12, 3, 25) {real, imag} */,
  {32'h41b30560, 32'hc1ccfaf7} /* (12, 3, 24) {real, imag} */,
  {32'h41c0d3d6, 32'h4089f5b6} /* (12, 3, 23) {real, imag} */,
  {32'h400f9476, 32'hc0f131d8} /* (12, 3, 22) {real, imag} */,
  {32'hc10648f9, 32'h40093eac} /* (12, 3, 21) {real, imag} */,
  {32'hc09c74ba, 32'h3f7e70c4} /* (12, 3, 20) {real, imag} */,
  {32'hc0b8b918, 32'hc0cad76c} /* (12, 3, 19) {real, imag} */,
  {32'hc131414e, 32'hc14da552} /* (12, 3, 18) {real, imag} */,
  {32'hbefd6064, 32'h4130ecf8} /* (12, 3, 17) {real, imag} */,
  {32'h3fab2892, 32'h4103207f} /* (12, 3, 16) {real, imag} */,
  {32'h3d26f400, 32'hc02872c3} /* (12, 3, 15) {real, imag} */,
  {32'h4140d174, 32'hc1b66366} /* (12, 3, 14) {real, imag} */,
  {32'h40e0bfcd, 32'h3f411428} /* (12, 3, 13) {real, imag} */,
  {32'hbf777728, 32'h41002321} /* (12, 3, 12) {real, imag} */,
  {32'h3e1b77f8, 32'h3ff0360a} /* (12, 3, 11) {real, imag} */,
  {32'h415aeefa, 32'hc0d73c36} /* (12, 3, 10) {real, imag} */,
  {32'hc0f32a41, 32'h3fa1388e} /* (12, 3, 9) {real, imag} */,
  {32'hc11f6a52, 32'h4191faf9} /* (12, 3, 8) {real, imag} */,
  {32'h41421172, 32'hc1840ec2} /* (12, 3, 7) {real, imag} */,
  {32'h41e0d454, 32'h41a74a15} /* (12, 3, 6) {real, imag} */,
  {32'h3f6fd260, 32'h420c5d78} /* (12, 3, 5) {real, imag} */,
  {32'hc1a7b10e, 32'h404836a2} /* (12, 3, 4) {real, imag} */,
  {32'hc1a2e696, 32'hc03b32f8} /* (12, 3, 3) {real, imag} */,
  {32'hc128edd3, 32'hc2cfd050} /* (12, 3, 2) {real, imag} */,
  {32'h4312a3e9, 32'h42ea5577} /* (12, 3, 1) {real, imag} */,
  {32'hc10d2149, 32'h40c7578c} /* (12, 3, 0) {real, imag} */,
  {32'hc497a83c, 32'hc178cf0d} /* (12, 2, 31) {real, imag} */,
  {32'h4410d81c, 32'hc31eaae8} /* (12, 2, 30) {real, imag} */,
  {32'h414652fa, 32'h41d9fe6a} /* (12, 2, 29) {real, imag} */,
  {32'hc1ddc005, 32'h4264f300} /* (12, 2, 28) {real, imag} */,
  {32'h420a77f5, 32'hc27ff0ed} /* (12, 2, 27) {real, imag} */,
  {32'h41c01a4f, 32'hc0038ca4} /* (12, 2, 26) {real, imag} */,
  {32'hc1a564aa, 32'h401e9024} /* (12, 2, 25) {real, imag} */,
  {32'h409fef56, 32'hc22d5feb} /* (12, 2, 24) {real, imag} */,
  {32'hc155106e, 32'h4062f3b2} /* (12, 2, 23) {real, imag} */,
  {32'hbf2616c0, 32'h411de8c6} /* (12, 2, 22) {real, imag} */,
  {32'h41982ee2, 32'hc0e80d46} /* (12, 2, 21) {real, imag} */,
  {32'hc18883d2, 32'h4024e536} /* (12, 2, 20) {real, imag} */,
  {32'h3e64a3a0, 32'h40c07170} /* (12, 2, 19) {real, imag} */,
  {32'h3f07fa99, 32'hc1956b41} /* (12, 2, 18) {real, imag} */,
  {32'hc1223768, 32'h411c3d1c} /* (12, 2, 17) {real, imag} */,
  {32'h402fd85c, 32'h405e13b1} /* (12, 2, 16) {real, imag} */,
  {32'hc1370633, 32'hc09610f8} /* (12, 2, 15) {real, imag} */,
  {32'h419fb44e, 32'h41b52066} /* (12, 2, 14) {real, imag} */,
  {32'h3f580674, 32'hc0876737} /* (12, 2, 13) {real, imag} */,
  {32'h40c9d1cf, 32'h417f73f2} /* (12, 2, 12) {real, imag} */,
  {32'h40035d5e, 32'h41d94946} /* (12, 2, 11) {real, imag} */,
  {32'hc09c5747, 32'hc003ad38} /* (12, 2, 10) {real, imag} */,
  {32'hc15da304, 32'hbfd6421c} /* (12, 2, 9) {real, imag} */,
  {32'h41923302, 32'h416edf45} /* (12, 2, 8) {real, imag} */,
  {32'hc1baad82, 32'hc0af3b90} /* (12, 2, 7) {real, imag} */,
  {32'h40d54688, 32'h41edd322} /* (12, 2, 6) {real, imag} */,
  {32'h421fe174, 32'h4294b361} /* (12, 2, 5) {real, imag} */,
  {32'hc2bf031d, 32'hc2613fe7} /* (12, 2, 4) {real, imag} */,
  {32'h416ad44f, 32'h404dec46} /* (12, 2, 3) {real, imag} */,
  {32'h43b3884d, 32'hc30b266a} /* (12, 2, 2) {real, imag} */,
  {32'hc4277074, 32'h429ec049} /* (12, 2, 1) {real, imag} */,
  {32'hc4170c5e, 32'hc2ae9758} /* (12, 2, 0) {real, imag} */,
  {32'h44c82ad4, 32'hc39e442a} /* (12, 1, 31) {real, imag} */,
  {32'hc3c996dd, 32'h419d7d75} /* (12, 1, 30) {real, imag} */,
  {32'h3ecc7e60, 32'h41d14ad1} /* (12, 1, 29) {real, imag} */,
  {32'h42a8dd31, 32'h4243f438} /* (12, 1, 28) {real, imag} */,
  {32'hc302d0df, 32'hc192267f} /* (12, 1, 27) {real, imag} */,
  {32'h4137bf7e, 32'hbfc3a2e8} /* (12, 1, 26) {real, imag} */,
  {32'h3ef52830, 32'hc0c3bb92} /* (12, 1, 25) {real, imag} */,
  {32'hc163a5e7, 32'hbfc53760} /* (12, 1, 24) {real, imag} */,
  {32'hc1870fa2, 32'hc0eff2d8} /* (12, 1, 23) {real, imag} */,
  {32'h41d95c2a, 32'h41d1dde3} /* (12, 1, 22) {real, imag} */,
  {32'hc1ba5049, 32'h41d08e26} /* (12, 1, 21) {real, imag} */,
  {32'hc1b4d5fa, 32'h40148662} /* (12, 1, 20) {real, imag} */,
  {32'hc0bb366d, 32'h413b3332} /* (12, 1, 19) {real, imag} */,
  {32'h418bc016, 32'h409f11d7} /* (12, 1, 18) {real, imag} */,
  {32'h4124ae14, 32'h411f5256} /* (12, 1, 17) {real, imag} */,
  {32'h3f1d3b54, 32'h40045edd} /* (12, 1, 16) {real, imag} */,
  {32'h410515ae, 32'h40d3341d} /* (12, 1, 15) {real, imag} */,
  {32'h40ca4ffc, 32'hc051755e} /* (12, 1, 14) {real, imag} */,
  {32'hc023e17f, 32'hc035f07d} /* (12, 1, 13) {real, imag} */,
  {32'h41091fa2, 32'hc16dba92} /* (12, 1, 12) {real, imag} */,
  {32'hbf86ff92, 32'hc1aca6b3} /* (12, 1, 11) {real, imag} */,
  {32'hc110a74c, 32'hc0627cf8} /* (12, 1, 10) {real, imag} */,
  {32'hc0818bd4, 32'hc0b55bcb} /* (12, 1, 9) {real, imag} */,
  {32'hc118265b, 32'hc22d55c8} /* (12, 1, 8) {real, imag} */,
  {32'h419c62ee, 32'h40fe0faa} /* (12, 1, 7) {real, imag} */,
  {32'hbfbdca10, 32'hc1f86efc} /* (12, 1, 6) {real, imag} */,
  {32'hc297b820, 32'hc1330fcc} /* (12, 1, 5) {real, imag} */,
  {32'hc1d5e5f8, 32'h428a5466} /* (12, 1, 4) {real, imag} */,
  {32'hc17c7a62, 32'hbeb1b2c0} /* (12, 1, 3) {real, imag} */,
  {32'hc4178599, 32'hc4040624} /* (12, 1, 2) {real, imag} */,
  {32'h450a1a57, 32'h44a42047} /* (12, 1, 1) {real, imag} */,
  {32'h45027137, 32'h42fc5dd8} /* (12, 1, 0) {real, imag} */,
  {32'h449cf0bc, 32'hc483701f} /* (12, 0, 31) {real, imag} */,
  {32'hc3430253, 32'h439168d5} /* (12, 0, 30) {real, imag} */,
  {32'hc23b3ad8, 32'h4154aeb0} /* (12, 0, 29) {real, imag} */,
  {32'h3fc0c4de, 32'h42336765} /* (12, 0, 28) {real, imag} */,
  {32'hc2542466, 32'h40806153} /* (12, 0, 27) {real, imag} */,
  {32'hc20cf3cc, 32'hc136a980} /* (12, 0, 26) {real, imag} */,
  {32'h3fc2a6f6, 32'hc1f96b02} /* (12, 0, 25) {real, imag} */,
  {32'hc08e3e02, 32'h41f1e5c6} /* (12, 0, 24) {real, imag} */,
  {32'hc06688be, 32'h41947590} /* (12, 0, 23) {real, imag} */,
  {32'hc1d69249, 32'h4157f8e4} /* (12, 0, 22) {real, imag} */,
  {32'hc058c978, 32'hc09d5898} /* (12, 0, 21) {real, imag} */,
  {32'hc0ef1c08, 32'hc01b6488} /* (12, 0, 20) {real, imag} */,
  {32'hbf05d79c, 32'h41356a60} /* (12, 0, 19) {real, imag} */,
  {32'hbee29920, 32'hc162bfce} /* (12, 0, 18) {real, imag} */,
  {32'hc0144bf5, 32'hc121eb9c} /* (12, 0, 17) {real, imag} */,
  {32'h404175e4, 32'h00000000} /* (12, 0, 16) {real, imag} */,
  {32'hc0144bf5, 32'h4121eb9c} /* (12, 0, 15) {real, imag} */,
  {32'hbee29920, 32'h4162bfce} /* (12, 0, 14) {real, imag} */,
  {32'hbf05d79c, 32'hc1356a60} /* (12, 0, 13) {real, imag} */,
  {32'hc0ef1c08, 32'h401b6488} /* (12, 0, 12) {real, imag} */,
  {32'hc058c978, 32'h409d5898} /* (12, 0, 11) {real, imag} */,
  {32'hc1d69249, 32'hc157f8e4} /* (12, 0, 10) {real, imag} */,
  {32'hc06688be, 32'hc1947590} /* (12, 0, 9) {real, imag} */,
  {32'hc08e3e02, 32'hc1f1e5c6} /* (12, 0, 8) {real, imag} */,
  {32'h3fc2a6f6, 32'h41f96b02} /* (12, 0, 7) {real, imag} */,
  {32'hc20cf3cc, 32'h4136a980} /* (12, 0, 6) {real, imag} */,
  {32'hc2542466, 32'hc0806153} /* (12, 0, 5) {real, imag} */,
  {32'h3fc0c4de, 32'hc2336765} /* (12, 0, 4) {real, imag} */,
  {32'hc23b3ad8, 32'hc154aeb0} /* (12, 0, 3) {real, imag} */,
  {32'hc3430253, 32'hc39168d5} /* (12, 0, 2) {real, imag} */,
  {32'h449cf0bc, 32'h4483701f} /* (12, 0, 1) {real, imag} */,
  {32'h44fee150, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h4519e3e7, 32'hc4afb621} /* (11, 31, 31) {real, imag} */,
  {32'hc423c4f9, 32'h4411f708} /* (11, 31, 30) {real, imag} */,
  {32'h419a8a95, 32'hc12f0cb7} /* (11, 31, 29) {real, imag} */,
  {32'hc1890778, 32'hc206aac5} /* (11, 31, 28) {real, imag} */,
  {32'hc2c977e0, 32'h41db971f} /* (11, 31, 27) {real, imag} */,
  {32'hc21ff0dc, 32'h419ed53d} /* (11, 31, 26) {real, imag} */,
  {32'h415375ce, 32'hc15247be} /* (11, 31, 25) {real, imag} */,
  {32'hc1adc14c, 32'h41d476fd} /* (11, 31, 24) {real, imag} */,
  {32'hc06a4a50, 32'hc149b67f} /* (11, 31, 23) {real, imag} */,
  {32'hc01b7a58, 32'h41cc444a} /* (11, 31, 22) {real, imag} */,
  {32'hc0be8105, 32'hc00599f8} /* (11, 31, 21) {real, imag} */,
  {32'h41010d18, 32'h3f2add90} /* (11, 31, 20) {real, imag} */,
  {32'h40aead9e, 32'h40d33833} /* (11, 31, 19) {real, imag} */,
  {32'h4064843e, 32'h41494fd0} /* (11, 31, 18) {real, imag} */,
  {32'h4082144c, 32'hc15e22b7} /* (11, 31, 17) {real, imag} */,
  {32'h408d58e0, 32'hc00b5178} /* (11, 31, 16) {real, imag} */,
  {32'h4062abba, 32'h40327d7b} /* (11, 31, 15) {real, imag} */,
  {32'h41492734, 32'hc0acc043} /* (11, 31, 14) {real, imag} */,
  {32'hc154bc87, 32'h41011ae7} /* (11, 31, 13) {real, imag} */,
  {32'hbef4ff30, 32'h40ebd418} /* (11, 31, 12) {real, imag} */,
  {32'hc1a4b3b3, 32'hc183fd85} /* (11, 31, 11) {real, imag} */,
  {32'h41b0ff67, 32'hc15d148e} /* (11, 31, 10) {real, imag} */,
  {32'hc0a78aaa, 32'hbf96b98c} /* (11, 31, 9) {real, imag} */,
  {32'hc1bbe2a0, 32'hc135c5c2} /* (11, 31, 8) {real, imag} */,
  {32'hbf1e8988, 32'h3f38fcc0} /* (11, 31, 7) {real, imag} */,
  {32'hc13e4c19, 32'h41179d96} /* (11, 31, 6) {real, imag} */,
  {32'hc2cbfb52, 32'h41c2caa2} /* (11, 31, 5) {real, imag} */,
  {32'h4292dd6a, 32'hc299fd52} /* (11, 31, 4) {real, imag} */,
  {32'hc2060f91, 32'hc1392c88} /* (11, 31, 3) {real, imag} */,
  {32'hc3d0f2a6, 32'hc22397b6} /* (11, 31, 2) {real, imag} */,
  {32'h44d828b8, 32'h43a8e473} /* (11, 31, 1) {real, imag} */,
  {32'h450eea0c, 32'hc30f22b4} /* (11, 31, 0) {real, imag} */,
  {32'hc4322ee0, 32'hc314410d} /* (11, 30, 31) {real, imag} */,
  {32'h43cfd23c, 32'h4314bb92} /* (11, 30, 30) {real, imag} */,
  {32'h41c20d4e, 32'hc1283537} /* (11, 30, 29) {real, imag} */,
  {32'hc2b8eb7c, 32'h4260db92} /* (11, 30, 28) {real, imag} */,
  {32'h4203386e, 32'hc2a7a44e} /* (11, 30, 27) {real, imag} */,
  {32'h40fd25a2, 32'hc1806988} /* (11, 30, 26) {real, imag} */,
  {32'h40fc800a, 32'h412df187} /* (11, 30, 25) {real, imag} */,
  {32'h41b9ea27, 32'h40bbcba8} /* (11, 30, 24) {real, imag} */,
  {32'hc09ec5e5, 32'hc03048d6} /* (11, 30, 23) {real, imag} */,
  {32'hc169774a, 32'hc15d6098} /* (11, 30, 22) {real, imag} */,
  {32'hc01d7fdb, 32'hc12a87b8} /* (11, 30, 21) {real, imag} */,
  {32'hc0a61eab, 32'hc11d2899} /* (11, 30, 20) {real, imag} */,
  {32'hc08631ae, 32'hc1372442} /* (11, 30, 19) {real, imag} */,
  {32'hc0f3e864, 32'hc1743ab2} /* (11, 30, 18) {real, imag} */,
  {32'hc052eabc, 32'h3f0399b4} /* (11, 30, 17) {real, imag} */,
  {32'h410832fd, 32'hc1146250} /* (11, 30, 16) {real, imag} */,
  {32'hc04e5bdc, 32'h3f1afbc8} /* (11, 30, 15) {real, imag} */,
  {32'h405b82a4, 32'h4024a3b0} /* (11, 30, 14) {real, imag} */,
  {32'h40c43f56, 32'h40a49ffc} /* (11, 30, 13) {real, imag} */,
  {32'h403c91c2, 32'h40ed56de} /* (11, 30, 12) {real, imag} */,
  {32'h40d4685b, 32'h4187d2e6} /* (11, 30, 11) {real, imag} */,
  {32'hc0b819b6, 32'hbfd7072e} /* (11, 30, 10) {real, imag} */,
  {32'hc144d794, 32'hbfdc5d61} /* (11, 30, 9) {real, imag} */,
  {32'h419d2549, 32'h41a8191e} /* (11, 30, 8) {real, imag} */,
  {32'h4007a0e0, 32'hc199f4ae} /* (11, 30, 7) {real, imag} */,
  {32'h41a733b4, 32'hbfae574c} /* (11, 30, 6) {real, imag} */,
  {32'h4265d2a9, 32'h4278bc99} /* (11, 30, 5) {real, imag} */,
  {32'hc19dab10, 32'hc295816a} /* (11, 30, 4) {real, imag} */,
  {32'h41663a8e, 32'hc18f9b23} /* (11, 30, 3) {real, imag} */,
  {32'h44146cf5, 32'h4329b6b9} /* (11, 30, 2) {real, imag} */,
  {32'hc4a2d3e7, 32'h42a5fec6} /* (11, 30, 1) {real, imag} */,
  {32'hc4305fe6, 32'h42b997dd} /* (11, 30, 0) {real, imag} */,
  {32'h42fa8474, 32'hc2b84752} /* (11, 29, 31) {real, imag} */,
  {32'h40ea39a6, 32'h42bf8072} /* (11, 29, 30) {real, imag} */,
  {32'hc1e791f8, 32'hc19ded94} /* (11, 29, 29) {real, imag} */,
  {32'hc1f0392a, 32'hc12a3156} /* (11, 29, 28) {real, imag} */,
  {32'hc0dc2517, 32'hc1845129} /* (11, 29, 27) {real, imag} */,
  {32'h412bb0d2, 32'hc1733f0e} /* (11, 29, 26) {real, imag} */,
  {32'h404ea700, 32'h416af6a7} /* (11, 29, 25) {real, imag} */,
  {32'h3e9138e0, 32'h40f0f7d0} /* (11, 29, 24) {real, imag} */,
  {32'hc0716e68, 32'hc041a13a} /* (11, 29, 23) {real, imag} */,
  {32'h3f9710a0, 32'hc0ed1b36} /* (11, 29, 22) {real, imag} */,
  {32'h4108b0bc, 32'hbd8c3880} /* (11, 29, 21) {real, imag} */,
  {32'hc1012b32, 32'hc06951ac} /* (11, 29, 20) {real, imag} */,
  {32'h40ecedaa, 32'h40886d88} /* (11, 29, 19) {real, imag} */,
  {32'h41676c87, 32'h41a51786} /* (11, 29, 18) {real, imag} */,
  {32'hc13b24df, 32'hc10e0241} /* (11, 29, 17) {real, imag} */,
  {32'h40bd5da3, 32'hc061fd4c} /* (11, 29, 16) {real, imag} */,
  {32'h40bd38b9, 32'hc1841238} /* (11, 29, 15) {real, imag} */,
  {32'h4134affd, 32'h4020026a} /* (11, 29, 14) {real, imag} */,
  {32'hc187b2e5, 32'h40814518} /* (11, 29, 13) {real, imag} */,
  {32'h4064c866, 32'hc0547bf8} /* (11, 29, 12) {real, imag} */,
  {32'h4122f6f6, 32'hc158ef20} /* (11, 29, 11) {real, imag} */,
  {32'hc0a4b3df, 32'hbfbcf700} /* (11, 29, 10) {real, imag} */,
  {32'h3f71a5d8, 32'h4194ef0d} /* (11, 29, 9) {real, imag} */,
  {32'h417b6f24, 32'h41054884} /* (11, 29, 8) {real, imag} */,
  {32'h4156db18, 32'hc154215b} /* (11, 29, 7) {real, imag} */,
  {32'h41768f00, 32'hc1be8ddb} /* (11, 29, 6) {real, imag} */,
  {32'hc21c72a8, 32'hc1ab8ddc} /* (11, 29, 5) {real, imag} */,
  {32'h421165ae, 32'hc223b7ce} /* (11, 29, 4) {real, imag} */,
  {32'hc184aeb0, 32'hc0715d71} /* (11, 29, 3) {real, imag} */,
  {32'h4275944e, 32'h4311ba98} /* (11, 29, 2) {real, imag} */,
  {32'hc30b19d8, 32'hc2a69cd3} /* (11, 29, 1) {real, imag} */,
  {32'h40d248fc, 32'hc14f0fc0} /* (11, 29, 0) {real, imag} */,
  {32'h43408df8, 32'hc21aa2ac} /* (11, 28, 31) {real, imag} */,
  {32'hc2a5b734, 32'h426af7c2} /* (11, 28, 30) {real, imag} */,
  {32'h41c4c972, 32'hbf8db810} /* (11, 28, 29) {real, imag} */,
  {32'h408864dc, 32'hc21d08d7} /* (11, 28, 28) {real, imag} */,
  {32'h41944aaa, 32'h41bd6c61} /* (11, 28, 27) {real, imag} */,
  {32'hc161ea33, 32'hc1ccde3e} /* (11, 28, 26) {real, imag} */,
  {32'h415d8def, 32'h4146b910} /* (11, 28, 25) {real, imag} */,
  {32'hc18470a1, 32'h419d0aa0} /* (11, 28, 24) {real, imag} */,
  {32'hc0efe966, 32'hc1202c9a} /* (11, 28, 23) {real, imag} */,
  {32'hc1ac3ae6, 32'h409685fd} /* (11, 28, 22) {real, imag} */,
  {32'h40261298, 32'h408a158f} /* (11, 28, 21) {real, imag} */,
  {32'h40974fb1, 32'hbfb6711f} /* (11, 28, 20) {real, imag} */,
  {32'hc03d8d3c, 32'hbf85ca08} /* (11, 28, 19) {real, imag} */,
  {32'h41347fd0, 32'h4154a1c6} /* (11, 28, 18) {real, imag} */,
  {32'hbfd4d751, 32'h400c8a8c} /* (11, 28, 17) {real, imag} */,
  {32'h3f5e33e4, 32'hc089c9a2} /* (11, 28, 16) {real, imag} */,
  {32'h40a20678, 32'hc09290b5} /* (11, 28, 15) {real, imag} */,
  {32'hc0d22f46, 32'h41a19aa7} /* (11, 28, 14) {real, imag} */,
  {32'h40bf2560, 32'hc0bcba06} /* (11, 28, 13) {real, imag} */,
  {32'h419d46bd, 32'hc10f87bd} /* (11, 28, 12) {real, imag} */,
  {32'hc160655e, 32'hc099afab} /* (11, 28, 11) {real, imag} */,
  {32'hc0f226ea, 32'h4080b536} /* (11, 28, 10) {real, imag} */,
  {32'h41947f2e, 32'h411ab064} /* (11, 28, 9) {real, imag} */,
  {32'hbf92162c, 32'h4107a07a} /* (11, 28, 8) {real, imag} */,
  {32'h41992fcc, 32'hc10f1535} /* (11, 28, 7) {real, imag} */,
  {32'hc0df84ac, 32'h40992348} /* (11, 28, 6) {real, imag} */,
  {32'hc0972a33, 32'hc1067687} /* (11, 28, 5) {real, imag} */,
  {32'h40acb6dd, 32'h3fcc8da0} /* (11, 28, 4) {real, imag} */,
  {32'hc12a0525, 32'h4156b3d5} /* (11, 28, 3) {real, imag} */,
  {32'hc2eacd1f, 32'h42aeaad3} /* (11, 28, 2) {real, imag} */,
  {32'h41f12752, 32'hc2b171a3} /* (11, 28, 1) {real, imag} */,
  {32'h42371a2a, 32'h3ed3c900} /* (11, 28, 0) {real, imag} */,
  {32'hc152afba, 32'h429b86e8} /* (11, 27, 31) {real, imag} */,
  {32'h419c603c, 32'hc1e2af0e} /* (11, 27, 30) {real, imag} */,
  {32'hc1e1aeae, 32'h411ab5d8} /* (11, 27, 29) {real, imag} */,
  {32'h40b385ed, 32'h410fdb2b} /* (11, 27, 28) {real, imag} */,
  {32'h420c3aec, 32'h3d65d000} /* (11, 27, 27) {real, imag} */,
  {32'hc206c45e, 32'h3f643060} /* (11, 27, 26) {real, imag} */,
  {32'h40c57cf0, 32'hc1266bd1} /* (11, 27, 25) {real, imag} */,
  {32'h41958817, 32'hc1b456b8} /* (11, 27, 24) {real, imag} */,
  {32'hc0d808dd, 32'h40f59015} /* (11, 27, 23) {real, imag} */,
  {32'hc16c06de, 32'hc13d5356} /* (11, 27, 22) {real, imag} */,
  {32'h41a7ecc2, 32'h4117f42c} /* (11, 27, 21) {real, imag} */,
  {32'h41199806, 32'hc1a1c47b} /* (11, 27, 20) {real, imag} */,
  {32'h41193244, 32'hc0d5e48a} /* (11, 27, 19) {real, imag} */,
  {32'hc0d68376, 32'hc0ddd840} /* (11, 27, 18) {real, imag} */,
  {32'h411ad574, 32'h40c69c88} /* (11, 27, 17) {real, imag} */,
  {32'hc0e6084e, 32'hc0532214} /* (11, 27, 16) {real, imag} */,
  {32'h3edb8f30, 32'hc00f20ed} /* (11, 27, 15) {real, imag} */,
  {32'hc0ec6be4, 32'hc0ae0a89} /* (11, 27, 14) {real, imag} */,
  {32'h4193b0f3, 32'hc152a230} /* (11, 27, 13) {real, imag} */,
  {32'h40dd3ebd, 32'hbe1af880} /* (11, 27, 12) {real, imag} */,
  {32'hc0bb3320, 32'h418b8876} /* (11, 27, 11) {real, imag} */,
  {32'h4072929e, 32'hc0bd5cf2} /* (11, 27, 10) {real, imag} */,
  {32'hc026fa62, 32'h410064bc} /* (11, 27, 9) {real, imag} */,
  {32'h416d21c6, 32'h42154064} /* (11, 27, 8) {real, imag} */,
  {32'h40a87fe2, 32'h404d7b0d} /* (11, 27, 7) {real, imag} */,
  {32'h4144eb58, 32'h4119232a} /* (11, 27, 6) {real, imag} */,
  {32'h413895f0, 32'hc19b62d4} /* (11, 27, 5) {real, imag} */,
  {32'hc17f6a43, 32'hc24c7d5a} /* (11, 27, 4) {real, imag} */,
  {32'hc1ac5d22, 32'hc0c05c8f} /* (11, 27, 3) {real, imag} */,
  {32'h41310ea8, 32'h3ec55ca0} /* (11, 27, 2) {real, imag} */,
  {32'hc2dd9576, 32'h40822142} /* (11, 27, 1) {real, imag} */,
  {32'hc26523e2, 32'h41b3bf32} /* (11, 27, 0) {real, imag} */,
  {32'h40c96e12, 32'hc07a914c} /* (11, 26, 31) {real, imag} */,
  {32'h41bd3b27, 32'hc02ec9d4} /* (11, 26, 30) {real, imag} */,
  {32'h412cf6ce, 32'hc13b53ce} /* (11, 26, 29) {real, imag} */,
  {32'h4057e907, 32'hbf8121ee} /* (11, 26, 28) {real, imag} */,
  {32'h405e31f8, 32'h40ff9437} /* (11, 26, 27) {real, imag} */,
  {32'h41678efc, 32'h41116e6f} /* (11, 26, 26) {real, imag} */,
  {32'h40b0c996, 32'hc0c38d3f} /* (11, 26, 25) {real, imag} */,
  {32'hc131b418, 32'h41a06d98} /* (11, 26, 24) {real, imag} */,
  {32'hc121182b, 32'h400bfc3c} /* (11, 26, 23) {real, imag} */,
  {32'hc03fbdf4, 32'hc0ce27d4} /* (11, 26, 22) {real, imag} */,
  {32'h3f928438, 32'h41977d73} /* (11, 26, 21) {real, imag} */,
  {32'hbfc4be28, 32'h413d48fb} /* (11, 26, 20) {real, imag} */,
  {32'h3f5834ba, 32'hc0f39882} /* (11, 26, 19) {real, imag} */,
  {32'hc0b887f2, 32'hc0a08380} /* (11, 26, 18) {real, imag} */,
  {32'hbfa420db, 32'hbf845aae} /* (11, 26, 17) {real, imag} */,
  {32'h409365f0, 32'hc0160636} /* (11, 26, 16) {real, imag} */,
  {32'h410eadfe, 32'h4153b2f1} /* (11, 26, 15) {real, imag} */,
  {32'hc0a8c3f6, 32'hc11c6a6e} /* (11, 26, 14) {real, imag} */,
  {32'hc0b4c180, 32'hc17721e5} /* (11, 26, 13) {real, imag} */,
  {32'h3f9137b0, 32'h40fd4931} /* (11, 26, 12) {real, imag} */,
  {32'h409dd059, 32'hc1202712} /* (11, 26, 11) {real, imag} */,
  {32'h41772a30, 32'hc1222b18} /* (11, 26, 10) {real, imag} */,
  {32'h40e4c837, 32'hc1a7a0c4} /* (11, 26, 9) {real, imag} */,
  {32'hc02f5070, 32'hc19b8af7} /* (11, 26, 8) {real, imag} */,
  {32'hc0b778a6, 32'h412446f7} /* (11, 26, 7) {real, imag} */,
  {32'h411ccf90, 32'hc1cd0c5c} /* (11, 26, 6) {real, imag} */,
  {32'h41a71be8, 32'hbf2172e0} /* (11, 26, 5) {real, imag} */,
  {32'h41713f90, 32'h4203cec3} /* (11, 26, 4) {real, imag} */,
  {32'h4091186f, 32'h4152a84f} /* (11, 26, 3) {real, imag} */,
  {32'h3f2ec7f0, 32'h419a41e2} /* (11, 26, 2) {real, imag} */,
  {32'h41f382c9, 32'h42232261} /* (11, 26, 1) {real, imag} */,
  {32'h4078911e, 32'hc199aa50} /* (11, 26, 0) {real, imag} */,
  {32'hc060d314, 32'hc116a4fc} /* (11, 25, 31) {real, imag} */,
  {32'hc06a312c, 32'hc078a121} /* (11, 25, 30) {real, imag} */,
  {32'h400b8ac8, 32'h406e98b8} /* (11, 25, 29) {real, imag} */,
  {32'h41ae6631, 32'hc0b3dd2e} /* (11, 25, 28) {real, imag} */,
  {32'hc1cb1748, 32'h40669f6a} /* (11, 25, 27) {real, imag} */,
  {32'h4111be26, 32'h42033c4d} /* (11, 25, 26) {real, imag} */,
  {32'h40e46a5a, 32'hc189aafa} /* (11, 25, 25) {real, imag} */,
  {32'h41776976, 32'h40805d6e} /* (11, 25, 24) {real, imag} */,
  {32'hc053c95a, 32'h3fa56820} /* (11, 25, 23) {real, imag} */,
  {32'h41514df9, 32'hc0d29eee} /* (11, 25, 22) {real, imag} */,
  {32'h411414b0, 32'h40714dfa} /* (11, 25, 21) {real, imag} */,
  {32'hc0c22bf9, 32'h407c8c97} /* (11, 25, 20) {real, imag} */,
  {32'hc0b237b0, 32'hc11fc0a6} /* (11, 25, 19) {real, imag} */,
  {32'hc0857f89, 32'h3fd06940} /* (11, 25, 18) {real, imag} */,
  {32'hc0692234, 32'hc0499aee} /* (11, 25, 17) {real, imag} */,
  {32'hc10c16fe, 32'hc14322db} /* (11, 25, 16) {real, imag} */,
  {32'hc099e815, 32'h411055f4} /* (11, 25, 15) {real, imag} */,
  {32'hc1236167, 32'hbf3ecba8} /* (11, 25, 14) {real, imag} */,
  {32'h419a8ff8, 32'hc203f69d} /* (11, 25, 13) {real, imag} */,
  {32'h408ee328, 32'hbfa431d7} /* (11, 25, 12) {real, imag} */,
  {32'h411e146e, 32'hc172cda1} /* (11, 25, 11) {real, imag} */,
  {32'hc0968f50, 32'hc1470a82} /* (11, 25, 10) {real, imag} */,
  {32'hc15f1173, 32'hc12355d0} /* (11, 25, 9) {real, imag} */,
  {32'hc1fd756e, 32'h414a1301} /* (11, 25, 8) {real, imag} */,
  {32'h419e7bb1, 32'h3e5fcf80} /* (11, 25, 7) {real, imag} */,
  {32'hc1212222, 32'h407766e0} /* (11, 25, 6) {real, imag} */,
  {32'h412651bb, 32'hc121b3fe} /* (11, 25, 5) {real, imag} */,
  {32'hc0af5151, 32'hc0deb02a} /* (11, 25, 4) {real, imag} */,
  {32'h416c3f48, 32'hc12d2d1a} /* (11, 25, 3) {real, imag} */,
  {32'hc10cbe28, 32'hbf9c4440} /* (11, 25, 2) {real, imag} */,
  {32'h41ad2a66, 32'hc11a4ffc} /* (11, 25, 1) {real, imag} */,
  {32'h411efa4e, 32'hc1015e98} /* (11, 25, 0) {real, imag} */,
  {32'hc204a9f2, 32'h413331fa} /* (11, 24, 31) {real, imag} */,
  {32'h42153914, 32'hc1adfb5d} /* (11, 24, 30) {real, imag} */,
  {32'hc070239e, 32'h40fc8c1d} /* (11, 24, 29) {real, imag} */,
  {32'hc200dcdc, 32'h40e926af} /* (11, 24, 28) {real, imag} */,
  {32'h3ff41750, 32'hc12874d9} /* (11, 24, 27) {real, imag} */,
  {32'h40ef565e, 32'hc15bfcbf} /* (11, 24, 26) {real, imag} */,
  {32'hc1a15946, 32'h411bf3ab} /* (11, 24, 25) {real, imag} */,
  {32'hc15dd500, 32'h402dc656} /* (11, 24, 24) {real, imag} */,
  {32'hc155ce7a, 32'h41811965} /* (11, 24, 23) {real, imag} */,
  {32'h40e3c7f9, 32'hc1647665} /* (11, 24, 22) {real, imag} */,
  {32'hc0c4d19c, 32'hc182e78f} /* (11, 24, 21) {real, imag} */,
  {32'h413833d1, 32'h417a3d9e} /* (11, 24, 20) {real, imag} */,
  {32'hc0cdceea, 32'h40b78920} /* (11, 24, 19) {real, imag} */,
  {32'h4153b056, 32'hc13773e8} /* (11, 24, 18) {real, imag} */,
  {32'hc18f04f8, 32'hc014091a} /* (11, 24, 17) {real, imag} */,
  {32'hbedec990, 32'hc02e279a} /* (11, 24, 16) {real, imag} */,
  {32'hc0452532, 32'hc0b95ec6} /* (11, 24, 15) {real, imag} */,
  {32'h4118ede9, 32'hbf8b25cc} /* (11, 24, 14) {real, imag} */,
  {32'hbf82f46f, 32'h3fd12ee8} /* (11, 24, 13) {real, imag} */,
  {32'h4185e238, 32'hc089b4d3} /* (11, 24, 12) {real, imag} */,
  {32'h40be4f85, 32'h40b6f008} /* (11, 24, 11) {real, imag} */,
  {32'h41a12279, 32'hc02445e2} /* (11, 24, 10) {real, imag} */,
  {32'h4081bd6e, 32'hbf086570} /* (11, 24, 9) {real, imag} */,
  {32'hc17e0448, 32'h412e5000} /* (11, 24, 8) {real, imag} */,
  {32'h41112d4e, 32'h41bef202} /* (11, 24, 7) {real, imag} */,
  {32'h3f8d93e8, 32'hc2238c64} /* (11, 24, 6) {real, imag} */,
  {32'h3f5aabb0, 32'h411da75e} /* (11, 24, 5) {real, imag} */,
  {32'h41476264, 32'hc11808f9} /* (11, 24, 4) {real, imag} */,
  {32'hc209217c, 32'hc06abc1e} /* (11, 24, 3) {real, imag} */,
  {32'h42098232, 32'h40e77cc2} /* (11, 24, 2) {real, imag} */,
  {32'hc25a8b79, 32'h41f51222} /* (11, 24, 1) {real, imag} */,
  {32'h3fd10ab4, 32'h419e97e1} /* (11, 24, 0) {real, imag} */,
  {32'h40f0aee9, 32'hc19c7f16} /* (11, 23, 31) {real, imag} */,
  {32'hc02c88ba, 32'h41ca0b98} /* (11, 23, 30) {real, imag} */,
  {32'h41369645, 32'h414a50e5} /* (11, 23, 29) {real, imag} */,
  {32'hc19b5f7a, 32'hbf46ec5c} /* (11, 23, 28) {real, imag} */,
  {32'h4040ac38, 32'hbfc02a8c} /* (11, 23, 27) {real, imag} */,
  {32'h403c9064, 32'hc02d84bc} /* (11, 23, 26) {real, imag} */,
  {32'hc05dc92d, 32'h419799ac} /* (11, 23, 25) {real, imag} */,
  {32'hc13e460c, 32'h418ec476} /* (11, 23, 24) {real, imag} */,
  {32'h4010ead4, 32'hc1bfa93a} /* (11, 23, 23) {real, imag} */,
  {32'hc128e8e6, 32'hc189faa8} /* (11, 23, 22) {real, imag} */,
  {32'hc101576e, 32'hbed522d0} /* (11, 23, 21) {real, imag} */,
  {32'h4134be96, 32'h41af811e} /* (11, 23, 20) {real, imag} */,
  {32'hc1bff504, 32'h4115b854} /* (11, 23, 19) {real, imag} */,
  {32'h3e88e448, 32'hbf8f42a4} /* (11, 23, 18) {real, imag} */,
  {32'hc04f503f, 32'hbd52cfc0} /* (11, 23, 17) {real, imag} */,
  {32'hc089bd6c, 32'h406ad762} /* (11, 23, 16) {real, imag} */,
  {32'hc042613f, 32'hc0a56aea} /* (11, 23, 15) {real, imag} */,
  {32'hbe097f40, 32'hc10dbfaa} /* (11, 23, 14) {real, imag} */,
  {32'h4206eaa8, 32'h41065e67} /* (11, 23, 13) {real, imag} */,
  {32'h408282d8, 32'hc14bb1ab} /* (11, 23, 12) {real, imag} */,
  {32'hc12ad22d, 32'h41418e8c} /* (11, 23, 11) {real, imag} */,
  {32'hc0a07753, 32'h41c4f3b6} /* (11, 23, 10) {real, imag} */,
  {32'hc087df60, 32'hc128f6ba} /* (11, 23, 9) {real, imag} */,
  {32'h40e07521, 32'hc17464f5} /* (11, 23, 8) {real, imag} */,
  {32'h3e5e8d80, 32'hc13241a2} /* (11, 23, 7) {real, imag} */,
  {32'h41786a6f, 32'h415de02e} /* (11, 23, 6) {real, imag} */,
  {32'hc10c7099, 32'hc00061ee} /* (11, 23, 5) {real, imag} */,
  {32'hc0895366, 32'h4078bf2c} /* (11, 23, 4) {real, imag} */,
  {32'h41101d72, 32'hbf9d8090} /* (11, 23, 3) {real, imag} */,
  {32'h414d0668, 32'h419ccfe2} /* (11, 23, 2) {real, imag} */,
  {32'hc2184f52, 32'hc184d277} /* (11, 23, 1) {real, imag} */,
  {32'h3fb538c0, 32'h3ff0d664} /* (11, 23, 0) {real, imag} */,
  {32'hc0a0c462, 32'hc1d37303} /* (11, 22, 31) {real, imag} */,
  {32'h4118ce9f, 32'h415f67af} /* (11, 22, 30) {real, imag} */,
  {32'h3fa2fa94, 32'hc17e02ba} /* (11, 22, 29) {real, imag} */,
  {32'h413dd00e, 32'hc1ddffd4} /* (11, 22, 28) {real, imag} */,
  {32'h41d3c16c, 32'h411bd967} /* (11, 22, 27) {real, imag} */,
  {32'h40fa3b61, 32'h41ae1520} /* (11, 22, 26) {real, imag} */,
  {32'hc0f268c6, 32'h4018f59f} /* (11, 22, 25) {real, imag} */,
  {32'hbf882b3e, 32'h40c8ed3e} /* (11, 22, 24) {real, imag} */,
  {32'h416af9ec, 32'hc1031f08} /* (11, 22, 23) {real, imag} */,
  {32'hbf86bd9c, 32'h419387fd} /* (11, 22, 22) {real, imag} */,
  {32'h3f22d1e0, 32'h3eea53ec} /* (11, 22, 21) {real, imag} */,
  {32'hbf8e4ae4, 32'h4009aee4} /* (11, 22, 20) {real, imag} */,
  {32'h403092fd, 32'hc11dc1d2} /* (11, 22, 19) {real, imag} */,
  {32'h40abbcd6, 32'h3c303700} /* (11, 22, 18) {real, imag} */,
  {32'hc0d3228e, 32'hc0da562f} /* (11, 22, 17) {real, imag} */,
  {32'hc1319682, 32'h4036da8c} /* (11, 22, 16) {real, imag} */,
  {32'h418e6d35, 32'hc18a5b19} /* (11, 22, 15) {real, imag} */,
  {32'h3e067e88, 32'h41848862} /* (11, 22, 14) {real, imag} */,
  {32'hc079ffba, 32'h40ca1133} /* (11, 22, 13) {real, imag} */,
  {32'hc02925b3, 32'hc10c407c} /* (11, 22, 12) {real, imag} */,
  {32'h409afe57, 32'hc03590ef} /* (11, 22, 11) {real, imag} */,
  {32'hc0552da9, 32'hc09b4a54} /* (11, 22, 10) {real, imag} */,
  {32'h407cda40, 32'hc15a0be4} /* (11, 22, 9) {real, imag} */,
  {32'hc095afdb, 32'h401b9178} /* (11, 22, 8) {real, imag} */,
  {32'hc0efc91f, 32'hc070e1aa} /* (11, 22, 7) {real, imag} */,
  {32'h40205897, 32'h40d150f6} /* (11, 22, 6) {real, imag} */,
  {32'hc1dc28b8, 32'h3fe52cf4} /* (11, 22, 5) {real, imag} */,
  {32'h419455c2, 32'h412f83a5} /* (11, 22, 4) {real, imag} */,
  {32'hc055a50f, 32'h412a051c} /* (11, 22, 3) {real, imag} */,
  {32'hc09f7792, 32'hbe9538c0} /* (11, 22, 2) {real, imag} */,
  {32'h3f6b9808, 32'hc1d21d4a} /* (11, 22, 1) {real, imag} */,
  {32'h41065a20, 32'h419f1d5c} /* (11, 22, 0) {real, imag} */,
  {32'hc012ec86, 32'h419039a0} /* (11, 21, 31) {real, imag} */,
  {32'hc138ee30, 32'hc21b35fa} /* (11, 21, 30) {real, imag} */,
  {32'hc0eb313e, 32'hc1b307cc} /* (11, 21, 29) {real, imag} */,
  {32'h41a3fbab, 32'h413d531d} /* (11, 21, 28) {real, imag} */,
  {32'h4094d8cc, 32'hc1945781} /* (11, 21, 27) {real, imag} */,
  {32'h41125f86, 32'h40e97029} /* (11, 21, 26) {real, imag} */,
  {32'hc165c47d, 32'hc1a89a4a} /* (11, 21, 25) {real, imag} */,
  {32'h412075c7, 32'hc054866c} /* (11, 21, 24) {real, imag} */,
  {32'h41d0c1f3, 32'h41284b4a} /* (11, 21, 23) {real, imag} */,
  {32'h3fd228dc, 32'h40ac909c} /* (11, 21, 22) {real, imag} */,
  {32'hc11e15db, 32'h400b6dbb} /* (11, 21, 21) {real, imag} */,
  {32'h401523e6, 32'h405734d8} /* (11, 21, 20) {real, imag} */,
  {32'hc0d389a6, 32'hc11e0c86} /* (11, 21, 19) {real, imag} */,
  {32'h402b0bda, 32'h40a80de6} /* (11, 21, 18) {real, imag} */,
  {32'hc0250bf2, 32'h40dc7f05} /* (11, 21, 17) {real, imag} */,
  {32'h4066e886, 32'hc12bbf1b} /* (11, 21, 16) {real, imag} */,
  {32'h404b7bc2, 32'h3f0a608c} /* (11, 21, 15) {real, imag} */,
  {32'hc09deea0, 32'hc167038a} /* (11, 21, 14) {real, imag} */,
  {32'hc13f1045, 32'hc1377c16} /* (11, 21, 13) {real, imag} */,
  {32'h413a9203, 32'hc07ffb18} /* (11, 21, 12) {real, imag} */,
  {32'h413ffb10, 32'hc04ce78f} /* (11, 21, 11) {real, imag} */,
  {32'hbf5e28d8, 32'h411b4528} /* (11, 21, 10) {real, imag} */,
  {32'hc175e3d4, 32'h41582d8b} /* (11, 21, 9) {real, imag} */,
  {32'h4133a3a4, 32'h40f12c23} /* (11, 21, 8) {real, imag} */,
  {32'h40832bbc, 32'hc18be722} /* (11, 21, 7) {real, imag} */,
  {32'hc15c2d73, 32'h4118c248} /* (11, 21, 6) {real, imag} */,
  {32'hbfc66ff4, 32'hc0be0c47} /* (11, 21, 5) {real, imag} */,
  {32'hc11de1f4, 32'hc14fe524} /* (11, 21, 4) {real, imag} */,
  {32'h4087ed19, 32'h40cf819d} /* (11, 21, 3) {real, imag} */,
  {32'h41f9d3a5, 32'h3f94ec22} /* (11, 21, 2) {real, imag} */,
  {32'hc03380c4, 32'h417b3e32} /* (11, 21, 1) {real, imag} */,
  {32'hc135545f, 32'h41a16ea7} /* (11, 21, 0) {real, imag} */,
  {32'hc063695b, 32'h4095891c} /* (11, 20, 31) {real, imag} */,
  {32'h4172e050, 32'hc18d7f35} /* (11, 20, 30) {real, imag} */,
  {32'h40a2d303, 32'hc093375d} /* (11, 20, 29) {real, imag} */,
  {32'h40f38eff, 32'h412772a9} /* (11, 20, 28) {real, imag} */,
  {32'hc08ffabb, 32'h416285c3} /* (11, 20, 27) {real, imag} */,
  {32'h40c1ffaf, 32'h411ab223} /* (11, 20, 26) {real, imag} */,
  {32'hbfeb6770, 32'h41cc102a} /* (11, 20, 25) {real, imag} */,
  {32'h40ef5be3, 32'hc11d7268} /* (11, 20, 24) {real, imag} */,
  {32'hc1a121f3, 32'h414a41b9} /* (11, 20, 23) {real, imag} */,
  {32'h40c52cd5, 32'h40d5974e} /* (11, 20, 22) {real, imag} */,
  {32'h3ed03760, 32'hc109f1bb} /* (11, 20, 21) {real, imag} */,
  {32'h40320812, 32'hc13841ec} /* (11, 20, 20) {real, imag} */,
  {32'hc0f66565, 32'hbfd37c0e} /* (11, 20, 19) {real, imag} */,
  {32'hc1078bea, 32'hbf83e6e8} /* (11, 20, 18) {real, imag} */,
  {32'h401e775d, 32'hbfa3f000} /* (11, 20, 17) {real, imag} */,
  {32'hbf4c20e0, 32'h41524812} /* (11, 20, 16) {real, imag} */,
  {32'hc087b7b6, 32'h3e01d900} /* (11, 20, 15) {real, imag} */,
  {32'hc1372d10, 32'h40d65268} /* (11, 20, 14) {real, imag} */,
  {32'h3f6afb29, 32'hc01bc556} /* (11, 20, 13) {real, imag} */,
  {32'hc06aa10f, 32'hc13fd042} /* (11, 20, 12) {real, imag} */,
  {32'hc1c4d284, 32'hc024c847} /* (11, 20, 11) {real, imag} */,
  {32'h412c6647, 32'h3e553848} /* (11, 20, 10) {real, imag} */,
  {32'hc106c1d8, 32'hc140a258} /* (11, 20, 9) {real, imag} */,
  {32'h41158ee5, 32'h3eb28be0} /* (11, 20, 8) {real, imag} */,
  {32'h40e5d586, 32'hc0bae68b} /* (11, 20, 7) {real, imag} */,
  {32'h40a57376, 32'hc18fdb31} /* (11, 20, 6) {real, imag} */,
  {32'hbeb53f78, 32'h4162c80d} /* (11, 20, 5) {real, imag} */,
  {32'hc0c39c81, 32'h40de2a18} /* (11, 20, 4) {real, imag} */,
  {32'hc0fdf11e, 32'hc1646e74} /* (11, 20, 3) {real, imag} */,
  {32'hc164309e, 32'h40be6c70} /* (11, 20, 2) {real, imag} */,
  {32'h40c672de, 32'hc184bc29} /* (11, 20, 1) {real, imag} */,
  {32'hc0e1425c, 32'hbed0e4b0} /* (11, 20, 0) {real, imag} */,
  {32'h3f95c668, 32'hc0111c0a} /* (11, 19, 31) {real, imag} */,
  {32'hc091c23a, 32'hc09daca4} /* (11, 19, 30) {real, imag} */,
  {32'hc0a4eb29, 32'h4081f15a} /* (11, 19, 29) {real, imag} */,
  {32'hbfd0df80, 32'hc12c2f2f} /* (11, 19, 28) {real, imag} */,
  {32'hc0c373d7, 32'h40dfb4b8} /* (11, 19, 27) {real, imag} */,
  {32'hc01a6f36, 32'h402ae0e8} /* (11, 19, 26) {real, imag} */,
  {32'h3f96e688, 32'hc085a003} /* (11, 19, 25) {real, imag} */,
  {32'hc0e21b77, 32'h404d0250} /* (11, 19, 24) {real, imag} */,
  {32'hc11230ce, 32'h3f8392b0} /* (11, 19, 23) {real, imag} */,
  {32'hc106a2ba, 32'hc0851f84} /* (11, 19, 22) {real, imag} */,
  {32'hc1017d07, 32'h4014afd8} /* (11, 19, 21) {real, imag} */,
  {32'hbe73b080, 32'h4140da66} /* (11, 19, 20) {real, imag} */,
  {32'h405805d4, 32'hc10c3366} /* (11, 19, 19) {real, imag} */,
  {32'h4010f658, 32'hc14be1c0} /* (11, 19, 18) {real, imag} */,
  {32'hbf41dc32, 32'h4152f052} /* (11, 19, 17) {real, imag} */,
  {32'hc13d39f7, 32'hc09a6498} /* (11, 19, 16) {real, imag} */,
  {32'hbf1baa30, 32'hbf5957c0} /* (11, 19, 15) {real, imag} */,
  {32'hc0b0363a, 32'h40861102} /* (11, 19, 14) {real, imag} */,
  {32'hbfee6358, 32'hc15b616f} /* (11, 19, 13) {real, imag} */,
  {32'hc17622fd, 32'h41d73804} /* (11, 19, 12) {real, imag} */,
  {32'h400ac154, 32'hc11d95f8} /* (11, 19, 11) {real, imag} */,
  {32'hc00c0820, 32'h40c362a9} /* (11, 19, 10) {real, imag} */,
  {32'h41ab6688, 32'hc0989d22} /* (11, 19, 9) {real, imag} */,
  {32'hbfcb059a, 32'h4156c84e} /* (11, 19, 8) {real, imag} */,
  {32'h40694022, 32'h41900edf} /* (11, 19, 7) {real, imag} */,
  {32'hc16889f8, 32'h40e36d4f} /* (11, 19, 6) {real, imag} */,
  {32'h40401413, 32'hbfd90f24} /* (11, 19, 5) {real, imag} */,
  {32'h4176718e, 32'hc12b1a06} /* (11, 19, 4) {real, imag} */,
  {32'h411e3c0c, 32'hbf9fc780} /* (11, 19, 3) {real, imag} */,
  {32'hc0542f68, 32'hc05facf6} /* (11, 19, 2) {real, imag} */,
  {32'hc0112bbe, 32'h4196aa90} /* (11, 19, 1) {real, imag} */,
  {32'h40a88106, 32'hc1142a72} /* (11, 19, 0) {real, imag} */,
  {32'h4015ef78, 32'h41b6066c} /* (11, 18, 31) {real, imag} */,
  {32'h41546afe, 32'hbfb5a16e} /* (11, 18, 30) {real, imag} */,
  {32'hc0cee6a6, 32'h410d9c2b} /* (11, 18, 29) {real, imag} */,
  {32'hc1421abb, 32'h40895554} /* (11, 18, 28) {real, imag} */,
  {32'h407a3fae, 32'hc0a02af8} /* (11, 18, 27) {real, imag} */,
  {32'hc0d78ec7, 32'hc061b9ea} /* (11, 18, 26) {real, imag} */,
  {32'hc0df56e1, 32'h402a17d7} /* (11, 18, 25) {real, imag} */,
  {32'h408f5067, 32'hc1111576} /* (11, 18, 24) {real, imag} */,
  {32'hc0409792, 32'hc0e391d0} /* (11, 18, 23) {real, imag} */,
  {32'h41a18260, 32'hc1e2ded8} /* (11, 18, 22) {real, imag} */,
  {32'hc0aa871c, 32'hc0d3b42c} /* (11, 18, 21) {real, imag} */,
  {32'hc1a0be93, 32'hbfbf45f0} /* (11, 18, 20) {real, imag} */,
  {32'h3f4554ba, 32'h3fcd2a28} /* (11, 18, 19) {real, imag} */,
  {32'h3fa56a10, 32'hbeafee50} /* (11, 18, 18) {real, imag} */,
  {32'hc08de419, 32'hc138bd86} /* (11, 18, 17) {real, imag} */,
  {32'hc1280a04, 32'hc03780e8} /* (11, 18, 16) {real, imag} */,
  {32'h41014dcc, 32'hc131108e} /* (11, 18, 15) {real, imag} */,
  {32'hc0ca3592, 32'h411d602a} /* (11, 18, 14) {real, imag} */,
  {32'h3f96892c, 32'h4145f1f9} /* (11, 18, 13) {real, imag} */,
  {32'hc101937c, 32'h40e00c7e} /* (11, 18, 12) {real, imag} */,
  {32'h41272d1c, 32'hc0ad5542} /* (11, 18, 11) {real, imag} */,
  {32'h3ffb0e5c, 32'hc0f06a8c} /* (11, 18, 10) {real, imag} */,
  {32'hbec01cf8, 32'h3ff466c6} /* (11, 18, 9) {real, imag} */,
  {32'hbeb8d630, 32'hbedc4af0} /* (11, 18, 8) {real, imag} */,
  {32'h4013bd2e, 32'h403662ba} /* (11, 18, 7) {real, imag} */,
  {32'hc0788ba6, 32'h4006c544} /* (11, 18, 6) {real, imag} */,
  {32'h3f85a945, 32'h416edaa0} /* (11, 18, 5) {real, imag} */,
  {32'hc13e4a8b, 32'hc152f601} /* (11, 18, 4) {real, imag} */,
  {32'hc109f2de, 32'hc1061db8} /* (11, 18, 3) {real, imag} */,
  {32'hc10451c0, 32'hc15e4891} /* (11, 18, 2) {real, imag} */,
  {32'hc123e667, 32'h410f57ad} /* (11, 18, 1) {real, imag} */,
  {32'hbee31000, 32'h4126cb40} /* (11, 18, 0) {real, imag} */,
  {32'hc0e7d8ea, 32'hc06f4b10} /* (11, 17, 31) {real, imag} */,
  {32'h411cb621, 32'h40dbb5ce} /* (11, 17, 30) {real, imag} */,
  {32'h4123adf0, 32'hbf42ec2c} /* (11, 17, 29) {real, imag} */,
  {32'hc19a87e6, 32'h40ee0ab2} /* (11, 17, 28) {real, imag} */,
  {32'hbfa7d0a8, 32'hc0baedf7} /* (11, 17, 27) {real, imag} */,
  {32'hbfbf304e, 32'hc01b66c2} /* (11, 17, 26) {real, imag} */,
  {32'h3f8fa0da, 32'h410dbeef} /* (11, 17, 25) {real, imag} */,
  {32'h415f3b0b, 32'hc0dda07c} /* (11, 17, 24) {real, imag} */,
  {32'hbf546b20, 32'hc1036108} /* (11, 17, 23) {real, imag} */,
  {32'hc11c8eea, 32'h3e17c360} /* (11, 17, 22) {real, imag} */,
  {32'hc1966a3b, 32'h40df9263} /* (11, 17, 21) {real, imag} */,
  {32'h40c47840, 32'h40f2808d} /* (11, 17, 20) {real, imag} */,
  {32'h40eac7d1, 32'hbf7d0278} /* (11, 17, 19) {real, imag} */,
  {32'h40ca2a56, 32'h4149b688} /* (11, 17, 18) {real, imag} */,
  {32'h404467b8, 32'hbfd70918} /* (11, 17, 17) {real, imag} */,
  {32'hc13ac271, 32'hc0ced706} /* (11, 17, 16) {real, imag} */,
  {32'h3f2c8b08, 32'hc091a62c} /* (11, 17, 15) {real, imag} */,
  {32'hc01648c8, 32'h3f0cf8c0} /* (11, 17, 14) {real, imag} */,
  {32'hc15019c3, 32'h4094c8d8} /* (11, 17, 13) {real, imag} */,
  {32'hc0b33a3e, 32'h41a6a527} /* (11, 17, 12) {real, imag} */,
  {32'hc08bbcbe, 32'h40ee97b9} /* (11, 17, 11) {real, imag} */,
  {32'hc173654e, 32'h40dc453b} /* (11, 17, 10) {real, imag} */,
  {32'hc0088dfb, 32'h3c18c400} /* (11, 17, 9) {real, imag} */,
  {32'hc01f7f29, 32'hc0fff7a0} /* (11, 17, 8) {real, imag} */,
  {32'hc15eb238, 32'hc036dd46} /* (11, 17, 7) {real, imag} */,
  {32'h41955488, 32'hc02694d9} /* (11, 17, 6) {real, imag} */,
  {32'hc0f909a4, 32'hc119c4c0} /* (11, 17, 5) {real, imag} */,
  {32'h413d2a3e, 32'hc0e8a866} /* (11, 17, 4) {real, imag} */,
  {32'h3f0f490c, 32'h402f6a65} /* (11, 17, 3) {real, imag} */,
  {32'h409e65d0, 32'hc00f4217} /* (11, 17, 2) {real, imag} */,
  {32'hc08aa525, 32'hc0d4fd9a} /* (11, 17, 1) {real, imag} */,
  {32'h4084a3d0, 32'hc0b8b3b6} /* (11, 17, 0) {real, imag} */,
  {32'hbf96f33c, 32'h406e0960} /* (11, 16, 31) {real, imag} */,
  {32'hc0b52dba, 32'h3d29de80} /* (11, 16, 30) {real, imag} */,
  {32'h40354424, 32'h4137a8d0} /* (11, 16, 29) {real, imag} */,
  {32'h3fff32f0, 32'h40b5080f} /* (11, 16, 28) {real, imag} */,
  {32'h40aace02, 32'hc0e83f19} /* (11, 16, 27) {real, imag} */,
  {32'h3dd5c140, 32'h3f80010a} /* (11, 16, 26) {real, imag} */,
  {32'h3f124c06, 32'hc084cfde} /* (11, 16, 25) {real, imag} */,
  {32'h4013e9a8, 32'hc0658e27} /* (11, 16, 24) {real, imag} */,
  {32'hc08e808d, 32'hc04d5fe9} /* (11, 16, 23) {real, imag} */,
  {32'h403594ee, 32'h3f668f1b} /* (11, 16, 22) {real, imag} */,
  {32'hc04bd210, 32'h3e9bdff4} /* (11, 16, 21) {real, imag} */,
  {32'h409a6da4, 32'h4192dd71} /* (11, 16, 20) {real, imag} */,
  {32'hc085af36, 32'h40c1d001} /* (11, 16, 19) {real, imag} */,
  {32'h40b264de, 32'h40b5fd6d} /* (11, 16, 18) {real, imag} */,
  {32'h403b9cae, 32'hc0d34d36} /* (11, 16, 17) {real, imag} */,
  {32'h408e5488, 32'h00000000} /* (11, 16, 16) {real, imag} */,
  {32'h403b9cae, 32'h40d34d36} /* (11, 16, 15) {real, imag} */,
  {32'h40b264de, 32'hc0b5fd6d} /* (11, 16, 14) {real, imag} */,
  {32'hc085af36, 32'hc0c1d001} /* (11, 16, 13) {real, imag} */,
  {32'h409a6da4, 32'hc192dd71} /* (11, 16, 12) {real, imag} */,
  {32'hc04bd210, 32'hbe9bdff4} /* (11, 16, 11) {real, imag} */,
  {32'h403594ee, 32'hbf668f1b} /* (11, 16, 10) {real, imag} */,
  {32'hc08e808d, 32'h404d5fe9} /* (11, 16, 9) {real, imag} */,
  {32'h4013e9a8, 32'h40658e27} /* (11, 16, 8) {real, imag} */,
  {32'h3f124c06, 32'h4084cfde} /* (11, 16, 7) {real, imag} */,
  {32'h3dd5c140, 32'hbf80010a} /* (11, 16, 6) {real, imag} */,
  {32'h40aace02, 32'h40e83f19} /* (11, 16, 5) {real, imag} */,
  {32'h3fff32f0, 32'hc0b5080f} /* (11, 16, 4) {real, imag} */,
  {32'h40354424, 32'hc137a8d0} /* (11, 16, 3) {real, imag} */,
  {32'hc0b52dba, 32'hbd29de80} /* (11, 16, 2) {real, imag} */,
  {32'hbf96f33c, 32'hc06e0960} /* (11, 16, 1) {real, imag} */,
  {32'hc06d7256, 32'h00000000} /* (11, 16, 0) {real, imag} */,
  {32'hc08aa525, 32'h40d4fd9a} /* (11, 15, 31) {real, imag} */,
  {32'h409e65d0, 32'h400f4217} /* (11, 15, 30) {real, imag} */,
  {32'h3f0f490c, 32'hc02f6a65} /* (11, 15, 29) {real, imag} */,
  {32'h413d2a3e, 32'h40e8a866} /* (11, 15, 28) {real, imag} */,
  {32'hc0f909a4, 32'h4119c4c0} /* (11, 15, 27) {real, imag} */,
  {32'h41955488, 32'h402694d9} /* (11, 15, 26) {real, imag} */,
  {32'hc15eb238, 32'h4036dd46} /* (11, 15, 25) {real, imag} */,
  {32'hc01f7f29, 32'h40fff7a0} /* (11, 15, 24) {real, imag} */,
  {32'hc0088dfb, 32'hbc18c400} /* (11, 15, 23) {real, imag} */,
  {32'hc173654e, 32'hc0dc453b} /* (11, 15, 22) {real, imag} */,
  {32'hc08bbcbe, 32'hc0ee97b9} /* (11, 15, 21) {real, imag} */,
  {32'hc0b33a3e, 32'hc1a6a527} /* (11, 15, 20) {real, imag} */,
  {32'hc15019c3, 32'hc094c8d8} /* (11, 15, 19) {real, imag} */,
  {32'hc01648c8, 32'hbf0cf8c0} /* (11, 15, 18) {real, imag} */,
  {32'h3f2c8b08, 32'h4091a62c} /* (11, 15, 17) {real, imag} */,
  {32'hc13ac271, 32'h40ced706} /* (11, 15, 16) {real, imag} */,
  {32'h404467b8, 32'h3fd70918} /* (11, 15, 15) {real, imag} */,
  {32'h40ca2a56, 32'hc149b688} /* (11, 15, 14) {real, imag} */,
  {32'h40eac7d1, 32'h3f7d0278} /* (11, 15, 13) {real, imag} */,
  {32'h40c47840, 32'hc0f2808d} /* (11, 15, 12) {real, imag} */,
  {32'hc1966a3b, 32'hc0df9263} /* (11, 15, 11) {real, imag} */,
  {32'hc11c8eea, 32'hbe17c360} /* (11, 15, 10) {real, imag} */,
  {32'hbf546b20, 32'h41036108} /* (11, 15, 9) {real, imag} */,
  {32'h415f3b0b, 32'h40dda07c} /* (11, 15, 8) {real, imag} */,
  {32'h3f8fa0da, 32'hc10dbeef} /* (11, 15, 7) {real, imag} */,
  {32'hbfbf304e, 32'h401b66c2} /* (11, 15, 6) {real, imag} */,
  {32'hbfa7d0a8, 32'h40baedf7} /* (11, 15, 5) {real, imag} */,
  {32'hc19a87e6, 32'hc0ee0ab2} /* (11, 15, 4) {real, imag} */,
  {32'h4123adf0, 32'h3f42ec2c} /* (11, 15, 3) {real, imag} */,
  {32'h411cb621, 32'hc0dbb5ce} /* (11, 15, 2) {real, imag} */,
  {32'hc0e7d8ea, 32'h406f4b10} /* (11, 15, 1) {real, imag} */,
  {32'h4084a3d0, 32'h40b8b3b6} /* (11, 15, 0) {real, imag} */,
  {32'hc123e667, 32'hc10f57ad} /* (11, 14, 31) {real, imag} */,
  {32'hc10451c0, 32'h415e4891} /* (11, 14, 30) {real, imag} */,
  {32'hc109f2de, 32'h41061db8} /* (11, 14, 29) {real, imag} */,
  {32'hc13e4a8b, 32'h4152f601} /* (11, 14, 28) {real, imag} */,
  {32'h3f85a945, 32'hc16edaa0} /* (11, 14, 27) {real, imag} */,
  {32'hc0788ba6, 32'hc006c544} /* (11, 14, 26) {real, imag} */,
  {32'h4013bd2e, 32'hc03662ba} /* (11, 14, 25) {real, imag} */,
  {32'hbeb8d630, 32'h3edc4af0} /* (11, 14, 24) {real, imag} */,
  {32'hbec01cf8, 32'hbff466c6} /* (11, 14, 23) {real, imag} */,
  {32'h3ffb0e5c, 32'h40f06a8c} /* (11, 14, 22) {real, imag} */,
  {32'h41272d1c, 32'h40ad5542} /* (11, 14, 21) {real, imag} */,
  {32'hc101937c, 32'hc0e00c7e} /* (11, 14, 20) {real, imag} */,
  {32'h3f96892c, 32'hc145f1f9} /* (11, 14, 19) {real, imag} */,
  {32'hc0ca3592, 32'hc11d602a} /* (11, 14, 18) {real, imag} */,
  {32'h41014dcc, 32'h4131108e} /* (11, 14, 17) {real, imag} */,
  {32'hc1280a04, 32'h403780e8} /* (11, 14, 16) {real, imag} */,
  {32'hc08de419, 32'h4138bd86} /* (11, 14, 15) {real, imag} */,
  {32'h3fa56a10, 32'h3eafee50} /* (11, 14, 14) {real, imag} */,
  {32'h3f4554ba, 32'hbfcd2a28} /* (11, 14, 13) {real, imag} */,
  {32'hc1a0be93, 32'h3fbf45f0} /* (11, 14, 12) {real, imag} */,
  {32'hc0aa871c, 32'h40d3b42c} /* (11, 14, 11) {real, imag} */,
  {32'h41a18260, 32'h41e2ded8} /* (11, 14, 10) {real, imag} */,
  {32'hc0409792, 32'h40e391d0} /* (11, 14, 9) {real, imag} */,
  {32'h408f5067, 32'h41111576} /* (11, 14, 8) {real, imag} */,
  {32'hc0df56e1, 32'hc02a17d7} /* (11, 14, 7) {real, imag} */,
  {32'hc0d78ec7, 32'h4061b9ea} /* (11, 14, 6) {real, imag} */,
  {32'h407a3fae, 32'h40a02af8} /* (11, 14, 5) {real, imag} */,
  {32'hc1421abb, 32'hc0895554} /* (11, 14, 4) {real, imag} */,
  {32'hc0cee6a6, 32'hc10d9c2b} /* (11, 14, 3) {real, imag} */,
  {32'h41546afe, 32'h3fb5a16e} /* (11, 14, 2) {real, imag} */,
  {32'h4015ef78, 32'hc1b6066c} /* (11, 14, 1) {real, imag} */,
  {32'hbee31000, 32'hc126cb40} /* (11, 14, 0) {real, imag} */,
  {32'hc0112bbe, 32'hc196aa90} /* (11, 13, 31) {real, imag} */,
  {32'hc0542f68, 32'h405facf6} /* (11, 13, 30) {real, imag} */,
  {32'h411e3c0c, 32'h3f9fc780} /* (11, 13, 29) {real, imag} */,
  {32'h4176718e, 32'h412b1a06} /* (11, 13, 28) {real, imag} */,
  {32'h40401413, 32'h3fd90f24} /* (11, 13, 27) {real, imag} */,
  {32'hc16889f8, 32'hc0e36d4f} /* (11, 13, 26) {real, imag} */,
  {32'h40694022, 32'hc1900edf} /* (11, 13, 25) {real, imag} */,
  {32'hbfcb059a, 32'hc156c84e} /* (11, 13, 24) {real, imag} */,
  {32'h41ab6688, 32'h40989d22} /* (11, 13, 23) {real, imag} */,
  {32'hc00c0820, 32'hc0c362a9} /* (11, 13, 22) {real, imag} */,
  {32'h400ac154, 32'h411d95f8} /* (11, 13, 21) {real, imag} */,
  {32'hc17622fd, 32'hc1d73804} /* (11, 13, 20) {real, imag} */,
  {32'hbfee6358, 32'h415b616f} /* (11, 13, 19) {real, imag} */,
  {32'hc0b0363a, 32'hc0861102} /* (11, 13, 18) {real, imag} */,
  {32'hbf1baa30, 32'h3f5957c0} /* (11, 13, 17) {real, imag} */,
  {32'hc13d39f7, 32'h409a6498} /* (11, 13, 16) {real, imag} */,
  {32'hbf41dc32, 32'hc152f052} /* (11, 13, 15) {real, imag} */,
  {32'h4010f658, 32'h414be1c0} /* (11, 13, 14) {real, imag} */,
  {32'h405805d4, 32'h410c3366} /* (11, 13, 13) {real, imag} */,
  {32'hbe73b080, 32'hc140da66} /* (11, 13, 12) {real, imag} */,
  {32'hc1017d07, 32'hc014afd8} /* (11, 13, 11) {real, imag} */,
  {32'hc106a2ba, 32'h40851f84} /* (11, 13, 10) {real, imag} */,
  {32'hc11230ce, 32'hbf8392b0} /* (11, 13, 9) {real, imag} */,
  {32'hc0e21b77, 32'hc04d0250} /* (11, 13, 8) {real, imag} */,
  {32'h3f96e688, 32'h4085a003} /* (11, 13, 7) {real, imag} */,
  {32'hc01a6f36, 32'hc02ae0e8} /* (11, 13, 6) {real, imag} */,
  {32'hc0c373d7, 32'hc0dfb4b8} /* (11, 13, 5) {real, imag} */,
  {32'hbfd0df80, 32'h412c2f2f} /* (11, 13, 4) {real, imag} */,
  {32'hc0a4eb29, 32'hc081f15a} /* (11, 13, 3) {real, imag} */,
  {32'hc091c23a, 32'h409daca4} /* (11, 13, 2) {real, imag} */,
  {32'h3f95c668, 32'h40111c0a} /* (11, 13, 1) {real, imag} */,
  {32'h40a88106, 32'h41142a72} /* (11, 13, 0) {real, imag} */,
  {32'h40c672de, 32'h4184bc29} /* (11, 12, 31) {real, imag} */,
  {32'hc164309e, 32'hc0be6c70} /* (11, 12, 30) {real, imag} */,
  {32'hc0fdf11e, 32'h41646e74} /* (11, 12, 29) {real, imag} */,
  {32'hc0c39c81, 32'hc0de2a18} /* (11, 12, 28) {real, imag} */,
  {32'hbeb53f78, 32'hc162c80d} /* (11, 12, 27) {real, imag} */,
  {32'h40a57376, 32'h418fdb31} /* (11, 12, 26) {real, imag} */,
  {32'h40e5d586, 32'h40bae68b} /* (11, 12, 25) {real, imag} */,
  {32'h41158ee5, 32'hbeb28be0} /* (11, 12, 24) {real, imag} */,
  {32'hc106c1d8, 32'h4140a258} /* (11, 12, 23) {real, imag} */,
  {32'h412c6647, 32'hbe553848} /* (11, 12, 22) {real, imag} */,
  {32'hc1c4d284, 32'h4024c847} /* (11, 12, 21) {real, imag} */,
  {32'hc06aa10f, 32'h413fd042} /* (11, 12, 20) {real, imag} */,
  {32'h3f6afb29, 32'h401bc556} /* (11, 12, 19) {real, imag} */,
  {32'hc1372d10, 32'hc0d65268} /* (11, 12, 18) {real, imag} */,
  {32'hc087b7b6, 32'hbe01d900} /* (11, 12, 17) {real, imag} */,
  {32'hbf4c20e0, 32'hc1524812} /* (11, 12, 16) {real, imag} */,
  {32'h401e775d, 32'h3fa3f000} /* (11, 12, 15) {real, imag} */,
  {32'hc1078bea, 32'h3f83e6e8} /* (11, 12, 14) {real, imag} */,
  {32'hc0f66565, 32'h3fd37c0e} /* (11, 12, 13) {real, imag} */,
  {32'h40320812, 32'h413841ec} /* (11, 12, 12) {real, imag} */,
  {32'h3ed03760, 32'h4109f1bb} /* (11, 12, 11) {real, imag} */,
  {32'h40c52cd5, 32'hc0d5974e} /* (11, 12, 10) {real, imag} */,
  {32'hc1a121f3, 32'hc14a41b9} /* (11, 12, 9) {real, imag} */,
  {32'h40ef5be3, 32'h411d7268} /* (11, 12, 8) {real, imag} */,
  {32'hbfeb6770, 32'hc1cc102a} /* (11, 12, 7) {real, imag} */,
  {32'h40c1ffaf, 32'hc11ab223} /* (11, 12, 6) {real, imag} */,
  {32'hc08ffabb, 32'hc16285c3} /* (11, 12, 5) {real, imag} */,
  {32'h40f38eff, 32'hc12772a9} /* (11, 12, 4) {real, imag} */,
  {32'h40a2d303, 32'h4093375d} /* (11, 12, 3) {real, imag} */,
  {32'h4172e050, 32'h418d7f35} /* (11, 12, 2) {real, imag} */,
  {32'hc063695b, 32'hc095891c} /* (11, 12, 1) {real, imag} */,
  {32'hc0e1425c, 32'h3ed0e4b0} /* (11, 12, 0) {real, imag} */,
  {32'hc03380c4, 32'hc17b3e32} /* (11, 11, 31) {real, imag} */,
  {32'h41f9d3a5, 32'hbf94ec22} /* (11, 11, 30) {real, imag} */,
  {32'h4087ed19, 32'hc0cf819d} /* (11, 11, 29) {real, imag} */,
  {32'hc11de1f4, 32'h414fe524} /* (11, 11, 28) {real, imag} */,
  {32'hbfc66ff4, 32'h40be0c47} /* (11, 11, 27) {real, imag} */,
  {32'hc15c2d73, 32'hc118c248} /* (11, 11, 26) {real, imag} */,
  {32'h40832bbc, 32'h418be722} /* (11, 11, 25) {real, imag} */,
  {32'h4133a3a4, 32'hc0f12c23} /* (11, 11, 24) {real, imag} */,
  {32'hc175e3d4, 32'hc1582d8b} /* (11, 11, 23) {real, imag} */,
  {32'hbf5e28d8, 32'hc11b4528} /* (11, 11, 22) {real, imag} */,
  {32'h413ffb10, 32'h404ce78f} /* (11, 11, 21) {real, imag} */,
  {32'h413a9203, 32'h407ffb18} /* (11, 11, 20) {real, imag} */,
  {32'hc13f1045, 32'h41377c16} /* (11, 11, 19) {real, imag} */,
  {32'hc09deea0, 32'h4167038a} /* (11, 11, 18) {real, imag} */,
  {32'h404b7bc2, 32'hbf0a608c} /* (11, 11, 17) {real, imag} */,
  {32'h4066e886, 32'h412bbf1b} /* (11, 11, 16) {real, imag} */,
  {32'hc0250bf2, 32'hc0dc7f05} /* (11, 11, 15) {real, imag} */,
  {32'h402b0bda, 32'hc0a80de6} /* (11, 11, 14) {real, imag} */,
  {32'hc0d389a6, 32'h411e0c86} /* (11, 11, 13) {real, imag} */,
  {32'h401523e6, 32'hc05734d8} /* (11, 11, 12) {real, imag} */,
  {32'hc11e15db, 32'hc00b6dbb} /* (11, 11, 11) {real, imag} */,
  {32'h3fd228dc, 32'hc0ac909c} /* (11, 11, 10) {real, imag} */,
  {32'h41d0c1f3, 32'hc1284b4a} /* (11, 11, 9) {real, imag} */,
  {32'h412075c7, 32'h4054866c} /* (11, 11, 8) {real, imag} */,
  {32'hc165c47d, 32'h41a89a4a} /* (11, 11, 7) {real, imag} */,
  {32'h41125f86, 32'hc0e97029} /* (11, 11, 6) {real, imag} */,
  {32'h4094d8cc, 32'h41945781} /* (11, 11, 5) {real, imag} */,
  {32'h41a3fbab, 32'hc13d531d} /* (11, 11, 4) {real, imag} */,
  {32'hc0eb313e, 32'h41b307cc} /* (11, 11, 3) {real, imag} */,
  {32'hc138ee30, 32'h421b35fa} /* (11, 11, 2) {real, imag} */,
  {32'hc012ec86, 32'hc19039a0} /* (11, 11, 1) {real, imag} */,
  {32'hc135545f, 32'hc1a16ea7} /* (11, 11, 0) {real, imag} */,
  {32'h3f6b9808, 32'h41d21d4a} /* (11, 10, 31) {real, imag} */,
  {32'hc09f7792, 32'h3e9538c0} /* (11, 10, 30) {real, imag} */,
  {32'hc055a50f, 32'hc12a051c} /* (11, 10, 29) {real, imag} */,
  {32'h419455c2, 32'hc12f83a5} /* (11, 10, 28) {real, imag} */,
  {32'hc1dc28b8, 32'hbfe52cf4} /* (11, 10, 27) {real, imag} */,
  {32'h40205897, 32'hc0d150f6} /* (11, 10, 26) {real, imag} */,
  {32'hc0efc91f, 32'h4070e1aa} /* (11, 10, 25) {real, imag} */,
  {32'hc095afdb, 32'hc01b9178} /* (11, 10, 24) {real, imag} */,
  {32'h407cda40, 32'h415a0be4} /* (11, 10, 23) {real, imag} */,
  {32'hc0552da9, 32'h409b4a54} /* (11, 10, 22) {real, imag} */,
  {32'h409afe57, 32'h403590ef} /* (11, 10, 21) {real, imag} */,
  {32'hc02925b3, 32'h410c407c} /* (11, 10, 20) {real, imag} */,
  {32'hc079ffba, 32'hc0ca1133} /* (11, 10, 19) {real, imag} */,
  {32'h3e067e88, 32'hc1848862} /* (11, 10, 18) {real, imag} */,
  {32'h418e6d35, 32'h418a5b19} /* (11, 10, 17) {real, imag} */,
  {32'hc1319682, 32'hc036da8c} /* (11, 10, 16) {real, imag} */,
  {32'hc0d3228e, 32'h40da562f} /* (11, 10, 15) {real, imag} */,
  {32'h40abbcd6, 32'hbc303700} /* (11, 10, 14) {real, imag} */,
  {32'h403092fd, 32'h411dc1d2} /* (11, 10, 13) {real, imag} */,
  {32'hbf8e4ae4, 32'hc009aee4} /* (11, 10, 12) {real, imag} */,
  {32'h3f22d1e0, 32'hbeea53ec} /* (11, 10, 11) {real, imag} */,
  {32'hbf86bd9c, 32'hc19387fd} /* (11, 10, 10) {real, imag} */,
  {32'h416af9ec, 32'h41031f08} /* (11, 10, 9) {real, imag} */,
  {32'hbf882b3e, 32'hc0c8ed3e} /* (11, 10, 8) {real, imag} */,
  {32'hc0f268c6, 32'hc018f59f} /* (11, 10, 7) {real, imag} */,
  {32'h40fa3b61, 32'hc1ae1520} /* (11, 10, 6) {real, imag} */,
  {32'h41d3c16c, 32'hc11bd967} /* (11, 10, 5) {real, imag} */,
  {32'h413dd00e, 32'h41ddffd4} /* (11, 10, 4) {real, imag} */,
  {32'h3fa2fa94, 32'h417e02ba} /* (11, 10, 3) {real, imag} */,
  {32'h4118ce9f, 32'hc15f67af} /* (11, 10, 2) {real, imag} */,
  {32'hc0a0c462, 32'h41d37303} /* (11, 10, 1) {real, imag} */,
  {32'h41065a20, 32'hc19f1d5c} /* (11, 10, 0) {real, imag} */,
  {32'hc2184f52, 32'h4184d277} /* (11, 9, 31) {real, imag} */,
  {32'h414d0668, 32'hc19ccfe2} /* (11, 9, 30) {real, imag} */,
  {32'h41101d72, 32'h3f9d8090} /* (11, 9, 29) {real, imag} */,
  {32'hc0895366, 32'hc078bf2c} /* (11, 9, 28) {real, imag} */,
  {32'hc10c7099, 32'h400061ee} /* (11, 9, 27) {real, imag} */,
  {32'h41786a6f, 32'hc15de02e} /* (11, 9, 26) {real, imag} */,
  {32'h3e5e8d80, 32'h413241a2} /* (11, 9, 25) {real, imag} */,
  {32'h40e07521, 32'h417464f5} /* (11, 9, 24) {real, imag} */,
  {32'hc087df60, 32'h4128f6ba} /* (11, 9, 23) {real, imag} */,
  {32'hc0a07753, 32'hc1c4f3b6} /* (11, 9, 22) {real, imag} */,
  {32'hc12ad22d, 32'hc1418e8c} /* (11, 9, 21) {real, imag} */,
  {32'h408282d8, 32'h414bb1ab} /* (11, 9, 20) {real, imag} */,
  {32'h4206eaa8, 32'hc1065e67} /* (11, 9, 19) {real, imag} */,
  {32'hbe097f40, 32'h410dbfaa} /* (11, 9, 18) {real, imag} */,
  {32'hc042613f, 32'h40a56aea} /* (11, 9, 17) {real, imag} */,
  {32'hc089bd6c, 32'hc06ad762} /* (11, 9, 16) {real, imag} */,
  {32'hc04f503f, 32'h3d52cfc0} /* (11, 9, 15) {real, imag} */,
  {32'h3e88e448, 32'h3f8f42a4} /* (11, 9, 14) {real, imag} */,
  {32'hc1bff504, 32'hc115b854} /* (11, 9, 13) {real, imag} */,
  {32'h4134be96, 32'hc1af811e} /* (11, 9, 12) {real, imag} */,
  {32'hc101576e, 32'h3ed522d0} /* (11, 9, 11) {real, imag} */,
  {32'hc128e8e6, 32'h4189faa8} /* (11, 9, 10) {real, imag} */,
  {32'h4010ead4, 32'h41bfa93a} /* (11, 9, 9) {real, imag} */,
  {32'hc13e460c, 32'hc18ec476} /* (11, 9, 8) {real, imag} */,
  {32'hc05dc92d, 32'hc19799ac} /* (11, 9, 7) {real, imag} */,
  {32'h403c9064, 32'h402d84bc} /* (11, 9, 6) {real, imag} */,
  {32'h4040ac38, 32'h3fc02a8c} /* (11, 9, 5) {real, imag} */,
  {32'hc19b5f7a, 32'h3f46ec5c} /* (11, 9, 4) {real, imag} */,
  {32'h41369645, 32'hc14a50e5} /* (11, 9, 3) {real, imag} */,
  {32'hc02c88ba, 32'hc1ca0b98} /* (11, 9, 2) {real, imag} */,
  {32'h40f0aee9, 32'h419c7f16} /* (11, 9, 1) {real, imag} */,
  {32'h3fb538c0, 32'hbff0d664} /* (11, 9, 0) {real, imag} */,
  {32'hc25a8b79, 32'hc1f51222} /* (11, 8, 31) {real, imag} */,
  {32'h42098232, 32'hc0e77cc2} /* (11, 8, 30) {real, imag} */,
  {32'hc209217c, 32'h406abc1e} /* (11, 8, 29) {real, imag} */,
  {32'h41476264, 32'h411808f9} /* (11, 8, 28) {real, imag} */,
  {32'h3f5aabb0, 32'hc11da75e} /* (11, 8, 27) {real, imag} */,
  {32'h3f8d93e8, 32'h42238c64} /* (11, 8, 26) {real, imag} */,
  {32'h41112d4e, 32'hc1bef202} /* (11, 8, 25) {real, imag} */,
  {32'hc17e0448, 32'hc12e5000} /* (11, 8, 24) {real, imag} */,
  {32'h4081bd6e, 32'h3f086570} /* (11, 8, 23) {real, imag} */,
  {32'h41a12279, 32'h402445e2} /* (11, 8, 22) {real, imag} */,
  {32'h40be4f85, 32'hc0b6f008} /* (11, 8, 21) {real, imag} */,
  {32'h4185e238, 32'h4089b4d3} /* (11, 8, 20) {real, imag} */,
  {32'hbf82f46f, 32'hbfd12ee8} /* (11, 8, 19) {real, imag} */,
  {32'h4118ede9, 32'h3f8b25cc} /* (11, 8, 18) {real, imag} */,
  {32'hc0452532, 32'h40b95ec6} /* (11, 8, 17) {real, imag} */,
  {32'hbedec990, 32'h402e279a} /* (11, 8, 16) {real, imag} */,
  {32'hc18f04f8, 32'h4014091a} /* (11, 8, 15) {real, imag} */,
  {32'h4153b056, 32'h413773e8} /* (11, 8, 14) {real, imag} */,
  {32'hc0cdceea, 32'hc0b78920} /* (11, 8, 13) {real, imag} */,
  {32'h413833d1, 32'hc17a3d9e} /* (11, 8, 12) {real, imag} */,
  {32'hc0c4d19c, 32'h4182e78f} /* (11, 8, 11) {real, imag} */,
  {32'h40e3c7f9, 32'h41647665} /* (11, 8, 10) {real, imag} */,
  {32'hc155ce7a, 32'hc1811965} /* (11, 8, 9) {real, imag} */,
  {32'hc15dd500, 32'hc02dc656} /* (11, 8, 8) {real, imag} */,
  {32'hc1a15946, 32'hc11bf3ab} /* (11, 8, 7) {real, imag} */,
  {32'h40ef565e, 32'h415bfcbf} /* (11, 8, 6) {real, imag} */,
  {32'h3ff41750, 32'h412874d9} /* (11, 8, 5) {real, imag} */,
  {32'hc200dcdc, 32'hc0e926af} /* (11, 8, 4) {real, imag} */,
  {32'hc070239e, 32'hc0fc8c1d} /* (11, 8, 3) {real, imag} */,
  {32'h42153914, 32'h41adfb5d} /* (11, 8, 2) {real, imag} */,
  {32'hc204a9f2, 32'hc13331fa} /* (11, 8, 1) {real, imag} */,
  {32'h3fd10ab4, 32'hc19e97e1} /* (11, 8, 0) {real, imag} */,
  {32'h41ad2a66, 32'h411a4ffc} /* (11, 7, 31) {real, imag} */,
  {32'hc10cbe28, 32'h3f9c4440} /* (11, 7, 30) {real, imag} */,
  {32'h416c3f48, 32'h412d2d1a} /* (11, 7, 29) {real, imag} */,
  {32'hc0af5151, 32'h40deb02a} /* (11, 7, 28) {real, imag} */,
  {32'h412651bb, 32'h4121b3fe} /* (11, 7, 27) {real, imag} */,
  {32'hc1212222, 32'hc07766e0} /* (11, 7, 26) {real, imag} */,
  {32'h419e7bb1, 32'hbe5fcf80} /* (11, 7, 25) {real, imag} */,
  {32'hc1fd756e, 32'hc14a1301} /* (11, 7, 24) {real, imag} */,
  {32'hc15f1173, 32'h412355d0} /* (11, 7, 23) {real, imag} */,
  {32'hc0968f50, 32'h41470a82} /* (11, 7, 22) {real, imag} */,
  {32'h411e146e, 32'h4172cda1} /* (11, 7, 21) {real, imag} */,
  {32'h408ee328, 32'h3fa431d7} /* (11, 7, 20) {real, imag} */,
  {32'h419a8ff8, 32'h4203f69d} /* (11, 7, 19) {real, imag} */,
  {32'hc1236167, 32'h3f3ecba8} /* (11, 7, 18) {real, imag} */,
  {32'hc099e815, 32'hc11055f4} /* (11, 7, 17) {real, imag} */,
  {32'hc10c16fe, 32'h414322db} /* (11, 7, 16) {real, imag} */,
  {32'hc0692234, 32'h40499aee} /* (11, 7, 15) {real, imag} */,
  {32'hc0857f89, 32'hbfd06940} /* (11, 7, 14) {real, imag} */,
  {32'hc0b237b0, 32'h411fc0a6} /* (11, 7, 13) {real, imag} */,
  {32'hc0c22bf9, 32'hc07c8c97} /* (11, 7, 12) {real, imag} */,
  {32'h411414b0, 32'hc0714dfa} /* (11, 7, 11) {real, imag} */,
  {32'h41514df9, 32'h40d29eee} /* (11, 7, 10) {real, imag} */,
  {32'hc053c95a, 32'hbfa56820} /* (11, 7, 9) {real, imag} */,
  {32'h41776976, 32'hc0805d6e} /* (11, 7, 8) {real, imag} */,
  {32'h40e46a5a, 32'h4189aafa} /* (11, 7, 7) {real, imag} */,
  {32'h4111be26, 32'hc2033c4d} /* (11, 7, 6) {real, imag} */,
  {32'hc1cb1748, 32'hc0669f6a} /* (11, 7, 5) {real, imag} */,
  {32'h41ae6631, 32'h40b3dd2e} /* (11, 7, 4) {real, imag} */,
  {32'h400b8ac8, 32'hc06e98b8} /* (11, 7, 3) {real, imag} */,
  {32'hc06a312c, 32'h4078a121} /* (11, 7, 2) {real, imag} */,
  {32'hc060d314, 32'h4116a4fc} /* (11, 7, 1) {real, imag} */,
  {32'h411efa4e, 32'h41015e98} /* (11, 7, 0) {real, imag} */,
  {32'h41f382c9, 32'hc2232261} /* (11, 6, 31) {real, imag} */,
  {32'h3f2ec7f0, 32'hc19a41e2} /* (11, 6, 30) {real, imag} */,
  {32'h4091186f, 32'hc152a84f} /* (11, 6, 29) {real, imag} */,
  {32'h41713f90, 32'hc203cec3} /* (11, 6, 28) {real, imag} */,
  {32'h41a71be8, 32'h3f2172e0} /* (11, 6, 27) {real, imag} */,
  {32'h411ccf90, 32'h41cd0c5c} /* (11, 6, 26) {real, imag} */,
  {32'hc0b778a6, 32'hc12446f7} /* (11, 6, 25) {real, imag} */,
  {32'hc02f5070, 32'h419b8af7} /* (11, 6, 24) {real, imag} */,
  {32'h40e4c837, 32'h41a7a0c4} /* (11, 6, 23) {real, imag} */,
  {32'h41772a30, 32'h41222b18} /* (11, 6, 22) {real, imag} */,
  {32'h409dd059, 32'h41202712} /* (11, 6, 21) {real, imag} */,
  {32'h3f9137b0, 32'hc0fd4931} /* (11, 6, 20) {real, imag} */,
  {32'hc0b4c180, 32'h417721e5} /* (11, 6, 19) {real, imag} */,
  {32'hc0a8c3f6, 32'h411c6a6e} /* (11, 6, 18) {real, imag} */,
  {32'h410eadfe, 32'hc153b2f1} /* (11, 6, 17) {real, imag} */,
  {32'h409365f0, 32'h40160636} /* (11, 6, 16) {real, imag} */,
  {32'hbfa420db, 32'h3f845aae} /* (11, 6, 15) {real, imag} */,
  {32'hc0b887f2, 32'h40a08380} /* (11, 6, 14) {real, imag} */,
  {32'h3f5834ba, 32'h40f39882} /* (11, 6, 13) {real, imag} */,
  {32'hbfc4be28, 32'hc13d48fb} /* (11, 6, 12) {real, imag} */,
  {32'h3f928438, 32'hc1977d73} /* (11, 6, 11) {real, imag} */,
  {32'hc03fbdf4, 32'h40ce27d4} /* (11, 6, 10) {real, imag} */,
  {32'hc121182b, 32'hc00bfc3c} /* (11, 6, 9) {real, imag} */,
  {32'hc131b418, 32'hc1a06d98} /* (11, 6, 8) {real, imag} */,
  {32'h40b0c996, 32'h40c38d3f} /* (11, 6, 7) {real, imag} */,
  {32'h41678efc, 32'hc1116e6f} /* (11, 6, 6) {real, imag} */,
  {32'h405e31f8, 32'hc0ff9437} /* (11, 6, 5) {real, imag} */,
  {32'h4057e907, 32'h3f8121ee} /* (11, 6, 4) {real, imag} */,
  {32'h412cf6ce, 32'h413b53ce} /* (11, 6, 3) {real, imag} */,
  {32'h41bd3b27, 32'h402ec9d4} /* (11, 6, 2) {real, imag} */,
  {32'h40c96e12, 32'h407a914c} /* (11, 6, 1) {real, imag} */,
  {32'h4078911e, 32'h4199aa50} /* (11, 6, 0) {real, imag} */,
  {32'hc2dd9576, 32'hc0822142} /* (11, 5, 31) {real, imag} */,
  {32'h41310ea8, 32'hbec55ca0} /* (11, 5, 30) {real, imag} */,
  {32'hc1ac5d22, 32'h40c05c8f} /* (11, 5, 29) {real, imag} */,
  {32'hc17f6a43, 32'h424c7d5a} /* (11, 5, 28) {real, imag} */,
  {32'h413895f0, 32'h419b62d4} /* (11, 5, 27) {real, imag} */,
  {32'h4144eb58, 32'hc119232a} /* (11, 5, 26) {real, imag} */,
  {32'h40a87fe2, 32'hc04d7b0d} /* (11, 5, 25) {real, imag} */,
  {32'h416d21c6, 32'hc2154064} /* (11, 5, 24) {real, imag} */,
  {32'hc026fa62, 32'hc10064bc} /* (11, 5, 23) {real, imag} */,
  {32'h4072929e, 32'h40bd5cf2} /* (11, 5, 22) {real, imag} */,
  {32'hc0bb3320, 32'hc18b8876} /* (11, 5, 21) {real, imag} */,
  {32'h40dd3ebd, 32'h3e1af880} /* (11, 5, 20) {real, imag} */,
  {32'h4193b0f3, 32'h4152a230} /* (11, 5, 19) {real, imag} */,
  {32'hc0ec6be4, 32'h40ae0a89} /* (11, 5, 18) {real, imag} */,
  {32'h3edb8f30, 32'h400f20ed} /* (11, 5, 17) {real, imag} */,
  {32'hc0e6084e, 32'h40532214} /* (11, 5, 16) {real, imag} */,
  {32'h411ad574, 32'hc0c69c88} /* (11, 5, 15) {real, imag} */,
  {32'hc0d68376, 32'h40ddd840} /* (11, 5, 14) {real, imag} */,
  {32'h41193244, 32'h40d5e48a} /* (11, 5, 13) {real, imag} */,
  {32'h41199806, 32'h41a1c47b} /* (11, 5, 12) {real, imag} */,
  {32'h41a7ecc2, 32'hc117f42c} /* (11, 5, 11) {real, imag} */,
  {32'hc16c06de, 32'h413d5356} /* (11, 5, 10) {real, imag} */,
  {32'hc0d808dd, 32'hc0f59015} /* (11, 5, 9) {real, imag} */,
  {32'h41958817, 32'h41b456b8} /* (11, 5, 8) {real, imag} */,
  {32'h40c57cf0, 32'h41266bd1} /* (11, 5, 7) {real, imag} */,
  {32'hc206c45e, 32'hbf643060} /* (11, 5, 6) {real, imag} */,
  {32'h420c3aec, 32'hbd65d000} /* (11, 5, 5) {real, imag} */,
  {32'h40b385ed, 32'hc10fdb2b} /* (11, 5, 4) {real, imag} */,
  {32'hc1e1aeae, 32'hc11ab5d8} /* (11, 5, 3) {real, imag} */,
  {32'h419c603c, 32'h41e2af0e} /* (11, 5, 2) {real, imag} */,
  {32'hc152afba, 32'hc29b86e8} /* (11, 5, 1) {real, imag} */,
  {32'hc26523e2, 32'hc1b3bf32} /* (11, 5, 0) {real, imag} */,
  {32'h41f12752, 32'h42b171a3} /* (11, 4, 31) {real, imag} */,
  {32'hc2eacd1f, 32'hc2aeaad3} /* (11, 4, 30) {real, imag} */,
  {32'hc12a0525, 32'hc156b3d5} /* (11, 4, 29) {real, imag} */,
  {32'h40acb6dd, 32'hbfcc8da0} /* (11, 4, 28) {real, imag} */,
  {32'hc0972a33, 32'h41067687} /* (11, 4, 27) {real, imag} */,
  {32'hc0df84ac, 32'hc0992348} /* (11, 4, 26) {real, imag} */,
  {32'h41992fcc, 32'h410f1535} /* (11, 4, 25) {real, imag} */,
  {32'hbf92162c, 32'hc107a07a} /* (11, 4, 24) {real, imag} */,
  {32'h41947f2e, 32'hc11ab064} /* (11, 4, 23) {real, imag} */,
  {32'hc0f226ea, 32'hc080b536} /* (11, 4, 22) {real, imag} */,
  {32'hc160655e, 32'h4099afab} /* (11, 4, 21) {real, imag} */,
  {32'h419d46bd, 32'h410f87bd} /* (11, 4, 20) {real, imag} */,
  {32'h40bf2560, 32'h40bcba06} /* (11, 4, 19) {real, imag} */,
  {32'hc0d22f46, 32'hc1a19aa7} /* (11, 4, 18) {real, imag} */,
  {32'h40a20678, 32'h409290b5} /* (11, 4, 17) {real, imag} */,
  {32'h3f5e33e4, 32'h4089c9a2} /* (11, 4, 16) {real, imag} */,
  {32'hbfd4d751, 32'hc00c8a8c} /* (11, 4, 15) {real, imag} */,
  {32'h41347fd0, 32'hc154a1c6} /* (11, 4, 14) {real, imag} */,
  {32'hc03d8d3c, 32'h3f85ca08} /* (11, 4, 13) {real, imag} */,
  {32'h40974fb1, 32'h3fb6711f} /* (11, 4, 12) {real, imag} */,
  {32'h40261298, 32'hc08a158f} /* (11, 4, 11) {real, imag} */,
  {32'hc1ac3ae6, 32'hc09685fd} /* (11, 4, 10) {real, imag} */,
  {32'hc0efe966, 32'h41202c9a} /* (11, 4, 9) {real, imag} */,
  {32'hc18470a1, 32'hc19d0aa0} /* (11, 4, 8) {real, imag} */,
  {32'h415d8def, 32'hc146b910} /* (11, 4, 7) {real, imag} */,
  {32'hc161ea33, 32'h41ccde3e} /* (11, 4, 6) {real, imag} */,
  {32'h41944aaa, 32'hc1bd6c61} /* (11, 4, 5) {real, imag} */,
  {32'h408864dc, 32'h421d08d7} /* (11, 4, 4) {real, imag} */,
  {32'h41c4c972, 32'h3f8db810} /* (11, 4, 3) {real, imag} */,
  {32'hc2a5b734, 32'hc26af7c2} /* (11, 4, 2) {real, imag} */,
  {32'h43408df8, 32'h421aa2ac} /* (11, 4, 1) {real, imag} */,
  {32'h42371a2a, 32'hbed3c900} /* (11, 4, 0) {real, imag} */,
  {32'hc30b19d8, 32'h42a69cd3} /* (11, 3, 31) {real, imag} */,
  {32'h4275944e, 32'hc311ba98} /* (11, 3, 30) {real, imag} */,
  {32'hc184aeb0, 32'h40715d71} /* (11, 3, 29) {real, imag} */,
  {32'h421165ae, 32'h4223b7ce} /* (11, 3, 28) {real, imag} */,
  {32'hc21c72a8, 32'h41ab8ddc} /* (11, 3, 27) {real, imag} */,
  {32'h41768f00, 32'h41be8ddb} /* (11, 3, 26) {real, imag} */,
  {32'h4156db18, 32'h4154215b} /* (11, 3, 25) {real, imag} */,
  {32'h417b6f24, 32'hc1054884} /* (11, 3, 24) {real, imag} */,
  {32'h3f71a5d8, 32'hc194ef0d} /* (11, 3, 23) {real, imag} */,
  {32'hc0a4b3df, 32'h3fbcf700} /* (11, 3, 22) {real, imag} */,
  {32'h4122f6f6, 32'h4158ef20} /* (11, 3, 21) {real, imag} */,
  {32'h4064c866, 32'h40547bf8} /* (11, 3, 20) {real, imag} */,
  {32'hc187b2e5, 32'hc0814518} /* (11, 3, 19) {real, imag} */,
  {32'h4134affd, 32'hc020026a} /* (11, 3, 18) {real, imag} */,
  {32'h40bd38b9, 32'h41841238} /* (11, 3, 17) {real, imag} */,
  {32'h40bd5da3, 32'h4061fd4c} /* (11, 3, 16) {real, imag} */,
  {32'hc13b24df, 32'h410e0241} /* (11, 3, 15) {real, imag} */,
  {32'h41676c87, 32'hc1a51786} /* (11, 3, 14) {real, imag} */,
  {32'h40ecedaa, 32'hc0886d88} /* (11, 3, 13) {real, imag} */,
  {32'hc1012b32, 32'h406951ac} /* (11, 3, 12) {real, imag} */,
  {32'h4108b0bc, 32'h3d8c3880} /* (11, 3, 11) {real, imag} */,
  {32'h3f9710a0, 32'h40ed1b36} /* (11, 3, 10) {real, imag} */,
  {32'hc0716e68, 32'h4041a13a} /* (11, 3, 9) {real, imag} */,
  {32'h3e9138e0, 32'hc0f0f7d0} /* (11, 3, 8) {real, imag} */,
  {32'h404ea700, 32'hc16af6a7} /* (11, 3, 7) {real, imag} */,
  {32'h412bb0d2, 32'h41733f0e} /* (11, 3, 6) {real, imag} */,
  {32'hc0dc2517, 32'h41845129} /* (11, 3, 5) {real, imag} */,
  {32'hc1f0392a, 32'h412a3156} /* (11, 3, 4) {real, imag} */,
  {32'hc1e791f8, 32'h419ded94} /* (11, 3, 3) {real, imag} */,
  {32'h40ea39a6, 32'hc2bf8072} /* (11, 3, 2) {real, imag} */,
  {32'h42fa8474, 32'h42b84752} /* (11, 3, 1) {real, imag} */,
  {32'h40d248fc, 32'h414f0fc0} /* (11, 3, 0) {real, imag} */,
  {32'hc4a2d3e7, 32'hc2a5fec6} /* (11, 2, 31) {real, imag} */,
  {32'h44146cf5, 32'hc329b6b9} /* (11, 2, 30) {real, imag} */,
  {32'h41663a8e, 32'h418f9b23} /* (11, 2, 29) {real, imag} */,
  {32'hc19dab10, 32'h4295816a} /* (11, 2, 28) {real, imag} */,
  {32'h4265d2a9, 32'hc278bc99} /* (11, 2, 27) {real, imag} */,
  {32'h41a733b4, 32'h3fae574c} /* (11, 2, 26) {real, imag} */,
  {32'h4007a0e0, 32'h4199f4ae} /* (11, 2, 25) {real, imag} */,
  {32'h419d2549, 32'hc1a8191e} /* (11, 2, 24) {real, imag} */,
  {32'hc144d794, 32'h3fdc5d61} /* (11, 2, 23) {real, imag} */,
  {32'hc0b819b6, 32'h3fd7072e} /* (11, 2, 22) {real, imag} */,
  {32'h40d4685b, 32'hc187d2e6} /* (11, 2, 21) {real, imag} */,
  {32'h403c91c2, 32'hc0ed56de} /* (11, 2, 20) {real, imag} */,
  {32'h40c43f56, 32'hc0a49ffc} /* (11, 2, 19) {real, imag} */,
  {32'h405b82a4, 32'hc024a3b0} /* (11, 2, 18) {real, imag} */,
  {32'hc04e5bdc, 32'hbf1afbc8} /* (11, 2, 17) {real, imag} */,
  {32'h410832fd, 32'h41146250} /* (11, 2, 16) {real, imag} */,
  {32'hc052eabc, 32'hbf0399b4} /* (11, 2, 15) {real, imag} */,
  {32'hc0f3e864, 32'h41743ab2} /* (11, 2, 14) {real, imag} */,
  {32'hc08631ae, 32'h41372442} /* (11, 2, 13) {real, imag} */,
  {32'hc0a61eab, 32'h411d2899} /* (11, 2, 12) {real, imag} */,
  {32'hc01d7fdb, 32'h412a87b8} /* (11, 2, 11) {real, imag} */,
  {32'hc169774a, 32'h415d6098} /* (11, 2, 10) {real, imag} */,
  {32'hc09ec5e5, 32'h403048d6} /* (11, 2, 9) {real, imag} */,
  {32'h41b9ea27, 32'hc0bbcba8} /* (11, 2, 8) {real, imag} */,
  {32'h40fc800a, 32'hc12df187} /* (11, 2, 7) {real, imag} */,
  {32'h40fd25a2, 32'h41806988} /* (11, 2, 6) {real, imag} */,
  {32'h4203386e, 32'h42a7a44e} /* (11, 2, 5) {real, imag} */,
  {32'hc2b8eb7c, 32'hc260db92} /* (11, 2, 4) {real, imag} */,
  {32'h41c20d4e, 32'h41283537} /* (11, 2, 3) {real, imag} */,
  {32'h43cfd23c, 32'hc314bb92} /* (11, 2, 2) {real, imag} */,
  {32'hc4322ee0, 32'h4314410d} /* (11, 2, 1) {real, imag} */,
  {32'hc4305fe6, 32'hc2b997dd} /* (11, 2, 0) {real, imag} */,
  {32'h44d828b8, 32'hc3a8e473} /* (11, 1, 31) {real, imag} */,
  {32'hc3d0f2a6, 32'h422397b6} /* (11, 1, 30) {real, imag} */,
  {32'hc2060f91, 32'h41392c88} /* (11, 1, 29) {real, imag} */,
  {32'h4292dd6a, 32'h4299fd52} /* (11, 1, 28) {real, imag} */,
  {32'hc2cbfb52, 32'hc1c2caa2} /* (11, 1, 27) {real, imag} */,
  {32'hc13e4c19, 32'hc1179d96} /* (11, 1, 26) {real, imag} */,
  {32'hbf1e8988, 32'hbf38fcc0} /* (11, 1, 25) {real, imag} */,
  {32'hc1bbe2a0, 32'h4135c5c2} /* (11, 1, 24) {real, imag} */,
  {32'hc0a78aaa, 32'h3f96b98c} /* (11, 1, 23) {real, imag} */,
  {32'h41b0ff67, 32'h415d148e} /* (11, 1, 22) {real, imag} */,
  {32'hc1a4b3b3, 32'h4183fd85} /* (11, 1, 21) {real, imag} */,
  {32'hbef4ff30, 32'hc0ebd418} /* (11, 1, 20) {real, imag} */,
  {32'hc154bc87, 32'hc1011ae7} /* (11, 1, 19) {real, imag} */,
  {32'h41492734, 32'h40acc043} /* (11, 1, 18) {real, imag} */,
  {32'h4062abba, 32'hc0327d7b} /* (11, 1, 17) {real, imag} */,
  {32'h408d58e0, 32'h400b5178} /* (11, 1, 16) {real, imag} */,
  {32'h4082144c, 32'h415e22b7} /* (11, 1, 15) {real, imag} */,
  {32'h4064843e, 32'hc1494fd0} /* (11, 1, 14) {real, imag} */,
  {32'h40aead9e, 32'hc0d33833} /* (11, 1, 13) {real, imag} */,
  {32'h41010d18, 32'hbf2add90} /* (11, 1, 12) {real, imag} */,
  {32'hc0be8105, 32'h400599f8} /* (11, 1, 11) {real, imag} */,
  {32'hc01b7a58, 32'hc1cc444a} /* (11, 1, 10) {real, imag} */,
  {32'hc06a4a50, 32'h4149b67f} /* (11, 1, 9) {real, imag} */,
  {32'hc1adc14c, 32'hc1d476fd} /* (11, 1, 8) {real, imag} */,
  {32'h415375ce, 32'h415247be} /* (11, 1, 7) {real, imag} */,
  {32'hc21ff0dc, 32'hc19ed53d} /* (11, 1, 6) {real, imag} */,
  {32'hc2c977e0, 32'hc1db971f} /* (11, 1, 5) {real, imag} */,
  {32'hc1890778, 32'h4206aac5} /* (11, 1, 4) {real, imag} */,
  {32'h419a8a95, 32'h412f0cb7} /* (11, 1, 3) {real, imag} */,
  {32'hc423c4f9, 32'hc411f708} /* (11, 1, 2) {real, imag} */,
  {32'h4519e3e7, 32'h44afb621} /* (11, 1, 1) {real, imag} */,
  {32'h450eea0c, 32'h430f22b4} /* (11, 1, 0) {real, imag} */,
  {32'h44af8898, 32'hc48f875f} /* (11, 0, 31) {real, imag} */,
  {32'hc35361cb, 32'h43993e16} /* (11, 0, 30) {real, imag} */,
  {32'hc2527aea, 32'h41627042} /* (11, 0, 29) {real, imag} */,
  {32'hc17fd20c, 32'h4207513c} /* (11, 0, 28) {real, imag} */,
  {32'hc23d83d5, 32'h422c4a98} /* (11, 0, 27) {real, imag} */,
  {32'hc0d424e8, 32'h40143660} /* (11, 0, 26) {real, imag} */,
  {32'h41b8b7ee, 32'hc138fe24} /* (11, 0, 25) {real, imag} */,
  {32'h41502eed, 32'h4148aa2a} /* (11, 0, 24) {real, imag} */,
  {32'hc11c6dd5, 32'h41997224} /* (11, 0, 23) {real, imag} */,
  {32'h413f3bdc, 32'h3fd2e7c4} /* (11, 0, 22) {real, imag} */,
  {32'hc11176a8, 32'h4110c282} /* (11, 0, 21) {real, imag} */,
  {32'hc09e8999, 32'hbfc8f784} /* (11, 0, 20) {real, imag} */,
  {32'hc0a231af, 32'hc0cc03cc} /* (11, 0, 19) {real, imag} */,
  {32'h410a32a0, 32'hc082c9d3} /* (11, 0, 18) {real, imag} */,
  {32'hc0047984, 32'hc0fab4f5} /* (11, 0, 17) {real, imag} */,
  {32'hc10f5536, 32'h00000000} /* (11, 0, 16) {real, imag} */,
  {32'hc0047984, 32'h40fab4f5} /* (11, 0, 15) {real, imag} */,
  {32'h410a32a0, 32'h4082c9d3} /* (11, 0, 14) {real, imag} */,
  {32'hc0a231af, 32'h40cc03cc} /* (11, 0, 13) {real, imag} */,
  {32'hc09e8999, 32'h3fc8f784} /* (11, 0, 12) {real, imag} */,
  {32'hc11176a8, 32'hc110c282} /* (11, 0, 11) {real, imag} */,
  {32'h413f3bdc, 32'hbfd2e7c4} /* (11, 0, 10) {real, imag} */,
  {32'hc11c6dd5, 32'hc1997224} /* (11, 0, 9) {real, imag} */,
  {32'h41502eed, 32'hc148aa2a} /* (11, 0, 8) {real, imag} */,
  {32'h41b8b7ee, 32'h4138fe24} /* (11, 0, 7) {real, imag} */,
  {32'hc0d424e8, 32'hc0143660} /* (11, 0, 6) {real, imag} */,
  {32'hc23d83d5, 32'hc22c4a98} /* (11, 0, 5) {real, imag} */,
  {32'hc17fd20c, 32'hc207513c} /* (11, 0, 4) {real, imag} */,
  {32'hc2527aea, 32'hc1627042} /* (11, 0, 3) {real, imag} */,
  {32'hc35361cb, 32'hc3993e16} /* (11, 0, 2) {real, imag} */,
  {32'h44af8898, 32'h448f875f} /* (11, 0, 1) {real, imag} */,
  {32'h4511a423, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h451efe91, 32'hc4aba8a3} /* (10, 31, 31) {real, imag} */,
  {32'hc426c6c3, 32'h441153f9} /* (10, 31, 30) {real, imag} */,
  {32'h413a26f6, 32'hc18fa254} /* (10, 31, 29) {real, imag} */,
  {32'h41ee46f0, 32'hc194ad6e} /* (10, 31, 28) {real, imag} */,
  {32'hc298ff05, 32'h422e35bf} /* (10, 31, 27) {real, imag} */,
  {32'hc1f2cde9, 32'h416495df} /* (10, 31, 26) {real, imag} */,
  {32'h41cbec46, 32'hc0585798} /* (10, 31, 25) {real, imag} */,
  {32'hc0cb65a5, 32'h421efba0} /* (10, 31, 24) {real, imag} */,
  {32'h415610f2, 32'hc1536679} /* (10, 31, 23) {real, imag} */,
  {32'hc1b840ff, 32'h41a64742} /* (10, 31, 22) {real, imag} */,
  {32'hc08245ae, 32'h41812527} /* (10, 31, 21) {real, imag} */,
  {32'hc0a09591, 32'h40b3e00a} /* (10, 31, 20) {real, imag} */,
  {32'h400bff88, 32'hc05fbd1d} /* (10, 31, 19) {real, imag} */,
  {32'hc1800dfd, 32'h40859b5b} /* (10, 31, 18) {real, imag} */,
  {32'h4051caf9, 32'hc0732b67} /* (10, 31, 17) {real, imag} */,
  {32'h40b83cba, 32'hc1152a10} /* (10, 31, 16) {real, imag} */,
  {32'h3f91158e, 32'hc04c2d37} /* (10, 31, 15) {real, imag} */,
  {32'hc090a2dc, 32'hc19a1f74} /* (10, 31, 14) {real, imag} */,
  {32'h412db4a1, 32'h40c40fd4} /* (10, 31, 13) {real, imag} */,
  {32'h4000cd76, 32'hc1a25556} /* (10, 31, 12) {real, imag} */,
  {32'hc1990ec6, 32'hc18a5b84} /* (10, 31, 11) {real, imag} */,
  {32'h417baf31, 32'hc0e19633} /* (10, 31, 10) {real, imag} */,
  {32'hc145b17c, 32'h409df8ba} /* (10, 31, 9) {real, imag} */,
  {32'hc1417d14, 32'hc17e305e} /* (10, 31, 8) {real, imag} */,
  {32'h419a37d0, 32'h40bdf30c} /* (10, 31, 7) {real, imag} */,
  {32'hc0c39d6c, 32'hc1a2217c} /* (10, 31, 6) {real, imag} */,
  {32'hc2ac58a1, 32'hc0b16332} /* (10, 31, 5) {real, imag} */,
  {32'h42a40b94, 32'hc2c8fb02} /* (10, 31, 4) {real, imag} */,
  {32'hc23f9288, 32'h4140efc8} /* (10, 31, 3) {real, imag} */,
  {32'hc3c8ff00, 32'hc2835e8e} /* (10, 31, 2) {real, imag} */,
  {32'h44dbfc61, 32'h43c114bf} /* (10, 31, 1) {real, imag} */,
  {32'h4513f624, 32'hc31af701} /* (10, 31, 0) {real, imag} */,
  {32'hc4396d1f, 32'hc3432882} /* (10, 30, 31) {real, imag} */,
  {32'h43d96382, 32'h42fb0336} /* (10, 30, 30) {real, imag} */,
  {32'h4118f22c, 32'hc1bbb3fa} /* (10, 30, 29) {real, imag} */,
  {32'hc2da8845, 32'h42234d5f} /* (10, 30, 28) {real, imag} */,
  {32'h41b8be07, 32'hc2a4d4b0} /* (10, 30, 27) {real, imag} */,
  {32'h4120cdd9, 32'h413c4cc4} /* (10, 30, 26) {real, imag} */,
  {32'hc0b0361a, 32'hc090cd6e} /* (10, 30, 25) {real, imag} */,
  {32'h411e3d37, 32'hc15981f6} /* (10, 30, 24) {real, imag} */,
  {32'h40a4d237, 32'hc116ef5e} /* (10, 30, 23) {real, imag} */,
  {32'hc105d3ce, 32'h411270b6} /* (10, 30, 22) {real, imag} */,
  {32'h40765eba, 32'hc174724e} /* (10, 30, 21) {real, imag} */,
  {32'h3eaf0bb0, 32'h40ba3025} /* (10, 30, 20) {real, imag} */,
  {32'hc1626ec2, 32'h3fcfc3ce} /* (10, 30, 19) {real, imag} */,
  {32'hc0de5ca0, 32'h40c7287e} /* (10, 30, 18) {real, imag} */,
  {32'h40b0702c, 32'h40596098} /* (10, 30, 17) {real, imag} */,
  {32'h3fc072d6, 32'h3e8ce4e4} /* (10, 30, 16) {real, imag} */,
  {32'hc11f4e31, 32'h40a609e4} /* (10, 30, 15) {real, imag} */,
  {32'h415c69c6, 32'h3ef554c0} /* (10, 30, 14) {real, imag} */,
  {32'hc11bee8f, 32'hc13b9980} /* (10, 30, 13) {real, imag} */,
  {32'hc0193ade, 32'hc164c944} /* (10, 30, 12) {real, imag} */,
  {32'h41025ba0, 32'h41cd0b2e} /* (10, 30, 11) {real, imag} */,
  {32'hc1be6041, 32'h406e3dcc} /* (10, 30, 10) {real, imag} */,
  {32'hc159558d, 32'hc17da11c} /* (10, 30, 9) {real, imag} */,
  {32'h41ffbe08, 32'h41be5976} /* (10, 30, 8) {real, imag} */,
  {32'hbfceed28, 32'hc104b9c6} /* (10, 30, 7) {real, imag} */,
  {32'h415b121c, 32'h4131844a} /* (10, 30, 6) {real, imag} */,
  {32'h426cdb99, 32'h4283366a} /* (10, 30, 5) {real, imag} */,
  {32'hc1d745ae, 32'hc297b2b2} /* (10, 30, 4) {real, imag} */,
  {32'h421c33fc, 32'hc179fe47} /* (10, 30, 3) {real, imag} */,
  {32'h441603b2, 32'h43375182} /* (10, 30, 2) {real, imag} */,
  {32'hc4a5fe8d, 32'h429c5516} /* (10, 30, 1) {real, imag} */,
  {32'hc43a787e, 32'h42c83579} /* (10, 30, 0) {real, imag} */,
  {32'h42e2072d, 32'hc2af14e8} /* (10, 29, 31) {real, imag} */,
  {32'hc109bafa, 32'h42bcc3f5} /* (10, 29, 30) {real, imag} */,
  {32'hc1e2777a, 32'hc1bf6ded} /* (10, 29, 29) {real, imag} */,
  {32'hc2008b65, 32'hc1421998} /* (10, 29, 28) {real, imag} */,
  {32'hc1641416, 32'hc0a3e9b0} /* (10, 29, 27) {real, imag} */,
  {32'hc0931ff0, 32'h4028e1e6} /* (10, 29, 26) {real, imag} */,
  {32'hc1b941ad, 32'hc05b583a} /* (10, 29, 25) {real, imag} */,
  {32'hc0a8a9cd, 32'hc14d286b} /* (10, 29, 24) {real, imag} */,
  {32'h40b0e5d8, 32'h40a71cfc} /* (10, 29, 23) {real, imag} */,
  {32'h4143d934, 32'hc18a43c2} /* (10, 29, 22) {real, imag} */,
  {32'h40c6ee46, 32'hc11d725a} /* (10, 29, 21) {real, imag} */,
  {32'h4102f34d, 32'h41744d4e} /* (10, 29, 20) {real, imag} */,
  {32'hc0793449, 32'h41023aba} /* (10, 29, 19) {real, imag} */,
  {32'h4037676e, 32'h4183083f} /* (10, 29, 18) {real, imag} */,
  {32'h414e35d1, 32'h4077aef0} /* (10, 29, 17) {real, imag} */,
  {32'h4100181d, 32'h41235781} /* (10, 29, 16) {real, imag} */,
  {32'h40f8e119, 32'h4127a2b7} /* (10, 29, 15) {real, imag} */,
  {32'h3e3f6c60, 32'h40e61e3c} /* (10, 29, 14) {real, imag} */,
  {32'hc050782a, 32'hc08ed0de} /* (10, 29, 13) {real, imag} */,
  {32'hc0c069a9, 32'h4063beb6} /* (10, 29, 12) {real, imag} */,
  {32'h4085c79c, 32'hc14b789a} /* (10, 29, 11) {real, imag} */,
  {32'hc1cfb06f, 32'h4101a298} /* (10, 29, 10) {real, imag} */,
  {32'hc125ea66, 32'hbff8f1ec} /* (10, 29, 9) {real, imag} */,
  {32'h414fb88f, 32'hbf1aa348} /* (10, 29, 8) {real, imag} */,
  {32'hc02912a0, 32'hc14d37e6} /* (10, 29, 7) {real, imag} */,
  {32'h4110f1bc, 32'hc14cc7d7} /* (10, 29, 6) {real, imag} */,
  {32'hc2250c8d, 32'hc118a6f2} /* (10, 29, 5) {real, imag} */,
  {32'h426266e6, 32'hc1f1744a} /* (10, 29, 4) {real, imag} */,
  {32'hc18d50d6, 32'h416aafbd} /* (10, 29, 3) {real, imag} */,
  {32'h428616b9, 32'h4306af0b} /* (10, 29, 2) {real, imag} */,
  {32'hc3132d8f, 32'hc2969b15} /* (10, 29, 1) {real, imag} */,
  {32'hc18b8942, 32'hc153d01e} /* (10, 29, 0) {real, imag} */,
  {32'h4320d659, 32'hc1f4a87c} /* (10, 28, 31) {real, imag} */,
  {32'hc2723e65, 32'h42867505} /* (10, 28, 30) {real, imag} */,
  {32'hc1be0e15, 32'hc1c8c00c} /* (10, 28, 29) {real, imag} */,
  {32'h4103c62a, 32'hc22d6279} /* (10, 28, 28) {real, imag} */,
  {32'h41bb4502, 32'h41ea884e} /* (10, 28, 27) {real, imag} */,
  {32'hc10e99b2, 32'hc0f08c46} /* (10, 28, 26) {real, imag} */,
  {32'hc08ea97a, 32'h4170f572} /* (10, 28, 25) {real, imag} */,
  {32'hc0fa4f8a, 32'h4195bba6} /* (10, 28, 24) {real, imag} */,
  {32'h4128f3dc, 32'hbf46fc50} /* (10, 28, 23) {real, imag} */,
  {32'h40c785c2, 32'hc0b6f94a} /* (10, 28, 22) {real, imag} */,
  {32'h412d264f, 32'h41a4f36a} /* (10, 28, 21) {real, imag} */,
  {32'hbfd5ee12, 32'hc100befa} /* (10, 28, 20) {real, imag} */,
  {32'h41198148, 32'h40b5d58a} /* (10, 28, 19) {real, imag} */,
  {32'h414b1034, 32'h40d1dd42} /* (10, 28, 18) {real, imag} */,
  {32'hc1715748, 32'hc042e7de} /* (10, 28, 17) {real, imag} */,
  {32'hc0c12340, 32'hc0be4c8e} /* (10, 28, 16) {real, imag} */,
  {32'hbf694099, 32'hc11789d1} /* (10, 28, 15) {real, imag} */,
  {32'hc17985ac, 32'h40d4fb4d} /* (10, 28, 14) {real, imag} */,
  {32'hc022d4be, 32'hc07e574f} /* (10, 28, 13) {real, imag} */,
  {32'hbfa6e504, 32'hc0a2caea} /* (10, 28, 12) {real, imag} */,
  {32'h401a743e, 32'h41484bda} /* (10, 28, 11) {real, imag} */,
  {32'hbffcab1e, 32'h414c7819} /* (10, 28, 10) {real, imag} */,
  {32'h42018976, 32'hc02a7794} /* (10, 28, 9) {real, imag} */,
  {32'h40fa51c2, 32'h41b2c919} /* (10, 28, 8) {real, imag} */,
  {32'h418a8bbe, 32'h412248d0} /* (10, 28, 7) {real, imag} */,
  {32'hc1c2a438, 32'hc1f64a91} /* (10, 28, 6) {real, imag} */,
  {32'hc1bdf03a, 32'h40374726} /* (10, 28, 5) {real, imag} */,
  {32'h41d9b136, 32'h3f9431c0} /* (10, 28, 4) {real, imag} */,
  {32'hc122bd6f, 32'h411e0276} /* (10, 28, 3) {real, imag} */,
  {32'hc2d31cbd, 32'h425e677d} /* (10, 28, 2) {real, imag} */,
  {32'h424fee04, 32'hc2c31e08} /* (10, 28, 1) {real, imag} */,
  {32'h420e4851, 32'hc1c8d2d6} /* (10, 28, 0) {real, imag} */,
  {32'hc1b97270, 32'h4296f74f} /* (10, 27, 31) {real, imag} */,
  {32'h40b58d21, 32'hc24f3922} /* (10, 27, 30) {real, imag} */,
  {32'hbf8781a6, 32'hc0e7cf3e} /* (10, 27, 29) {real, imag} */,
  {32'hc1498c26, 32'h406c0e60} /* (10, 27, 28) {real, imag} */,
  {32'h416b48f2, 32'hc04a52fc} /* (10, 27, 27) {real, imag} */,
  {32'hc142a20a, 32'hc0b6320f} /* (10, 27, 26) {real, imag} */,
  {32'h40e1c7d1, 32'h416cdcec} /* (10, 27, 25) {real, imag} */,
  {32'h4093ef7c, 32'hc1a614c8} /* (10, 27, 24) {real, imag} */,
  {32'h408065c7, 32'h3fcb01ae} /* (10, 27, 23) {real, imag} */,
  {32'hc04c3ce4, 32'hc0f836f4} /* (10, 27, 22) {real, imag} */,
  {32'hc13e69ec, 32'h403b47d4} /* (10, 27, 21) {real, imag} */,
  {32'h41304136, 32'h3f558a98} /* (10, 27, 20) {real, imag} */,
  {32'h41704e62, 32'hc045caa6} /* (10, 27, 19) {real, imag} */,
  {32'h3fd0c5a8, 32'hc18303a3} /* (10, 27, 18) {real, imag} */,
  {32'hc14c0665, 32'hc138def2} /* (10, 27, 17) {real, imag} */,
  {32'hc1365de8, 32'h3e7428e0} /* (10, 27, 16) {real, imag} */,
  {32'h40072c74, 32'h414ef872} /* (10, 27, 15) {real, imag} */,
  {32'hc1346b8a, 32'h4188a1de} /* (10, 27, 14) {real, imag} */,
  {32'hc0a51228, 32'h41147946} /* (10, 27, 13) {real, imag} */,
  {32'h3f4b6310, 32'h40889820} /* (10, 27, 12) {real, imag} */,
  {32'h413941ec, 32'h418fbac8} /* (10, 27, 11) {real, imag} */,
  {32'hbf708d80, 32'h4186e724} /* (10, 27, 10) {real, imag} */,
  {32'hc0fc6160, 32'hc1abe7ec} /* (10, 27, 9) {real, imag} */,
  {32'hc0fd51ed, 32'h41ce30a1} /* (10, 27, 8) {real, imag} */,
  {32'hc10b137d, 32'hc12aa6b6} /* (10, 27, 7) {real, imag} */,
  {32'h3f96d8a6, 32'h40accbba} /* (10, 27, 6) {real, imag} */,
  {32'hbf2065c0, 32'hc1889e1a} /* (10, 27, 5) {real, imag} */,
  {32'hc198c64c, 32'hc224a9bc} /* (10, 27, 4) {real, imag} */,
  {32'h40e32c50, 32'h40ae0a9c} /* (10, 27, 3) {real, imag} */,
  {32'h41a62202, 32'hbfb336e4} /* (10, 27, 2) {real, imag} */,
  {32'hc2eabc8a, 32'h420d0e4b} /* (10, 27, 1) {real, imag} */,
  {32'hc27fea3c, 32'h41af539a} /* (10, 27, 0) {real, imag} */,
  {32'h4092ea6f, 32'hc060ba35} /* (10, 26, 31) {real, imag} */,
  {32'h40b40756, 32'h41e53a70} /* (10, 26, 30) {real, imag} */,
  {32'hc18660e2, 32'hc119004f} /* (10, 26, 29) {real, imag} */,
  {32'hc170f791, 32'hc0adc047} /* (10, 26, 28) {real, imag} */,
  {32'h41751b72, 32'hc190de38} /* (10, 26, 27) {real, imag} */,
  {32'h41080f86, 32'hc0f865d0} /* (10, 26, 26) {real, imag} */,
  {32'h40db68c6, 32'hbf1a1a74} /* (10, 26, 25) {real, imag} */,
  {32'h4132085c, 32'h414d03a0} /* (10, 26, 24) {real, imag} */,
  {32'hc0d75db9, 32'h412da22c} /* (10, 26, 23) {real, imag} */,
  {32'hc12864fe, 32'h418a5a38} /* (10, 26, 22) {real, imag} */,
  {32'hbfc15018, 32'h403b5f55} /* (10, 26, 21) {real, imag} */,
  {32'h40bc5ec8, 32'hbfb5c8d8} /* (10, 26, 20) {real, imag} */,
  {32'h40d75e53, 32'hbe985e58} /* (10, 26, 19) {real, imag} */,
  {32'h40960ce0, 32'hc098a832} /* (10, 26, 18) {real, imag} */,
  {32'hc10d7742, 32'h4124c742} /* (10, 26, 17) {real, imag} */,
  {32'hc0ce252f, 32'hc0b410c8} /* (10, 26, 16) {real, imag} */,
  {32'hc0cf61ad, 32'hc1307e25} /* (10, 26, 15) {real, imag} */,
  {32'h415c0d4e, 32'hc0a28c80} /* (10, 26, 14) {real, imag} */,
  {32'h407485ac, 32'hc10f34d3} /* (10, 26, 13) {real, imag} */,
  {32'h40b07835, 32'h402cd542} /* (10, 26, 12) {real, imag} */,
  {32'h4184eafa, 32'hc047a064} /* (10, 26, 11) {real, imag} */,
  {32'hc149291f, 32'h411e04d6} /* (10, 26, 10) {real, imag} */,
  {32'h419723af, 32'hc1baa62b} /* (10, 26, 9) {real, imag} */,
  {32'hc18733ec, 32'h401e231a} /* (10, 26, 8) {real, imag} */,
  {32'h4069f31a, 32'hbfbea0aa} /* (10, 26, 7) {real, imag} */,
  {32'h418ce352, 32'h40480454} /* (10, 26, 6) {real, imag} */,
  {32'hc0734e34, 32'h41826ce0} /* (10, 26, 5) {real, imag} */,
  {32'h41855990, 32'h41745ae2} /* (10, 26, 4) {real, imag} */,
  {32'h413775b0, 32'hc0e30794} /* (10, 26, 3) {real, imag} */,
  {32'h40b3ca98, 32'h41979fa5} /* (10, 26, 2) {real, imag} */,
  {32'h40d830fb, 32'h41efaceb} /* (10, 26, 1) {real, imag} */,
  {32'h41769ea5, 32'hc2090978} /* (10, 26, 0) {real, imag} */,
  {32'h4111935c, 32'hc2049c11} /* (10, 25, 31) {real, imag} */,
  {32'hc1ef7fec, 32'hc0afa876} /* (10, 25, 30) {real, imag} */,
  {32'h40ad01ea, 32'hbf1be220} /* (10, 25, 29) {real, imag} */,
  {32'h41099ee6, 32'h3fd119ac} /* (10, 25, 28) {real, imag} */,
  {32'hc13c49d7, 32'h41734e13} /* (10, 25, 27) {real, imag} */,
  {32'h41ad079d, 32'h4147d92e} /* (10, 25, 26) {real, imag} */,
  {32'h3f23ec04, 32'hc0ca5ba0} /* (10, 25, 25) {real, imag} */,
  {32'hc0ea2445, 32'h4078ea24} /* (10, 25, 24) {real, imag} */,
  {32'h40f8411d, 32'hc0eb41af} /* (10, 25, 23) {real, imag} */,
  {32'hc1112bac, 32'h418bc44e} /* (10, 25, 22) {real, imag} */,
  {32'h41047a21, 32'hc008cd62} /* (10, 25, 21) {real, imag} */,
  {32'hc04daff6, 32'h40f992ea} /* (10, 25, 20) {real, imag} */,
  {32'hc091c783, 32'hc18c4352} /* (10, 25, 19) {real, imag} */,
  {32'hc0af21c1, 32'hc0b7241a} /* (10, 25, 18) {real, imag} */,
  {32'hc0649754, 32'hc042f983} /* (10, 25, 17) {real, imag} */,
  {32'h40ac5d66, 32'hc09f3b01} /* (10, 25, 16) {real, imag} */,
  {32'hc11373db, 32'hbf2716b4} /* (10, 25, 15) {real, imag} */,
  {32'h408dbfbd, 32'hbf85f2dc} /* (10, 25, 14) {real, imag} */,
  {32'h4114a0c8, 32'h3efd6268} /* (10, 25, 13) {real, imag} */,
  {32'hc184d64e, 32'h4114327a} /* (10, 25, 12) {real, imag} */,
  {32'h415bf115, 32'hc0dc1bf8} /* (10, 25, 11) {real, imag} */,
  {32'h40ba942b, 32'h4003dab0} /* (10, 25, 10) {real, imag} */,
  {32'hc186f702, 32'h4169e925} /* (10, 25, 9) {real, imag} */,
  {32'hc1a46fb4, 32'hc021a142} /* (10, 25, 8) {real, imag} */,
  {32'h40f63c32, 32'h411856da} /* (10, 25, 7) {real, imag} */,
  {32'h3f9aec8c, 32'hbed979c0} /* (10, 25, 6) {real, imag} */,
  {32'hc10c15e7, 32'hc0b1358c} /* (10, 25, 5) {real, imag} */,
  {32'h3fe60260, 32'hc0fd965e} /* (10, 25, 4) {real, imag} */,
  {32'hc1c36b20, 32'hc1ff86b0} /* (10, 25, 3) {real, imag} */,
  {32'hc14bf404, 32'h41cc03fe} /* (10, 25, 2) {real, imag} */,
  {32'h41b45426, 32'hc1b3471e} /* (10, 25, 1) {real, imag} */,
  {32'h409304cd, 32'h40d6311a} /* (10, 25, 0) {real, imag} */,
  {32'hc1ad2c34, 32'h41a0f196} /* (10, 24, 31) {real, imag} */,
  {32'h41e6be6d, 32'hc1210aa6} /* (10, 24, 30) {real, imag} */,
  {32'hbfe9c1f0, 32'hc0044dea} /* (10, 24, 29) {real, imag} */,
  {32'hc198bc52, 32'h3fcfee58} /* (10, 24, 28) {real, imag} */,
  {32'h41545845, 32'h4132d86a} /* (10, 24, 27) {real, imag} */,
  {32'h413d43ec, 32'hc0c6fdc7} /* (10, 24, 26) {real, imag} */,
  {32'h41d2ab84, 32'hc0f806b1} /* (10, 24, 25) {real, imag} */,
  {32'h40e87609, 32'hc01fe71c} /* (10, 24, 24) {real, imag} */,
  {32'hc138d2d8, 32'hc13c13a2} /* (10, 24, 23) {real, imag} */,
  {32'h40b573bc, 32'hc10ba8b5} /* (10, 24, 22) {real, imag} */,
  {32'h41007f1a, 32'hc0be2169} /* (10, 24, 21) {real, imag} */,
  {32'h4171e022, 32'hbec96a18} /* (10, 24, 20) {real, imag} */,
  {32'hc1888a74, 32'hc04a7901} /* (10, 24, 19) {real, imag} */,
  {32'h40df11f0, 32'h410ae8e6} /* (10, 24, 18) {real, imag} */,
  {32'hc0c97abf, 32'h3f43a9f2} /* (10, 24, 17) {real, imag} */,
  {32'h40c4da08, 32'hc018bed6} /* (10, 24, 16) {real, imag} */,
  {32'h3dda7270, 32'h404904d4} /* (10, 24, 15) {real, imag} */,
  {32'h40daee5c, 32'h3f8d43ac} /* (10, 24, 14) {real, imag} */,
  {32'h40af29d7, 32'h40a352b2} /* (10, 24, 13) {real, imag} */,
  {32'hc0ceebb0, 32'hc17d0eab} /* (10, 24, 12) {real, imag} */,
  {32'hc1c3b31c, 32'hc14361e6} /* (10, 24, 11) {real, imag} */,
  {32'h412944f4, 32'hc1822d24} /* (10, 24, 10) {real, imag} */,
  {32'h3c402e00, 32'h409fece4} /* (10, 24, 9) {real, imag} */,
  {32'h40ebd6da, 32'hc02cd5d8} /* (10, 24, 8) {real, imag} */,
  {32'h40e6b0ee, 32'h409f6f35} /* (10, 24, 7) {real, imag} */,
  {32'hc0baa38a, 32'hbe681530} /* (10, 24, 6) {real, imag} */,
  {32'h4123aa99, 32'hc1a579c8} /* (10, 24, 5) {real, imag} */,
  {32'h4014b4e0, 32'hc16822cc} /* (10, 24, 4) {real, imag} */,
  {32'hc1cfcd71, 32'h4131a35c} /* (10, 24, 3) {real, imag} */,
  {32'h41d18910, 32'h40d37ba4} /* (10, 24, 2) {real, imag} */,
  {32'hc2324ca9, 32'h4115a032} /* (10, 24, 1) {real, imag} */,
  {32'hc0f07ef0, 32'h400f89fc} /* (10, 24, 0) {real, imag} */,
  {32'hc12d7b7c, 32'hc0bde6b8} /* (10, 23, 31) {real, imag} */,
  {32'h411e96bb, 32'h3f4981d0} /* (10, 23, 30) {real, imag} */,
  {32'h415da0d6, 32'hc0cf3848} /* (10, 23, 29) {real, imag} */,
  {32'hc186fc80, 32'h40a9addd} /* (10, 23, 28) {real, imag} */,
  {32'hc1d22072, 32'hc157c20d} /* (10, 23, 27) {real, imag} */,
  {32'h41689094, 32'h40dc2979} /* (10, 23, 26) {real, imag} */,
  {32'hc1122fa2, 32'hc14efc3d} /* (10, 23, 25) {real, imag} */,
  {32'hc135bec8, 32'hc1009cb6} /* (10, 23, 24) {real, imag} */,
  {32'hbf729870, 32'h40887d20} /* (10, 23, 23) {real, imag} */,
  {32'h40d73946, 32'h4131deb1} /* (10, 23, 22) {real, imag} */,
  {32'h41472496, 32'h40abf07f} /* (10, 23, 21) {real, imag} */,
  {32'hc145b78c, 32'hc05e6720} /* (10, 23, 20) {real, imag} */,
  {32'h4061e7b6, 32'h411fb2e6} /* (10, 23, 19) {real, imag} */,
  {32'hc03635f4, 32'h403c833a} /* (10, 23, 18) {real, imag} */,
  {32'hbf2f4150, 32'hc12f4e2e} /* (10, 23, 17) {real, imag} */,
  {32'h40879d7f, 32'hc07dba8f} /* (10, 23, 16) {real, imag} */,
  {32'hc1282b3c, 32'hc1823df6} /* (10, 23, 15) {real, imag} */,
  {32'h3fccee5c, 32'h41312e48} /* (10, 23, 14) {real, imag} */,
  {32'h406b7ec2, 32'h410cd24a} /* (10, 23, 13) {real, imag} */,
  {32'h40c9da7e, 32'h410c08d7} /* (10, 23, 12) {real, imag} */,
  {32'hc0053802, 32'h3f236c64} /* (10, 23, 11) {real, imag} */,
  {32'hc19427e9, 32'hc102f0e6} /* (10, 23, 10) {real, imag} */,
  {32'h4011e82e, 32'hc14f8337} /* (10, 23, 9) {real, imag} */,
  {32'hbf96f18c, 32'h40b60382} /* (10, 23, 8) {real, imag} */,
  {32'hc12dcd50, 32'hc18190c1} /* (10, 23, 7) {real, imag} */,
  {32'hbf7179d0, 32'hc05685ff} /* (10, 23, 6) {real, imag} */,
  {32'h418f3cf5, 32'h4167d96e} /* (10, 23, 5) {real, imag} */,
  {32'h4194934c, 32'h41829b66} /* (10, 23, 4) {real, imag} */,
  {32'h403fb233, 32'hc18e6b00} /* (10, 23, 3) {real, imag} */,
  {32'h401dce12, 32'h409385a6} /* (10, 23, 2) {real, imag} */,
  {32'hc0e5a079, 32'hc15b8d0e} /* (10, 23, 1) {real, imag} */,
  {32'h40b517b8, 32'hc0d6c3dc} /* (10, 23, 0) {real, imag} */,
  {32'h40d9c25e, 32'h41908b20} /* (10, 22, 31) {real, imag} */,
  {32'h413895e7, 32'h40993912} /* (10, 22, 30) {real, imag} */,
  {32'h418d75af, 32'hc1068f18} /* (10, 22, 29) {real, imag} */,
  {32'h401825ee, 32'hbe9b75d0} /* (10, 22, 28) {real, imag} */,
  {32'hc02b4a98, 32'hc0d7adaa} /* (10, 22, 27) {real, imag} */,
  {32'h40283776, 32'hc1f67f42} /* (10, 22, 26) {real, imag} */,
  {32'hc0d804ea, 32'h40bea2dc} /* (10, 22, 25) {real, imag} */,
  {32'h412e088a, 32'hc0cf30ef} /* (10, 22, 24) {real, imag} */,
  {32'hbf005a22, 32'hc1581694} /* (10, 22, 23) {real, imag} */,
  {32'hc190f4c0, 32'hc110c952} /* (10, 22, 22) {real, imag} */,
  {32'hbee3c410, 32'hbe80e9b0} /* (10, 22, 21) {real, imag} */,
  {32'h3f891e00, 32'h404a9fc3} /* (10, 22, 20) {real, imag} */,
  {32'h409003ce, 32'hc105c85e} /* (10, 22, 19) {real, imag} */,
  {32'hc1161929, 32'h41a87432} /* (10, 22, 18) {real, imag} */,
  {32'hc0994ae7, 32'h4017c988} /* (10, 22, 17) {real, imag} */,
  {32'h41168a7a, 32'hbf2d6051} /* (10, 22, 16) {real, imag} */,
  {32'h405ec206, 32'hc0d138ca} /* (10, 22, 15) {real, imag} */,
  {32'hc13bf96e, 32'hc173cac3} /* (10, 22, 14) {real, imag} */,
  {32'hc1c98cd9, 32'hc091347f} /* (10, 22, 13) {real, imag} */,
  {32'hc0dbbeca, 32'h41246791} /* (10, 22, 12) {real, imag} */,
  {32'hbf6dc230, 32'hc0132a68} /* (10, 22, 11) {real, imag} */,
  {32'h418e6c07, 32'hc0edadd4} /* (10, 22, 10) {real, imag} */,
  {32'h421a1203, 32'h41a2080c} /* (10, 22, 9) {real, imag} */,
  {32'h3f52c518, 32'hc15996de} /* (10, 22, 8) {real, imag} */,
  {32'hc1826acb, 32'h408b28e0} /* (10, 22, 7) {real, imag} */,
  {32'hc123ff92, 32'hc048b41c} /* (10, 22, 6) {real, imag} */,
  {32'h41263e9d, 32'h3f7eaff0} /* (10, 22, 5) {real, imag} */,
  {32'hc157ba32, 32'h415cc7e4} /* (10, 22, 4) {real, imag} */,
  {32'hc18609a1, 32'hc18f223e} /* (10, 22, 3) {real, imag} */,
  {32'hc182c7f1, 32'h412b0303} /* (10, 22, 2) {real, imag} */,
  {32'h415d45b6, 32'hc1bacea2} /* (10, 22, 1) {real, imag} */,
  {32'h40e13321, 32'h414b08e4} /* (10, 22, 0) {real, imag} */,
  {32'h405d58c0, 32'h41e19644} /* (10, 21, 31) {real, imag} */,
  {32'h414dcae8, 32'hc1ea414a} /* (10, 21, 30) {real, imag} */,
  {32'h41093868, 32'h415120c0} /* (10, 21, 29) {real, imag} */,
  {32'hc09f56df, 32'hbfca6b50} /* (10, 21, 28) {real, imag} */,
  {32'hc09ff534, 32'h40a80f58} /* (10, 21, 27) {real, imag} */,
  {32'hc1433582, 32'hbe99f688} /* (10, 21, 26) {real, imag} */,
  {32'h413a55ca, 32'h3da46ec0} /* (10, 21, 25) {real, imag} */,
  {32'hc04b67e1, 32'hc08cbced} /* (10, 21, 24) {real, imag} */,
  {32'h3fe526d8, 32'hc07e96a8} /* (10, 21, 23) {real, imag} */,
  {32'h40a2dfa0, 32'hc16ba651} /* (10, 21, 22) {real, imag} */,
  {32'h40073354, 32'h4157ca2c} /* (10, 21, 21) {real, imag} */,
  {32'h40e7de01, 32'h40429630} /* (10, 21, 20) {real, imag} */,
  {32'h4103ec10, 32'hc01fe034} /* (10, 21, 19) {real, imag} */,
  {32'hbf694eb0, 32'hc0c48978} /* (10, 21, 18) {real, imag} */,
  {32'hbf8cab43, 32'h408a2d41} /* (10, 21, 17) {real, imag} */,
  {32'h3fde7fe8, 32'h40af9a24} /* (10, 21, 16) {real, imag} */,
  {32'hbfa14410, 32'hc00fefb8} /* (10, 21, 15) {real, imag} */,
  {32'h3fe16fd0, 32'hc0d51636} /* (10, 21, 14) {real, imag} */,
  {32'h410fb54c, 32'h412d9d10} /* (10, 21, 13) {real, imag} */,
  {32'hc0ce49e6, 32'hbfa90bbc} /* (10, 21, 12) {real, imag} */,
  {32'hc03c2e66, 32'h4040431c} /* (10, 21, 11) {real, imag} */,
  {32'hc0b53044, 32'h411066e5} /* (10, 21, 10) {real, imag} */,
  {32'hc04bd6b4, 32'h41459990} /* (10, 21, 9) {real, imag} */,
  {32'h4122f08e, 32'h40e9b0ca} /* (10, 21, 8) {real, imag} */,
  {32'h3f6adecc, 32'h401e0f44} /* (10, 21, 7) {real, imag} */,
  {32'h3ffda398, 32'h41495140} /* (10, 21, 6) {real, imag} */,
  {32'hc098f5cc, 32'hc1bb91f0} /* (10, 21, 5) {real, imag} */,
  {32'hc0ed3def, 32'hc11922e0} /* (10, 21, 4) {real, imag} */,
  {32'h40870ad0, 32'hc0c82455} /* (10, 21, 3) {real, imag} */,
  {32'h41886ff5, 32'h4150a396} /* (10, 21, 2) {real, imag} */,
  {32'hc1b54e9f, 32'h41d6649e} /* (10, 21, 1) {real, imag} */,
  {32'hc10117b3, 32'h411bf5fa} /* (10, 21, 0) {real, imag} */,
  {32'h3fb63077, 32'h41317e1a} /* (10, 20, 31) {real, imag} */,
  {32'h409e5fac, 32'hbfa73846} /* (10, 20, 30) {real, imag} */,
  {32'h3d00cbc0, 32'h3f7db7b8} /* (10, 20, 29) {real, imag} */,
  {32'h3fe26a58, 32'h3e6f53c0} /* (10, 20, 28) {real, imag} */,
  {32'h3fb58808, 32'hc09997ae} /* (10, 20, 27) {real, imag} */,
  {32'hc093d743, 32'hc11b6d45} /* (10, 20, 26) {real, imag} */,
  {32'h405d3a60, 32'h3fb5a350} /* (10, 20, 25) {real, imag} */,
  {32'h413def97, 32'h4127fe78} /* (10, 20, 24) {real, imag} */,
  {32'hc0af8391, 32'h412e4d25} /* (10, 20, 23) {real, imag} */,
  {32'h403f504a, 32'hc18adf40} /* (10, 20, 22) {real, imag} */,
  {32'h413733ec, 32'h4111b54c} /* (10, 20, 21) {real, imag} */,
  {32'h40f5f3a3, 32'hc1eced0c} /* (10, 20, 20) {real, imag} */,
  {32'h40ba8f47, 32'hc02021fe} /* (10, 20, 19) {real, imag} */,
  {32'hbf1c8914, 32'hbe475dc0} /* (10, 20, 18) {real, imag} */,
  {32'hbf0172fa, 32'hc0d9c364} /* (10, 20, 17) {real, imag} */,
  {32'h40b54b75, 32'h4165d598} /* (10, 20, 16) {real, imag} */,
  {32'h419ab58a, 32'h40a96599} /* (10, 20, 15) {real, imag} */,
  {32'h41afb95c, 32'hc1592250} /* (10, 20, 14) {real, imag} */,
  {32'h414c2470, 32'hbef779b0} /* (10, 20, 13) {real, imag} */,
  {32'h4152590b, 32'h415ba271} /* (10, 20, 12) {real, imag} */,
  {32'hc0b25d14, 32'hc196fb79} /* (10, 20, 11) {real, imag} */,
  {32'hc0875636, 32'hc1995dfc} /* (10, 20, 10) {real, imag} */,
  {32'hc1676069, 32'hc0af3fc4} /* (10, 20, 9) {real, imag} */,
  {32'hc1b2548e, 32'h4190ad5c} /* (10, 20, 8) {real, imag} */,
  {32'h3d4f3c00, 32'h410f4533} /* (10, 20, 7) {real, imag} */,
  {32'h3f10fbce, 32'hc00159b1} /* (10, 20, 6) {real, imag} */,
  {32'hc1798fe0, 32'hbfa95612} /* (10, 20, 5) {real, imag} */,
  {32'h4198d651, 32'hc160cd8e} /* (10, 20, 4) {real, imag} */,
  {32'hc05af31c, 32'hc0efe81a} /* (10, 20, 3) {real, imag} */,
  {32'hbfaea8d4, 32'h40a095f6} /* (10, 20, 2) {real, imag} */,
  {32'h400bf65c, 32'h407497fc} /* (10, 20, 1) {real, imag} */,
  {32'h4168350e, 32'h400c8508} /* (10, 20, 0) {real, imag} */,
  {32'h40b23490, 32'hc1663914} /* (10, 19, 31) {real, imag} */,
  {32'hbe8a9490, 32'hc065422e} /* (10, 19, 30) {real, imag} */,
  {32'hc12d8fbf, 32'h40f2091a} /* (10, 19, 29) {real, imag} */,
  {32'hc12e5727, 32'hc019a04c} /* (10, 19, 28) {real, imag} */,
  {32'h40c99f61, 32'hbf9af158} /* (10, 19, 27) {real, imag} */,
  {32'h419c23d8, 32'h40c505f7} /* (10, 19, 26) {real, imag} */,
  {32'hc1ac7dc0, 32'hbf73c0ca} /* (10, 19, 25) {real, imag} */,
  {32'hc0340354, 32'h410d177e} /* (10, 19, 24) {real, imag} */,
  {32'hc1b660cc, 32'h3f1663b0} /* (10, 19, 23) {real, imag} */,
  {32'h40df9149, 32'hc118da90} /* (10, 19, 22) {real, imag} */,
  {32'hc0f896e7, 32'h3ff89f4c} /* (10, 19, 21) {real, imag} */,
  {32'hc116b404, 32'hc1c20a74} /* (10, 19, 20) {real, imag} */,
  {32'h4154107a, 32'hc12d62a8} /* (10, 19, 19) {real, imag} */,
  {32'h41680b84, 32'hbfbaedd6} /* (10, 19, 18) {real, imag} */,
  {32'hc08c162a, 32'hc07a210e} /* (10, 19, 17) {real, imag} */,
  {32'h40af03d6, 32'h407c8cda} /* (10, 19, 16) {real, imag} */,
  {32'h405edb84, 32'h418ae738} /* (10, 19, 15) {real, imag} */,
  {32'hc0cc3f0a, 32'h40569af3} /* (10, 19, 14) {real, imag} */,
  {32'h3ecaf8c0, 32'hc17c77d8} /* (10, 19, 13) {real, imag} */,
  {32'hc1969dd6, 32'h4095e2fa} /* (10, 19, 12) {real, imag} */,
  {32'h411cd426, 32'h41193716} /* (10, 19, 11) {real, imag} */,
  {32'hc0e22446, 32'hc148f396} /* (10, 19, 10) {real, imag} */,
  {32'hc01cc818, 32'hc0d4d5bc} /* (10, 19, 9) {real, imag} */,
  {32'h418111f8, 32'h410cf746} /* (10, 19, 8) {real, imag} */,
  {32'h411dead6, 32'hc0090416} /* (10, 19, 7) {real, imag} */,
  {32'hc1132130, 32'h41219e85} /* (10, 19, 6) {real, imag} */,
  {32'hbf194300, 32'h3ede28a0} /* (10, 19, 5) {real, imag} */,
  {32'hc1ab81e9, 32'hc0ae1866} /* (10, 19, 4) {real, imag} */,
  {32'hc03ae008, 32'h4147b4ee} /* (10, 19, 3) {real, imag} */,
  {32'h41228d1b, 32'hc014a478} /* (10, 19, 2) {real, imag} */,
  {32'h408747f5, 32'h406f4240} /* (10, 19, 1) {real, imag} */,
  {32'hc107d3e4, 32'h40861249} /* (10, 19, 0) {real, imag} */,
  {32'hc0cb93d4, 32'h41384052} /* (10, 18, 31) {real, imag} */,
  {32'hc160aa65, 32'hc112c846} /* (10, 18, 30) {real, imag} */,
  {32'h406fd0c1, 32'hc0f3f306} /* (10, 18, 29) {real, imag} */,
  {32'hc0e4ea3c, 32'h407b6aad} /* (10, 18, 28) {real, imag} */,
  {32'hc14c9a3d, 32'hc0627354} /* (10, 18, 27) {real, imag} */,
  {32'hc10fb9c9, 32'hc169e6c8} /* (10, 18, 26) {real, imag} */,
  {32'h3f8c5564, 32'hc0e7fa78} /* (10, 18, 25) {real, imag} */,
  {32'h3fa314e8, 32'hbeab1246} /* (10, 18, 24) {real, imag} */,
  {32'h409cb73e, 32'h40e70cf2} /* (10, 18, 23) {real, imag} */,
  {32'hbfdcc1ac, 32'hc0c935a2} /* (10, 18, 22) {real, imag} */,
  {32'hc10282fd, 32'hc1335619} /* (10, 18, 21) {real, imag} */,
  {32'hc0802586, 32'h409a33f8} /* (10, 18, 20) {real, imag} */,
  {32'hbfa475ec, 32'h40e19900} /* (10, 18, 19) {real, imag} */,
  {32'hc1a69095, 32'hc10886d4} /* (10, 18, 18) {real, imag} */,
  {32'hc0c89a27, 32'h41110f98} /* (10, 18, 17) {real, imag} */,
  {32'hc1229c90, 32'h3fcbee20} /* (10, 18, 16) {real, imag} */,
  {32'hc09ebb90, 32'hc07ca7f7} /* (10, 18, 15) {real, imag} */,
  {32'hc175dc4c, 32'hbf845bb6} /* (10, 18, 14) {real, imag} */,
  {32'hc0bf9eac, 32'hc092f9cf} /* (10, 18, 13) {real, imag} */,
  {32'h41431bd0, 32'hbfa973f8} /* (10, 18, 12) {real, imag} */,
  {32'hc13c7bc3, 32'hbc62e580} /* (10, 18, 11) {real, imag} */,
  {32'h417a794a, 32'hc0e1b230} /* (10, 18, 10) {real, imag} */,
  {32'hc12dd784, 32'h3f1d87c8} /* (10, 18, 9) {real, imag} */,
  {32'h408b06ce, 32'hbf512674} /* (10, 18, 8) {real, imag} */,
  {32'h40e8882c, 32'hbe94e880} /* (10, 18, 7) {real, imag} */,
  {32'h3fd03c48, 32'hc00e8f8a} /* (10, 18, 6) {real, imag} */,
  {32'h408da36a, 32'hc12789a6} /* (10, 18, 5) {real, imag} */,
  {32'hbf0fafa4, 32'h4198f33e} /* (10, 18, 4) {real, imag} */,
  {32'hbff283b4, 32'hc1405b34} /* (10, 18, 3) {real, imag} */,
  {32'h4121f970, 32'hc0035f1a} /* (10, 18, 2) {real, imag} */,
  {32'hc07c3d54, 32'h406fd73c} /* (10, 18, 1) {real, imag} */,
  {32'h40b817ae, 32'hbd3f4500} /* (10, 18, 0) {real, imag} */,
  {32'h3eba0ab0, 32'h40192a1e} /* (10, 17, 31) {real, imag} */,
  {32'h4130822e, 32'h3fb8a801} /* (10, 17, 30) {real, imag} */,
  {32'h40997e5f, 32'h3f8d814c} /* (10, 17, 29) {real, imag} */,
  {32'hc088bbd0, 32'h3e8cf420} /* (10, 17, 28) {real, imag} */,
  {32'hbfcea818, 32'hc107a424} /* (10, 17, 27) {real, imag} */,
  {32'hc051947f, 32'hc14285c1} /* (10, 17, 26) {real, imag} */,
  {32'hc0099612, 32'hc09bfdbb} /* (10, 17, 25) {real, imag} */,
  {32'h4059ede6, 32'hc05ee504} /* (10, 17, 24) {real, imag} */,
  {32'h40f444c5, 32'h3fa6f574} /* (10, 17, 23) {real, imag} */,
  {32'hc08165e2, 32'hc1244cc3} /* (10, 17, 22) {real, imag} */,
  {32'h4110b14c, 32'hbfd00dc0} /* (10, 17, 21) {real, imag} */,
  {32'hbf3ee0c0, 32'h3fe653cb} /* (10, 17, 20) {real, imag} */,
  {32'h410e1378, 32'h4161c03a} /* (10, 17, 19) {real, imag} */,
  {32'h40922540, 32'h40a2ac6c} /* (10, 17, 18) {real, imag} */,
  {32'hbfc81c40, 32'h4123ba62} /* (10, 17, 17) {real, imag} */,
  {32'hbfca1a4d, 32'h40598e40} /* (10, 17, 16) {real, imag} */,
  {32'h400b0468, 32'hbf8166ac} /* (10, 17, 15) {real, imag} */,
  {32'h3f3da87d, 32'hc03ea20c} /* (10, 17, 14) {real, imag} */,
  {32'h40e1be9c, 32'hc1314358} /* (10, 17, 13) {real, imag} */,
  {32'hbff1bebc, 32'hc047a6fa} /* (10, 17, 12) {real, imag} */,
  {32'hc0e17af8, 32'hc14422e6} /* (10, 17, 11) {real, imag} */,
  {32'hc15bcf1f, 32'hbfd5be90} /* (10, 17, 10) {real, imag} */,
  {32'h4003ee6a, 32'h40e5a8fc} /* (10, 17, 9) {real, imag} */,
  {32'hc0bf516a, 32'h3f9370ef} /* (10, 17, 8) {real, imag} */,
  {32'h4128045a, 32'hc08c9e97} /* (10, 17, 7) {real, imag} */,
  {32'h3fd3490d, 32'hc13a02aa} /* (10, 17, 6) {real, imag} */,
  {32'hbf75c7f8, 32'h4012d3fa} /* (10, 17, 5) {real, imag} */,
  {32'h408e4152, 32'hc09a45a4} /* (10, 17, 4) {real, imag} */,
  {32'hc028f10e, 32'h41234b36} /* (10, 17, 3) {real, imag} */,
  {32'h3f08b810, 32'h413d5f0c} /* (10, 17, 2) {real, imag} */,
  {32'hc111233c, 32'hc12ee632} /* (10, 17, 1) {real, imag} */,
  {32'hbfe4cf9e, 32'h3f857ca2} /* (10, 17, 0) {real, imag} */,
  {32'h40a0a4de, 32'h4093ad0a} /* (10, 16, 31) {real, imag} */,
  {32'h41152492, 32'h3f48019c} /* (10, 16, 30) {real, imag} */,
  {32'hc09cb169, 32'h407ba4c1} /* (10, 16, 29) {real, imag} */,
  {32'hbd8e80e0, 32'h410b8c0c} /* (10, 16, 28) {real, imag} */,
  {32'h3ffe8f82, 32'h40478213} /* (10, 16, 27) {real, imag} */,
  {32'h40a7d178, 32'h4020b31e} /* (10, 16, 26) {real, imag} */,
  {32'hc0bf5ce9, 32'h408a15d2} /* (10, 16, 25) {real, imag} */,
  {32'hc1458213, 32'hbfd4d3cc} /* (10, 16, 24) {real, imag} */,
  {32'hc0906e0e, 32'hc0abffa1} /* (10, 16, 23) {real, imag} */,
  {32'h40cb6be0, 32'h3d341c00} /* (10, 16, 22) {real, imag} */,
  {32'hc0dd8390, 32'hc1603c63} /* (10, 16, 21) {real, imag} */,
  {32'hbf7d9048, 32'hc0669390} /* (10, 16, 20) {real, imag} */,
  {32'h4071d3a7, 32'hc112e71c} /* (10, 16, 19) {real, imag} */,
  {32'h408165b9, 32'hc14fa58c} /* (10, 16, 18) {real, imag} */,
  {32'h4135cee0, 32'hbfc73f12} /* (10, 16, 17) {real, imag} */,
  {32'hc0f29103, 32'h00000000} /* (10, 16, 16) {real, imag} */,
  {32'h4135cee0, 32'h3fc73f12} /* (10, 16, 15) {real, imag} */,
  {32'h408165b9, 32'h414fa58c} /* (10, 16, 14) {real, imag} */,
  {32'h4071d3a7, 32'h4112e71c} /* (10, 16, 13) {real, imag} */,
  {32'hbf7d9048, 32'h40669390} /* (10, 16, 12) {real, imag} */,
  {32'hc0dd8390, 32'h41603c63} /* (10, 16, 11) {real, imag} */,
  {32'h40cb6be0, 32'hbd341c00} /* (10, 16, 10) {real, imag} */,
  {32'hc0906e0e, 32'h40abffa1} /* (10, 16, 9) {real, imag} */,
  {32'hc1458213, 32'h3fd4d3cc} /* (10, 16, 8) {real, imag} */,
  {32'hc0bf5ce9, 32'hc08a15d2} /* (10, 16, 7) {real, imag} */,
  {32'h40a7d178, 32'hc020b31e} /* (10, 16, 6) {real, imag} */,
  {32'h3ffe8f82, 32'hc0478213} /* (10, 16, 5) {real, imag} */,
  {32'hbd8e80e0, 32'hc10b8c0c} /* (10, 16, 4) {real, imag} */,
  {32'hc09cb169, 32'hc07ba4c1} /* (10, 16, 3) {real, imag} */,
  {32'h41152492, 32'hbf48019c} /* (10, 16, 2) {real, imag} */,
  {32'h40a0a4de, 32'hc093ad0a} /* (10, 16, 1) {real, imag} */,
  {32'hc0061760, 32'h00000000} /* (10, 16, 0) {real, imag} */,
  {32'hc111233c, 32'h412ee632} /* (10, 15, 31) {real, imag} */,
  {32'h3f08b810, 32'hc13d5f0c} /* (10, 15, 30) {real, imag} */,
  {32'hc028f10e, 32'hc1234b36} /* (10, 15, 29) {real, imag} */,
  {32'h408e4152, 32'h409a45a4} /* (10, 15, 28) {real, imag} */,
  {32'hbf75c7f8, 32'hc012d3fa} /* (10, 15, 27) {real, imag} */,
  {32'h3fd3490d, 32'h413a02aa} /* (10, 15, 26) {real, imag} */,
  {32'h4128045a, 32'h408c9e97} /* (10, 15, 25) {real, imag} */,
  {32'hc0bf516a, 32'hbf9370ef} /* (10, 15, 24) {real, imag} */,
  {32'h4003ee6a, 32'hc0e5a8fc} /* (10, 15, 23) {real, imag} */,
  {32'hc15bcf1f, 32'h3fd5be90} /* (10, 15, 22) {real, imag} */,
  {32'hc0e17af8, 32'h414422e6} /* (10, 15, 21) {real, imag} */,
  {32'hbff1bebc, 32'h4047a6fa} /* (10, 15, 20) {real, imag} */,
  {32'h40e1be9c, 32'h41314358} /* (10, 15, 19) {real, imag} */,
  {32'h3f3da87d, 32'h403ea20c} /* (10, 15, 18) {real, imag} */,
  {32'h400b0468, 32'h3f8166ac} /* (10, 15, 17) {real, imag} */,
  {32'hbfca1a4d, 32'hc0598e40} /* (10, 15, 16) {real, imag} */,
  {32'hbfc81c40, 32'hc123ba62} /* (10, 15, 15) {real, imag} */,
  {32'h40922540, 32'hc0a2ac6c} /* (10, 15, 14) {real, imag} */,
  {32'h410e1378, 32'hc161c03a} /* (10, 15, 13) {real, imag} */,
  {32'hbf3ee0c0, 32'hbfe653cb} /* (10, 15, 12) {real, imag} */,
  {32'h4110b14c, 32'h3fd00dc0} /* (10, 15, 11) {real, imag} */,
  {32'hc08165e2, 32'h41244cc3} /* (10, 15, 10) {real, imag} */,
  {32'h40f444c5, 32'hbfa6f574} /* (10, 15, 9) {real, imag} */,
  {32'h4059ede6, 32'h405ee504} /* (10, 15, 8) {real, imag} */,
  {32'hc0099612, 32'h409bfdbb} /* (10, 15, 7) {real, imag} */,
  {32'hc051947f, 32'h414285c1} /* (10, 15, 6) {real, imag} */,
  {32'hbfcea818, 32'h4107a424} /* (10, 15, 5) {real, imag} */,
  {32'hc088bbd0, 32'hbe8cf420} /* (10, 15, 4) {real, imag} */,
  {32'h40997e5f, 32'hbf8d814c} /* (10, 15, 3) {real, imag} */,
  {32'h4130822e, 32'hbfb8a801} /* (10, 15, 2) {real, imag} */,
  {32'h3eba0ab0, 32'hc0192a1e} /* (10, 15, 1) {real, imag} */,
  {32'hbfe4cf9e, 32'hbf857ca2} /* (10, 15, 0) {real, imag} */,
  {32'hc07c3d54, 32'hc06fd73c} /* (10, 14, 31) {real, imag} */,
  {32'h4121f970, 32'h40035f1a} /* (10, 14, 30) {real, imag} */,
  {32'hbff283b4, 32'h41405b34} /* (10, 14, 29) {real, imag} */,
  {32'hbf0fafa4, 32'hc198f33e} /* (10, 14, 28) {real, imag} */,
  {32'h408da36a, 32'h412789a6} /* (10, 14, 27) {real, imag} */,
  {32'h3fd03c48, 32'h400e8f8a} /* (10, 14, 26) {real, imag} */,
  {32'h40e8882c, 32'h3e94e880} /* (10, 14, 25) {real, imag} */,
  {32'h408b06ce, 32'h3f512674} /* (10, 14, 24) {real, imag} */,
  {32'hc12dd784, 32'hbf1d87c8} /* (10, 14, 23) {real, imag} */,
  {32'h417a794a, 32'h40e1b230} /* (10, 14, 22) {real, imag} */,
  {32'hc13c7bc3, 32'h3c62e580} /* (10, 14, 21) {real, imag} */,
  {32'h41431bd0, 32'h3fa973f8} /* (10, 14, 20) {real, imag} */,
  {32'hc0bf9eac, 32'h4092f9cf} /* (10, 14, 19) {real, imag} */,
  {32'hc175dc4c, 32'h3f845bb6} /* (10, 14, 18) {real, imag} */,
  {32'hc09ebb90, 32'h407ca7f7} /* (10, 14, 17) {real, imag} */,
  {32'hc1229c90, 32'hbfcbee20} /* (10, 14, 16) {real, imag} */,
  {32'hc0c89a27, 32'hc1110f98} /* (10, 14, 15) {real, imag} */,
  {32'hc1a69095, 32'h410886d4} /* (10, 14, 14) {real, imag} */,
  {32'hbfa475ec, 32'hc0e19900} /* (10, 14, 13) {real, imag} */,
  {32'hc0802586, 32'hc09a33f8} /* (10, 14, 12) {real, imag} */,
  {32'hc10282fd, 32'h41335619} /* (10, 14, 11) {real, imag} */,
  {32'hbfdcc1ac, 32'h40c935a2} /* (10, 14, 10) {real, imag} */,
  {32'h409cb73e, 32'hc0e70cf2} /* (10, 14, 9) {real, imag} */,
  {32'h3fa314e8, 32'h3eab1246} /* (10, 14, 8) {real, imag} */,
  {32'h3f8c5564, 32'h40e7fa78} /* (10, 14, 7) {real, imag} */,
  {32'hc10fb9c9, 32'h4169e6c8} /* (10, 14, 6) {real, imag} */,
  {32'hc14c9a3d, 32'h40627354} /* (10, 14, 5) {real, imag} */,
  {32'hc0e4ea3c, 32'hc07b6aad} /* (10, 14, 4) {real, imag} */,
  {32'h406fd0c1, 32'h40f3f306} /* (10, 14, 3) {real, imag} */,
  {32'hc160aa65, 32'h4112c846} /* (10, 14, 2) {real, imag} */,
  {32'hc0cb93d4, 32'hc1384052} /* (10, 14, 1) {real, imag} */,
  {32'h40b817ae, 32'h3d3f4500} /* (10, 14, 0) {real, imag} */,
  {32'h408747f5, 32'hc06f4240} /* (10, 13, 31) {real, imag} */,
  {32'h41228d1b, 32'h4014a478} /* (10, 13, 30) {real, imag} */,
  {32'hc03ae008, 32'hc147b4ee} /* (10, 13, 29) {real, imag} */,
  {32'hc1ab81e9, 32'h40ae1866} /* (10, 13, 28) {real, imag} */,
  {32'hbf194300, 32'hbede28a0} /* (10, 13, 27) {real, imag} */,
  {32'hc1132130, 32'hc1219e85} /* (10, 13, 26) {real, imag} */,
  {32'h411dead6, 32'h40090416} /* (10, 13, 25) {real, imag} */,
  {32'h418111f8, 32'hc10cf746} /* (10, 13, 24) {real, imag} */,
  {32'hc01cc818, 32'h40d4d5bc} /* (10, 13, 23) {real, imag} */,
  {32'hc0e22446, 32'h4148f396} /* (10, 13, 22) {real, imag} */,
  {32'h411cd426, 32'hc1193716} /* (10, 13, 21) {real, imag} */,
  {32'hc1969dd6, 32'hc095e2fa} /* (10, 13, 20) {real, imag} */,
  {32'h3ecaf8c0, 32'h417c77d8} /* (10, 13, 19) {real, imag} */,
  {32'hc0cc3f0a, 32'hc0569af3} /* (10, 13, 18) {real, imag} */,
  {32'h405edb84, 32'hc18ae738} /* (10, 13, 17) {real, imag} */,
  {32'h40af03d6, 32'hc07c8cda} /* (10, 13, 16) {real, imag} */,
  {32'hc08c162a, 32'h407a210e} /* (10, 13, 15) {real, imag} */,
  {32'h41680b84, 32'h3fbaedd6} /* (10, 13, 14) {real, imag} */,
  {32'h4154107a, 32'h412d62a8} /* (10, 13, 13) {real, imag} */,
  {32'hc116b404, 32'h41c20a74} /* (10, 13, 12) {real, imag} */,
  {32'hc0f896e7, 32'hbff89f4c} /* (10, 13, 11) {real, imag} */,
  {32'h40df9149, 32'h4118da90} /* (10, 13, 10) {real, imag} */,
  {32'hc1b660cc, 32'hbf1663b0} /* (10, 13, 9) {real, imag} */,
  {32'hc0340354, 32'hc10d177e} /* (10, 13, 8) {real, imag} */,
  {32'hc1ac7dc0, 32'h3f73c0ca} /* (10, 13, 7) {real, imag} */,
  {32'h419c23d8, 32'hc0c505f7} /* (10, 13, 6) {real, imag} */,
  {32'h40c99f61, 32'h3f9af158} /* (10, 13, 5) {real, imag} */,
  {32'hc12e5727, 32'h4019a04c} /* (10, 13, 4) {real, imag} */,
  {32'hc12d8fbf, 32'hc0f2091a} /* (10, 13, 3) {real, imag} */,
  {32'hbe8a9490, 32'h4065422e} /* (10, 13, 2) {real, imag} */,
  {32'h40b23490, 32'h41663914} /* (10, 13, 1) {real, imag} */,
  {32'hc107d3e4, 32'hc0861249} /* (10, 13, 0) {real, imag} */,
  {32'h400bf65c, 32'hc07497fc} /* (10, 12, 31) {real, imag} */,
  {32'hbfaea8d4, 32'hc0a095f6} /* (10, 12, 30) {real, imag} */,
  {32'hc05af31c, 32'h40efe81a} /* (10, 12, 29) {real, imag} */,
  {32'h4198d651, 32'h4160cd8e} /* (10, 12, 28) {real, imag} */,
  {32'hc1798fe0, 32'h3fa95612} /* (10, 12, 27) {real, imag} */,
  {32'h3f10fbce, 32'h400159b1} /* (10, 12, 26) {real, imag} */,
  {32'h3d4f3c00, 32'hc10f4533} /* (10, 12, 25) {real, imag} */,
  {32'hc1b2548e, 32'hc190ad5c} /* (10, 12, 24) {real, imag} */,
  {32'hc1676069, 32'h40af3fc4} /* (10, 12, 23) {real, imag} */,
  {32'hc0875636, 32'h41995dfc} /* (10, 12, 22) {real, imag} */,
  {32'hc0b25d14, 32'h4196fb79} /* (10, 12, 21) {real, imag} */,
  {32'h4152590b, 32'hc15ba271} /* (10, 12, 20) {real, imag} */,
  {32'h414c2470, 32'h3ef779b0} /* (10, 12, 19) {real, imag} */,
  {32'h41afb95c, 32'h41592250} /* (10, 12, 18) {real, imag} */,
  {32'h419ab58a, 32'hc0a96599} /* (10, 12, 17) {real, imag} */,
  {32'h40b54b75, 32'hc165d598} /* (10, 12, 16) {real, imag} */,
  {32'hbf0172fa, 32'h40d9c364} /* (10, 12, 15) {real, imag} */,
  {32'hbf1c8914, 32'h3e475dc0} /* (10, 12, 14) {real, imag} */,
  {32'h40ba8f47, 32'h402021fe} /* (10, 12, 13) {real, imag} */,
  {32'h40f5f3a3, 32'h41eced0c} /* (10, 12, 12) {real, imag} */,
  {32'h413733ec, 32'hc111b54c} /* (10, 12, 11) {real, imag} */,
  {32'h403f504a, 32'h418adf40} /* (10, 12, 10) {real, imag} */,
  {32'hc0af8391, 32'hc12e4d25} /* (10, 12, 9) {real, imag} */,
  {32'h413def97, 32'hc127fe78} /* (10, 12, 8) {real, imag} */,
  {32'h405d3a60, 32'hbfb5a350} /* (10, 12, 7) {real, imag} */,
  {32'hc093d743, 32'h411b6d45} /* (10, 12, 6) {real, imag} */,
  {32'h3fb58808, 32'h409997ae} /* (10, 12, 5) {real, imag} */,
  {32'h3fe26a58, 32'hbe6f53c0} /* (10, 12, 4) {real, imag} */,
  {32'h3d00cbc0, 32'hbf7db7b8} /* (10, 12, 3) {real, imag} */,
  {32'h409e5fac, 32'h3fa73846} /* (10, 12, 2) {real, imag} */,
  {32'h3fb63077, 32'hc1317e1a} /* (10, 12, 1) {real, imag} */,
  {32'h4168350e, 32'hc00c8508} /* (10, 12, 0) {real, imag} */,
  {32'hc1b54e9f, 32'hc1d6649e} /* (10, 11, 31) {real, imag} */,
  {32'h41886ff5, 32'hc150a396} /* (10, 11, 30) {real, imag} */,
  {32'h40870ad0, 32'h40c82455} /* (10, 11, 29) {real, imag} */,
  {32'hc0ed3def, 32'h411922e0} /* (10, 11, 28) {real, imag} */,
  {32'hc098f5cc, 32'h41bb91f0} /* (10, 11, 27) {real, imag} */,
  {32'h3ffda398, 32'hc1495140} /* (10, 11, 26) {real, imag} */,
  {32'h3f6adecc, 32'hc01e0f44} /* (10, 11, 25) {real, imag} */,
  {32'h4122f08e, 32'hc0e9b0ca} /* (10, 11, 24) {real, imag} */,
  {32'hc04bd6b4, 32'hc1459990} /* (10, 11, 23) {real, imag} */,
  {32'hc0b53044, 32'hc11066e5} /* (10, 11, 22) {real, imag} */,
  {32'hc03c2e66, 32'hc040431c} /* (10, 11, 21) {real, imag} */,
  {32'hc0ce49e6, 32'h3fa90bbc} /* (10, 11, 20) {real, imag} */,
  {32'h410fb54c, 32'hc12d9d10} /* (10, 11, 19) {real, imag} */,
  {32'h3fe16fd0, 32'h40d51636} /* (10, 11, 18) {real, imag} */,
  {32'hbfa14410, 32'h400fefb8} /* (10, 11, 17) {real, imag} */,
  {32'h3fde7fe8, 32'hc0af9a24} /* (10, 11, 16) {real, imag} */,
  {32'hbf8cab43, 32'hc08a2d41} /* (10, 11, 15) {real, imag} */,
  {32'hbf694eb0, 32'h40c48978} /* (10, 11, 14) {real, imag} */,
  {32'h4103ec10, 32'h401fe034} /* (10, 11, 13) {real, imag} */,
  {32'h40e7de01, 32'hc0429630} /* (10, 11, 12) {real, imag} */,
  {32'h40073354, 32'hc157ca2c} /* (10, 11, 11) {real, imag} */,
  {32'h40a2dfa0, 32'h416ba651} /* (10, 11, 10) {real, imag} */,
  {32'h3fe526d8, 32'h407e96a8} /* (10, 11, 9) {real, imag} */,
  {32'hc04b67e1, 32'h408cbced} /* (10, 11, 8) {real, imag} */,
  {32'h413a55ca, 32'hbda46ec0} /* (10, 11, 7) {real, imag} */,
  {32'hc1433582, 32'h3e99f688} /* (10, 11, 6) {real, imag} */,
  {32'hc09ff534, 32'hc0a80f58} /* (10, 11, 5) {real, imag} */,
  {32'hc09f56df, 32'h3fca6b50} /* (10, 11, 4) {real, imag} */,
  {32'h41093868, 32'hc15120c0} /* (10, 11, 3) {real, imag} */,
  {32'h414dcae8, 32'h41ea414a} /* (10, 11, 2) {real, imag} */,
  {32'h405d58c0, 32'hc1e19644} /* (10, 11, 1) {real, imag} */,
  {32'hc10117b3, 32'hc11bf5fa} /* (10, 11, 0) {real, imag} */,
  {32'h415d45b6, 32'h41bacea2} /* (10, 10, 31) {real, imag} */,
  {32'hc182c7f1, 32'hc12b0303} /* (10, 10, 30) {real, imag} */,
  {32'hc18609a1, 32'h418f223e} /* (10, 10, 29) {real, imag} */,
  {32'hc157ba32, 32'hc15cc7e4} /* (10, 10, 28) {real, imag} */,
  {32'h41263e9d, 32'hbf7eaff0} /* (10, 10, 27) {real, imag} */,
  {32'hc123ff92, 32'h4048b41c} /* (10, 10, 26) {real, imag} */,
  {32'hc1826acb, 32'hc08b28e0} /* (10, 10, 25) {real, imag} */,
  {32'h3f52c518, 32'h415996de} /* (10, 10, 24) {real, imag} */,
  {32'h421a1203, 32'hc1a2080c} /* (10, 10, 23) {real, imag} */,
  {32'h418e6c07, 32'h40edadd4} /* (10, 10, 22) {real, imag} */,
  {32'hbf6dc230, 32'h40132a68} /* (10, 10, 21) {real, imag} */,
  {32'hc0dbbeca, 32'hc1246791} /* (10, 10, 20) {real, imag} */,
  {32'hc1c98cd9, 32'h4091347f} /* (10, 10, 19) {real, imag} */,
  {32'hc13bf96e, 32'h4173cac3} /* (10, 10, 18) {real, imag} */,
  {32'h405ec206, 32'h40d138ca} /* (10, 10, 17) {real, imag} */,
  {32'h41168a7a, 32'h3f2d6051} /* (10, 10, 16) {real, imag} */,
  {32'hc0994ae7, 32'hc017c988} /* (10, 10, 15) {real, imag} */,
  {32'hc1161929, 32'hc1a87432} /* (10, 10, 14) {real, imag} */,
  {32'h409003ce, 32'h4105c85e} /* (10, 10, 13) {real, imag} */,
  {32'h3f891e00, 32'hc04a9fc3} /* (10, 10, 12) {real, imag} */,
  {32'hbee3c410, 32'h3e80e9b0} /* (10, 10, 11) {real, imag} */,
  {32'hc190f4c0, 32'h4110c952} /* (10, 10, 10) {real, imag} */,
  {32'hbf005a22, 32'h41581694} /* (10, 10, 9) {real, imag} */,
  {32'h412e088a, 32'h40cf30ef} /* (10, 10, 8) {real, imag} */,
  {32'hc0d804ea, 32'hc0bea2dc} /* (10, 10, 7) {real, imag} */,
  {32'h40283776, 32'h41f67f42} /* (10, 10, 6) {real, imag} */,
  {32'hc02b4a98, 32'h40d7adaa} /* (10, 10, 5) {real, imag} */,
  {32'h401825ee, 32'h3e9b75d0} /* (10, 10, 4) {real, imag} */,
  {32'h418d75af, 32'h41068f18} /* (10, 10, 3) {real, imag} */,
  {32'h413895e7, 32'hc0993912} /* (10, 10, 2) {real, imag} */,
  {32'h40d9c25e, 32'hc1908b20} /* (10, 10, 1) {real, imag} */,
  {32'h40e13321, 32'hc14b08e4} /* (10, 10, 0) {real, imag} */,
  {32'hc0e5a079, 32'h415b8d0e} /* (10, 9, 31) {real, imag} */,
  {32'h401dce12, 32'hc09385a6} /* (10, 9, 30) {real, imag} */,
  {32'h403fb233, 32'h418e6b00} /* (10, 9, 29) {real, imag} */,
  {32'h4194934c, 32'hc1829b66} /* (10, 9, 28) {real, imag} */,
  {32'h418f3cf5, 32'hc167d96e} /* (10, 9, 27) {real, imag} */,
  {32'hbf7179d0, 32'h405685ff} /* (10, 9, 26) {real, imag} */,
  {32'hc12dcd50, 32'h418190c1} /* (10, 9, 25) {real, imag} */,
  {32'hbf96f18c, 32'hc0b60382} /* (10, 9, 24) {real, imag} */,
  {32'h4011e82e, 32'h414f8337} /* (10, 9, 23) {real, imag} */,
  {32'hc19427e9, 32'h4102f0e6} /* (10, 9, 22) {real, imag} */,
  {32'hc0053802, 32'hbf236c64} /* (10, 9, 21) {real, imag} */,
  {32'h40c9da7e, 32'hc10c08d7} /* (10, 9, 20) {real, imag} */,
  {32'h406b7ec2, 32'hc10cd24a} /* (10, 9, 19) {real, imag} */,
  {32'h3fccee5c, 32'hc1312e48} /* (10, 9, 18) {real, imag} */,
  {32'hc1282b3c, 32'h41823df6} /* (10, 9, 17) {real, imag} */,
  {32'h40879d7f, 32'h407dba8f} /* (10, 9, 16) {real, imag} */,
  {32'hbf2f4150, 32'h412f4e2e} /* (10, 9, 15) {real, imag} */,
  {32'hc03635f4, 32'hc03c833a} /* (10, 9, 14) {real, imag} */,
  {32'h4061e7b6, 32'hc11fb2e6} /* (10, 9, 13) {real, imag} */,
  {32'hc145b78c, 32'h405e6720} /* (10, 9, 12) {real, imag} */,
  {32'h41472496, 32'hc0abf07f} /* (10, 9, 11) {real, imag} */,
  {32'h40d73946, 32'hc131deb1} /* (10, 9, 10) {real, imag} */,
  {32'hbf729870, 32'hc0887d20} /* (10, 9, 9) {real, imag} */,
  {32'hc135bec8, 32'h41009cb6} /* (10, 9, 8) {real, imag} */,
  {32'hc1122fa2, 32'h414efc3d} /* (10, 9, 7) {real, imag} */,
  {32'h41689094, 32'hc0dc2979} /* (10, 9, 6) {real, imag} */,
  {32'hc1d22072, 32'h4157c20d} /* (10, 9, 5) {real, imag} */,
  {32'hc186fc80, 32'hc0a9addd} /* (10, 9, 4) {real, imag} */,
  {32'h415da0d6, 32'h40cf3848} /* (10, 9, 3) {real, imag} */,
  {32'h411e96bb, 32'hbf4981d0} /* (10, 9, 2) {real, imag} */,
  {32'hc12d7b7c, 32'h40bde6b8} /* (10, 9, 1) {real, imag} */,
  {32'h40b517b8, 32'h40d6c3dc} /* (10, 9, 0) {real, imag} */,
  {32'hc2324ca9, 32'hc115a032} /* (10, 8, 31) {real, imag} */,
  {32'h41d18910, 32'hc0d37ba4} /* (10, 8, 30) {real, imag} */,
  {32'hc1cfcd71, 32'hc131a35c} /* (10, 8, 29) {real, imag} */,
  {32'h4014b4e0, 32'h416822cc} /* (10, 8, 28) {real, imag} */,
  {32'h4123aa99, 32'h41a579c8} /* (10, 8, 27) {real, imag} */,
  {32'hc0baa38a, 32'h3e681530} /* (10, 8, 26) {real, imag} */,
  {32'h40e6b0ee, 32'hc09f6f35} /* (10, 8, 25) {real, imag} */,
  {32'h40ebd6da, 32'h402cd5d8} /* (10, 8, 24) {real, imag} */,
  {32'h3c402e00, 32'hc09fece4} /* (10, 8, 23) {real, imag} */,
  {32'h412944f4, 32'h41822d24} /* (10, 8, 22) {real, imag} */,
  {32'hc1c3b31c, 32'h414361e6} /* (10, 8, 21) {real, imag} */,
  {32'hc0ceebb0, 32'h417d0eab} /* (10, 8, 20) {real, imag} */,
  {32'h40af29d7, 32'hc0a352b2} /* (10, 8, 19) {real, imag} */,
  {32'h40daee5c, 32'hbf8d43ac} /* (10, 8, 18) {real, imag} */,
  {32'h3dda7270, 32'hc04904d4} /* (10, 8, 17) {real, imag} */,
  {32'h40c4da08, 32'h4018bed6} /* (10, 8, 16) {real, imag} */,
  {32'hc0c97abf, 32'hbf43a9f2} /* (10, 8, 15) {real, imag} */,
  {32'h40df11f0, 32'hc10ae8e6} /* (10, 8, 14) {real, imag} */,
  {32'hc1888a74, 32'h404a7901} /* (10, 8, 13) {real, imag} */,
  {32'h4171e022, 32'h3ec96a18} /* (10, 8, 12) {real, imag} */,
  {32'h41007f1a, 32'h40be2169} /* (10, 8, 11) {real, imag} */,
  {32'h40b573bc, 32'h410ba8b5} /* (10, 8, 10) {real, imag} */,
  {32'hc138d2d8, 32'h413c13a2} /* (10, 8, 9) {real, imag} */,
  {32'h40e87609, 32'h401fe71c} /* (10, 8, 8) {real, imag} */,
  {32'h41d2ab84, 32'h40f806b1} /* (10, 8, 7) {real, imag} */,
  {32'h413d43ec, 32'h40c6fdc7} /* (10, 8, 6) {real, imag} */,
  {32'h41545845, 32'hc132d86a} /* (10, 8, 5) {real, imag} */,
  {32'hc198bc52, 32'hbfcfee58} /* (10, 8, 4) {real, imag} */,
  {32'hbfe9c1f0, 32'h40044dea} /* (10, 8, 3) {real, imag} */,
  {32'h41e6be6d, 32'h41210aa6} /* (10, 8, 2) {real, imag} */,
  {32'hc1ad2c34, 32'hc1a0f196} /* (10, 8, 1) {real, imag} */,
  {32'hc0f07ef0, 32'hc00f89fc} /* (10, 8, 0) {real, imag} */,
  {32'h41b45426, 32'h41b3471e} /* (10, 7, 31) {real, imag} */,
  {32'hc14bf404, 32'hc1cc03fe} /* (10, 7, 30) {real, imag} */,
  {32'hc1c36b20, 32'h41ff86b0} /* (10, 7, 29) {real, imag} */,
  {32'h3fe60260, 32'h40fd965e} /* (10, 7, 28) {real, imag} */,
  {32'hc10c15e7, 32'h40b1358c} /* (10, 7, 27) {real, imag} */,
  {32'h3f9aec8c, 32'h3ed979c0} /* (10, 7, 26) {real, imag} */,
  {32'h40f63c32, 32'hc11856da} /* (10, 7, 25) {real, imag} */,
  {32'hc1a46fb4, 32'h4021a142} /* (10, 7, 24) {real, imag} */,
  {32'hc186f702, 32'hc169e925} /* (10, 7, 23) {real, imag} */,
  {32'h40ba942b, 32'hc003dab0} /* (10, 7, 22) {real, imag} */,
  {32'h415bf115, 32'h40dc1bf8} /* (10, 7, 21) {real, imag} */,
  {32'hc184d64e, 32'hc114327a} /* (10, 7, 20) {real, imag} */,
  {32'h4114a0c8, 32'hbefd6268} /* (10, 7, 19) {real, imag} */,
  {32'h408dbfbd, 32'h3f85f2dc} /* (10, 7, 18) {real, imag} */,
  {32'hc11373db, 32'h3f2716b4} /* (10, 7, 17) {real, imag} */,
  {32'h40ac5d66, 32'h409f3b01} /* (10, 7, 16) {real, imag} */,
  {32'hc0649754, 32'h4042f983} /* (10, 7, 15) {real, imag} */,
  {32'hc0af21c1, 32'h40b7241a} /* (10, 7, 14) {real, imag} */,
  {32'hc091c783, 32'h418c4352} /* (10, 7, 13) {real, imag} */,
  {32'hc04daff6, 32'hc0f992ea} /* (10, 7, 12) {real, imag} */,
  {32'h41047a21, 32'h4008cd62} /* (10, 7, 11) {real, imag} */,
  {32'hc1112bac, 32'hc18bc44e} /* (10, 7, 10) {real, imag} */,
  {32'h40f8411d, 32'h40eb41af} /* (10, 7, 9) {real, imag} */,
  {32'hc0ea2445, 32'hc078ea24} /* (10, 7, 8) {real, imag} */,
  {32'h3f23ec04, 32'h40ca5ba0} /* (10, 7, 7) {real, imag} */,
  {32'h41ad079d, 32'hc147d92e} /* (10, 7, 6) {real, imag} */,
  {32'hc13c49d7, 32'hc1734e13} /* (10, 7, 5) {real, imag} */,
  {32'h41099ee6, 32'hbfd119ac} /* (10, 7, 4) {real, imag} */,
  {32'h40ad01ea, 32'h3f1be220} /* (10, 7, 3) {real, imag} */,
  {32'hc1ef7fec, 32'h40afa876} /* (10, 7, 2) {real, imag} */,
  {32'h4111935c, 32'h42049c11} /* (10, 7, 1) {real, imag} */,
  {32'h409304cd, 32'hc0d6311a} /* (10, 7, 0) {real, imag} */,
  {32'h40d830fb, 32'hc1efaceb} /* (10, 6, 31) {real, imag} */,
  {32'h40b3ca98, 32'hc1979fa5} /* (10, 6, 30) {real, imag} */,
  {32'h413775b0, 32'h40e30794} /* (10, 6, 29) {real, imag} */,
  {32'h41855990, 32'hc1745ae2} /* (10, 6, 28) {real, imag} */,
  {32'hc0734e34, 32'hc1826ce0} /* (10, 6, 27) {real, imag} */,
  {32'h418ce352, 32'hc0480454} /* (10, 6, 26) {real, imag} */,
  {32'h4069f31a, 32'h3fbea0aa} /* (10, 6, 25) {real, imag} */,
  {32'hc18733ec, 32'hc01e231a} /* (10, 6, 24) {real, imag} */,
  {32'h419723af, 32'h41baa62b} /* (10, 6, 23) {real, imag} */,
  {32'hc149291f, 32'hc11e04d6} /* (10, 6, 22) {real, imag} */,
  {32'h4184eafa, 32'h4047a064} /* (10, 6, 21) {real, imag} */,
  {32'h40b07835, 32'hc02cd542} /* (10, 6, 20) {real, imag} */,
  {32'h407485ac, 32'h410f34d3} /* (10, 6, 19) {real, imag} */,
  {32'h415c0d4e, 32'h40a28c80} /* (10, 6, 18) {real, imag} */,
  {32'hc0cf61ad, 32'h41307e25} /* (10, 6, 17) {real, imag} */,
  {32'hc0ce252f, 32'h40b410c8} /* (10, 6, 16) {real, imag} */,
  {32'hc10d7742, 32'hc124c742} /* (10, 6, 15) {real, imag} */,
  {32'h40960ce0, 32'h4098a832} /* (10, 6, 14) {real, imag} */,
  {32'h40d75e53, 32'h3e985e58} /* (10, 6, 13) {real, imag} */,
  {32'h40bc5ec8, 32'h3fb5c8d8} /* (10, 6, 12) {real, imag} */,
  {32'hbfc15018, 32'hc03b5f55} /* (10, 6, 11) {real, imag} */,
  {32'hc12864fe, 32'hc18a5a38} /* (10, 6, 10) {real, imag} */,
  {32'hc0d75db9, 32'hc12da22c} /* (10, 6, 9) {real, imag} */,
  {32'h4132085c, 32'hc14d03a0} /* (10, 6, 8) {real, imag} */,
  {32'h40db68c6, 32'h3f1a1a74} /* (10, 6, 7) {real, imag} */,
  {32'h41080f86, 32'h40f865d0} /* (10, 6, 6) {real, imag} */,
  {32'h41751b72, 32'h4190de38} /* (10, 6, 5) {real, imag} */,
  {32'hc170f791, 32'h40adc047} /* (10, 6, 4) {real, imag} */,
  {32'hc18660e2, 32'h4119004f} /* (10, 6, 3) {real, imag} */,
  {32'h40b40756, 32'hc1e53a70} /* (10, 6, 2) {real, imag} */,
  {32'h4092ea6f, 32'h4060ba35} /* (10, 6, 1) {real, imag} */,
  {32'h41769ea5, 32'h42090978} /* (10, 6, 0) {real, imag} */,
  {32'hc2eabc8a, 32'hc20d0e4b} /* (10, 5, 31) {real, imag} */,
  {32'h41a62202, 32'h3fb336e4} /* (10, 5, 30) {real, imag} */,
  {32'h40e32c50, 32'hc0ae0a9c} /* (10, 5, 29) {real, imag} */,
  {32'hc198c64c, 32'h4224a9bc} /* (10, 5, 28) {real, imag} */,
  {32'hbf2065c0, 32'h41889e1a} /* (10, 5, 27) {real, imag} */,
  {32'h3f96d8a6, 32'hc0accbba} /* (10, 5, 26) {real, imag} */,
  {32'hc10b137d, 32'h412aa6b6} /* (10, 5, 25) {real, imag} */,
  {32'hc0fd51ed, 32'hc1ce30a1} /* (10, 5, 24) {real, imag} */,
  {32'hc0fc6160, 32'h41abe7ec} /* (10, 5, 23) {real, imag} */,
  {32'hbf708d80, 32'hc186e724} /* (10, 5, 22) {real, imag} */,
  {32'h413941ec, 32'hc18fbac8} /* (10, 5, 21) {real, imag} */,
  {32'h3f4b6310, 32'hc0889820} /* (10, 5, 20) {real, imag} */,
  {32'hc0a51228, 32'hc1147946} /* (10, 5, 19) {real, imag} */,
  {32'hc1346b8a, 32'hc188a1de} /* (10, 5, 18) {real, imag} */,
  {32'h40072c74, 32'hc14ef872} /* (10, 5, 17) {real, imag} */,
  {32'hc1365de8, 32'hbe7428e0} /* (10, 5, 16) {real, imag} */,
  {32'hc14c0665, 32'h4138def2} /* (10, 5, 15) {real, imag} */,
  {32'h3fd0c5a8, 32'h418303a3} /* (10, 5, 14) {real, imag} */,
  {32'h41704e62, 32'h4045caa6} /* (10, 5, 13) {real, imag} */,
  {32'h41304136, 32'hbf558a98} /* (10, 5, 12) {real, imag} */,
  {32'hc13e69ec, 32'hc03b47d4} /* (10, 5, 11) {real, imag} */,
  {32'hc04c3ce4, 32'h40f836f4} /* (10, 5, 10) {real, imag} */,
  {32'h408065c7, 32'hbfcb01ae} /* (10, 5, 9) {real, imag} */,
  {32'h4093ef7c, 32'h41a614c8} /* (10, 5, 8) {real, imag} */,
  {32'h40e1c7d1, 32'hc16cdcec} /* (10, 5, 7) {real, imag} */,
  {32'hc142a20a, 32'h40b6320f} /* (10, 5, 6) {real, imag} */,
  {32'h416b48f2, 32'h404a52fc} /* (10, 5, 5) {real, imag} */,
  {32'hc1498c26, 32'hc06c0e60} /* (10, 5, 4) {real, imag} */,
  {32'hbf8781a6, 32'h40e7cf3e} /* (10, 5, 3) {real, imag} */,
  {32'h40b58d21, 32'h424f3922} /* (10, 5, 2) {real, imag} */,
  {32'hc1b97270, 32'hc296f74f} /* (10, 5, 1) {real, imag} */,
  {32'hc27fea3c, 32'hc1af539a} /* (10, 5, 0) {real, imag} */,
  {32'h424fee04, 32'h42c31e08} /* (10, 4, 31) {real, imag} */,
  {32'hc2d31cbd, 32'hc25e677d} /* (10, 4, 30) {real, imag} */,
  {32'hc122bd6f, 32'hc11e0276} /* (10, 4, 29) {real, imag} */,
  {32'h41d9b136, 32'hbf9431c0} /* (10, 4, 28) {real, imag} */,
  {32'hc1bdf03a, 32'hc0374726} /* (10, 4, 27) {real, imag} */,
  {32'hc1c2a438, 32'h41f64a91} /* (10, 4, 26) {real, imag} */,
  {32'h418a8bbe, 32'hc12248d0} /* (10, 4, 25) {real, imag} */,
  {32'h40fa51c2, 32'hc1b2c919} /* (10, 4, 24) {real, imag} */,
  {32'h42018976, 32'h402a7794} /* (10, 4, 23) {real, imag} */,
  {32'hbffcab1e, 32'hc14c7819} /* (10, 4, 22) {real, imag} */,
  {32'h401a743e, 32'hc1484bda} /* (10, 4, 21) {real, imag} */,
  {32'hbfa6e504, 32'h40a2caea} /* (10, 4, 20) {real, imag} */,
  {32'hc022d4be, 32'h407e574f} /* (10, 4, 19) {real, imag} */,
  {32'hc17985ac, 32'hc0d4fb4d} /* (10, 4, 18) {real, imag} */,
  {32'hbf694099, 32'h411789d1} /* (10, 4, 17) {real, imag} */,
  {32'hc0c12340, 32'h40be4c8e} /* (10, 4, 16) {real, imag} */,
  {32'hc1715748, 32'h4042e7de} /* (10, 4, 15) {real, imag} */,
  {32'h414b1034, 32'hc0d1dd42} /* (10, 4, 14) {real, imag} */,
  {32'h41198148, 32'hc0b5d58a} /* (10, 4, 13) {real, imag} */,
  {32'hbfd5ee12, 32'h4100befa} /* (10, 4, 12) {real, imag} */,
  {32'h412d264f, 32'hc1a4f36a} /* (10, 4, 11) {real, imag} */,
  {32'h40c785c2, 32'h40b6f94a} /* (10, 4, 10) {real, imag} */,
  {32'h4128f3dc, 32'h3f46fc50} /* (10, 4, 9) {real, imag} */,
  {32'hc0fa4f8a, 32'hc195bba6} /* (10, 4, 8) {real, imag} */,
  {32'hc08ea97a, 32'hc170f572} /* (10, 4, 7) {real, imag} */,
  {32'hc10e99b2, 32'h40f08c46} /* (10, 4, 6) {real, imag} */,
  {32'h41bb4502, 32'hc1ea884e} /* (10, 4, 5) {real, imag} */,
  {32'h4103c62a, 32'h422d6279} /* (10, 4, 4) {real, imag} */,
  {32'hc1be0e15, 32'h41c8c00c} /* (10, 4, 3) {real, imag} */,
  {32'hc2723e65, 32'hc2867505} /* (10, 4, 2) {real, imag} */,
  {32'h4320d659, 32'h41f4a87c} /* (10, 4, 1) {real, imag} */,
  {32'h420e4851, 32'h41c8d2d6} /* (10, 4, 0) {real, imag} */,
  {32'hc3132d8f, 32'h42969b15} /* (10, 3, 31) {real, imag} */,
  {32'h428616b9, 32'hc306af0b} /* (10, 3, 30) {real, imag} */,
  {32'hc18d50d6, 32'hc16aafbd} /* (10, 3, 29) {real, imag} */,
  {32'h426266e6, 32'h41f1744a} /* (10, 3, 28) {real, imag} */,
  {32'hc2250c8d, 32'h4118a6f2} /* (10, 3, 27) {real, imag} */,
  {32'h4110f1bc, 32'h414cc7d7} /* (10, 3, 26) {real, imag} */,
  {32'hc02912a0, 32'h414d37e6} /* (10, 3, 25) {real, imag} */,
  {32'h414fb88f, 32'h3f1aa348} /* (10, 3, 24) {real, imag} */,
  {32'hc125ea66, 32'h3ff8f1ec} /* (10, 3, 23) {real, imag} */,
  {32'hc1cfb06f, 32'hc101a298} /* (10, 3, 22) {real, imag} */,
  {32'h4085c79c, 32'h414b789a} /* (10, 3, 21) {real, imag} */,
  {32'hc0c069a9, 32'hc063beb6} /* (10, 3, 20) {real, imag} */,
  {32'hc050782a, 32'h408ed0de} /* (10, 3, 19) {real, imag} */,
  {32'h3e3f6c60, 32'hc0e61e3c} /* (10, 3, 18) {real, imag} */,
  {32'h40f8e119, 32'hc127a2b7} /* (10, 3, 17) {real, imag} */,
  {32'h4100181d, 32'hc1235781} /* (10, 3, 16) {real, imag} */,
  {32'h414e35d1, 32'hc077aef0} /* (10, 3, 15) {real, imag} */,
  {32'h4037676e, 32'hc183083f} /* (10, 3, 14) {real, imag} */,
  {32'hc0793449, 32'hc1023aba} /* (10, 3, 13) {real, imag} */,
  {32'h4102f34d, 32'hc1744d4e} /* (10, 3, 12) {real, imag} */,
  {32'h40c6ee46, 32'h411d725a} /* (10, 3, 11) {real, imag} */,
  {32'h4143d934, 32'h418a43c2} /* (10, 3, 10) {real, imag} */,
  {32'h40b0e5d8, 32'hc0a71cfc} /* (10, 3, 9) {real, imag} */,
  {32'hc0a8a9cd, 32'h414d286b} /* (10, 3, 8) {real, imag} */,
  {32'hc1b941ad, 32'h405b583a} /* (10, 3, 7) {real, imag} */,
  {32'hc0931ff0, 32'hc028e1e6} /* (10, 3, 6) {real, imag} */,
  {32'hc1641416, 32'h40a3e9b0} /* (10, 3, 5) {real, imag} */,
  {32'hc2008b65, 32'h41421998} /* (10, 3, 4) {real, imag} */,
  {32'hc1e2777a, 32'h41bf6ded} /* (10, 3, 3) {real, imag} */,
  {32'hc109bafa, 32'hc2bcc3f5} /* (10, 3, 2) {real, imag} */,
  {32'h42e2072d, 32'h42af14e8} /* (10, 3, 1) {real, imag} */,
  {32'hc18b8942, 32'h4153d01e} /* (10, 3, 0) {real, imag} */,
  {32'hc4a5fe8d, 32'hc29c5516} /* (10, 2, 31) {real, imag} */,
  {32'h441603b2, 32'hc3375182} /* (10, 2, 30) {real, imag} */,
  {32'h421c33fc, 32'h4179fe47} /* (10, 2, 29) {real, imag} */,
  {32'hc1d745ae, 32'h4297b2b2} /* (10, 2, 28) {real, imag} */,
  {32'h426cdb99, 32'hc283366a} /* (10, 2, 27) {real, imag} */,
  {32'h415b121c, 32'hc131844a} /* (10, 2, 26) {real, imag} */,
  {32'hbfceed28, 32'h4104b9c6} /* (10, 2, 25) {real, imag} */,
  {32'h41ffbe08, 32'hc1be5976} /* (10, 2, 24) {real, imag} */,
  {32'hc159558d, 32'h417da11c} /* (10, 2, 23) {real, imag} */,
  {32'hc1be6041, 32'hc06e3dcc} /* (10, 2, 22) {real, imag} */,
  {32'h41025ba0, 32'hc1cd0b2e} /* (10, 2, 21) {real, imag} */,
  {32'hc0193ade, 32'h4164c944} /* (10, 2, 20) {real, imag} */,
  {32'hc11bee8f, 32'h413b9980} /* (10, 2, 19) {real, imag} */,
  {32'h415c69c6, 32'hbef554c0} /* (10, 2, 18) {real, imag} */,
  {32'hc11f4e31, 32'hc0a609e4} /* (10, 2, 17) {real, imag} */,
  {32'h3fc072d6, 32'hbe8ce4e4} /* (10, 2, 16) {real, imag} */,
  {32'h40b0702c, 32'hc0596098} /* (10, 2, 15) {real, imag} */,
  {32'hc0de5ca0, 32'hc0c7287e} /* (10, 2, 14) {real, imag} */,
  {32'hc1626ec2, 32'hbfcfc3ce} /* (10, 2, 13) {real, imag} */,
  {32'h3eaf0bb0, 32'hc0ba3025} /* (10, 2, 12) {real, imag} */,
  {32'h40765eba, 32'h4174724e} /* (10, 2, 11) {real, imag} */,
  {32'hc105d3ce, 32'hc11270b6} /* (10, 2, 10) {real, imag} */,
  {32'h40a4d237, 32'h4116ef5e} /* (10, 2, 9) {real, imag} */,
  {32'h411e3d37, 32'h415981f6} /* (10, 2, 8) {real, imag} */,
  {32'hc0b0361a, 32'h4090cd6e} /* (10, 2, 7) {real, imag} */,
  {32'h4120cdd9, 32'hc13c4cc4} /* (10, 2, 6) {real, imag} */,
  {32'h41b8be07, 32'h42a4d4b0} /* (10, 2, 5) {real, imag} */,
  {32'hc2da8845, 32'hc2234d5f} /* (10, 2, 4) {real, imag} */,
  {32'h4118f22c, 32'h41bbb3fa} /* (10, 2, 3) {real, imag} */,
  {32'h43d96382, 32'hc2fb0336} /* (10, 2, 2) {real, imag} */,
  {32'hc4396d1f, 32'h43432882} /* (10, 2, 1) {real, imag} */,
  {32'hc43a787e, 32'hc2c83579} /* (10, 2, 0) {real, imag} */,
  {32'h44dbfc61, 32'hc3c114bf} /* (10, 1, 31) {real, imag} */,
  {32'hc3c8ff00, 32'h42835e8e} /* (10, 1, 30) {real, imag} */,
  {32'hc23f9288, 32'hc140efc8} /* (10, 1, 29) {real, imag} */,
  {32'h42a40b94, 32'h42c8fb02} /* (10, 1, 28) {real, imag} */,
  {32'hc2ac58a1, 32'h40b16332} /* (10, 1, 27) {real, imag} */,
  {32'hc0c39d6c, 32'h41a2217c} /* (10, 1, 26) {real, imag} */,
  {32'h419a37d0, 32'hc0bdf30c} /* (10, 1, 25) {real, imag} */,
  {32'hc1417d14, 32'h417e305e} /* (10, 1, 24) {real, imag} */,
  {32'hc145b17c, 32'hc09df8ba} /* (10, 1, 23) {real, imag} */,
  {32'h417baf31, 32'h40e19633} /* (10, 1, 22) {real, imag} */,
  {32'hc1990ec6, 32'h418a5b84} /* (10, 1, 21) {real, imag} */,
  {32'h4000cd76, 32'h41a25556} /* (10, 1, 20) {real, imag} */,
  {32'h412db4a1, 32'hc0c40fd4} /* (10, 1, 19) {real, imag} */,
  {32'hc090a2dc, 32'h419a1f74} /* (10, 1, 18) {real, imag} */,
  {32'h3f91158e, 32'h404c2d37} /* (10, 1, 17) {real, imag} */,
  {32'h40b83cba, 32'h41152a10} /* (10, 1, 16) {real, imag} */,
  {32'h4051caf9, 32'h40732b67} /* (10, 1, 15) {real, imag} */,
  {32'hc1800dfd, 32'hc0859b5b} /* (10, 1, 14) {real, imag} */,
  {32'h400bff88, 32'h405fbd1d} /* (10, 1, 13) {real, imag} */,
  {32'hc0a09591, 32'hc0b3e00a} /* (10, 1, 12) {real, imag} */,
  {32'hc08245ae, 32'hc1812527} /* (10, 1, 11) {real, imag} */,
  {32'hc1b840ff, 32'hc1a64742} /* (10, 1, 10) {real, imag} */,
  {32'h415610f2, 32'h41536679} /* (10, 1, 9) {real, imag} */,
  {32'hc0cb65a5, 32'hc21efba0} /* (10, 1, 8) {real, imag} */,
  {32'h41cbec46, 32'h40585798} /* (10, 1, 7) {real, imag} */,
  {32'hc1f2cde9, 32'hc16495df} /* (10, 1, 6) {real, imag} */,
  {32'hc298ff05, 32'hc22e35bf} /* (10, 1, 5) {real, imag} */,
  {32'h41ee46f0, 32'h4194ad6e} /* (10, 1, 4) {real, imag} */,
  {32'h413a26f6, 32'h418fa254} /* (10, 1, 3) {real, imag} */,
  {32'hc426c6c3, 32'hc41153f9} /* (10, 1, 2) {real, imag} */,
  {32'h451efe91, 32'h44aba8a3} /* (10, 1, 1) {real, imag} */,
  {32'h4513f624, 32'h431af701} /* (10, 1, 0) {real, imag} */,
  {32'h44b62b0a, 32'hc4930090} /* (10, 0, 31) {real, imag} */,
  {32'hc34a9d4c, 32'h43afe09a} /* (10, 0, 30) {real, imag} */,
  {32'hc2817688, 32'h4182c4d1} /* (10, 0, 29) {real, imag} */,
  {32'hc144c8d5, 32'h41cc18e6} /* (10, 0, 28) {real, imag} */,
  {32'hc26dba18, 32'h41dbe344} /* (10, 0, 27) {real, imag} */,
  {32'hbef87650, 32'h40b0d6e8} /* (10, 0, 26) {real, imag} */,
  {32'h41137829, 32'hc155b1c4} /* (10, 0, 25) {real, imag} */,
  {32'hc082dc94, 32'h42126efa} /* (10, 0, 24) {real, imag} */,
  {32'h40d33a04, 32'hc063b507} /* (10, 0, 23) {real, imag} */,
  {32'h4106aa57, 32'h40154caa} /* (10, 0, 22) {real, imag} */,
  {32'h3fcbadf6, 32'h414472e2} /* (10, 0, 21) {real, imag} */,
  {32'hbf8569cc, 32'hbeee6f18} /* (10, 0, 20) {real, imag} */,
  {32'hc074a4ee, 32'hc19b686a} /* (10, 0, 19) {real, imag} */,
  {32'h4058b5f0, 32'hc0cc7708} /* (10, 0, 18) {real, imag} */,
  {32'hbff78be0, 32'h3f9be7bc} /* (10, 0, 17) {real, imag} */,
  {32'hc15a7012, 32'h00000000} /* (10, 0, 16) {real, imag} */,
  {32'hbff78be0, 32'hbf9be7bc} /* (10, 0, 15) {real, imag} */,
  {32'h4058b5f0, 32'h40cc7708} /* (10, 0, 14) {real, imag} */,
  {32'hc074a4ee, 32'h419b686a} /* (10, 0, 13) {real, imag} */,
  {32'hbf8569cc, 32'h3eee6f18} /* (10, 0, 12) {real, imag} */,
  {32'h3fcbadf6, 32'hc14472e2} /* (10, 0, 11) {real, imag} */,
  {32'h4106aa57, 32'hc0154caa} /* (10, 0, 10) {real, imag} */,
  {32'h40d33a04, 32'h4063b507} /* (10, 0, 9) {real, imag} */,
  {32'hc082dc94, 32'hc2126efa} /* (10, 0, 8) {real, imag} */,
  {32'h41137829, 32'h4155b1c4} /* (10, 0, 7) {real, imag} */,
  {32'hbef87650, 32'hc0b0d6e8} /* (10, 0, 6) {real, imag} */,
  {32'hc26dba18, 32'hc1dbe344} /* (10, 0, 5) {real, imag} */,
  {32'hc144c8d5, 32'hc1cc18e6} /* (10, 0, 4) {real, imag} */,
  {32'hc2817688, 32'hc182c4d1} /* (10, 0, 3) {real, imag} */,
  {32'hc34a9d4c, 32'hc3afe09a} /* (10, 0, 2) {real, imag} */,
  {32'h44b62b0a, 32'h44930090} /* (10, 0, 1) {real, imag} */,
  {32'h4519ca44, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h4519b1b4, 32'hc4a09d10} /* (9, 31, 31) {real, imag} */,
  {32'hc41b750a, 32'h440b2cf5} /* (9, 31, 30) {real, imag} */,
  {32'hc1775210, 32'hc16dedac} /* (9, 31, 29) {real, imag} */,
  {32'h428c7824, 32'hc1210898} /* (9, 31, 28) {real, imag} */,
  {32'hc2b88f86, 32'h41b5d8cf} /* (9, 31, 27) {real, imag} */,
  {32'hc21272ca, 32'h415bcfb1} /* (9, 31, 26) {real, imag} */,
  {32'h4187fa93, 32'h40bfd081} /* (9, 31, 25) {real, imag} */,
  {32'hc112a991, 32'h41d873d2} /* (9, 31, 24) {real, imag} */,
  {32'h3ec65ae0, 32'hc1377dbe} /* (9, 31, 23) {real, imag} */,
  {32'hc1a6cade, 32'h4173b006} /* (9, 31, 22) {real, imag} */,
  {32'h404ec3a4, 32'h41a40c9a} /* (9, 31, 21) {real, imag} */,
  {32'h40fcdd38, 32'h418a3c1d} /* (9, 31, 20) {real, imag} */,
  {32'h4148b3bf, 32'h3f636a60} /* (9, 31, 19) {real, imag} */,
  {32'h405ad65a, 32'h4110be98} /* (9, 31, 18) {real, imag} */,
  {32'hc15aedf0, 32'hc08217d0} /* (9, 31, 17) {real, imag} */,
  {32'hc010715f, 32'hc0fc766a} /* (9, 31, 16) {real, imag} */,
  {32'h3e961ec4, 32'hbfc0c49c} /* (9, 31, 15) {real, imag} */,
  {32'hc1830a4a, 32'hc1c43cca} /* (9, 31, 14) {real, imag} */,
  {32'h40898cc8, 32'h4123a916} /* (9, 31, 13) {real, imag} */,
  {32'h4124890c, 32'hc10d52f6} /* (9, 31, 12) {real, imag} */,
  {32'hc1dd6582, 32'hc134f38a} /* (9, 31, 11) {real, imag} */,
  {32'hc05acc0c, 32'hc0aadedc} /* (9, 31, 10) {real, imag} */,
  {32'h414aca9c, 32'hbf245c50} /* (9, 31, 9) {real, imag} */,
  {32'hc1e9ef22, 32'hc071dc1c} /* (9, 31, 8) {real, imag} */,
  {32'h42167626, 32'h41b868f7} /* (9, 31, 7) {real, imag} */,
  {32'hc1a08e7c, 32'h41389bdc} /* (9, 31, 6) {real, imag} */,
  {32'hc2a95a45, 32'h41dc97f4} /* (9, 31, 5) {real, imag} */,
  {32'h429d877b, 32'hc2c0738a} /* (9, 31, 4) {real, imag} */,
  {32'hc2336371, 32'h41a2051b} /* (9, 31, 3) {real, imag} */,
  {32'hc3bbee4a, 32'hc28e708b} /* (9, 31, 2) {real, imag} */,
  {32'h44d2283a, 32'h43d3f00b} /* (9, 31, 1) {real, imag} */,
  {32'h45105eca, 32'hc35c289a} /* (9, 31, 0) {real, imag} */,
  {32'hc432a101, 32'hc3446f42} /* (9, 30, 31) {real, imag} */,
  {32'h43d8527b, 32'h42ec34d2} /* (9, 30, 30) {real, imag} */,
  {32'hc18dac46, 32'hc12f5658} /* (9, 30, 29) {real, imag} */,
  {32'hc2b8aad1, 32'h424ab37a} /* (9, 30, 28) {real, imag} */,
  {32'h42390c3a, 32'hc231fd35} /* (9, 30, 27) {real, imag} */,
  {32'h4182dcee, 32'h41337d9d} /* (9, 30, 26) {real, imag} */,
  {32'hc1df366c, 32'h3f8f0c70} /* (9, 30, 25) {real, imag} */,
  {32'h4190afbf, 32'hc11f2e7b} /* (9, 30, 24) {real, imag} */,
  {32'h411d899e, 32'hc134fd31} /* (9, 30, 23) {real, imag} */,
  {32'hc17fd13e, 32'h41470152} /* (9, 30, 22) {real, imag} */,
  {32'h410e2894, 32'hc127577c} /* (9, 30, 21) {real, imag} */,
  {32'h411d3200, 32'h40bca626} /* (9, 30, 20) {real, imag} */,
  {32'h4047ec5c, 32'h3f1b9480} /* (9, 30, 19) {real, imag} */,
  {32'hc02ec384, 32'hc0b2e074} /* (9, 30, 18) {real, imag} */,
  {32'hc03a2220, 32'h412c8000} /* (9, 30, 17) {real, imag} */,
  {32'h40deddd0, 32'h409b5aa5} /* (9, 30, 16) {real, imag} */,
  {32'hc0930a8a, 32'hbfc7aecc} /* (9, 30, 15) {real, imag} */,
  {32'hbff7cdf2, 32'h41e3eb3d} /* (9, 30, 14) {real, imag} */,
  {32'h40c26e5c, 32'h40937cb0} /* (9, 30, 13) {real, imag} */,
  {32'hc03b6334, 32'hc0aabf42} /* (9, 30, 12) {real, imag} */,
  {32'hc0fb4764, 32'hbcc078c0} /* (9, 30, 11) {real, imag} */,
  {32'h3f838d64, 32'hc0619436} /* (9, 30, 10) {real, imag} */,
  {32'h4135e4b7, 32'hc190bdaf} /* (9, 30, 9) {real, imag} */,
  {32'h41effc58, 32'h4196d7ef} /* (9, 30, 8) {real, imag} */,
  {32'hc119d8cb, 32'h40cb52c9} /* (9, 30, 7) {real, imag} */,
  {32'h41540f24, 32'h419890a7} /* (9, 30, 6) {real, imag} */,
  {32'h42abba8f, 32'h420fb289} /* (9, 30, 5) {real, imag} */,
  {32'hc186c26b, 32'hc292eebb} /* (9, 30, 4) {real, imag} */,
  {32'h419a4284, 32'hc230401d} /* (9, 30, 3) {real, imag} */,
  {32'h440f54ac, 32'h433538f6} /* (9, 30, 2) {real, imag} */,
  {32'hc4a2fd64, 32'h4242606e} /* (9, 30, 1) {real, imag} */,
  {32'hc42ff663, 32'h4300b112} /* (9, 30, 0) {real, imag} */,
  {32'h42c52f9a, 32'hc2d115a2} /* (9, 29, 31) {real, imag} */,
  {32'hbf5755c0, 32'h42ca9267} /* (9, 29, 30) {real, imag} */,
  {32'hc1f177e0, 32'hc108571a} /* (9, 29, 29) {real, imag} */,
  {32'hc22221b2, 32'hc07ff548} /* (9, 29, 28) {real, imag} */,
  {32'hc0d9758c, 32'hc0782040} /* (9, 29, 27) {real, imag} */,
  {32'hbf12e8c0, 32'hc1a8b76b} /* (9, 29, 26) {real, imag} */,
  {32'hc103746e, 32'h40b77d52} /* (9, 29, 25) {real, imag} */,
  {32'hc1cb02f4, 32'hc1248d92} /* (9, 29, 24) {real, imag} */,
  {32'hbdec5a10, 32'hc0c0f446} /* (9, 29, 23) {real, imag} */,
  {32'hc13cffc4, 32'hc1562576} /* (9, 29, 22) {real, imag} */,
  {32'hc045076c, 32'h3f965254} /* (9, 29, 21) {real, imag} */,
  {32'h41601a8e, 32'hc0d0f065} /* (9, 29, 20) {real, imag} */,
  {32'hc04b693a, 32'hc0eca620} /* (9, 29, 19) {real, imag} */,
  {32'hc0af22ad, 32'hc0b4f981} /* (9, 29, 18) {real, imag} */,
  {32'h411df930, 32'hc1096487} /* (9, 29, 17) {real, imag} */,
  {32'h404f2860, 32'h40cc41ff} /* (9, 29, 16) {real, imag} */,
  {32'h40a98de0, 32'h413cb9e8} /* (9, 29, 15) {real, imag} */,
  {32'h4119840e, 32'hc09a57d2} /* (9, 29, 14) {real, imag} */,
  {32'h412ac4d1, 32'h40068634} /* (9, 29, 13) {real, imag} */,
  {32'h40b5d577, 32'hc03ea28a} /* (9, 29, 12) {real, imag} */,
  {32'hc09bd94e, 32'h4135716c} /* (9, 29, 11) {real, imag} */,
  {32'hc13fc771, 32'hbf543014} /* (9, 29, 10) {real, imag} */,
  {32'hc0dacbc2, 32'hc10e4e75} /* (9, 29, 9) {real, imag} */,
  {32'h418ce24b, 32'h4190014e} /* (9, 29, 8) {real, imag} */,
  {32'hc1922f2b, 32'h40c2ea38} /* (9, 29, 7) {real, imag} */,
  {32'h3f94d3d8, 32'hc15a4ed6} /* (9, 29, 6) {real, imag} */,
  {32'hc224ce6e, 32'h413a1917} /* (9, 29, 5) {real, imag} */,
  {32'h41ef50c3, 32'hc081faa6} /* (9, 29, 4) {real, imag} */,
  {32'h3fd336b4, 32'hc1eb199d} /* (9, 29, 3) {real, imag} */,
  {32'h428a0160, 32'h432a8cc7} /* (9, 29, 2) {real, imag} */,
  {32'hc2feea4c, 32'hc2278557} /* (9, 29, 1) {real, imag} */,
  {32'hc120eb90, 32'h41e257cc} /* (9, 29, 0) {real, imag} */,
  {32'h430dff05, 32'hc2094c94} /* (9, 28, 31) {real, imag} */,
  {32'hc24694f6, 32'h42a88ca7} /* (9, 28, 30) {real, imag} */,
  {32'hc21c4e87, 32'hc2532e9c} /* (9, 28, 29) {real, imag} */,
  {32'h416aa38e, 32'hc19dab8d} /* (9, 28, 28) {real, imag} */,
  {32'hc0d00e40, 32'h41d059f2} /* (9, 28, 27) {real, imag} */,
  {32'h41bd1858, 32'h401e1364} /* (9, 28, 26) {real, imag} */,
  {32'hbfdeb5e0, 32'h417fa0e4} /* (9, 28, 25) {real, imag} */,
  {32'hc115bbe0, 32'h411c68a3} /* (9, 28, 24) {real, imag} */,
  {32'h40b25510, 32'h408f40c4} /* (9, 28, 23) {real, imag} */,
  {32'h411ae7a4, 32'hc08fb2c9} /* (9, 28, 22) {real, imag} */,
  {32'h40da790f, 32'h412d6fdd} /* (9, 28, 21) {real, imag} */,
  {32'hc1d897d5, 32'hc10eb4ec} /* (9, 28, 20) {real, imag} */,
  {32'hc08c0e3e, 32'h40afb75a} /* (9, 28, 19) {real, imag} */,
  {32'h3fad2042, 32'h40bdc6a5} /* (9, 28, 18) {real, imag} */,
  {32'h40a2a01a, 32'hc080f911} /* (9, 28, 17) {real, imag} */,
  {32'hc0c7b2e5, 32'hbfdba0e2} /* (9, 28, 16) {real, imag} */,
  {32'h4118a53c, 32'h40a1dc22} /* (9, 28, 15) {real, imag} */,
  {32'hc107a3f4, 32'h401d2ee4} /* (9, 28, 14) {real, imag} */,
  {32'hc15f7d20, 32'h41824abc} /* (9, 28, 13) {real, imag} */,
  {32'h4174b962, 32'h40112bfa} /* (9, 28, 12) {real, imag} */,
  {32'hc0238ece, 32'hc1b2aba0} /* (9, 28, 11) {real, imag} */,
  {32'hc0df5969, 32'h408ba6f6} /* (9, 28, 10) {real, imag} */,
  {32'h4165f52a, 32'h400ffaf8} /* (9, 28, 9) {real, imag} */,
  {32'h40816374, 32'h414259ce} /* (9, 28, 8) {real, imag} */,
  {32'h405b1766, 32'hc18c45ad} /* (9, 28, 7) {real, imag} */,
  {32'hc15d4d0a, 32'hc128cd71} /* (9, 28, 6) {real, imag} */,
  {32'hc1af5c3e, 32'h41be297f} /* (9, 28, 5) {real, imag} */,
  {32'h4203af83, 32'hc0b7006e} /* (9, 28, 4) {real, imag} */,
  {32'hc1535150, 32'h411a7a75} /* (9, 28, 3) {real, imag} */,
  {32'hc2bb769c, 32'h4298c6ae} /* (9, 28, 2) {real, imag} */,
  {32'h41b382f6, 32'hc2cc40c4} /* (9, 28, 1) {real, imag} */,
  {32'h4214a618, 32'hc1c19450} /* (9, 28, 0) {real, imag} */,
  {32'hc20e53da, 32'h42983dde} /* (9, 27, 31) {real, imag} */,
  {32'h41faff09, 32'hc21ee39a} /* (9, 27, 30) {real, imag} */,
  {32'hc1edfd25, 32'h4141ee4b} /* (9, 27, 29) {real, imag} */,
  {32'hc130a827, 32'h409f1190} /* (9, 27, 28) {real, imag} */,
  {32'h421b9724, 32'hc13d4d47} /* (9, 27, 27) {real, imag} */,
  {32'hc09e2312, 32'hc12b7902} /* (9, 27, 26) {real, imag} */,
  {32'hc0832666, 32'h416c7b3a} /* (9, 27, 25) {real, imag} */,
  {32'hbe003680, 32'h3fc9e728} /* (9, 27, 24) {real, imag} */,
  {32'h40a298c5, 32'h40c41566} /* (9, 27, 23) {real, imag} */,
  {32'h400fa0ac, 32'hc1e81e0d} /* (9, 27, 22) {real, imag} */,
  {32'hc00cb252, 32'hc18f4ff0} /* (9, 27, 21) {real, imag} */,
  {32'hbf9b9978, 32'hbfa2a30f} /* (9, 27, 20) {real, imag} */,
  {32'hc0284551, 32'hbff54bd0} /* (9, 27, 19) {real, imag} */,
  {32'h411496c4, 32'h3f5ce59c} /* (9, 27, 18) {real, imag} */,
  {32'h40d26ddc, 32'hbee436b4} /* (9, 27, 17) {real, imag} */,
  {32'h413dd0d8, 32'hbebd9e50} /* (9, 27, 16) {real, imag} */,
  {32'hc067b16a, 32'hc0eed38f} /* (9, 27, 15) {real, imag} */,
  {32'h3fd9e90c, 32'h4007e700} /* (9, 27, 14) {real, imag} */,
  {32'hc15efd1a, 32'hc128249b} /* (9, 27, 13) {real, imag} */,
  {32'hc11141a3, 32'h407477c2} /* (9, 27, 12) {real, imag} */,
  {32'h412b022b, 32'hc00c35a6} /* (9, 27, 11) {real, imag} */,
  {32'hc1b3b325, 32'h3e4d0100} /* (9, 27, 10) {real, imag} */,
  {32'h411501cb, 32'hbf3aa684} /* (9, 27, 9) {real, imag} */,
  {32'h413d15c2, 32'h40089c91} /* (9, 27, 8) {real, imag} */,
  {32'hc0ac7bdc, 32'hc1a11e4b} /* (9, 27, 7) {real, imag} */,
  {32'h412c16aa, 32'hc1c38d36} /* (9, 27, 6) {real, imag} */,
  {32'hc07b17c8, 32'hc1109960} /* (9, 27, 5) {real, imag} */,
  {32'hc105b0bb, 32'hbfbb7200} /* (9, 27, 4) {real, imag} */,
  {32'h419c6dff, 32'hc145efd5} /* (9, 27, 3) {real, imag} */,
  {32'h41848bb4, 32'h4107af27} /* (9, 27, 2) {real, imag} */,
  {32'hc2d1ec08, 32'h4081e296} /* (9, 27, 1) {real, imag} */,
  {32'hc259bfcc, 32'h41efe0a2} /* (9, 27, 0) {real, imag} */,
  {32'h41290938, 32'hc11a57f6} /* (9, 26, 31) {real, imag} */,
  {32'hc1dffff6, 32'h41c0c6d2} /* (9, 26, 30) {real, imag} */,
  {32'hc0e07254, 32'h40cd7805} /* (9, 26, 29) {real, imag} */,
  {32'h413292da, 32'h3fc10dc0} /* (9, 26, 28) {real, imag} */,
  {32'h40e7392e, 32'h3e56fd80} /* (9, 26, 27) {real, imag} */,
  {32'h4156bd63, 32'hc1006a9d} /* (9, 26, 26) {real, imag} */,
  {32'h40c2633a, 32'hc0b02450} /* (9, 26, 25) {real, imag} */,
  {32'h40dd23a8, 32'h41234e5d} /* (9, 26, 24) {real, imag} */,
  {32'hbfe8a5fc, 32'hc06432de} /* (9, 26, 23) {real, imag} */,
  {32'hc05745cc, 32'hc1a96a98} /* (9, 26, 22) {real, imag} */,
  {32'h415ff534, 32'hc1b1599c} /* (9, 26, 21) {real, imag} */,
  {32'hc182cfed, 32'hc14014dc} /* (9, 26, 20) {real, imag} */,
  {32'hbec60770, 32'hbff850f4} /* (9, 26, 19) {real, imag} */,
  {32'hc09861d8, 32'h40a31c67} /* (9, 26, 18) {real, imag} */,
  {32'h411278fa, 32'hc088cb0a} /* (9, 26, 17) {real, imag} */,
  {32'hc1297b59, 32'h40171e7e} /* (9, 26, 16) {real, imag} */,
  {32'hc0bc3bb4, 32'hc0f3f20d} /* (9, 26, 15) {real, imag} */,
  {32'h404e8858, 32'hc1247d7c} /* (9, 26, 14) {real, imag} */,
  {32'h40d7ff22, 32'h410faeaa} /* (9, 26, 13) {real, imag} */,
  {32'h3f3c3738, 32'hc062e628} /* (9, 26, 12) {real, imag} */,
  {32'h4103c4a6, 32'hc1146f09} /* (9, 26, 11) {real, imag} */,
  {32'h40d95fcf, 32'h4142d8b2} /* (9, 26, 10) {real, imag} */,
  {32'h40c95adb, 32'hc13dbd84} /* (9, 26, 9) {real, imag} */,
  {32'hc0918b75, 32'hc041bd62} /* (9, 26, 8) {real, imag} */,
  {32'hc121ca64, 32'hbf9de6e6} /* (9, 26, 7) {real, imag} */,
  {32'h41b1d271, 32'hc1a78c22} /* (9, 26, 6) {real, imag} */,
  {32'hc0adf51d, 32'h407f1a2c} /* (9, 26, 5) {real, imag} */,
  {32'h41b9c2ba, 32'h41a820c9} /* (9, 26, 4) {real, imag} */,
  {32'hbcf10200, 32'hc15c52b8} /* (9, 26, 3) {real, imag} */,
  {32'h410c098d, 32'hc0a5c617} /* (9, 26, 2) {real, imag} */,
  {32'h40106338, 32'hc16c182d} /* (9, 26, 1) {real, imag} */,
  {32'h401f004c, 32'hc19194ac} /* (9, 26, 0) {real, imag} */,
  {32'h3e28d720, 32'hc1b46930} /* (9, 25, 31) {real, imag} */,
  {32'hc1154f9d, 32'h41d0af36} /* (9, 25, 30) {real, imag} */,
  {32'hbff318cc, 32'hc0a4c9dc} /* (9, 25, 29) {real, imag} */,
  {32'h4026d8df, 32'hc1180da2} /* (9, 25, 28) {real, imag} */,
  {32'h41ae0abc, 32'hc081ccb5} /* (9, 25, 27) {real, imag} */,
  {32'h3f6893f0, 32'h411cf9f4} /* (9, 25, 26) {real, imag} */,
  {32'h40fc3dca, 32'h41365872} /* (9, 25, 25) {real, imag} */,
  {32'hc1337814, 32'hc0bb3a40} /* (9, 25, 24) {real, imag} */,
  {32'h40fd5ab0, 32'hc18c4f5b} /* (9, 25, 23) {real, imag} */,
  {32'h41278658, 32'h40e51bba} /* (9, 25, 22) {real, imag} */,
  {32'h40ce1327, 32'hc098c76a} /* (9, 25, 21) {real, imag} */,
  {32'hc10702ef, 32'hbf9d1b9a} /* (9, 25, 20) {real, imag} */,
  {32'h40d1304a, 32'h41aa97e8} /* (9, 25, 19) {real, imag} */,
  {32'hc18d5daf, 32'hc027a090} /* (9, 25, 18) {real, imag} */,
  {32'hc144446e, 32'hc08ac34c} /* (9, 25, 17) {real, imag} */,
  {32'hc010a314, 32'h4034c2ca} /* (9, 25, 16) {real, imag} */,
  {32'h412eb7af, 32'hc00ed740} /* (9, 25, 15) {real, imag} */,
  {32'h4025c396, 32'h40ea10f6} /* (9, 25, 14) {real, imag} */,
  {32'h41320fea, 32'hc12917ba} /* (9, 25, 13) {real, imag} */,
  {32'h40efbfe4, 32'hc1356422} /* (9, 25, 12) {real, imag} */,
  {32'hc10f11e6, 32'h4069ed31} /* (9, 25, 11) {real, imag} */,
  {32'h408fe90a, 32'hc134339a} /* (9, 25, 10) {real, imag} */,
  {32'hc1bf03b2, 32'h4024b61c} /* (9, 25, 9) {real, imag} */,
  {32'hbfa03af8, 32'h41a9dd94} /* (9, 25, 8) {real, imag} */,
  {32'hc095c019, 32'h415a9bc7} /* (9, 25, 7) {real, imag} */,
  {32'hc01429f6, 32'hc00b1ec8} /* (9, 25, 6) {real, imag} */,
  {32'hc1a64e32, 32'hc11998ba} /* (9, 25, 5) {real, imag} */,
  {32'hc105b476, 32'h40dcacf0} /* (9, 25, 4) {real, imag} */,
  {32'hc100d1fe, 32'hc1008979} /* (9, 25, 3) {real, imag} */,
  {32'h3f3320f0, 32'h41c56090} /* (9, 25, 2) {real, imag} */,
  {32'h418d0f0b, 32'hc14206ed} /* (9, 25, 1) {real, imag} */,
  {32'hc093b8dd, 32'hc0b92cb6} /* (9, 25, 0) {real, imag} */,
  {32'hc0c09db9, 32'h418e2ef2} /* (9, 24, 31) {real, imag} */,
  {32'h40db9691, 32'h4126c05a} /* (9, 24, 30) {real, imag} */,
  {32'hbf34bb00, 32'hc137909a} /* (9, 24, 29) {real, imag} */,
  {32'h40e59cee, 32'hc0604ecc} /* (9, 24, 28) {real, imag} */,
  {32'h41a1bb48, 32'h402a1284} /* (9, 24, 27) {real, imag} */,
  {32'hc0b35e82, 32'hbf9467ec} /* (9, 24, 26) {real, imag} */,
  {32'h41687c3a, 32'hc207439c} /* (9, 24, 25) {real, imag} */,
  {32'hc156b7f6, 32'hc193374b} /* (9, 24, 24) {real, imag} */,
  {32'h405726ba, 32'hc138668b} /* (9, 24, 23) {real, imag} */,
  {32'hc0cd28c2, 32'hc06d0bb8} /* (9, 24, 22) {real, imag} */,
  {32'hc0a638de, 32'h40491660} /* (9, 24, 21) {real, imag} */,
  {32'hc142ac24, 32'h4014dad1} /* (9, 24, 20) {real, imag} */,
  {32'h400e1b4c, 32'h40d31e45} /* (9, 24, 19) {real, imag} */,
  {32'hc0b60709, 32'hc130e052} /* (9, 24, 18) {real, imag} */,
  {32'hc1055741, 32'hbdbde780} /* (9, 24, 17) {real, imag} */,
  {32'h41284177, 32'hc008d2f0} /* (9, 24, 16) {real, imag} */,
  {32'hc11cf51d, 32'h4187981c} /* (9, 24, 15) {real, imag} */,
  {32'h40b43d0d, 32'hc0f1d7cb} /* (9, 24, 14) {real, imag} */,
  {32'hbf5575a0, 32'hc09d2aef} /* (9, 24, 13) {real, imag} */,
  {32'h3f76592c, 32'h40638db1} /* (9, 24, 12) {real, imag} */,
  {32'hc06f0b20, 32'hc16af8cc} /* (9, 24, 11) {real, imag} */,
  {32'hc105869f, 32'hc11d33b8} /* (9, 24, 10) {real, imag} */,
  {32'hc1c4f950, 32'h40a151ce} /* (9, 24, 9) {real, imag} */,
  {32'hc0101b68, 32'h412be38c} /* (9, 24, 8) {real, imag} */,
  {32'h40d15f48, 32'h4082ce15} /* (9, 24, 7) {real, imag} */,
  {32'h409461b4, 32'h418e0432} /* (9, 24, 6) {real, imag} */,
  {32'h40065b38, 32'h3f1a3428} /* (9, 24, 5) {real, imag} */,
  {32'h41079894, 32'hc1f35b23} /* (9, 24, 4) {real, imag} */,
  {32'h4010dde7, 32'h4163fc8c} /* (9, 24, 3) {real, imag} */,
  {32'h41f9c2d7, 32'hc115260e} /* (9, 24, 2) {real, imag} */,
  {32'hc22b9308, 32'h41b21bbd} /* (9, 24, 1) {real, imag} */,
  {32'hc20b388c, 32'h4141f294} /* (9, 24, 0) {real, imag} */,
  {32'h41d1964f, 32'h4107fbde} /* (9, 23, 31) {real, imag} */,
  {32'h4168f3cc, 32'h413b5eb7} /* (9, 23, 30) {real, imag} */,
  {32'h41290906, 32'hc13ff948} /* (9, 23, 29) {real, imag} */,
  {32'hc1939144, 32'hc1481848} /* (9, 23, 28) {real, imag} */,
  {32'hc1948df5, 32'h403c8e90} /* (9, 23, 27) {real, imag} */,
  {32'hc115a206, 32'hc14027aa} /* (9, 23, 26) {real, imag} */,
  {32'hc0ebc9de, 32'hc18f8dec} /* (9, 23, 25) {real, imag} */,
  {32'h413fc2e9, 32'h418a8aa8} /* (9, 23, 24) {real, imag} */,
  {32'hc12b39a1, 32'h404f7b6e} /* (9, 23, 23) {real, imag} */,
  {32'h41c839b3, 32'hc12276db} /* (9, 23, 22) {real, imag} */,
  {32'hbf769a34, 32'h4113a178} /* (9, 23, 21) {real, imag} */,
  {32'hc136e39d, 32'hbf8e6c98} /* (9, 23, 20) {real, imag} */,
  {32'hc0f8d97a, 32'hc1391768} /* (9, 23, 19) {real, imag} */,
  {32'h3feab22c, 32'hbf847d0a} /* (9, 23, 18) {real, imag} */,
  {32'h406513d3, 32'h41468d6e} /* (9, 23, 17) {real, imag} */,
  {32'h412d974e, 32'hbfcffaca} /* (9, 23, 16) {real, imag} */,
  {32'hbfbaa008, 32'hc0c22151} /* (9, 23, 15) {real, imag} */,
  {32'h40d511a0, 32'hbf40d170} /* (9, 23, 14) {real, imag} */,
  {32'hc18e3a41, 32'hc1b287f4} /* (9, 23, 13) {real, imag} */,
  {32'hc04dde10, 32'hc0158a28} /* (9, 23, 12) {real, imag} */,
  {32'hc13f1268, 32'h406e6bd5} /* (9, 23, 11) {real, imag} */,
  {32'h40a63dcc, 32'h4134c2ee} /* (9, 23, 10) {real, imag} */,
  {32'h404aad82, 32'h40cde7fe} /* (9, 23, 9) {real, imag} */,
  {32'hc13ae645, 32'h410b0e76} /* (9, 23, 8) {real, imag} */,
  {32'h40ea2840, 32'h4013f88f} /* (9, 23, 7) {real, imag} */,
  {32'hc088eafd, 32'h3ff8cb20} /* (9, 23, 6) {real, imag} */,
  {32'hc0721c05, 32'hc1497cd5} /* (9, 23, 5) {real, imag} */,
  {32'hc08fa26c, 32'hc00d6e22} /* (9, 23, 4) {real, imag} */,
  {32'h413408a2, 32'hc0ea9ccc} /* (9, 23, 3) {real, imag} */,
  {32'hc0fd5536, 32'h41b01132} /* (9, 23, 2) {real, imag} */,
  {32'hc110f302, 32'hc18b683c} /* (9, 23, 1) {real, imag} */,
  {32'h41081a94, 32'h41820bc7} /* (9, 23, 0) {real, imag} */,
  {32'h41233d98, 32'hc1732f6d} /* (9, 22, 31) {real, imag} */,
  {32'h402215a1, 32'hbf95223e} /* (9, 22, 30) {real, imag} */,
  {32'h418c27ef, 32'h3edb2690} /* (9, 22, 29) {real, imag} */,
  {32'hc15fd0b2, 32'hbf7c0638} /* (9, 22, 28) {real, imag} */,
  {32'hc114ceee, 32'h414e3614} /* (9, 22, 27) {real, imag} */,
  {32'h40740717, 32'hbe5282e0} /* (9, 22, 26) {real, imag} */,
  {32'h416ec109, 32'h418b2f41} /* (9, 22, 25) {real, imag} */,
  {32'h411bd2ab, 32'hc0cb51fd} /* (9, 22, 24) {real, imag} */,
  {32'h3f0a3250, 32'h41931044} /* (9, 22, 23) {real, imag} */,
  {32'hc1cf2a5b, 32'hbecae300} /* (9, 22, 22) {real, imag} */,
  {32'h40d00520, 32'h410d35cc} /* (9, 22, 21) {real, imag} */,
  {32'hc0b2f56f, 32'h40104ae2} /* (9, 22, 20) {real, imag} */,
  {32'hc1258c60, 32'h417ed0e6} /* (9, 22, 19) {real, imag} */,
  {32'h41b400d4, 32'hc189e9f0} /* (9, 22, 18) {real, imag} */,
  {32'hc006e7d6, 32'h409eccc1} /* (9, 22, 17) {real, imag} */,
  {32'hc0b79a71, 32'h3f2849d0} /* (9, 22, 16) {real, imag} */,
  {32'h3f28b8bc, 32'h40f79e3b} /* (9, 22, 15) {real, imag} */,
  {32'hc18de962, 32'h410427ab} /* (9, 22, 14) {real, imag} */,
  {32'hc1a496b2, 32'h4094d05a} /* (9, 22, 13) {real, imag} */,
  {32'hbf615188, 32'hc141fef4} /* (9, 22, 12) {real, imag} */,
  {32'h41616c4a, 32'hc097a936} /* (9, 22, 11) {real, imag} */,
  {32'h40cf4308, 32'h41237fa5} /* (9, 22, 10) {real, imag} */,
  {32'hbf62ec48, 32'h4136caa0} /* (9, 22, 9) {real, imag} */,
  {32'h40ffa908, 32'hc024b358} /* (9, 22, 8) {real, imag} */,
  {32'hc1153db3, 32'hc0509d0e} /* (9, 22, 7) {real, imag} */,
  {32'h41038eeb, 32'h40469cf6} /* (9, 22, 6) {real, imag} */,
  {32'hc080da64, 32'h3f970de8} /* (9, 22, 5) {real, imag} */,
  {32'hc1274539, 32'h40b51160} /* (9, 22, 4) {real, imag} */,
  {32'hbfe3c370, 32'hc1302d04} /* (9, 22, 3) {real, imag} */,
  {32'h3fb6182e, 32'h40e3a9f0} /* (9, 22, 2) {real, imag} */,
  {32'h4190603d, 32'h41202b35} /* (9, 22, 1) {real, imag} */,
  {32'hc19d7a93, 32'hc0c2dd4d} /* (9, 22, 0) {real, imag} */,
  {32'hc0e57d9a, 32'h41729ca6} /* (9, 21, 31) {real, imag} */,
  {32'h4063d485, 32'h3fad276c} /* (9, 21, 30) {real, imag} */,
  {32'h4128dac4, 32'hc1434522} /* (9, 21, 29) {real, imag} */,
  {32'hc192aa7e, 32'h40cc5c3a} /* (9, 21, 28) {real, imag} */,
  {32'h3fdb916c, 32'hc0ac8542} /* (9, 21, 27) {real, imag} */,
  {32'h40bd3c41, 32'h40e499dd} /* (9, 21, 26) {real, imag} */,
  {32'hc0a71438, 32'hc082fca2} /* (9, 21, 25) {real, imag} */,
  {32'h3ee0aec0, 32'hc136c532} /* (9, 21, 24) {real, imag} */,
  {32'hc1176cb5, 32'hbfd5a670} /* (9, 21, 23) {real, imag} */,
  {32'hc0dc36e2, 32'hc037dd8a} /* (9, 21, 22) {real, imag} */,
  {32'hc11f4117, 32'hc16cdde4} /* (9, 21, 21) {real, imag} */,
  {32'h3f49d8f8, 32'h40cad478} /* (9, 21, 20) {real, imag} */,
  {32'h40c45724, 32'h4185862d} /* (9, 21, 19) {real, imag} */,
  {32'h3e586c00, 32'h41f0445d} /* (9, 21, 18) {real, imag} */,
  {32'h405d8ca2, 32'hc0e71420} /* (9, 21, 17) {real, imag} */,
  {32'h40cf5b26, 32'hc1183972} /* (9, 21, 16) {real, imag} */,
  {32'hc149ee60, 32'h3f9f090b} /* (9, 21, 15) {real, imag} */,
  {32'h3f3e5aa0, 32'h407ab20c} /* (9, 21, 14) {real, imag} */,
  {32'hc1981146, 32'hc09d84ed} /* (9, 21, 13) {real, imag} */,
  {32'hc10f9c8c, 32'h4132e161} /* (9, 21, 12) {real, imag} */,
  {32'h412f3a78, 32'hc172a8d5} /* (9, 21, 11) {real, imag} */,
  {32'hbf825360, 32'hc1907dd4} /* (9, 21, 10) {real, imag} */,
  {32'h3f4b4390, 32'h4099fbe2} /* (9, 21, 9) {real, imag} */,
  {32'h40fc2b0e, 32'hc1449334} /* (9, 21, 8) {real, imag} */,
  {32'hc0dd9477, 32'h40aa72a6} /* (9, 21, 7) {real, imag} */,
  {32'hc097c05a, 32'h3fa81e30} /* (9, 21, 6) {real, imag} */,
  {32'h415c0d49, 32'hc0c795b8} /* (9, 21, 5) {real, imag} */,
  {32'h4121d3e2, 32'h4178e4d4} /* (9, 21, 4) {real, imag} */,
  {32'hbf021080, 32'hc1982141} /* (9, 21, 3) {real, imag} */,
  {32'h407df1b8, 32'hc08735ab} /* (9, 21, 2) {real, imag} */,
  {32'hc1a247c5, 32'h41688766} /* (9, 21, 1) {real, imag} */,
  {32'hc1be043d, 32'h408cd588} /* (9, 21, 0) {real, imag} */,
  {32'h3fd60cd4, 32'h41831d6e} /* (9, 20, 31) {real, imag} */,
  {32'h411092e7, 32'h40a6c0a6} /* (9, 20, 30) {real, imag} */,
  {32'hc1a1b6f6, 32'h410abe67} /* (9, 20, 29) {real, imag} */,
  {32'h41529958, 32'hc07a9a4f} /* (9, 20, 28) {real, imag} */,
  {32'h413a84b7, 32'hc14be5c5} /* (9, 20, 27) {real, imag} */,
  {32'h402a00a1, 32'hc0aabea6} /* (9, 20, 26) {real, imag} */,
  {32'hc1e01c02, 32'h4135a725} /* (9, 20, 25) {real, imag} */,
  {32'hc14c63c6, 32'h41a1d086} /* (9, 20, 24) {real, imag} */,
  {32'h4065c818, 32'hbe7cf830} /* (9, 20, 23) {real, imag} */,
  {32'hbfb0a1f2, 32'h416b157b} /* (9, 20, 22) {real, imag} */,
  {32'h3e9b220c, 32'h412be35e} /* (9, 20, 21) {real, imag} */,
  {32'hc03e7ef6, 32'h3fa41738} /* (9, 20, 20) {real, imag} */,
  {32'hc0aaf2cb, 32'h414c5bae} /* (9, 20, 19) {real, imag} */,
  {32'hc0ebbbce, 32'h4138770c} /* (9, 20, 18) {real, imag} */,
  {32'h40bf0496, 32'hc12116fa} /* (9, 20, 17) {real, imag} */,
  {32'h3f4f6218, 32'hc14e49be} /* (9, 20, 16) {real, imag} */,
  {32'h3ec44378, 32'h40c13296} /* (9, 20, 15) {real, imag} */,
  {32'h41a4fdbe, 32'h41100fef} /* (9, 20, 14) {real, imag} */,
  {32'hc127c7be, 32'h3ff4e84c} /* (9, 20, 13) {real, imag} */,
  {32'h40a5920b, 32'hc0299d92} /* (9, 20, 12) {real, imag} */,
  {32'h403cc150, 32'h4007208a} /* (9, 20, 11) {real, imag} */,
  {32'h409011d6, 32'h413d90d3} /* (9, 20, 10) {real, imag} */,
  {32'h40c406eb, 32'h414c2cac} /* (9, 20, 9) {real, imag} */,
  {32'hc1b97102, 32'hc0c5f8e8} /* (9, 20, 8) {real, imag} */,
  {32'h419ac234, 32'h41397f2a} /* (9, 20, 7) {real, imag} */,
  {32'hc16265ca, 32'hc046abaf} /* (9, 20, 6) {real, imag} */,
  {32'h4116701f, 32'h407e2ba0} /* (9, 20, 5) {real, imag} */,
  {32'h4105d2f1, 32'hc0a6581b} /* (9, 20, 4) {real, imag} */,
  {32'hc10f87ad, 32'hc0e23f7c} /* (9, 20, 3) {real, imag} */,
  {32'h41165e62, 32'h40b80b10} /* (9, 20, 2) {real, imag} */,
  {32'h40a708ef, 32'h410b862d} /* (9, 20, 1) {real, imag} */,
  {32'h4003d0ff, 32'hc1224e9a} /* (9, 20, 0) {real, imag} */,
  {32'hbf014318, 32'h3f2e6ea0} /* (9, 19, 31) {real, imag} */,
  {32'h407ce838, 32'hbe928740} /* (9, 19, 30) {real, imag} */,
  {32'hbfce3dfe, 32'h3fd12d54} /* (9, 19, 29) {real, imag} */,
  {32'h3f5a5726, 32'hc0db7154} /* (9, 19, 28) {real, imag} */,
  {32'h409517bb, 32'h3f0cadec} /* (9, 19, 27) {real, imag} */,
  {32'hc065278a, 32'h410152e3} /* (9, 19, 26) {real, imag} */,
  {32'hc07fe130, 32'h4148f194} /* (9, 19, 25) {real, imag} */,
  {32'h4089b365, 32'hbf01b7d0} /* (9, 19, 24) {real, imag} */,
  {32'hc04385a7, 32'hc1102ba8} /* (9, 19, 23) {real, imag} */,
  {32'h4159abb0, 32'h4064a862} /* (9, 19, 22) {real, imag} */,
  {32'hc16f50db, 32'h3ebc2ef8} /* (9, 19, 21) {real, imag} */,
  {32'hc0d09110, 32'h4123fc48} /* (9, 19, 20) {real, imag} */,
  {32'h3f7c719a, 32'h419a9fe2} /* (9, 19, 19) {real, imag} */,
  {32'h3fad6ea8, 32'hc00407a4} /* (9, 19, 18) {real, imag} */,
  {32'h40ca72ac, 32'hc1337377} /* (9, 19, 17) {real, imag} */,
  {32'hc11bdd34, 32'h40a3021a} /* (9, 19, 16) {real, imag} */,
  {32'h4085e81a, 32'hc0fe6164} /* (9, 19, 15) {real, imag} */,
  {32'hc0d69992, 32'hc13ff6a9} /* (9, 19, 14) {real, imag} */,
  {32'h41068832, 32'h403fce79} /* (9, 19, 13) {real, imag} */,
  {32'hc135a3f8, 32'hc11e9e92} /* (9, 19, 12) {real, imag} */,
  {32'h41083dcf, 32'h41290f2b} /* (9, 19, 11) {real, imag} */,
  {32'h40a2c20e, 32'h3fd5160c} /* (9, 19, 10) {real, imag} */,
  {32'h3f81a880, 32'hc1a51a62} /* (9, 19, 9) {real, imag} */,
  {32'hbfbbbcb9, 32'h40a66348} /* (9, 19, 8) {real, imag} */,
  {32'hbfb85982, 32'h40a5a5ff} /* (9, 19, 7) {real, imag} */,
  {32'h418892e1, 32'h40c65662} /* (9, 19, 6) {real, imag} */,
  {32'h4123bb86, 32'h408c42ac} /* (9, 19, 5) {real, imag} */,
  {32'hc189dbf3, 32'hbf887192} /* (9, 19, 4) {real, imag} */,
  {32'hc0d48223, 32'hc0260bc6} /* (9, 19, 3) {real, imag} */,
  {32'h3f411f30, 32'hc1202ff0} /* (9, 19, 2) {real, imag} */,
  {32'hbf918aa0, 32'h4077d528} /* (9, 19, 1) {real, imag} */,
  {32'hc0161680, 32'h41295179} /* (9, 19, 0) {real, imag} */,
  {32'h3e985538, 32'h41416020} /* (9, 18, 31) {real, imag} */,
  {32'hbf095dc0, 32'h40addac8} /* (9, 18, 30) {real, imag} */,
  {32'hc0d0ef0a, 32'h41975d2d} /* (9, 18, 29) {real, imag} */,
  {32'h40941e55, 32'h40814b97} /* (9, 18, 28) {real, imag} */,
  {32'hc0a0826d, 32'h40393c2a} /* (9, 18, 27) {real, imag} */,
  {32'hbf1fb7c8, 32'h3f820574} /* (9, 18, 26) {real, imag} */,
  {32'h40514bfb, 32'h40ec2fd2} /* (9, 18, 25) {real, imag} */,
  {32'hbff24638, 32'hc065b09e} /* (9, 18, 24) {real, imag} */,
  {32'h3ef850aa, 32'h413d3f9b} /* (9, 18, 23) {real, imag} */,
  {32'h3fcaf9d8, 32'h3ffea744} /* (9, 18, 22) {real, imag} */,
  {32'hc1213f18, 32'h41041a31} /* (9, 18, 21) {real, imag} */,
  {32'h400b56be, 32'hc04a17d8} /* (9, 18, 20) {real, imag} */,
  {32'hc0c29c40, 32'hbff05144} /* (9, 18, 19) {real, imag} */,
  {32'hbfc34798, 32'h3fcd7216} /* (9, 18, 18) {real, imag} */,
  {32'h3eec9a80, 32'hc08a37c1} /* (9, 18, 17) {real, imag} */,
  {32'h419fcc36, 32'h40c25145} /* (9, 18, 16) {real, imag} */,
  {32'hc108d54a, 32'hc0464c2a} /* (9, 18, 15) {real, imag} */,
  {32'h415e9881, 32'hc1229d08} /* (9, 18, 14) {real, imag} */,
  {32'hc063dd9c, 32'hc09b673b} /* (9, 18, 13) {real, imag} */,
  {32'hc0a397f9, 32'h41255073} /* (9, 18, 12) {real, imag} */,
  {32'h41608b89, 32'hc011fc4a} /* (9, 18, 11) {real, imag} */,
  {32'h40cca8d2, 32'h41450ed4} /* (9, 18, 10) {real, imag} */,
  {32'hc1104790, 32'h41242777} /* (9, 18, 9) {real, imag} */,
  {32'h41996520, 32'h40c46606} /* (9, 18, 8) {real, imag} */,
  {32'h4119fd0e, 32'hbfe5045d} /* (9, 18, 7) {real, imag} */,
  {32'h3fffab80, 32'h4145fd48} /* (9, 18, 6) {real, imag} */,
  {32'h41160144, 32'hc184d019} /* (9, 18, 5) {real, imag} */,
  {32'h40a6af1d, 32'h418ff41c} /* (9, 18, 4) {real, imag} */,
  {32'h4021380a, 32'hc0a7399f} /* (9, 18, 3) {real, imag} */,
  {32'h413b4179, 32'h4097e474} /* (9, 18, 2) {real, imag} */,
  {32'hbf8c0e90, 32'h3ebbbc60} /* (9, 18, 1) {real, imag} */,
  {32'hc0637268, 32'h403ac67c} /* (9, 18, 0) {real, imag} */,
  {32'h3f2796b0, 32'hc09aaf44} /* (9, 17, 31) {real, imag} */,
  {32'h400978fc, 32'h408f60da} /* (9, 17, 30) {real, imag} */,
  {32'h40e6fa50, 32'h400b008f} /* (9, 17, 29) {real, imag} */,
  {32'hc01f8094, 32'hbf5beff8} /* (9, 17, 28) {real, imag} */,
  {32'hbffc3dba, 32'hc0e104cc} /* (9, 17, 27) {real, imag} */,
  {32'h40b65e4c, 32'hc0f0c9c8} /* (9, 17, 26) {real, imag} */,
  {32'h410991a1, 32'hc0e9294e} /* (9, 17, 25) {real, imag} */,
  {32'hc1058377, 32'hc13de941} /* (9, 17, 24) {real, imag} */,
  {32'h40aa521a, 32'hc18c442e} /* (9, 17, 23) {real, imag} */,
  {32'hc148e88e, 32'h408fd35e} /* (9, 17, 22) {real, imag} */,
  {32'hc050ecc6, 32'h412fd43e} /* (9, 17, 21) {real, imag} */,
  {32'hbf725c58, 32'h40347c3d} /* (9, 17, 20) {real, imag} */,
  {32'hc17ff72b, 32'h4002957f} /* (9, 17, 19) {real, imag} */,
  {32'h4102e48d, 32'hc10bc63e} /* (9, 17, 18) {real, imag} */,
  {32'hc127d660, 32'h41020f6d} /* (9, 17, 17) {real, imag} */,
  {32'hbfa522a2, 32'h4149e0ae} /* (9, 17, 16) {real, imag} */,
  {32'h40994c50, 32'h3f283448} /* (9, 17, 15) {real, imag} */,
  {32'h408221fb, 32'h3ed7b660} /* (9, 17, 14) {real, imag} */,
  {32'h412d267f, 32'h40c80a22} /* (9, 17, 13) {real, imag} */,
  {32'h3ebec248, 32'h40e59767} /* (9, 17, 12) {real, imag} */,
  {32'hc094dc14, 32'h3f9e84e4} /* (9, 17, 11) {real, imag} */,
  {32'hc0b0fa66, 32'h3f85aed8} /* (9, 17, 10) {real, imag} */,
  {32'hc0add149, 32'hc0d99b4c} /* (9, 17, 9) {real, imag} */,
  {32'h400b7e08, 32'hc0a08d36} /* (9, 17, 8) {real, imag} */,
  {32'h408c981f, 32'hbf9fe508} /* (9, 17, 7) {real, imag} */,
  {32'hc0fb69c1, 32'h41487038} /* (9, 17, 6) {real, imag} */,
  {32'hbfaf5ea2, 32'hbfb495fa} /* (9, 17, 5) {real, imag} */,
  {32'h40230b2b, 32'hc08ee1e6} /* (9, 17, 4) {real, imag} */,
  {32'h405d3deb, 32'h406c32e9} /* (9, 17, 3) {real, imag} */,
  {32'hbddd3200, 32'h41512753} /* (9, 17, 2) {real, imag} */,
  {32'hbfc1e1fc, 32'hbff29520} /* (9, 17, 1) {real, imag} */,
  {32'hc11b1a58, 32'hbe2cae00} /* (9, 17, 0) {real, imag} */,
  {32'hc0334c11, 32'h412231cd} /* (9, 16, 31) {real, imag} */,
  {32'hc110aa3c, 32'hc0f76e1a} /* (9, 16, 30) {real, imag} */,
  {32'h40a9cdf6, 32'h405c1184} /* (9, 16, 29) {real, imag} */,
  {32'h405c25a0, 32'hc10c1626} /* (9, 16, 28) {real, imag} */,
  {32'hc0feb055, 32'hc1180731} /* (9, 16, 27) {real, imag} */,
  {32'hc03b5791, 32'h3ec38c30} /* (9, 16, 26) {real, imag} */,
  {32'h408105b2, 32'hbf740510} /* (9, 16, 25) {real, imag} */,
  {32'h400716d4, 32'hc1215a09} /* (9, 16, 24) {real, imag} */,
  {32'hbf8f4316, 32'h3f530130} /* (9, 16, 23) {real, imag} */,
  {32'hc09b4fa0, 32'h4158dfc6} /* (9, 16, 22) {real, imag} */,
  {32'hc09175c4, 32'hc09faa8c} /* (9, 16, 21) {real, imag} */,
  {32'h414c489e, 32'hc0db9380} /* (9, 16, 20) {real, imag} */,
  {32'h412c45ca, 32'hc187ed7a} /* (9, 16, 19) {real, imag} */,
  {32'hc0c0f9ca, 32'hc02b1351} /* (9, 16, 18) {real, imag} */,
  {32'h3e9bd754, 32'h4125bc1e} /* (9, 16, 17) {real, imag} */,
  {32'h40ad2dc8, 32'h00000000} /* (9, 16, 16) {real, imag} */,
  {32'h3e9bd754, 32'hc125bc1e} /* (9, 16, 15) {real, imag} */,
  {32'hc0c0f9ca, 32'h402b1351} /* (9, 16, 14) {real, imag} */,
  {32'h412c45ca, 32'h4187ed7a} /* (9, 16, 13) {real, imag} */,
  {32'h414c489e, 32'h40db9380} /* (9, 16, 12) {real, imag} */,
  {32'hc09175c4, 32'h409faa8c} /* (9, 16, 11) {real, imag} */,
  {32'hc09b4fa0, 32'hc158dfc6} /* (9, 16, 10) {real, imag} */,
  {32'hbf8f4316, 32'hbf530130} /* (9, 16, 9) {real, imag} */,
  {32'h400716d4, 32'h41215a09} /* (9, 16, 8) {real, imag} */,
  {32'h408105b2, 32'h3f740510} /* (9, 16, 7) {real, imag} */,
  {32'hc03b5791, 32'hbec38c30} /* (9, 16, 6) {real, imag} */,
  {32'hc0feb055, 32'h41180731} /* (9, 16, 5) {real, imag} */,
  {32'h405c25a0, 32'h410c1626} /* (9, 16, 4) {real, imag} */,
  {32'h40a9cdf6, 32'hc05c1184} /* (9, 16, 3) {real, imag} */,
  {32'hc110aa3c, 32'h40f76e1a} /* (9, 16, 2) {real, imag} */,
  {32'hc0334c11, 32'hc12231cd} /* (9, 16, 1) {real, imag} */,
  {32'h409aab86, 32'h00000000} /* (9, 16, 0) {real, imag} */,
  {32'hbfc1e1fc, 32'h3ff29520} /* (9, 15, 31) {real, imag} */,
  {32'hbddd3200, 32'hc1512753} /* (9, 15, 30) {real, imag} */,
  {32'h405d3deb, 32'hc06c32e9} /* (9, 15, 29) {real, imag} */,
  {32'h40230b2b, 32'h408ee1e6} /* (9, 15, 28) {real, imag} */,
  {32'hbfaf5ea2, 32'h3fb495fa} /* (9, 15, 27) {real, imag} */,
  {32'hc0fb69c1, 32'hc1487038} /* (9, 15, 26) {real, imag} */,
  {32'h408c981f, 32'h3f9fe508} /* (9, 15, 25) {real, imag} */,
  {32'h400b7e08, 32'h40a08d36} /* (9, 15, 24) {real, imag} */,
  {32'hc0add149, 32'h40d99b4c} /* (9, 15, 23) {real, imag} */,
  {32'hc0b0fa66, 32'hbf85aed8} /* (9, 15, 22) {real, imag} */,
  {32'hc094dc14, 32'hbf9e84e4} /* (9, 15, 21) {real, imag} */,
  {32'h3ebec248, 32'hc0e59767} /* (9, 15, 20) {real, imag} */,
  {32'h412d267f, 32'hc0c80a22} /* (9, 15, 19) {real, imag} */,
  {32'h408221fb, 32'hbed7b660} /* (9, 15, 18) {real, imag} */,
  {32'h40994c50, 32'hbf283448} /* (9, 15, 17) {real, imag} */,
  {32'hbfa522a2, 32'hc149e0ae} /* (9, 15, 16) {real, imag} */,
  {32'hc127d660, 32'hc1020f6d} /* (9, 15, 15) {real, imag} */,
  {32'h4102e48d, 32'h410bc63e} /* (9, 15, 14) {real, imag} */,
  {32'hc17ff72b, 32'hc002957f} /* (9, 15, 13) {real, imag} */,
  {32'hbf725c58, 32'hc0347c3d} /* (9, 15, 12) {real, imag} */,
  {32'hc050ecc6, 32'hc12fd43e} /* (9, 15, 11) {real, imag} */,
  {32'hc148e88e, 32'hc08fd35e} /* (9, 15, 10) {real, imag} */,
  {32'h40aa521a, 32'h418c442e} /* (9, 15, 9) {real, imag} */,
  {32'hc1058377, 32'h413de941} /* (9, 15, 8) {real, imag} */,
  {32'h410991a1, 32'h40e9294e} /* (9, 15, 7) {real, imag} */,
  {32'h40b65e4c, 32'h40f0c9c8} /* (9, 15, 6) {real, imag} */,
  {32'hbffc3dba, 32'h40e104cc} /* (9, 15, 5) {real, imag} */,
  {32'hc01f8094, 32'h3f5beff8} /* (9, 15, 4) {real, imag} */,
  {32'h40e6fa50, 32'hc00b008f} /* (9, 15, 3) {real, imag} */,
  {32'h400978fc, 32'hc08f60da} /* (9, 15, 2) {real, imag} */,
  {32'h3f2796b0, 32'h409aaf44} /* (9, 15, 1) {real, imag} */,
  {32'hc11b1a58, 32'h3e2cae00} /* (9, 15, 0) {real, imag} */,
  {32'hbf8c0e90, 32'hbebbbc60} /* (9, 14, 31) {real, imag} */,
  {32'h413b4179, 32'hc097e474} /* (9, 14, 30) {real, imag} */,
  {32'h4021380a, 32'h40a7399f} /* (9, 14, 29) {real, imag} */,
  {32'h40a6af1d, 32'hc18ff41c} /* (9, 14, 28) {real, imag} */,
  {32'h41160144, 32'h4184d019} /* (9, 14, 27) {real, imag} */,
  {32'h3fffab80, 32'hc145fd48} /* (9, 14, 26) {real, imag} */,
  {32'h4119fd0e, 32'h3fe5045d} /* (9, 14, 25) {real, imag} */,
  {32'h41996520, 32'hc0c46606} /* (9, 14, 24) {real, imag} */,
  {32'hc1104790, 32'hc1242777} /* (9, 14, 23) {real, imag} */,
  {32'h40cca8d2, 32'hc1450ed4} /* (9, 14, 22) {real, imag} */,
  {32'h41608b89, 32'h4011fc4a} /* (9, 14, 21) {real, imag} */,
  {32'hc0a397f9, 32'hc1255073} /* (9, 14, 20) {real, imag} */,
  {32'hc063dd9c, 32'h409b673b} /* (9, 14, 19) {real, imag} */,
  {32'h415e9881, 32'h41229d08} /* (9, 14, 18) {real, imag} */,
  {32'hc108d54a, 32'h40464c2a} /* (9, 14, 17) {real, imag} */,
  {32'h419fcc36, 32'hc0c25145} /* (9, 14, 16) {real, imag} */,
  {32'h3eec9a80, 32'h408a37c1} /* (9, 14, 15) {real, imag} */,
  {32'hbfc34798, 32'hbfcd7216} /* (9, 14, 14) {real, imag} */,
  {32'hc0c29c40, 32'h3ff05144} /* (9, 14, 13) {real, imag} */,
  {32'h400b56be, 32'h404a17d8} /* (9, 14, 12) {real, imag} */,
  {32'hc1213f18, 32'hc1041a31} /* (9, 14, 11) {real, imag} */,
  {32'h3fcaf9d8, 32'hbffea744} /* (9, 14, 10) {real, imag} */,
  {32'h3ef850aa, 32'hc13d3f9b} /* (9, 14, 9) {real, imag} */,
  {32'hbff24638, 32'h4065b09e} /* (9, 14, 8) {real, imag} */,
  {32'h40514bfb, 32'hc0ec2fd2} /* (9, 14, 7) {real, imag} */,
  {32'hbf1fb7c8, 32'hbf820574} /* (9, 14, 6) {real, imag} */,
  {32'hc0a0826d, 32'hc0393c2a} /* (9, 14, 5) {real, imag} */,
  {32'h40941e55, 32'hc0814b97} /* (9, 14, 4) {real, imag} */,
  {32'hc0d0ef0a, 32'hc1975d2d} /* (9, 14, 3) {real, imag} */,
  {32'hbf095dc0, 32'hc0addac8} /* (9, 14, 2) {real, imag} */,
  {32'h3e985538, 32'hc1416020} /* (9, 14, 1) {real, imag} */,
  {32'hc0637268, 32'hc03ac67c} /* (9, 14, 0) {real, imag} */,
  {32'hbf918aa0, 32'hc077d528} /* (9, 13, 31) {real, imag} */,
  {32'h3f411f30, 32'h41202ff0} /* (9, 13, 30) {real, imag} */,
  {32'hc0d48223, 32'h40260bc6} /* (9, 13, 29) {real, imag} */,
  {32'hc189dbf3, 32'h3f887192} /* (9, 13, 28) {real, imag} */,
  {32'h4123bb86, 32'hc08c42ac} /* (9, 13, 27) {real, imag} */,
  {32'h418892e1, 32'hc0c65662} /* (9, 13, 26) {real, imag} */,
  {32'hbfb85982, 32'hc0a5a5ff} /* (9, 13, 25) {real, imag} */,
  {32'hbfbbbcb9, 32'hc0a66348} /* (9, 13, 24) {real, imag} */,
  {32'h3f81a880, 32'h41a51a62} /* (9, 13, 23) {real, imag} */,
  {32'h40a2c20e, 32'hbfd5160c} /* (9, 13, 22) {real, imag} */,
  {32'h41083dcf, 32'hc1290f2b} /* (9, 13, 21) {real, imag} */,
  {32'hc135a3f8, 32'h411e9e92} /* (9, 13, 20) {real, imag} */,
  {32'h41068832, 32'hc03fce79} /* (9, 13, 19) {real, imag} */,
  {32'hc0d69992, 32'h413ff6a9} /* (9, 13, 18) {real, imag} */,
  {32'h4085e81a, 32'h40fe6164} /* (9, 13, 17) {real, imag} */,
  {32'hc11bdd34, 32'hc0a3021a} /* (9, 13, 16) {real, imag} */,
  {32'h40ca72ac, 32'h41337377} /* (9, 13, 15) {real, imag} */,
  {32'h3fad6ea8, 32'h400407a4} /* (9, 13, 14) {real, imag} */,
  {32'h3f7c719a, 32'hc19a9fe2} /* (9, 13, 13) {real, imag} */,
  {32'hc0d09110, 32'hc123fc48} /* (9, 13, 12) {real, imag} */,
  {32'hc16f50db, 32'hbebc2ef8} /* (9, 13, 11) {real, imag} */,
  {32'h4159abb0, 32'hc064a862} /* (9, 13, 10) {real, imag} */,
  {32'hc04385a7, 32'h41102ba8} /* (9, 13, 9) {real, imag} */,
  {32'h4089b365, 32'h3f01b7d0} /* (9, 13, 8) {real, imag} */,
  {32'hc07fe130, 32'hc148f194} /* (9, 13, 7) {real, imag} */,
  {32'hc065278a, 32'hc10152e3} /* (9, 13, 6) {real, imag} */,
  {32'h409517bb, 32'hbf0cadec} /* (9, 13, 5) {real, imag} */,
  {32'h3f5a5726, 32'h40db7154} /* (9, 13, 4) {real, imag} */,
  {32'hbfce3dfe, 32'hbfd12d54} /* (9, 13, 3) {real, imag} */,
  {32'h407ce838, 32'h3e928740} /* (9, 13, 2) {real, imag} */,
  {32'hbf014318, 32'hbf2e6ea0} /* (9, 13, 1) {real, imag} */,
  {32'hc0161680, 32'hc1295179} /* (9, 13, 0) {real, imag} */,
  {32'h40a708ef, 32'hc10b862d} /* (9, 12, 31) {real, imag} */,
  {32'h41165e62, 32'hc0b80b10} /* (9, 12, 30) {real, imag} */,
  {32'hc10f87ad, 32'h40e23f7c} /* (9, 12, 29) {real, imag} */,
  {32'h4105d2f1, 32'h40a6581b} /* (9, 12, 28) {real, imag} */,
  {32'h4116701f, 32'hc07e2ba0} /* (9, 12, 27) {real, imag} */,
  {32'hc16265ca, 32'h4046abaf} /* (9, 12, 26) {real, imag} */,
  {32'h419ac234, 32'hc1397f2a} /* (9, 12, 25) {real, imag} */,
  {32'hc1b97102, 32'h40c5f8e8} /* (9, 12, 24) {real, imag} */,
  {32'h40c406eb, 32'hc14c2cac} /* (9, 12, 23) {real, imag} */,
  {32'h409011d6, 32'hc13d90d3} /* (9, 12, 22) {real, imag} */,
  {32'h403cc150, 32'hc007208a} /* (9, 12, 21) {real, imag} */,
  {32'h40a5920b, 32'h40299d92} /* (9, 12, 20) {real, imag} */,
  {32'hc127c7be, 32'hbff4e84c} /* (9, 12, 19) {real, imag} */,
  {32'h41a4fdbe, 32'hc1100fef} /* (9, 12, 18) {real, imag} */,
  {32'h3ec44378, 32'hc0c13296} /* (9, 12, 17) {real, imag} */,
  {32'h3f4f6218, 32'h414e49be} /* (9, 12, 16) {real, imag} */,
  {32'h40bf0496, 32'h412116fa} /* (9, 12, 15) {real, imag} */,
  {32'hc0ebbbce, 32'hc138770c} /* (9, 12, 14) {real, imag} */,
  {32'hc0aaf2cb, 32'hc14c5bae} /* (9, 12, 13) {real, imag} */,
  {32'hc03e7ef6, 32'hbfa41738} /* (9, 12, 12) {real, imag} */,
  {32'h3e9b220c, 32'hc12be35e} /* (9, 12, 11) {real, imag} */,
  {32'hbfb0a1f2, 32'hc16b157b} /* (9, 12, 10) {real, imag} */,
  {32'h4065c818, 32'h3e7cf830} /* (9, 12, 9) {real, imag} */,
  {32'hc14c63c6, 32'hc1a1d086} /* (9, 12, 8) {real, imag} */,
  {32'hc1e01c02, 32'hc135a725} /* (9, 12, 7) {real, imag} */,
  {32'h402a00a1, 32'h40aabea6} /* (9, 12, 6) {real, imag} */,
  {32'h413a84b7, 32'h414be5c5} /* (9, 12, 5) {real, imag} */,
  {32'h41529958, 32'h407a9a4f} /* (9, 12, 4) {real, imag} */,
  {32'hc1a1b6f6, 32'hc10abe67} /* (9, 12, 3) {real, imag} */,
  {32'h411092e7, 32'hc0a6c0a6} /* (9, 12, 2) {real, imag} */,
  {32'h3fd60cd4, 32'hc1831d6e} /* (9, 12, 1) {real, imag} */,
  {32'h4003d0ff, 32'h41224e9a} /* (9, 12, 0) {real, imag} */,
  {32'hc1a247c5, 32'hc1688766} /* (9, 11, 31) {real, imag} */,
  {32'h407df1b8, 32'h408735ab} /* (9, 11, 30) {real, imag} */,
  {32'hbf021080, 32'h41982141} /* (9, 11, 29) {real, imag} */,
  {32'h4121d3e2, 32'hc178e4d4} /* (9, 11, 28) {real, imag} */,
  {32'h415c0d49, 32'h40c795b8} /* (9, 11, 27) {real, imag} */,
  {32'hc097c05a, 32'hbfa81e30} /* (9, 11, 26) {real, imag} */,
  {32'hc0dd9477, 32'hc0aa72a6} /* (9, 11, 25) {real, imag} */,
  {32'h40fc2b0e, 32'h41449334} /* (9, 11, 24) {real, imag} */,
  {32'h3f4b4390, 32'hc099fbe2} /* (9, 11, 23) {real, imag} */,
  {32'hbf825360, 32'h41907dd4} /* (9, 11, 22) {real, imag} */,
  {32'h412f3a78, 32'h4172a8d5} /* (9, 11, 21) {real, imag} */,
  {32'hc10f9c8c, 32'hc132e161} /* (9, 11, 20) {real, imag} */,
  {32'hc1981146, 32'h409d84ed} /* (9, 11, 19) {real, imag} */,
  {32'h3f3e5aa0, 32'hc07ab20c} /* (9, 11, 18) {real, imag} */,
  {32'hc149ee60, 32'hbf9f090b} /* (9, 11, 17) {real, imag} */,
  {32'h40cf5b26, 32'h41183972} /* (9, 11, 16) {real, imag} */,
  {32'h405d8ca2, 32'h40e71420} /* (9, 11, 15) {real, imag} */,
  {32'h3e586c00, 32'hc1f0445d} /* (9, 11, 14) {real, imag} */,
  {32'h40c45724, 32'hc185862d} /* (9, 11, 13) {real, imag} */,
  {32'h3f49d8f8, 32'hc0cad478} /* (9, 11, 12) {real, imag} */,
  {32'hc11f4117, 32'h416cdde4} /* (9, 11, 11) {real, imag} */,
  {32'hc0dc36e2, 32'h4037dd8a} /* (9, 11, 10) {real, imag} */,
  {32'hc1176cb5, 32'h3fd5a670} /* (9, 11, 9) {real, imag} */,
  {32'h3ee0aec0, 32'h4136c532} /* (9, 11, 8) {real, imag} */,
  {32'hc0a71438, 32'h4082fca2} /* (9, 11, 7) {real, imag} */,
  {32'h40bd3c41, 32'hc0e499dd} /* (9, 11, 6) {real, imag} */,
  {32'h3fdb916c, 32'h40ac8542} /* (9, 11, 5) {real, imag} */,
  {32'hc192aa7e, 32'hc0cc5c3a} /* (9, 11, 4) {real, imag} */,
  {32'h4128dac4, 32'h41434522} /* (9, 11, 3) {real, imag} */,
  {32'h4063d485, 32'hbfad276c} /* (9, 11, 2) {real, imag} */,
  {32'hc0e57d9a, 32'hc1729ca6} /* (9, 11, 1) {real, imag} */,
  {32'hc1be043d, 32'hc08cd588} /* (9, 11, 0) {real, imag} */,
  {32'h4190603d, 32'hc1202b35} /* (9, 10, 31) {real, imag} */,
  {32'h3fb6182e, 32'hc0e3a9f0} /* (9, 10, 30) {real, imag} */,
  {32'hbfe3c370, 32'h41302d04} /* (9, 10, 29) {real, imag} */,
  {32'hc1274539, 32'hc0b51160} /* (9, 10, 28) {real, imag} */,
  {32'hc080da64, 32'hbf970de8} /* (9, 10, 27) {real, imag} */,
  {32'h41038eeb, 32'hc0469cf6} /* (9, 10, 26) {real, imag} */,
  {32'hc1153db3, 32'h40509d0e} /* (9, 10, 25) {real, imag} */,
  {32'h40ffa908, 32'h4024b358} /* (9, 10, 24) {real, imag} */,
  {32'hbf62ec48, 32'hc136caa0} /* (9, 10, 23) {real, imag} */,
  {32'h40cf4308, 32'hc1237fa5} /* (9, 10, 22) {real, imag} */,
  {32'h41616c4a, 32'h4097a936} /* (9, 10, 21) {real, imag} */,
  {32'hbf615188, 32'h4141fef4} /* (9, 10, 20) {real, imag} */,
  {32'hc1a496b2, 32'hc094d05a} /* (9, 10, 19) {real, imag} */,
  {32'hc18de962, 32'hc10427ab} /* (9, 10, 18) {real, imag} */,
  {32'h3f28b8bc, 32'hc0f79e3b} /* (9, 10, 17) {real, imag} */,
  {32'hc0b79a71, 32'hbf2849d0} /* (9, 10, 16) {real, imag} */,
  {32'hc006e7d6, 32'hc09eccc1} /* (9, 10, 15) {real, imag} */,
  {32'h41b400d4, 32'h4189e9f0} /* (9, 10, 14) {real, imag} */,
  {32'hc1258c60, 32'hc17ed0e6} /* (9, 10, 13) {real, imag} */,
  {32'hc0b2f56f, 32'hc0104ae2} /* (9, 10, 12) {real, imag} */,
  {32'h40d00520, 32'hc10d35cc} /* (9, 10, 11) {real, imag} */,
  {32'hc1cf2a5b, 32'h3ecae300} /* (9, 10, 10) {real, imag} */,
  {32'h3f0a3250, 32'hc1931044} /* (9, 10, 9) {real, imag} */,
  {32'h411bd2ab, 32'h40cb51fd} /* (9, 10, 8) {real, imag} */,
  {32'h416ec109, 32'hc18b2f41} /* (9, 10, 7) {real, imag} */,
  {32'h40740717, 32'h3e5282e0} /* (9, 10, 6) {real, imag} */,
  {32'hc114ceee, 32'hc14e3614} /* (9, 10, 5) {real, imag} */,
  {32'hc15fd0b2, 32'h3f7c0638} /* (9, 10, 4) {real, imag} */,
  {32'h418c27ef, 32'hbedb2690} /* (9, 10, 3) {real, imag} */,
  {32'h402215a1, 32'h3f95223e} /* (9, 10, 2) {real, imag} */,
  {32'h41233d98, 32'h41732f6d} /* (9, 10, 1) {real, imag} */,
  {32'hc19d7a93, 32'h40c2dd4d} /* (9, 10, 0) {real, imag} */,
  {32'hc110f302, 32'h418b683c} /* (9, 9, 31) {real, imag} */,
  {32'hc0fd5536, 32'hc1b01132} /* (9, 9, 30) {real, imag} */,
  {32'h413408a2, 32'h40ea9ccc} /* (9, 9, 29) {real, imag} */,
  {32'hc08fa26c, 32'h400d6e22} /* (9, 9, 28) {real, imag} */,
  {32'hc0721c05, 32'h41497cd5} /* (9, 9, 27) {real, imag} */,
  {32'hc088eafd, 32'hbff8cb20} /* (9, 9, 26) {real, imag} */,
  {32'h40ea2840, 32'hc013f88f} /* (9, 9, 25) {real, imag} */,
  {32'hc13ae645, 32'hc10b0e76} /* (9, 9, 24) {real, imag} */,
  {32'h404aad82, 32'hc0cde7fe} /* (9, 9, 23) {real, imag} */,
  {32'h40a63dcc, 32'hc134c2ee} /* (9, 9, 22) {real, imag} */,
  {32'hc13f1268, 32'hc06e6bd5} /* (9, 9, 21) {real, imag} */,
  {32'hc04dde10, 32'h40158a28} /* (9, 9, 20) {real, imag} */,
  {32'hc18e3a41, 32'h41b287f4} /* (9, 9, 19) {real, imag} */,
  {32'h40d511a0, 32'h3f40d170} /* (9, 9, 18) {real, imag} */,
  {32'hbfbaa008, 32'h40c22151} /* (9, 9, 17) {real, imag} */,
  {32'h412d974e, 32'h3fcffaca} /* (9, 9, 16) {real, imag} */,
  {32'h406513d3, 32'hc1468d6e} /* (9, 9, 15) {real, imag} */,
  {32'h3feab22c, 32'h3f847d0a} /* (9, 9, 14) {real, imag} */,
  {32'hc0f8d97a, 32'h41391768} /* (9, 9, 13) {real, imag} */,
  {32'hc136e39d, 32'h3f8e6c98} /* (9, 9, 12) {real, imag} */,
  {32'hbf769a34, 32'hc113a178} /* (9, 9, 11) {real, imag} */,
  {32'h41c839b3, 32'h412276db} /* (9, 9, 10) {real, imag} */,
  {32'hc12b39a1, 32'hc04f7b6e} /* (9, 9, 9) {real, imag} */,
  {32'h413fc2e9, 32'hc18a8aa8} /* (9, 9, 8) {real, imag} */,
  {32'hc0ebc9de, 32'h418f8dec} /* (9, 9, 7) {real, imag} */,
  {32'hc115a206, 32'h414027aa} /* (9, 9, 6) {real, imag} */,
  {32'hc1948df5, 32'hc03c8e90} /* (9, 9, 5) {real, imag} */,
  {32'hc1939144, 32'h41481848} /* (9, 9, 4) {real, imag} */,
  {32'h41290906, 32'h413ff948} /* (9, 9, 3) {real, imag} */,
  {32'h4168f3cc, 32'hc13b5eb7} /* (9, 9, 2) {real, imag} */,
  {32'h41d1964f, 32'hc107fbde} /* (9, 9, 1) {real, imag} */,
  {32'h41081a94, 32'hc1820bc7} /* (9, 9, 0) {real, imag} */,
  {32'hc22b9308, 32'hc1b21bbd} /* (9, 8, 31) {real, imag} */,
  {32'h41f9c2d7, 32'h4115260e} /* (9, 8, 30) {real, imag} */,
  {32'h4010dde7, 32'hc163fc8c} /* (9, 8, 29) {real, imag} */,
  {32'h41079894, 32'h41f35b23} /* (9, 8, 28) {real, imag} */,
  {32'h40065b38, 32'hbf1a3428} /* (9, 8, 27) {real, imag} */,
  {32'h409461b4, 32'hc18e0432} /* (9, 8, 26) {real, imag} */,
  {32'h40d15f48, 32'hc082ce15} /* (9, 8, 25) {real, imag} */,
  {32'hc0101b68, 32'hc12be38c} /* (9, 8, 24) {real, imag} */,
  {32'hc1c4f950, 32'hc0a151ce} /* (9, 8, 23) {real, imag} */,
  {32'hc105869f, 32'h411d33b8} /* (9, 8, 22) {real, imag} */,
  {32'hc06f0b20, 32'h416af8cc} /* (9, 8, 21) {real, imag} */,
  {32'h3f76592c, 32'hc0638db1} /* (9, 8, 20) {real, imag} */,
  {32'hbf5575a0, 32'h409d2aef} /* (9, 8, 19) {real, imag} */,
  {32'h40b43d0d, 32'h40f1d7cb} /* (9, 8, 18) {real, imag} */,
  {32'hc11cf51d, 32'hc187981c} /* (9, 8, 17) {real, imag} */,
  {32'h41284177, 32'h4008d2f0} /* (9, 8, 16) {real, imag} */,
  {32'hc1055741, 32'h3dbde780} /* (9, 8, 15) {real, imag} */,
  {32'hc0b60709, 32'h4130e052} /* (9, 8, 14) {real, imag} */,
  {32'h400e1b4c, 32'hc0d31e45} /* (9, 8, 13) {real, imag} */,
  {32'hc142ac24, 32'hc014dad1} /* (9, 8, 12) {real, imag} */,
  {32'hc0a638de, 32'hc0491660} /* (9, 8, 11) {real, imag} */,
  {32'hc0cd28c2, 32'h406d0bb8} /* (9, 8, 10) {real, imag} */,
  {32'h405726ba, 32'h4138668b} /* (9, 8, 9) {real, imag} */,
  {32'hc156b7f6, 32'h4193374b} /* (9, 8, 8) {real, imag} */,
  {32'h41687c3a, 32'h4207439c} /* (9, 8, 7) {real, imag} */,
  {32'hc0b35e82, 32'h3f9467ec} /* (9, 8, 6) {real, imag} */,
  {32'h41a1bb48, 32'hc02a1284} /* (9, 8, 5) {real, imag} */,
  {32'h40e59cee, 32'h40604ecc} /* (9, 8, 4) {real, imag} */,
  {32'hbf34bb00, 32'h4137909a} /* (9, 8, 3) {real, imag} */,
  {32'h40db9691, 32'hc126c05a} /* (9, 8, 2) {real, imag} */,
  {32'hc0c09db9, 32'hc18e2ef2} /* (9, 8, 1) {real, imag} */,
  {32'hc20b388c, 32'hc141f294} /* (9, 8, 0) {real, imag} */,
  {32'h418d0f0b, 32'h414206ed} /* (9, 7, 31) {real, imag} */,
  {32'h3f3320f0, 32'hc1c56090} /* (9, 7, 30) {real, imag} */,
  {32'hc100d1fe, 32'h41008979} /* (9, 7, 29) {real, imag} */,
  {32'hc105b476, 32'hc0dcacf0} /* (9, 7, 28) {real, imag} */,
  {32'hc1a64e32, 32'h411998ba} /* (9, 7, 27) {real, imag} */,
  {32'hc01429f6, 32'h400b1ec8} /* (9, 7, 26) {real, imag} */,
  {32'hc095c019, 32'hc15a9bc7} /* (9, 7, 25) {real, imag} */,
  {32'hbfa03af8, 32'hc1a9dd94} /* (9, 7, 24) {real, imag} */,
  {32'hc1bf03b2, 32'hc024b61c} /* (9, 7, 23) {real, imag} */,
  {32'h408fe90a, 32'h4134339a} /* (9, 7, 22) {real, imag} */,
  {32'hc10f11e6, 32'hc069ed31} /* (9, 7, 21) {real, imag} */,
  {32'h40efbfe4, 32'h41356422} /* (9, 7, 20) {real, imag} */,
  {32'h41320fea, 32'h412917ba} /* (9, 7, 19) {real, imag} */,
  {32'h4025c396, 32'hc0ea10f6} /* (9, 7, 18) {real, imag} */,
  {32'h412eb7af, 32'h400ed740} /* (9, 7, 17) {real, imag} */,
  {32'hc010a314, 32'hc034c2ca} /* (9, 7, 16) {real, imag} */,
  {32'hc144446e, 32'h408ac34c} /* (9, 7, 15) {real, imag} */,
  {32'hc18d5daf, 32'h4027a090} /* (9, 7, 14) {real, imag} */,
  {32'h40d1304a, 32'hc1aa97e8} /* (9, 7, 13) {real, imag} */,
  {32'hc10702ef, 32'h3f9d1b9a} /* (9, 7, 12) {real, imag} */,
  {32'h40ce1327, 32'h4098c76a} /* (9, 7, 11) {real, imag} */,
  {32'h41278658, 32'hc0e51bba} /* (9, 7, 10) {real, imag} */,
  {32'h40fd5ab0, 32'h418c4f5b} /* (9, 7, 9) {real, imag} */,
  {32'hc1337814, 32'h40bb3a40} /* (9, 7, 8) {real, imag} */,
  {32'h40fc3dca, 32'hc1365872} /* (9, 7, 7) {real, imag} */,
  {32'h3f6893f0, 32'hc11cf9f4} /* (9, 7, 6) {real, imag} */,
  {32'h41ae0abc, 32'h4081ccb5} /* (9, 7, 5) {real, imag} */,
  {32'h4026d8df, 32'h41180da2} /* (9, 7, 4) {real, imag} */,
  {32'hbff318cc, 32'h40a4c9dc} /* (9, 7, 3) {real, imag} */,
  {32'hc1154f9d, 32'hc1d0af36} /* (9, 7, 2) {real, imag} */,
  {32'h3e28d720, 32'h41b46930} /* (9, 7, 1) {real, imag} */,
  {32'hc093b8dd, 32'h40b92cb6} /* (9, 7, 0) {real, imag} */,
  {32'h40106338, 32'h416c182d} /* (9, 6, 31) {real, imag} */,
  {32'h410c098d, 32'h40a5c617} /* (9, 6, 30) {real, imag} */,
  {32'hbcf10200, 32'h415c52b8} /* (9, 6, 29) {real, imag} */,
  {32'h41b9c2ba, 32'hc1a820c9} /* (9, 6, 28) {real, imag} */,
  {32'hc0adf51d, 32'hc07f1a2c} /* (9, 6, 27) {real, imag} */,
  {32'h41b1d271, 32'h41a78c22} /* (9, 6, 26) {real, imag} */,
  {32'hc121ca64, 32'h3f9de6e6} /* (9, 6, 25) {real, imag} */,
  {32'hc0918b75, 32'h4041bd62} /* (9, 6, 24) {real, imag} */,
  {32'h40c95adb, 32'h413dbd84} /* (9, 6, 23) {real, imag} */,
  {32'h40d95fcf, 32'hc142d8b2} /* (9, 6, 22) {real, imag} */,
  {32'h4103c4a6, 32'h41146f09} /* (9, 6, 21) {real, imag} */,
  {32'h3f3c3738, 32'h4062e628} /* (9, 6, 20) {real, imag} */,
  {32'h40d7ff22, 32'hc10faeaa} /* (9, 6, 19) {real, imag} */,
  {32'h404e8858, 32'h41247d7c} /* (9, 6, 18) {real, imag} */,
  {32'hc0bc3bb4, 32'h40f3f20d} /* (9, 6, 17) {real, imag} */,
  {32'hc1297b59, 32'hc0171e7e} /* (9, 6, 16) {real, imag} */,
  {32'h411278fa, 32'h4088cb0a} /* (9, 6, 15) {real, imag} */,
  {32'hc09861d8, 32'hc0a31c67} /* (9, 6, 14) {real, imag} */,
  {32'hbec60770, 32'h3ff850f4} /* (9, 6, 13) {real, imag} */,
  {32'hc182cfed, 32'h414014dc} /* (9, 6, 12) {real, imag} */,
  {32'h415ff534, 32'h41b1599c} /* (9, 6, 11) {real, imag} */,
  {32'hc05745cc, 32'h41a96a98} /* (9, 6, 10) {real, imag} */,
  {32'hbfe8a5fc, 32'h406432de} /* (9, 6, 9) {real, imag} */,
  {32'h40dd23a8, 32'hc1234e5d} /* (9, 6, 8) {real, imag} */,
  {32'h40c2633a, 32'h40b02450} /* (9, 6, 7) {real, imag} */,
  {32'h4156bd63, 32'h41006a9d} /* (9, 6, 6) {real, imag} */,
  {32'h40e7392e, 32'hbe56fd80} /* (9, 6, 5) {real, imag} */,
  {32'h413292da, 32'hbfc10dc0} /* (9, 6, 4) {real, imag} */,
  {32'hc0e07254, 32'hc0cd7805} /* (9, 6, 3) {real, imag} */,
  {32'hc1dffff6, 32'hc1c0c6d2} /* (9, 6, 2) {real, imag} */,
  {32'h41290938, 32'h411a57f6} /* (9, 6, 1) {real, imag} */,
  {32'h401f004c, 32'h419194ac} /* (9, 6, 0) {real, imag} */,
  {32'hc2d1ec08, 32'hc081e296} /* (9, 5, 31) {real, imag} */,
  {32'h41848bb4, 32'hc107af27} /* (9, 5, 30) {real, imag} */,
  {32'h419c6dff, 32'h4145efd5} /* (9, 5, 29) {real, imag} */,
  {32'hc105b0bb, 32'h3fbb7200} /* (9, 5, 28) {real, imag} */,
  {32'hc07b17c8, 32'h41109960} /* (9, 5, 27) {real, imag} */,
  {32'h412c16aa, 32'h41c38d36} /* (9, 5, 26) {real, imag} */,
  {32'hc0ac7bdc, 32'h41a11e4b} /* (9, 5, 25) {real, imag} */,
  {32'h413d15c2, 32'hc0089c91} /* (9, 5, 24) {real, imag} */,
  {32'h411501cb, 32'h3f3aa684} /* (9, 5, 23) {real, imag} */,
  {32'hc1b3b325, 32'hbe4d0100} /* (9, 5, 22) {real, imag} */,
  {32'h412b022b, 32'h400c35a6} /* (9, 5, 21) {real, imag} */,
  {32'hc11141a3, 32'hc07477c2} /* (9, 5, 20) {real, imag} */,
  {32'hc15efd1a, 32'h4128249b} /* (9, 5, 19) {real, imag} */,
  {32'h3fd9e90c, 32'hc007e700} /* (9, 5, 18) {real, imag} */,
  {32'hc067b16a, 32'h40eed38f} /* (9, 5, 17) {real, imag} */,
  {32'h413dd0d8, 32'h3ebd9e50} /* (9, 5, 16) {real, imag} */,
  {32'h40d26ddc, 32'h3ee436b4} /* (9, 5, 15) {real, imag} */,
  {32'h411496c4, 32'hbf5ce59c} /* (9, 5, 14) {real, imag} */,
  {32'hc0284551, 32'h3ff54bd0} /* (9, 5, 13) {real, imag} */,
  {32'hbf9b9978, 32'h3fa2a30f} /* (9, 5, 12) {real, imag} */,
  {32'hc00cb252, 32'h418f4ff0} /* (9, 5, 11) {real, imag} */,
  {32'h400fa0ac, 32'h41e81e0d} /* (9, 5, 10) {real, imag} */,
  {32'h40a298c5, 32'hc0c41566} /* (9, 5, 9) {real, imag} */,
  {32'hbe003680, 32'hbfc9e728} /* (9, 5, 8) {real, imag} */,
  {32'hc0832666, 32'hc16c7b3a} /* (9, 5, 7) {real, imag} */,
  {32'hc09e2312, 32'h412b7902} /* (9, 5, 6) {real, imag} */,
  {32'h421b9724, 32'h413d4d47} /* (9, 5, 5) {real, imag} */,
  {32'hc130a827, 32'hc09f1190} /* (9, 5, 4) {real, imag} */,
  {32'hc1edfd25, 32'hc141ee4b} /* (9, 5, 3) {real, imag} */,
  {32'h41faff09, 32'h421ee39a} /* (9, 5, 2) {real, imag} */,
  {32'hc20e53da, 32'hc2983dde} /* (9, 5, 1) {real, imag} */,
  {32'hc259bfcc, 32'hc1efe0a2} /* (9, 5, 0) {real, imag} */,
  {32'h41b382f6, 32'h42cc40c4} /* (9, 4, 31) {real, imag} */,
  {32'hc2bb769c, 32'hc298c6ae} /* (9, 4, 30) {real, imag} */,
  {32'hc1535150, 32'hc11a7a75} /* (9, 4, 29) {real, imag} */,
  {32'h4203af83, 32'h40b7006e} /* (9, 4, 28) {real, imag} */,
  {32'hc1af5c3e, 32'hc1be297f} /* (9, 4, 27) {real, imag} */,
  {32'hc15d4d0a, 32'h4128cd71} /* (9, 4, 26) {real, imag} */,
  {32'h405b1766, 32'h418c45ad} /* (9, 4, 25) {real, imag} */,
  {32'h40816374, 32'hc14259ce} /* (9, 4, 24) {real, imag} */,
  {32'h4165f52a, 32'hc00ffaf8} /* (9, 4, 23) {real, imag} */,
  {32'hc0df5969, 32'hc08ba6f6} /* (9, 4, 22) {real, imag} */,
  {32'hc0238ece, 32'h41b2aba0} /* (9, 4, 21) {real, imag} */,
  {32'h4174b962, 32'hc0112bfa} /* (9, 4, 20) {real, imag} */,
  {32'hc15f7d20, 32'hc1824abc} /* (9, 4, 19) {real, imag} */,
  {32'hc107a3f4, 32'hc01d2ee4} /* (9, 4, 18) {real, imag} */,
  {32'h4118a53c, 32'hc0a1dc22} /* (9, 4, 17) {real, imag} */,
  {32'hc0c7b2e5, 32'h3fdba0e2} /* (9, 4, 16) {real, imag} */,
  {32'h40a2a01a, 32'h4080f911} /* (9, 4, 15) {real, imag} */,
  {32'h3fad2042, 32'hc0bdc6a5} /* (9, 4, 14) {real, imag} */,
  {32'hc08c0e3e, 32'hc0afb75a} /* (9, 4, 13) {real, imag} */,
  {32'hc1d897d5, 32'h410eb4ec} /* (9, 4, 12) {real, imag} */,
  {32'h40da790f, 32'hc12d6fdd} /* (9, 4, 11) {real, imag} */,
  {32'h411ae7a4, 32'h408fb2c9} /* (9, 4, 10) {real, imag} */,
  {32'h40b25510, 32'hc08f40c4} /* (9, 4, 9) {real, imag} */,
  {32'hc115bbe0, 32'hc11c68a3} /* (9, 4, 8) {real, imag} */,
  {32'hbfdeb5e0, 32'hc17fa0e4} /* (9, 4, 7) {real, imag} */,
  {32'h41bd1858, 32'hc01e1364} /* (9, 4, 6) {real, imag} */,
  {32'hc0d00e40, 32'hc1d059f2} /* (9, 4, 5) {real, imag} */,
  {32'h416aa38e, 32'h419dab8d} /* (9, 4, 4) {real, imag} */,
  {32'hc21c4e87, 32'h42532e9c} /* (9, 4, 3) {real, imag} */,
  {32'hc24694f6, 32'hc2a88ca7} /* (9, 4, 2) {real, imag} */,
  {32'h430dff05, 32'h42094c94} /* (9, 4, 1) {real, imag} */,
  {32'h4214a618, 32'h41c19450} /* (9, 4, 0) {real, imag} */,
  {32'hc2feea4c, 32'h42278557} /* (9, 3, 31) {real, imag} */,
  {32'h428a0160, 32'hc32a8cc7} /* (9, 3, 30) {real, imag} */,
  {32'h3fd336b4, 32'h41eb199d} /* (9, 3, 29) {real, imag} */,
  {32'h41ef50c3, 32'h4081faa6} /* (9, 3, 28) {real, imag} */,
  {32'hc224ce6e, 32'hc13a1917} /* (9, 3, 27) {real, imag} */,
  {32'h3f94d3d8, 32'h415a4ed6} /* (9, 3, 26) {real, imag} */,
  {32'hc1922f2b, 32'hc0c2ea38} /* (9, 3, 25) {real, imag} */,
  {32'h418ce24b, 32'hc190014e} /* (9, 3, 24) {real, imag} */,
  {32'hc0dacbc2, 32'h410e4e75} /* (9, 3, 23) {real, imag} */,
  {32'hc13fc771, 32'h3f543014} /* (9, 3, 22) {real, imag} */,
  {32'hc09bd94e, 32'hc135716c} /* (9, 3, 21) {real, imag} */,
  {32'h40b5d577, 32'h403ea28a} /* (9, 3, 20) {real, imag} */,
  {32'h412ac4d1, 32'hc0068634} /* (9, 3, 19) {real, imag} */,
  {32'h4119840e, 32'h409a57d2} /* (9, 3, 18) {real, imag} */,
  {32'h40a98de0, 32'hc13cb9e8} /* (9, 3, 17) {real, imag} */,
  {32'h404f2860, 32'hc0cc41ff} /* (9, 3, 16) {real, imag} */,
  {32'h411df930, 32'h41096487} /* (9, 3, 15) {real, imag} */,
  {32'hc0af22ad, 32'h40b4f981} /* (9, 3, 14) {real, imag} */,
  {32'hc04b693a, 32'h40eca620} /* (9, 3, 13) {real, imag} */,
  {32'h41601a8e, 32'h40d0f065} /* (9, 3, 12) {real, imag} */,
  {32'hc045076c, 32'hbf965254} /* (9, 3, 11) {real, imag} */,
  {32'hc13cffc4, 32'h41562576} /* (9, 3, 10) {real, imag} */,
  {32'hbdec5a10, 32'h40c0f446} /* (9, 3, 9) {real, imag} */,
  {32'hc1cb02f4, 32'h41248d92} /* (9, 3, 8) {real, imag} */,
  {32'hc103746e, 32'hc0b77d52} /* (9, 3, 7) {real, imag} */,
  {32'hbf12e8c0, 32'h41a8b76b} /* (9, 3, 6) {real, imag} */,
  {32'hc0d9758c, 32'h40782040} /* (9, 3, 5) {real, imag} */,
  {32'hc22221b2, 32'h407ff548} /* (9, 3, 4) {real, imag} */,
  {32'hc1f177e0, 32'h4108571a} /* (9, 3, 3) {real, imag} */,
  {32'hbf5755c0, 32'hc2ca9267} /* (9, 3, 2) {real, imag} */,
  {32'h42c52f9a, 32'h42d115a2} /* (9, 3, 1) {real, imag} */,
  {32'hc120eb90, 32'hc1e257cc} /* (9, 3, 0) {real, imag} */,
  {32'hc4a2fd64, 32'hc242606e} /* (9, 2, 31) {real, imag} */,
  {32'h440f54ac, 32'hc33538f6} /* (9, 2, 30) {real, imag} */,
  {32'h419a4284, 32'h4230401d} /* (9, 2, 29) {real, imag} */,
  {32'hc186c26b, 32'h4292eebb} /* (9, 2, 28) {real, imag} */,
  {32'h42abba8f, 32'hc20fb289} /* (9, 2, 27) {real, imag} */,
  {32'h41540f24, 32'hc19890a7} /* (9, 2, 26) {real, imag} */,
  {32'hc119d8cb, 32'hc0cb52c9} /* (9, 2, 25) {real, imag} */,
  {32'h41effc58, 32'hc196d7ef} /* (9, 2, 24) {real, imag} */,
  {32'h4135e4b7, 32'h4190bdaf} /* (9, 2, 23) {real, imag} */,
  {32'h3f838d64, 32'h40619436} /* (9, 2, 22) {real, imag} */,
  {32'hc0fb4764, 32'h3cc078c0} /* (9, 2, 21) {real, imag} */,
  {32'hc03b6334, 32'h40aabf42} /* (9, 2, 20) {real, imag} */,
  {32'h40c26e5c, 32'hc0937cb0} /* (9, 2, 19) {real, imag} */,
  {32'hbff7cdf2, 32'hc1e3eb3d} /* (9, 2, 18) {real, imag} */,
  {32'hc0930a8a, 32'h3fc7aecc} /* (9, 2, 17) {real, imag} */,
  {32'h40deddd0, 32'hc09b5aa5} /* (9, 2, 16) {real, imag} */,
  {32'hc03a2220, 32'hc12c8000} /* (9, 2, 15) {real, imag} */,
  {32'hc02ec384, 32'h40b2e074} /* (9, 2, 14) {real, imag} */,
  {32'h4047ec5c, 32'hbf1b9480} /* (9, 2, 13) {real, imag} */,
  {32'h411d3200, 32'hc0bca626} /* (9, 2, 12) {real, imag} */,
  {32'h410e2894, 32'h4127577c} /* (9, 2, 11) {real, imag} */,
  {32'hc17fd13e, 32'hc1470152} /* (9, 2, 10) {real, imag} */,
  {32'h411d899e, 32'h4134fd31} /* (9, 2, 9) {real, imag} */,
  {32'h4190afbf, 32'h411f2e7b} /* (9, 2, 8) {real, imag} */,
  {32'hc1df366c, 32'hbf8f0c70} /* (9, 2, 7) {real, imag} */,
  {32'h4182dcee, 32'hc1337d9d} /* (9, 2, 6) {real, imag} */,
  {32'h42390c3a, 32'h4231fd35} /* (9, 2, 5) {real, imag} */,
  {32'hc2b8aad1, 32'hc24ab37a} /* (9, 2, 4) {real, imag} */,
  {32'hc18dac46, 32'h412f5658} /* (9, 2, 3) {real, imag} */,
  {32'h43d8527b, 32'hc2ec34d2} /* (9, 2, 2) {real, imag} */,
  {32'hc432a101, 32'h43446f42} /* (9, 2, 1) {real, imag} */,
  {32'hc42ff663, 32'hc300b112} /* (9, 2, 0) {real, imag} */,
  {32'h44d2283a, 32'hc3d3f00b} /* (9, 1, 31) {real, imag} */,
  {32'hc3bbee4a, 32'h428e708b} /* (9, 1, 30) {real, imag} */,
  {32'hc2336371, 32'hc1a2051b} /* (9, 1, 29) {real, imag} */,
  {32'h429d877b, 32'h42c0738a} /* (9, 1, 28) {real, imag} */,
  {32'hc2a95a45, 32'hc1dc97f4} /* (9, 1, 27) {real, imag} */,
  {32'hc1a08e7c, 32'hc1389bdc} /* (9, 1, 26) {real, imag} */,
  {32'h42167626, 32'hc1b868f7} /* (9, 1, 25) {real, imag} */,
  {32'hc1e9ef22, 32'h4071dc1c} /* (9, 1, 24) {real, imag} */,
  {32'h414aca9c, 32'h3f245c50} /* (9, 1, 23) {real, imag} */,
  {32'hc05acc0c, 32'h40aadedc} /* (9, 1, 22) {real, imag} */,
  {32'hc1dd6582, 32'h4134f38a} /* (9, 1, 21) {real, imag} */,
  {32'h4124890c, 32'h410d52f6} /* (9, 1, 20) {real, imag} */,
  {32'h40898cc8, 32'hc123a916} /* (9, 1, 19) {real, imag} */,
  {32'hc1830a4a, 32'h41c43cca} /* (9, 1, 18) {real, imag} */,
  {32'h3e961ec4, 32'h3fc0c49c} /* (9, 1, 17) {real, imag} */,
  {32'hc010715f, 32'h40fc766a} /* (9, 1, 16) {real, imag} */,
  {32'hc15aedf0, 32'h408217d0} /* (9, 1, 15) {real, imag} */,
  {32'h405ad65a, 32'hc110be98} /* (9, 1, 14) {real, imag} */,
  {32'h4148b3bf, 32'hbf636a60} /* (9, 1, 13) {real, imag} */,
  {32'h40fcdd38, 32'hc18a3c1d} /* (9, 1, 12) {real, imag} */,
  {32'h404ec3a4, 32'hc1a40c9a} /* (9, 1, 11) {real, imag} */,
  {32'hc1a6cade, 32'hc173b006} /* (9, 1, 10) {real, imag} */,
  {32'h3ec65ae0, 32'h41377dbe} /* (9, 1, 9) {real, imag} */,
  {32'hc112a991, 32'hc1d873d2} /* (9, 1, 8) {real, imag} */,
  {32'h4187fa93, 32'hc0bfd081} /* (9, 1, 7) {real, imag} */,
  {32'hc21272ca, 32'hc15bcfb1} /* (9, 1, 6) {real, imag} */,
  {32'hc2b88f86, 32'hc1b5d8cf} /* (9, 1, 5) {real, imag} */,
  {32'h428c7824, 32'h41210898} /* (9, 1, 4) {real, imag} */,
  {32'hc1775210, 32'h416dedac} /* (9, 1, 3) {real, imag} */,
  {32'hc41b750a, 32'hc40b2cf5} /* (9, 1, 2) {real, imag} */,
  {32'h4519b1b4, 32'h44a09d10} /* (9, 1, 1) {real, imag} */,
  {32'h45105eca, 32'h435c289a} /* (9, 1, 0) {real, imag} */,
  {32'h44b18a4e, 32'hc4902210} /* (9, 0, 31) {real, imag} */,
  {32'hc33ae13a, 32'h43bc3442} /* (9, 0, 30) {real, imag} */,
  {32'hc253a414, 32'h41dcb57c} /* (9, 0, 29) {real, imag} */,
  {32'hc10003ec, 32'h404d0380} /* (9, 0, 28) {real, imag} */,
  {32'hc26b67c0, 32'hc07d899a} /* (9, 0, 27) {real, imag} */,
  {32'h410a8180, 32'hc0d28827} /* (9, 0, 26) {real, imag} */,
  {32'h412e9e63, 32'h4021af90} /* (9, 0, 25) {real, imag} */,
  {32'h41221586, 32'h4231fbf0} /* (9, 0, 24) {real, imag} */,
  {32'hbf0879f0, 32'hc15ca9bf} /* (9, 0, 23) {real, imag} */,
  {32'h414c5986, 32'h419ee578} /* (9, 0, 22) {real, imag} */,
  {32'hc1618145, 32'hc1522b5c} /* (9, 0, 21) {real, imag} */,
  {32'h40c8c07d, 32'hc05e21d0} /* (9, 0, 20) {real, imag} */,
  {32'h410e02ac, 32'hc16be810} /* (9, 0, 19) {real, imag} */,
  {32'h3f06d4b4, 32'h4152962c} /* (9, 0, 18) {real, imag} */,
  {32'hc14a8a4a, 32'hc0770406} /* (9, 0, 17) {real, imag} */,
  {32'h40c1a47e, 32'h00000000} /* (9, 0, 16) {real, imag} */,
  {32'hc14a8a4a, 32'h40770406} /* (9, 0, 15) {real, imag} */,
  {32'h3f06d4b4, 32'hc152962c} /* (9, 0, 14) {real, imag} */,
  {32'h410e02ac, 32'h416be810} /* (9, 0, 13) {real, imag} */,
  {32'h40c8c07d, 32'h405e21d0} /* (9, 0, 12) {real, imag} */,
  {32'hc1618145, 32'h41522b5c} /* (9, 0, 11) {real, imag} */,
  {32'h414c5986, 32'hc19ee578} /* (9, 0, 10) {real, imag} */,
  {32'hbf0879f0, 32'h415ca9bf} /* (9, 0, 9) {real, imag} */,
  {32'h41221586, 32'hc231fbf0} /* (9, 0, 8) {real, imag} */,
  {32'h412e9e63, 32'hc021af90} /* (9, 0, 7) {real, imag} */,
  {32'h410a8180, 32'h40d28827} /* (9, 0, 6) {real, imag} */,
  {32'hc26b67c0, 32'h407d899a} /* (9, 0, 5) {real, imag} */,
  {32'hc10003ec, 32'hc04d0380} /* (9, 0, 4) {real, imag} */,
  {32'hc253a414, 32'hc1dcb57c} /* (9, 0, 3) {real, imag} */,
  {32'hc33ae13a, 32'hc3bc3442} /* (9, 0, 2) {real, imag} */,
  {32'h44b18a4e, 32'h44902210} /* (9, 0, 1) {real, imag} */,
  {32'h45166e52, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h450bb595, 32'hc48a3849} /* (8, 31, 31) {real, imag} */,
  {32'hc40af8a8, 32'h4401b2e0} /* (8, 31, 30) {real, imag} */,
  {32'hc21060a1, 32'h42435b96} /* (8, 31, 29) {real, imag} */,
  {32'h42699c56, 32'h41835cb3} /* (8, 31, 28) {real, imag} */,
  {32'hc29f7400, 32'h41a6fb00} /* (8, 31, 27) {real, imag} */,
  {32'hc1d6180e, 32'h4069fab4} /* (8, 31, 26) {real, imag} */,
  {32'h412e5da6, 32'hc149af36} /* (8, 31, 25) {real, imag} */,
  {32'hc01f0128, 32'h41e99d99} /* (8, 31, 24) {real, imag} */,
  {32'hc109eb2a, 32'h418b9a8a} /* (8, 31, 23) {real, imag} */,
  {32'hc1bdb8a6, 32'h40cda082} /* (8, 31, 22) {real, imag} */,
  {32'hc1114d2c, 32'h41aec71a} /* (8, 31, 21) {real, imag} */,
  {32'h3fbe162c, 32'h419ccdf0} /* (8, 31, 20) {real, imag} */,
  {32'h40670ff6, 32'h3f8e4e50} /* (8, 31, 19) {real, imag} */,
  {32'h40e556b2, 32'h418606e2} /* (8, 31, 18) {real, imag} */,
  {32'h4087c8b9, 32'hc11b5098} /* (8, 31, 17) {real, imag} */,
  {32'h409f1e63, 32'hbf77e51e} /* (8, 31, 16) {real, imag} */,
  {32'hc01f94a6, 32'hbf31bf3c} /* (8, 31, 15) {real, imag} */,
  {32'hc12a4c87, 32'hc1989ca2} /* (8, 31, 14) {real, imag} */,
  {32'hc03c7b21, 32'h409ef37c} /* (8, 31, 13) {real, imag} */,
  {32'h414e6234, 32'h41a20ee9} /* (8, 31, 12) {real, imag} */,
  {32'hc22e581e, 32'hc0c9eff2} /* (8, 31, 11) {real, imag} */,
  {32'h400cc0b8, 32'hc0dbd85f} /* (8, 31, 10) {real, imag} */,
  {32'h40933ae0, 32'hc15d209e} /* (8, 31, 9) {real, imag} */,
  {32'hc211bc7d, 32'h3ea24140} /* (8, 31, 8) {real, imag} */,
  {32'h4195d823, 32'h415cee22} /* (8, 31, 7) {real, imag} */,
  {32'hc19807b8, 32'hc12ed425} /* (8, 31, 6) {real, imag} */,
  {32'hc2b5cc2c, 32'h4123a32d} /* (8, 31, 5) {real, imag} */,
  {32'h428394cd, 32'hc2a07ef2} /* (8, 31, 4) {real, imag} */,
  {32'hc100a106, 32'h40fe2978} /* (8, 31, 3) {real, imag} */,
  {32'hc3ab8065, 32'hc2969374} /* (8, 31, 2) {real, imag} */,
  {32'h44c3e72d, 32'h43c6ca94} /* (8, 31, 1) {real, imag} */,
  {32'h4504ce84, 32'hc36653ae} /* (8, 31, 0) {real, imag} */,
  {32'hc4203dbc, 32'hc3212c7c} /* (8, 30, 31) {real, imag} */,
  {32'h43cce94e, 32'h42ad8e00} /* (8, 30, 30) {real, imag} */,
  {32'hc1e50215, 32'hc0602560} /* (8, 30, 29) {real, imag} */,
  {32'hc2d758c2, 32'h41c3bede} /* (8, 30, 28) {real, imag} */,
  {32'h428c6076, 32'hc1dbbdea} /* (8, 30, 27) {real, imag} */,
  {32'h3fe42078, 32'hc0e0be35} /* (8, 30, 26) {real, imag} */,
  {32'hc190a884, 32'h42039adc} /* (8, 30, 25) {real, imag} */,
  {32'hc08f4426, 32'hc0018f42} /* (8, 30, 24) {real, imag} */,
  {32'h416c9750, 32'hc0e19701} /* (8, 30, 23) {real, imag} */,
  {32'hc0bbccc2, 32'h3f6216b0} /* (8, 30, 22) {real, imag} */,
  {32'hbfda6a86, 32'hc15848fc} /* (8, 30, 21) {real, imag} */,
  {32'h4153a7cb, 32'h4131c74c} /* (8, 30, 20) {real, imag} */,
  {32'h411e21f4, 32'h40e13645} /* (8, 30, 19) {real, imag} */,
  {32'hc0fced45, 32'hc1075247} /* (8, 30, 18) {real, imag} */,
  {32'hc148bf24, 32'hc0d7b4b5} /* (8, 30, 17) {real, imag} */,
  {32'hc121e42e, 32'hc11acf0c} /* (8, 30, 16) {real, imag} */,
  {32'h418739ba, 32'hc11d214c} /* (8, 30, 15) {real, imag} */,
  {32'hc11a609b, 32'h3ea83950} /* (8, 30, 14) {real, imag} */,
  {32'h3f0e9734, 32'h4130bbed} /* (8, 30, 13) {real, imag} */,
  {32'h4178535d, 32'h41cf1b82} /* (8, 30, 12) {real, imag} */,
  {32'hc107f4f8, 32'h40fc9800} /* (8, 30, 11) {real, imag} */,
  {32'hc1152825, 32'h406b0078} /* (8, 30, 10) {real, imag} */,
  {32'hc10e917f, 32'h401d929a} /* (8, 30, 9) {real, imag} */,
  {32'h41958887, 32'hbd0cca00} /* (8, 30, 8) {real, imag} */,
  {32'h41b7d1e8, 32'hc17e53be} /* (8, 30, 7) {real, imag} */,
  {32'h41a6cd38, 32'h413f15dd} /* (8, 30, 6) {real, imag} */,
  {32'h42a003a0, 32'h421caf60} /* (8, 30, 5) {real, imag} */,
  {32'hc1ff7fdc, 32'hc28ed330} /* (8, 30, 4) {real, imag} */,
  {32'hc1fb0fdb, 32'hc2920442} /* (8, 30, 3) {real, imag} */,
  {32'h440a3d64, 32'h4319eda6} /* (8, 30, 2) {real, imag} */,
  {32'hc498727c, 32'h41ffb2f2} /* (8, 30, 1) {real, imag} */,
  {32'hc41b20e7, 32'h43158d32} /* (8, 30, 0) {real, imag} */,
  {32'h42e35e97, 32'hc2cfbbd8} /* (8, 29, 31) {real, imag} */,
  {32'h41088d04, 32'h42afbae0} /* (8, 29, 30) {real, imag} */,
  {32'hc19fe610, 32'hc1096a58} /* (8, 29, 29) {real, imag} */,
  {32'hc25a96f3, 32'hc1c322c6} /* (8, 29, 28) {real, imag} */,
  {32'h4104af16, 32'hc1d7e300} /* (8, 29, 27) {real, imag} */,
  {32'hc0e275de, 32'hc072ee5c} /* (8, 29, 26) {real, imag} */,
  {32'hc1c471b5, 32'hc0348a10} /* (8, 29, 25) {real, imag} */,
  {32'h40539718, 32'hc157fcbc} /* (8, 29, 24) {real, imag} */,
  {32'h3f175ec0, 32'hc0ad7edd} /* (8, 29, 23) {real, imag} */,
  {32'hc10ab030, 32'hbee74d38} /* (8, 29, 22) {real, imag} */,
  {32'h40cfac72, 32'h406f0eaf} /* (8, 29, 21) {real, imag} */,
  {32'h413e90cb, 32'h40527004} /* (8, 29, 20) {real, imag} */,
  {32'hc03ae50c, 32'h40408295} /* (8, 29, 19) {real, imag} */,
  {32'hc072e101, 32'h412a0b76} /* (8, 29, 18) {real, imag} */,
  {32'hc18d1aa0, 32'hc05a01d8} /* (8, 29, 17) {real, imag} */,
  {32'hc16f6542, 32'hc12959d7} /* (8, 29, 16) {real, imag} */,
  {32'h41017329, 32'h3e050ff0} /* (8, 29, 15) {real, imag} */,
  {32'hc0cbf336, 32'h4119a022} /* (8, 29, 14) {real, imag} */,
  {32'h414214fb, 32'hc1875f48} /* (8, 29, 13) {real, imag} */,
  {32'h40b4b810, 32'hc00f69e6} /* (8, 29, 12) {real, imag} */,
  {32'h3f9272ea, 32'hc1107c32} /* (8, 29, 11) {real, imag} */,
  {32'h41b014cf, 32'hc114608e} /* (8, 29, 10) {real, imag} */,
  {32'h3ef3f120, 32'h41120a8a} /* (8, 29, 9) {real, imag} */,
  {32'hc1c19c86, 32'h41dee8f4} /* (8, 29, 8) {real, imag} */,
  {32'hc1c5f9d7, 32'hc1b3ce37} /* (8, 29, 7) {real, imag} */,
  {32'hc1377f2f, 32'hbfb4a574} /* (8, 29, 6) {real, imag} */,
  {32'hc22c0982, 32'h40c53252} /* (8, 29, 5) {real, imag} */,
  {32'h4206a215, 32'hc0b00a0c} /* (8, 29, 4) {real, imag} */,
  {32'h4114dccb, 32'hc20a6de0} /* (8, 29, 3) {real, imag} */,
  {32'h42894744, 32'h43190739} /* (8, 29, 2) {real, imag} */,
  {32'hc3093e46, 32'hc23626fc} /* (8, 29, 1) {real, imag} */,
  {32'h418dfd16, 32'h42084645} /* (8, 29, 0) {real, imag} */,
  {32'h431b5363, 32'hc28fdba4} /* (8, 28, 31) {real, imag} */,
  {32'hc2d2d024, 32'h428dc6d8} /* (8, 28, 30) {real, imag} */,
  {32'hc23f514c, 32'hc1ef7074} /* (8, 28, 29) {real, imag} */,
  {32'h41600eac, 32'hc04f0ee8} /* (8, 28, 28) {real, imag} */,
  {32'hc073e91d, 32'h421139ed} /* (8, 28, 27) {real, imag} */,
  {32'h41f62477, 32'h4064245c} /* (8, 28, 26) {real, imag} */,
  {32'h4092b5da, 32'h3fd4d568} /* (8, 28, 25) {real, imag} */,
  {32'h4148bd09, 32'h4224d9bc} /* (8, 28, 24) {real, imag} */,
  {32'hc0d0dfe5, 32'hc091c0a3} /* (8, 28, 23) {real, imag} */,
  {32'hc119e39d, 32'hc09558cb} /* (8, 28, 22) {real, imag} */,
  {32'h4194bde1, 32'hc072f5fa} /* (8, 28, 21) {real, imag} */,
  {32'h3fa32af4, 32'hc05b2d12} /* (8, 28, 20) {real, imag} */,
  {32'hbe9c3290, 32'hc1a7fdbe} /* (8, 28, 19) {real, imag} */,
  {32'h40d0ba30, 32'h411b4534} /* (8, 28, 18) {real, imag} */,
  {32'hc0d7fe1a, 32'h410b5554} /* (8, 28, 17) {real, imag} */,
  {32'h41418759, 32'h3f6c4b78} /* (8, 28, 16) {real, imag} */,
  {32'hc1096498, 32'h3ed20fe0} /* (8, 28, 15) {real, imag} */,
  {32'h3f7887d8, 32'h414984c5} /* (8, 28, 14) {real, imag} */,
  {32'hc04f186e, 32'hc0759e8d} /* (8, 28, 13) {real, imag} */,
  {32'h4064a5ae, 32'hc08acd0c} /* (8, 28, 12) {real, imag} */,
  {32'hbf85bf0c, 32'hc1622b63} /* (8, 28, 11) {real, imag} */,
  {32'h413c69c6, 32'h41694c04} /* (8, 28, 10) {real, imag} */,
  {32'h41b4e8f0, 32'h4083a134} /* (8, 28, 9) {real, imag} */,
  {32'hc1266fa4, 32'h415f1371} /* (8, 28, 8) {real, imag} */,
  {32'h40f9daf2, 32'hc0d571dc} /* (8, 28, 7) {real, imag} */,
  {32'hc102be28, 32'hc109bfce} /* (8, 28, 6) {real, imag} */,
  {32'hc18e30f6, 32'h4175b074} /* (8, 28, 5) {real, imag} */,
  {32'h41b762c1, 32'hc193291a} /* (8, 28, 4) {real, imag} */,
  {32'hc1bd52fa, 32'h40a1fec8} /* (8, 28, 3) {real, imag} */,
  {32'hc2ac3a41, 32'h42a30b6d} /* (8, 28, 2) {real, imag} */,
  {32'h41cd1bda, 32'hc2c3a0d8} /* (8, 28, 1) {real, imag} */,
  {32'h425cba62, 32'hc1cb1984} /* (8, 28, 0) {real, imag} */,
  {32'hc1e1dd3a, 32'h42803406} /* (8, 27, 31) {real, imag} */,
  {32'h41c4c139, 32'hc235c15c} /* (8, 27, 30) {real, imag} */,
  {32'hc17f891e, 32'h3ed0c570} /* (8, 27, 29) {real, imag} */,
  {32'hc199a4ea, 32'h41110346} /* (8, 27, 28) {real, imag} */,
  {32'h4241590c, 32'hc20f191d} /* (8, 27, 27) {real, imag} */,
  {32'hc050a0d8, 32'hc155a3bd} /* (8, 27, 26) {real, imag} */,
  {32'hc1347a94, 32'h411fbe62} /* (8, 27, 25) {real, imag} */,
  {32'h41956503, 32'h408601c4} /* (8, 27, 24) {real, imag} */,
  {32'hc04d9140, 32'hc117b90d} /* (8, 27, 23) {real, imag} */,
  {32'h40e158e9, 32'hc002028c} /* (8, 27, 22) {real, imag} */,
  {32'h411b0683, 32'h41971048} /* (8, 27, 21) {real, imag} */,
  {32'h4121277a, 32'h40d823c2} /* (8, 27, 20) {real, imag} */,
  {32'hc104c9f6, 32'hc06c48ec} /* (8, 27, 19) {real, imag} */,
  {32'hc12746a6, 32'hc1b27688} /* (8, 27, 18) {real, imag} */,
  {32'h414ca738, 32'hbf8f37a4} /* (8, 27, 17) {real, imag} */,
  {32'h410314b3, 32'hc0263d22} /* (8, 27, 16) {real, imag} */,
  {32'hc0a1ecfa, 32'h4020f380} /* (8, 27, 15) {real, imag} */,
  {32'hc0f480f6, 32'h405d50da} /* (8, 27, 14) {real, imag} */,
  {32'h41147cb8, 32'hc0c2c4a4} /* (8, 27, 13) {real, imag} */,
  {32'hc135eb5a, 32'h414210f2} /* (8, 27, 12) {real, imag} */,
  {32'h3f11f7f0, 32'h41af835c} /* (8, 27, 11) {real, imag} */,
  {32'h41046867, 32'h3fdb52a8} /* (8, 27, 10) {real, imag} */,
  {32'hbf59211c, 32'hc12f0302} /* (8, 27, 9) {real, imag} */,
  {32'h41675f10, 32'h419b53a4} /* (8, 27, 8) {real, imag} */,
  {32'h404812b8, 32'hc1377a2e} /* (8, 27, 7) {real, imag} */,
  {32'hc17fec05, 32'hc1ecd200} /* (8, 27, 6) {real, imag} */,
  {32'hc0af85c8, 32'h40dc86c0} /* (8, 27, 5) {real, imag} */,
  {32'h3fec1680, 32'h40b27da9} /* (8, 27, 4) {real, imag} */,
  {32'h41b96cb6, 32'hc05ccd84} /* (8, 27, 3) {real, imag} */,
  {32'h42139c8f, 32'h41cf5082} /* (8, 27, 2) {real, imag} */,
  {32'hc2a45f32, 32'h41268117} /* (8, 27, 1) {real, imag} */,
  {32'hc285626f, 32'h41af64cd} /* (8, 27, 0) {real, imag} */,
  {32'hc141a9e0, 32'h4140adb2} /* (8, 26, 31) {real, imag} */,
  {32'hc2026050, 32'h4163b8b4} /* (8, 26, 30) {real, imag} */,
  {32'h408c642c, 32'hc0aa9c49} /* (8, 26, 29) {real, imag} */,
  {32'h41729525, 32'h414f2690} /* (8, 26, 28) {real, imag} */,
  {32'h400b4c4c, 32'h4092a7a7} /* (8, 26, 27) {real, imag} */,
  {32'h412525d6, 32'hc1102f8f} /* (8, 26, 26) {real, imag} */,
  {32'hc1078555, 32'hc2132adc} /* (8, 26, 25) {real, imag} */,
  {32'h40317a9a, 32'hc0e7cab1} /* (8, 26, 24) {real, imag} */,
  {32'hc0fe0c32, 32'hbf62edb8} /* (8, 26, 23) {real, imag} */,
  {32'h416c69ea, 32'hc110c792} /* (8, 26, 22) {real, imag} */,
  {32'h41453715, 32'h4173b089} /* (8, 26, 21) {real, imag} */,
  {32'h41066f9f, 32'hc115083d} /* (8, 26, 20) {real, imag} */,
  {32'h412c16ae, 32'h4081eea8} /* (8, 26, 19) {real, imag} */,
  {32'h4103ab2e, 32'hc02bbf04} /* (8, 26, 18) {real, imag} */,
  {32'h409cd784, 32'h40f33dc2} /* (8, 26, 17) {real, imag} */,
  {32'hc0dfc13c, 32'h4046a443} /* (8, 26, 16) {real, imag} */,
  {32'h4081d552, 32'h4102b2b7} /* (8, 26, 15) {real, imag} */,
  {32'h41014c70, 32'h41281e2f} /* (8, 26, 14) {real, imag} */,
  {32'hc08cda54, 32'hc12d1013} /* (8, 26, 13) {real, imag} */,
  {32'hc19c9498, 32'h41ba7193} /* (8, 26, 12) {real, imag} */,
  {32'h4138a24b, 32'h3f62e78c} /* (8, 26, 11) {real, imag} */,
  {32'h416db58a, 32'h407ae31e} /* (8, 26, 10) {real, imag} */,
  {32'h418d37be, 32'hc146f048} /* (8, 26, 9) {real, imag} */,
  {32'h3eac5cd8, 32'h40b22f40} /* (8, 26, 8) {real, imag} */,
  {32'h3e839ff8, 32'hc006ad42} /* (8, 26, 7) {real, imag} */,
  {32'hc1596dca, 32'hc14e255c} /* (8, 26, 6) {real, imag} */,
  {32'h41255606, 32'hc1827fcf} /* (8, 26, 5) {real, imag} */,
  {32'hc02b32e4, 32'h40faf4b7} /* (8, 26, 4) {real, imag} */,
  {32'h404391bc, 32'hc0d19c6e} /* (8, 26, 3) {real, imag} */,
  {32'hbe223fc0, 32'hc04a774a} /* (8, 26, 2) {real, imag} */,
  {32'hc113337e, 32'h411d0403} /* (8, 26, 1) {real, imag} */,
  {32'hc128f784, 32'hc16d50a2} /* (8, 26, 0) {real, imag} */,
  {32'h4147b797, 32'hc1c725cf} /* (8, 25, 31) {real, imag} */,
  {32'hbfba0994, 32'h421b4ef0} /* (8, 25, 30) {real, imag} */,
  {32'hc1f9ef90, 32'hc1ccd28a} /* (8, 25, 29) {real, imag} */,
  {32'hc143ff04, 32'hbfa4ccc9} /* (8, 25, 28) {real, imag} */,
  {32'h410860d2, 32'hc092faa6} /* (8, 25, 27) {real, imag} */,
  {32'hc114a574, 32'h40c06b47} /* (8, 25, 26) {real, imag} */,
  {32'h4111d480, 32'h4119ba82} /* (8, 25, 25) {real, imag} */,
  {32'h40e466f4, 32'hc136c616} /* (8, 25, 24) {real, imag} */,
  {32'hc0e091b0, 32'hc1714b59} /* (8, 25, 23) {real, imag} */,
  {32'hc0204e30, 32'h3fb8f2b0} /* (8, 25, 22) {real, imag} */,
  {32'h418371a9, 32'hc04c8b86} /* (8, 25, 21) {real, imag} */,
  {32'hc1496cbe, 32'h40df5733} /* (8, 25, 20) {real, imag} */,
  {32'hc173a30a, 32'hbfab1194} /* (8, 25, 19) {real, imag} */,
  {32'h414f910f, 32'hc0610a3a} /* (8, 25, 18) {real, imag} */,
  {32'h40d78e06, 32'h41494efe} /* (8, 25, 17) {real, imag} */,
  {32'h405ab75e, 32'h3e8c5a30} /* (8, 25, 16) {real, imag} */,
  {32'h4080da92, 32'h40c12dcd} /* (8, 25, 15) {real, imag} */,
  {32'h41422796, 32'h41362cdc} /* (8, 25, 14) {real, imag} */,
  {32'h4119e5c6, 32'h4079f117} /* (8, 25, 13) {real, imag} */,
  {32'h4105e7e7, 32'hc0531ec0} /* (8, 25, 12) {real, imag} */,
  {32'hbff19858, 32'hc09bf2a8} /* (8, 25, 11) {real, imag} */,
  {32'hbf20a856, 32'hc14ea660} /* (8, 25, 10) {real, imag} */,
  {32'hc161dde2, 32'hc0598f37} /* (8, 25, 9) {real, imag} */,
  {32'h405272c6, 32'h40d4e389} /* (8, 25, 8) {real, imag} */,
  {32'hc1105f5e, 32'hc0bd15d5} /* (8, 25, 7) {real, imag} */,
  {32'h411c9b49, 32'h40bfe0a8} /* (8, 25, 6) {real, imag} */,
  {32'hc08e45ce, 32'hbe74b720} /* (8, 25, 5) {real, imag} */,
  {32'hc118ba23, 32'hc153e79f} /* (8, 25, 4) {real, imag} */,
  {32'h400bb6b6, 32'h41172242} /* (8, 25, 3) {real, imag} */,
  {32'h3f12f940, 32'h4160713a} /* (8, 25, 2) {real, imag} */,
  {32'hc0947a74, 32'h40e6c954} /* (8, 25, 1) {real, imag} */,
  {32'h419f600c, 32'hc10ba742} /* (8, 25, 0) {real, imag} */,
  {32'hc1c71e19, 32'h4175166e} /* (8, 24, 31) {real, imag} */,
  {32'h41c4b48c, 32'h3ded9780} /* (8, 24, 30) {real, imag} */,
  {32'h401ebc3c, 32'hc11e50d4} /* (8, 24, 29) {real, imag} */,
  {32'hc06fa31a, 32'h4194aa26} /* (8, 24, 28) {real, imag} */,
  {32'h411cd322, 32'hc0201c7e} /* (8, 24, 27) {real, imag} */,
  {32'hbfd327c0, 32'h4195483c} /* (8, 24, 26) {real, imag} */,
  {32'hc152cfeb, 32'hc1c0a1ed} /* (8, 24, 25) {real, imag} */,
  {32'hc0c2fbc4, 32'h414e4b69} /* (8, 24, 24) {real, imag} */,
  {32'h3e1893e0, 32'hc1391f5d} /* (8, 24, 23) {real, imag} */,
  {32'h418f8dbb, 32'hc10ea5bd} /* (8, 24, 22) {real, imag} */,
  {32'h40d910ca, 32'hbe59d600} /* (8, 24, 21) {real, imag} */,
  {32'h41200028, 32'h3ea488c8} /* (8, 24, 20) {real, imag} */,
  {32'h402d6963, 32'h412cf958} /* (8, 24, 19) {real, imag} */,
  {32'hc1573482, 32'hc0e75785} /* (8, 24, 18) {real, imag} */,
  {32'hbeb18a10, 32'hc02e8d62} /* (8, 24, 17) {real, imag} */,
  {32'h40cba8de, 32'hc08ad055} /* (8, 24, 16) {real, imag} */,
  {32'h40c37693, 32'hc128a6b2} /* (8, 24, 15) {real, imag} */,
  {32'hc0ffacf9, 32'h413d1d44} /* (8, 24, 14) {real, imag} */,
  {32'hc0df9239, 32'h405e8d58} /* (8, 24, 13) {real, imag} */,
  {32'h4055a426, 32'hc170035b} /* (8, 24, 12) {real, imag} */,
  {32'h3fac2baa, 32'hc03ae2c4} /* (8, 24, 11) {real, imag} */,
  {32'hbf60ae0b, 32'h3fbfc020} /* (8, 24, 10) {real, imag} */,
  {32'h404d317c, 32'h40bdb690} /* (8, 24, 9) {real, imag} */,
  {32'hbf43dca8, 32'h41707c13} /* (8, 24, 8) {real, imag} */,
  {32'hc034541c, 32'hc1554ef3} /* (8, 24, 7) {real, imag} */,
  {32'h418e7085, 32'h40a12d66} /* (8, 24, 6) {real, imag} */,
  {32'h4175b960, 32'h41036f92} /* (8, 24, 5) {real, imag} */,
  {32'h41e01a48, 32'h3c9b8f80} /* (8, 24, 4) {real, imag} */,
  {32'h408d2346, 32'hbfa8f49a} /* (8, 24, 3) {real, imag} */,
  {32'h41d9f388, 32'h402f43d6} /* (8, 24, 2) {real, imag} */,
  {32'hc22b588b, 32'h41f37c8e} /* (8, 24, 1) {real, imag} */,
  {32'hc1936038, 32'hbf1c9980} /* (8, 24, 0) {real, imag} */,
  {32'h40ae3e34, 32'hbf8722d4} /* (8, 23, 31) {real, imag} */,
  {32'hc057e46f, 32'h4183bd80} /* (8, 23, 30) {real, imag} */,
  {32'hbfefbaca, 32'h40cfcd6b} /* (8, 23, 29) {real, imag} */,
  {32'h4015ba23, 32'hc09322b6} /* (8, 23, 28) {real, imag} */,
  {32'hc0227b2c, 32'h41197c32} /* (8, 23, 27) {real, imag} */,
  {32'hc1308120, 32'h4045997a} /* (8, 23, 26) {real, imag} */,
  {32'hc0c90e47, 32'hc11f85ba} /* (8, 23, 25) {real, imag} */,
  {32'hc09b03f5, 32'h3f1a4628} /* (8, 23, 24) {real, imag} */,
  {32'hc153f2af, 32'hc18018ce} /* (8, 23, 23) {real, imag} */,
  {32'hc0c11e19, 32'hc0e63bff} /* (8, 23, 22) {real, imag} */,
  {32'h4075311c, 32'h3fc20a96} /* (8, 23, 21) {real, imag} */,
  {32'h41a8f4ea, 32'h4149c5c7} /* (8, 23, 20) {real, imag} */,
  {32'h3faa1ac8, 32'h41765ef1} /* (8, 23, 19) {real, imag} */,
  {32'h3fbc5d70, 32'hc105b13e} /* (8, 23, 18) {real, imag} */,
  {32'hc0f2c9bc, 32'hc15e0108} /* (8, 23, 17) {real, imag} */,
  {32'h4002d384, 32'hc0be27b1} /* (8, 23, 16) {real, imag} */,
  {32'hc01b7c33, 32'h408e8632} /* (8, 23, 15) {real, imag} */,
  {32'hc0e51436, 32'hc02c8e8e} /* (8, 23, 14) {real, imag} */,
  {32'hc0d363be, 32'h4106977a} /* (8, 23, 13) {real, imag} */,
  {32'h416c6859, 32'hc0b61877} /* (8, 23, 12) {real, imag} */,
  {32'h40b222a0, 32'hc1d4de4c} /* (8, 23, 11) {real, imag} */,
  {32'h411cdd0c, 32'h40e9511c} /* (8, 23, 10) {real, imag} */,
  {32'hbf3d1fe0, 32'hc0ffe028} /* (8, 23, 9) {real, imag} */,
  {32'hc0a93a42, 32'hc0de5bd6} /* (8, 23, 8) {real, imag} */,
  {32'hbf79a7f4, 32'h419895d0} /* (8, 23, 7) {real, imag} */,
  {32'hc0322c92, 32'h41673680} /* (8, 23, 6) {real, imag} */,
  {32'hc18ff435, 32'h401502f0} /* (8, 23, 5) {real, imag} */,
  {32'hc19a9344, 32'h3f5ea538} /* (8, 23, 4) {real, imag} */,
  {32'h40c40757, 32'hbf237808} /* (8, 23, 3) {real, imag} */,
  {32'h41801be1, 32'h41c82d02} /* (8, 23, 2) {real, imag} */,
  {32'hc1b75939, 32'hc1aed1db} /* (8, 23, 1) {real, imag} */,
  {32'hc1bf00d0, 32'h41d687ce} /* (8, 23, 0) {real, imag} */,
  {32'hc0ad8c29, 32'h404a7a20} /* (8, 22, 31) {real, imag} */,
  {32'h414a5af5, 32'hc0bfcc9a} /* (8, 22, 30) {real, imag} */,
  {32'hc13b5051, 32'hbf6c78da} /* (8, 22, 29) {real, imag} */,
  {32'h413f70de, 32'hc10ac131} /* (8, 22, 28) {real, imag} */,
  {32'hc14315e2, 32'h40506771} /* (8, 22, 27) {real, imag} */,
  {32'hc1a7dd91, 32'h3f2beaf8} /* (8, 22, 26) {real, imag} */,
  {32'h40cdfa1c, 32'h4115ff91} /* (8, 22, 25) {real, imag} */,
  {32'hbf7d9608, 32'hc0ed07b5} /* (8, 22, 24) {real, imag} */,
  {32'h41a562d9, 32'h40cb6f1b} /* (8, 22, 23) {real, imag} */,
  {32'h4093403a, 32'h40f5245a} /* (8, 22, 22) {real, imag} */,
  {32'h3d240b00, 32'hc0b6ad7c} /* (8, 22, 21) {real, imag} */,
  {32'h412e1097, 32'h40973398} /* (8, 22, 20) {real, imag} */,
  {32'h40135819, 32'hc1323515} /* (8, 22, 19) {real, imag} */,
  {32'hc0484b42, 32'h405d3018} /* (8, 22, 18) {real, imag} */,
  {32'h3fc7fd52, 32'hc1069a98} /* (8, 22, 17) {real, imag} */,
  {32'hc0e9f8aa, 32'hc051bed6} /* (8, 22, 16) {real, imag} */,
  {32'h4107b5ef, 32'h405b90a8} /* (8, 22, 15) {real, imag} */,
  {32'h3f722020, 32'h4080fdc8} /* (8, 22, 14) {real, imag} */,
  {32'h41394fca, 32'hc105d9a4} /* (8, 22, 13) {real, imag} */,
  {32'h411d7941, 32'h3f3b224c} /* (8, 22, 12) {real, imag} */,
  {32'h412a4f8a, 32'hc11e9dbc} /* (8, 22, 11) {real, imag} */,
  {32'hc0073572, 32'h40ac138b} /* (8, 22, 10) {real, imag} */,
  {32'hc1686a9b, 32'h40ee3314} /* (8, 22, 9) {real, imag} */,
  {32'hc0c067f1, 32'h413b7f13} /* (8, 22, 8) {real, imag} */,
  {32'hc18ec2d2, 32'h40372eea} /* (8, 22, 7) {real, imag} */,
  {32'hc153bc4d, 32'hc0cd4586} /* (8, 22, 6) {real, imag} */,
  {32'h4052d82c, 32'hc0e9bf85} /* (8, 22, 5) {real, imag} */,
  {32'h41a9b56d, 32'h3ffb3d02} /* (8, 22, 4) {real, imag} */,
  {32'hbe35b3c0, 32'h409983d6} /* (8, 22, 3) {real, imag} */,
  {32'hc120172c, 32'h400884f8} /* (8, 22, 2) {real, imag} */,
  {32'h3e832b70, 32'h3fe17bc8} /* (8, 22, 1) {real, imag} */,
  {32'hc0fa5f81, 32'hc11d3b3a} /* (8, 22, 0) {real, imag} */,
  {32'hc06ffe40, 32'h416dc1f0} /* (8, 21, 31) {real, imag} */,
  {32'h41140654, 32'hc1262ab4} /* (8, 21, 30) {real, imag} */,
  {32'hbfdb6708, 32'hc105d7ee} /* (8, 21, 29) {real, imag} */,
  {32'h41405847, 32'h40204283} /* (8, 21, 28) {real, imag} */,
  {32'hc1d5675d, 32'h4051725d} /* (8, 21, 27) {real, imag} */,
  {32'h406f1ea0, 32'hbfbae576} /* (8, 21, 26) {real, imag} */,
  {32'hc0e5c5c7, 32'h4091e722} /* (8, 21, 25) {real, imag} */,
  {32'hc1594768, 32'h41823c90} /* (8, 21, 24) {real, imag} */,
  {32'h4153a870, 32'h3f6f63f0} /* (8, 21, 23) {real, imag} */,
  {32'hc1ad1132, 32'hc209808d} /* (8, 21, 22) {real, imag} */,
  {32'h405aa7eb, 32'hc0b61875} /* (8, 21, 21) {real, imag} */,
  {32'hc13b9580, 32'h40d529b4} /* (8, 21, 20) {real, imag} */,
  {32'hc21a57ec, 32'hc0c217a2} /* (8, 21, 19) {real, imag} */,
  {32'h40724476, 32'h4045c6de} /* (8, 21, 18) {real, imag} */,
  {32'h408c9fca, 32'h3f9e3f94} /* (8, 21, 17) {real, imag} */,
  {32'h3f5f0d10, 32'h40e1f965} /* (8, 21, 16) {real, imag} */,
  {32'h3ed31500, 32'hc15b2730} /* (8, 21, 15) {real, imag} */,
  {32'hbeae9c68, 32'h41080698} /* (8, 21, 14) {real, imag} */,
  {32'h3fc1f4f6, 32'h40f666f6} /* (8, 21, 13) {real, imag} */,
  {32'h416e6cb2, 32'hc1280ce9} /* (8, 21, 12) {real, imag} */,
  {32'h4111e5b4, 32'h412629f5} /* (8, 21, 11) {real, imag} */,
  {32'hc12809dd, 32'h40080f88} /* (8, 21, 10) {real, imag} */,
  {32'hc0962e51, 32'hbf9c200a} /* (8, 21, 9) {real, imag} */,
  {32'hc07316e6, 32'h4000e447} /* (8, 21, 8) {real, imag} */,
  {32'hc09a6464, 32'h406eb3aa} /* (8, 21, 7) {real, imag} */,
  {32'h405299e0, 32'h41171ca4} /* (8, 21, 6) {real, imag} */,
  {32'h41a41030, 32'hc019b1ba} /* (8, 21, 5) {real, imag} */,
  {32'h40999a44, 32'hc16a3174} /* (8, 21, 4) {real, imag} */,
  {32'hc0249d82, 32'h4023a120} /* (8, 21, 3) {real, imag} */,
  {32'h407c0f6c, 32'hc1603e2a} /* (8, 21, 2) {real, imag} */,
  {32'h40fdfe98, 32'hc027f2ca} /* (8, 21, 1) {real, imag} */,
  {32'hc1de58f0, 32'h41f19ffb} /* (8, 21, 0) {real, imag} */,
  {32'h41164e44, 32'hc0a767df} /* (8, 20, 31) {real, imag} */,
  {32'hc0cf9ebc, 32'hc1844609} /* (8, 20, 30) {real, imag} */,
  {32'h409690b5, 32'h415008e3} /* (8, 20, 29) {real, imag} */,
  {32'hc0abb416, 32'h403c0d68} /* (8, 20, 28) {real, imag} */,
  {32'h41b31400, 32'hc1498edf} /* (8, 20, 27) {real, imag} */,
  {32'h40ac6c5d, 32'h3fbea744} /* (8, 20, 26) {real, imag} */,
  {32'hc13c7917, 32'hc01626de} /* (8, 20, 25) {real, imag} */,
  {32'hc06aa95c, 32'hc1bcc3af} /* (8, 20, 24) {real, imag} */,
  {32'h4182d65b, 32'h411e3488} /* (8, 20, 23) {real, imag} */,
  {32'hc03f40d0, 32'hbee8ac20} /* (8, 20, 22) {real, imag} */,
  {32'hc08b7635, 32'h40a29e51} /* (8, 20, 21) {real, imag} */,
  {32'h41667d72, 32'h4106a9d9} /* (8, 20, 20) {real, imag} */,
  {32'hc1a5fd20, 32'hbf2eaa56} /* (8, 20, 19) {real, imag} */,
  {32'hc032a3cf, 32'hc104ae1c} /* (8, 20, 18) {real, imag} */,
  {32'hbe8e81a0, 32'h41370b26} /* (8, 20, 17) {real, imag} */,
  {32'hc0411a54, 32'h3fa4a7fb} /* (8, 20, 16) {real, imag} */,
  {32'hbe856ee0, 32'hc09df81c} /* (8, 20, 15) {real, imag} */,
  {32'hc18f969b, 32'hc0c33a74} /* (8, 20, 14) {real, imag} */,
  {32'hc117baba, 32'hc0e30d05} /* (8, 20, 13) {real, imag} */,
  {32'hc1342018, 32'h41ae2721} /* (8, 20, 12) {real, imag} */,
  {32'h3f1eabb0, 32'hc11b6490} /* (8, 20, 11) {real, imag} */,
  {32'h41a54578, 32'hc1438cf4} /* (8, 20, 10) {real, imag} */,
  {32'hc13740dd, 32'h40d7cb75} /* (8, 20, 9) {real, imag} */,
  {32'hbfd47254, 32'hc0ac0f58} /* (8, 20, 8) {real, imag} */,
  {32'h411bdbd0, 32'hc14d104e} /* (8, 20, 7) {real, imag} */,
  {32'hc11fa9a6, 32'h419922f0} /* (8, 20, 6) {real, imag} */,
  {32'hc00cf69e, 32'h41771a44} /* (8, 20, 5) {real, imag} */,
  {32'hc0f1c692, 32'h4094ec5a} /* (8, 20, 4) {real, imag} */,
  {32'h40fb81ee, 32'hc0844b1c} /* (8, 20, 3) {real, imag} */,
  {32'h401d0cf0, 32'h40b1f03c} /* (8, 20, 2) {real, imag} */,
  {32'h40357610, 32'h41256b63} /* (8, 20, 1) {real, imag} */,
  {32'h40cdc9ca, 32'hc1a4456d} /* (8, 20, 0) {real, imag} */,
  {32'hbfd60340, 32'hc1df2a90} /* (8, 19, 31) {real, imag} */,
  {32'h415f8476, 32'h4086bf90} /* (8, 19, 30) {real, imag} */,
  {32'h41470a8a, 32'hc0c60a50} /* (8, 19, 29) {real, imag} */,
  {32'hc0cb0e2a, 32'hbfa4fce8} /* (8, 19, 28) {real, imag} */,
  {32'h40b18cee, 32'h40a1d524} /* (8, 19, 27) {real, imag} */,
  {32'h41435672, 32'hbfb97b96} /* (8, 19, 26) {real, imag} */,
  {32'h4187d2ae, 32'hc08118e3} /* (8, 19, 25) {real, imag} */,
  {32'h41709d9e, 32'h416100cc} /* (8, 19, 24) {real, imag} */,
  {32'hc061841e, 32'h4170edfd} /* (8, 19, 23) {real, imag} */,
  {32'h418754ba, 32'h405b34a1} /* (8, 19, 22) {real, imag} */,
  {32'hc0234285, 32'h417796d4} /* (8, 19, 21) {real, imag} */,
  {32'h409de766, 32'h3facb26e} /* (8, 19, 20) {real, imag} */,
  {32'hc01bf15e, 32'hc1531dab} /* (8, 19, 19) {real, imag} */,
  {32'h40f02d84, 32'h40ef9274} /* (8, 19, 18) {real, imag} */,
  {32'hc0cbd461, 32'h418324c6} /* (8, 19, 17) {real, imag} */,
  {32'hc0d46d20, 32'hc07051fc} /* (8, 19, 16) {real, imag} */,
  {32'hc0a3d86a, 32'h3fa95134} /* (8, 19, 15) {real, imag} */,
  {32'h3effaf78, 32'h3fd8aad2} /* (8, 19, 14) {real, imag} */,
  {32'h40322354, 32'hc0ab7052} /* (8, 19, 13) {real, imag} */,
  {32'h40e20512, 32'hc0d4add5} /* (8, 19, 12) {real, imag} */,
  {32'h3ef38708, 32'h413266ea} /* (8, 19, 11) {real, imag} */,
  {32'hc197b72e, 32'hbf8d4124} /* (8, 19, 10) {real, imag} */,
  {32'hbe83c000, 32'hc066dccf} /* (8, 19, 9) {real, imag} */,
  {32'h412198f4, 32'hc06e8b9d} /* (8, 19, 8) {real, imag} */,
  {32'h40da69d9, 32'hc0f7b405} /* (8, 19, 7) {real, imag} */,
  {32'hbfb02a70, 32'hc15bd2ba} /* (8, 19, 6) {real, imag} */,
  {32'h3da7c080, 32'hc0c69d80} /* (8, 19, 5) {real, imag} */,
  {32'h413c6651, 32'hc0e98e8c} /* (8, 19, 4) {real, imag} */,
  {32'h40bee376, 32'hc197228e} /* (8, 19, 3) {real, imag} */,
  {32'hc09dd4cc, 32'hc0f58c77} /* (8, 19, 2) {real, imag} */,
  {32'hc0c8bcfe, 32'hbf877c8c} /* (8, 19, 1) {real, imag} */,
  {32'h4124106c, 32'hbfe7d78c} /* (8, 19, 0) {real, imag} */,
  {32'h4153cbfc, 32'h413e0170} /* (8, 18, 31) {real, imag} */,
  {32'h40de92e4, 32'h3f4e3590} /* (8, 18, 30) {real, imag} */,
  {32'hbfb468ae, 32'hc0c22841} /* (8, 18, 29) {real, imag} */,
  {32'hc0093222, 32'hc0319555} /* (8, 18, 28) {real, imag} */,
  {32'hbfcbf918, 32'hc0962fc3} /* (8, 18, 27) {real, imag} */,
  {32'hc0cd9866, 32'h40bb6f6b} /* (8, 18, 26) {real, imag} */,
  {32'hc102d1bb, 32'h40a486a8} /* (8, 18, 25) {real, imag} */,
  {32'h40ae1984, 32'hc0389546} /* (8, 18, 24) {real, imag} */,
  {32'h402d071c, 32'h4119f14b} /* (8, 18, 23) {real, imag} */,
  {32'hc1b5da82, 32'hc11a5929} /* (8, 18, 22) {real, imag} */,
  {32'h3f2cc550, 32'hc139f222} /* (8, 18, 21) {real, imag} */,
  {32'h3f97e292, 32'h409677bf} /* (8, 18, 20) {real, imag} */,
  {32'h41059c40, 32'hbfeb6bb4} /* (8, 18, 19) {real, imag} */,
  {32'h411dd618, 32'hc1268fc6} /* (8, 18, 18) {real, imag} */,
  {32'h411217a2, 32'h4126007e} /* (8, 18, 17) {real, imag} */,
  {32'hc18b1ffe, 32'h400c377c} /* (8, 18, 16) {real, imag} */,
  {32'hbf4ad3cc, 32'hc13fefff} /* (8, 18, 15) {real, imag} */,
  {32'h40c06da6, 32'hc19681eb} /* (8, 18, 14) {real, imag} */,
  {32'h4178a3fa, 32'h41ade270} /* (8, 18, 13) {real, imag} */,
  {32'hbc964c80, 32'hbfec8ea0} /* (8, 18, 12) {real, imag} */,
  {32'h4101ae28, 32'hc0d4a2f5} /* (8, 18, 11) {real, imag} */,
  {32'hc0efcd54, 32'hc07b8b1e} /* (8, 18, 10) {real, imag} */,
  {32'h40c5076d, 32'hc18b0d72} /* (8, 18, 9) {real, imag} */,
  {32'h415291d2, 32'hc1228c56} /* (8, 18, 8) {real, imag} */,
  {32'h40f9f6af, 32'hbf66ef0a} /* (8, 18, 7) {real, imag} */,
  {32'hc183255f, 32'hc0448660} /* (8, 18, 6) {real, imag} */,
  {32'hc0958731, 32'h4138ac37} /* (8, 18, 5) {real, imag} */,
  {32'hbf8a8f68, 32'h416625a4} /* (8, 18, 4) {real, imag} */,
  {32'hc12df0c4, 32'h4173deb8} /* (8, 18, 3) {real, imag} */,
  {32'h4170c486, 32'hc13c062e} /* (8, 18, 2) {real, imag} */,
  {32'hc1062702, 32'h4126ea14} /* (8, 18, 1) {real, imag} */,
  {32'h3f0ca660, 32'h402bf25a} /* (8, 18, 0) {real, imag} */,
  {32'h3f8e012d, 32'hc133a4ea} /* (8, 17, 31) {real, imag} */,
  {32'h410c50c6, 32'h409cfc3b} /* (8, 17, 30) {real, imag} */,
  {32'hc02b26d9, 32'h40dfb314} /* (8, 17, 29) {real, imag} */,
  {32'hc15946f0, 32'h4087ec6e} /* (8, 17, 28) {real, imag} */,
  {32'hc08ca3c6, 32'h409a15b2} /* (8, 17, 27) {real, imag} */,
  {32'h40fac458, 32'h402669fc} /* (8, 17, 26) {real, imag} */,
  {32'hc0cc4750, 32'hc1896a83} /* (8, 17, 25) {real, imag} */,
  {32'hc0c6a24e, 32'h415a9349} /* (8, 17, 24) {real, imag} */,
  {32'hc16ca334, 32'h41668d29} /* (8, 17, 23) {real, imag} */,
  {32'hc0338cf8, 32'h40d9e5ee} /* (8, 17, 22) {real, imag} */,
  {32'h40706822, 32'h3fae9684} /* (8, 17, 21) {real, imag} */,
  {32'hc0d47a24, 32'h411bbb61} /* (8, 17, 20) {real, imag} */,
  {32'h4139af5d, 32'h40c57532} /* (8, 17, 19) {real, imag} */,
  {32'h40d9f8e6, 32'hc0133b6a} /* (8, 17, 18) {real, imag} */,
  {32'h40823d30, 32'hc0ba3d87} /* (8, 17, 17) {real, imag} */,
  {32'h3fde628a, 32'hc0f1ee05} /* (8, 17, 16) {real, imag} */,
  {32'h40094588, 32'hc11614e8} /* (8, 17, 15) {real, imag} */,
  {32'h409b4bc4, 32'h402486b5} /* (8, 17, 14) {real, imag} */,
  {32'hc017cf07, 32'hbf98820d} /* (8, 17, 13) {real, imag} */,
  {32'h3ecae3e8, 32'hc0b7ed34} /* (8, 17, 12) {real, imag} */,
  {32'hc137caba, 32'h40c3dd1d} /* (8, 17, 11) {real, imag} */,
  {32'hc155a555, 32'h4122f15a} /* (8, 17, 10) {real, imag} */,
  {32'h40cc4202, 32'h416928ce} /* (8, 17, 9) {real, imag} */,
  {32'h41117906, 32'h404245a0} /* (8, 17, 8) {real, imag} */,
  {32'hc000e1bc, 32'h40a641bc} /* (8, 17, 7) {real, imag} */,
  {32'h4124e711, 32'hc11a6108} /* (8, 17, 6) {real, imag} */,
  {32'h401ccc46, 32'h3b527400} /* (8, 17, 5) {real, imag} */,
  {32'h41196059, 32'hbfbab5dd} /* (8, 17, 4) {real, imag} */,
  {32'hc129a8a8, 32'hc106613c} /* (8, 17, 3) {real, imag} */,
  {32'hc037b425, 32'hc0de7c51} /* (8, 17, 2) {real, imag} */,
  {32'hc0323438, 32'hc08f1eba} /* (8, 17, 1) {real, imag} */,
  {32'hc03391aa, 32'h400b89ec} /* (8, 17, 0) {real, imag} */,
  {32'hc071a164, 32'hc03d0f4b} /* (8, 16, 31) {real, imag} */,
  {32'h3f515d20, 32'h40ddf9d8} /* (8, 16, 30) {real, imag} */,
  {32'hc14ec1f0, 32'h40e3ae31} /* (8, 16, 29) {real, imag} */,
  {32'hc042d52a, 32'hbf6642b4} /* (8, 16, 28) {real, imag} */,
  {32'h3fae27a4, 32'hc03f2e16} /* (8, 16, 27) {real, imag} */,
  {32'h3f576894, 32'h41152469} /* (8, 16, 26) {real, imag} */,
  {32'hc077881e, 32'h3e15c4c0} /* (8, 16, 25) {real, imag} */,
  {32'hc10d6653, 32'h40811a58} /* (8, 16, 24) {real, imag} */,
  {32'hc189dcba, 32'hc129071c} /* (8, 16, 23) {real, imag} */,
  {32'hc07633f4, 32'hc13660f1} /* (8, 16, 22) {real, imag} */,
  {32'h41045d9c, 32'hc08bc16b} /* (8, 16, 21) {real, imag} */,
  {32'h3eb61460, 32'hc0739e24} /* (8, 16, 20) {real, imag} */,
  {32'hc007c45e, 32'hc081fba8} /* (8, 16, 19) {real, imag} */,
  {32'hc1946b04, 32'hbfe6915f} /* (8, 16, 18) {real, imag} */,
  {32'h406c8df0, 32'hc04bea1b} /* (8, 16, 17) {real, imag} */,
  {32'h414c5874, 32'h00000000} /* (8, 16, 16) {real, imag} */,
  {32'h406c8df0, 32'h404bea1b} /* (8, 16, 15) {real, imag} */,
  {32'hc1946b04, 32'h3fe6915f} /* (8, 16, 14) {real, imag} */,
  {32'hc007c45e, 32'h4081fba8} /* (8, 16, 13) {real, imag} */,
  {32'h3eb61460, 32'h40739e24} /* (8, 16, 12) {real, imag} */,
  {32'h41045d9c, 32'h408bc16b} /* (8, 16, 11) {real, imag} */,
  {32'hc07633f4, 32'h413660f1} /* (8, 16, 10) {real, imag} */,
  {32'hc189dcba, 32'h4129071c} /* (8, 16, 9) {real, imag} */,
  {32'hc10d6653, 32'hc0811a58} /* (8, 16, 8) {real, imag} */,
  {32'hc077881e, 32'hbe15c4c0} /* (8, 16, 7) {real, imag} */,
  {32'h3f576894, 32'hc1152469} /* (8, 16, 6) {real, imag} */,
  {32'h3fae27a4, 32'h403f2e16} /* (8, 16, 5) {real, imag} */,
  {32'hc042d52a, 32'h3f6642b4} /* (8, 16, 4) {real, imag} */,
  {32'hc14ec1f0, 32'hc0e3ae31} /* (8, 16, 3) {real, imag} */,
  {32'h3f515d20, 32'hc0ddf9d8} /* (8, 16, 2) {real, imag} */,
  {32'hc071a164, 32'h403d0f4b} /* (8, 16, 1) {real, imag} */,
  {32'h40fd9edc, 32'h00000000} /* (8, 16, 0) {real, imag} */,
  {32'hc0323438, 32'h408f1eba} /* (8, 15, 31) {real, imag} */,
  {32'hc037b425, 32'h40de7c51} /* (8, 15, 30) {real, imag} */,
  {32'hc129a8a8, 32'h4106613c} /* (8, 15, 29) {real, imag} */,
  {32'h41196059, 32'h3fbab5dd} /* (8, 15, 28) {real, imag} */,
  {32'h401ccc46, 32'hbb527400} /* (8, 15, 27) {real, imag} */,
  {32'h4124e711, 32'h411a6108} /* (8, 15, 26) {real, imag} */,
  {32'hc000e1bc, 32'hc0a641bc} /* (8, 15, 25) {real, imag} */,
  {32'h41117906, 32'hc04245a0} /* (8, 15, 24) {real, imag} */,
  {32'h40cc4202, 32'hc16928ce} /* (8, 15, 23) {real, imag} */,
  {32'hc155a555, 32'hc122f15a} /* (8, 15, 22) {real, imag} */,
  {32'hc137caba, 32'hc0c3dd1d} /* (8, 15, 21) {real, imag} */,
  {32'h3ecae3e8, 32'h40b7ed34} /* (8, 15, 20) {real, imag} */,
  {32'hc017cf07, 32'h3f98820d} /* (8, 15, 19) {real, imag} */,
  {32'h409b4bc4, 32'hc02486b5} /* (8, 15, 18) {real, imag} */,
  {32'h40094588, 32'h411614e8} /* (8, 15, 17) {real, imag} */,
  {32'h3fde628a, 32'h40f1ee05} /* (8, 15, 16) {real, imag} */,
  {32'h40823d30, 32'h40ba3d87} /* (8, 15, 15) {real, imag} */,
  {32'h40d9f8e6, 32'h40133b6a} /* (8, 15, 14) {real, imag} */,
  {32'h4139af5d, 32'hc0c57532} /* (8, 15, 13) {real, imag} */,
  {32'hc0d47a24, 32'hc11bbb61} /* (8, 15, 12) {real, imag} */,
  {32'h40706822, 32'hbfae9684} /* (8, 15, 11) {real, imag} */,
  {32'hc0338cf8, 32'hc0d9e5ee} /* (8, 15, 10) {real, imag} */,
  {32'hc16ca334, 32'hc1668d29} /* (8, 15, 9) {real, imag} */,
  {32'hc0c6a24e, 32'hc15a9349} /* (8, 15, 8) {real, imag} */,
  {32'hc0cc4750, 32'h41896a83} /* (8, 15, 7) {real, imag} */,
  {32'h40fac458, 32'hc02669fc} /* (8, 15, 6) {real, imag} */,
  {32'hc08ca3c6, 32'hc09a15b2} /* (8, 15, 5) {real, imag} */,
  {32'hc15946f0, 32'hc087ec6e} /* (8, 15, 4) {real, imag} */,
  {32'hc02b26d9, 32'hc0dfb314} /* (8, 15, 3) {real, imag} */,
  {32'h410c50c6, 32'hc09cfc3b} /* (8, 15, 2) {real, imag} */,
  {32'h3f8e012d, 32'h4133a4ea} /* (8, 15, 1) {real, imag} */,
  {32'hc03391aa, 32'hc00b89ec} /* (8, 15, 0) {real, imag} */,
  {32'hc1062702, 32'hc126ea14} /* (8, 14, 31) {real, imag} */,
  {32'h4170c486, 32'h413c062e} /* (8, 14, 30) {real, imag} */,
  {32'hc12df0c4, 32'hc173deb8} /* (8, 14, 29) {real, imag} */,
  {32'hbf8a8f68, 32'hc16625a4} /* (8, 14, 28) {real, imag} */,
  {32'hc0958731, 32'hc138ac37} /* (8, 14, 27) {real, imag} */,
  {32'hc183255f, 32'h40448660} /* (8, 14, 26) {real, imag} */,
  {32'h40f9f6af, 32'h3f66ef0a} /* (8, 14, 25) {real, imag} */,
  {32'h415291d2, 32'h41228c56} /* (8, 14, 24) {real, imag} */,
  {32'h40c5076d, 32'h418b0d72} /* (8, 14, 23) {real, imag} */,
  {32'hc0efcd54, 32'h407b8b1e} /* (8, 14, 22) {real, imag} */,
  {32'h4101ae28, 32'h40d4a2f5} /* (8, 14, 21) {real, imag} */,
  {32'hbc964c80, 32'h3fec8ea0} /* (8, 14, 20) {real, imag} */,
  {32'h4178a3fa, 32'hc1ade270} /* (8, 14, 19) {real, imag} */,
  {32'h40c06da6, 32'h419681eb} /* (8, 14, 18) {real, imag} */,
  {32'hbf4ad3cc, 32'h413fefff} /* (8, 14, 17) {real, imag} */,
  {32'hc18b1ffe, 32'hc00c377c} /* (8, 14, 16) {real, imag} */,
  {32'h411217a2, 32'hc126007e} /* (8, 14, 15) {real, imag} */,
  {32'h411dd618, 32'h41268fc6} /* (8, 14, 14) {real, imag} */,
  {32'h41059c40, 32'h3feb6bb4} /* (8, 14, 13) {real, imag} */,
  {32'h3f97e292, 32'hc09677bf} /* (8, 14, 12) {real, imag} */,
  {32'h3f2cc550, 32'h4139f222} /* (8, 14, 11) {real, imag} */,
  {32'hc1b5da82, 32'h411a5929} /* (8, 14, 10) {real, imag} */,
  {32'h402d071c, 32'hc119f14b} /* (8, 14, 9) {real, imag} */,
  {32'h40ae1984, 32'h40389546} /* (8, 14, 8) {real, imag} */,
  {32'hc102d1bb, 32'hc0a486a8} /* (8, 14, 7) {real, imag} */,
  {32'hc0cd9866, 32'hc0bb6f6b} /* (8, 14, 6) {real, imag} */,
  {32'hbfcbf918, 32'h40962fc3} /* (8, 14, 5) {real, imag} */,
  {32'hc0093222, 32'h40319555} /* (8, 14, 4) {real, imag} */,
  {32'hbfb468ae, 32'h40c22841} /* (8, 14, 3) {real, imag} */,
  {32'h40de92e4, 32'hbf4e3590} /* (8, 14, 2) {real, imag} */,
  {32'h4153cbfc, 32'hc13e0170} /* (8, 14, 1) {real, imag} */,
  {32'h3f0ca660, 32'hc02bf25a} /* (8, 14, 0) {real, imag} */,
  {32'hc0c8bcfe, 32'h3f877c8c} /* (8, 13, 31) {real, imag} */,
  {32'hc09dd4cc, 32'h40f58c77} /* (8, 13, 30) {real, imag} */,
  {32'h40bee376, 32'h4197228e} /* (8, 13, 29) {real, imag} */,
  {32'h413c6651, 32'h40e98e8c} /* (8, 13, 28) {real, imag} */,
  {32'h3da7c080, 32'h40c69d80} /* (8, 13, 27) {real, imag} */,
  {32'hbfb02a70, 32'h415bd2ba} /* (8, 13, 26) {real, imag} */,
  {32'h40da69d9, 32'h40f7b405} /* (8, 13, 25) {real, imag} */,
  {32'h412198f4, 32'h406e8b9d} /* (8, 13, 24) {real, imag} */,
  {32'hbe83c000, 32'h4066dccf} /* (8, 13, 23) {real, imag} */,
  {32'hc197b72e, 32'h3f8d4124} /* (8, 13, 22) {real, imag} */,
  {32'h3ef38708, 32'hc13266ea} /* (8, 13, 21) {real, imag} */,
  {32'h40e20512, 32'h40d4add5} /* (8, 13, 20) {real, imag} */,
  {32'h40322354, 32'h40ab7052} /* (8, 13, 19) {real, imag} */,
  {32'h3effaf78, 32'hbfd8aad2} /* (8, 13, 18) {real, imag} */,
  {32'hc0a3d86a, 32'hbfa95134} /* (8, 13, 17) {real, imag} */,
  {32'hc0d46d20, 32'h407051fc} /* (8, 13, 16) {real, imag} */,
  {32'hc0cbd461, 32'hc18324c6} /* (8, 13, 15) {real, imag} */,
  {32'h40f02d84, 32'hc0ef9274} /* (8, 13, 14) {real, imag} */,
  {32'hc01bf15e, 32'h41531dab} /* (8, 13, 13) {real, imag} */,
  {32'h409de766, 32'hbfacb26e} /* (8, 13, 12) {real, imag} */,
  {32'hc0234285, 32'hc17796d4} /* (8, 13, 11) {real, imag} */,
  {32'h418754ba, 32'hc05b34a1} /* (8, 13, 10) {real, imag} */,
  {32'hc061841e, 32'hc170edfd} /* (8, 13, 9) {real, imag} */,
  {32'h41709d9e, 32'hc16100cc} /* (8, 13, 8) {real, imag} */,
  {32'h4187d2ae, 32'h408118e3} /* (8, 13, 7) {real, imag} */,
  {32'h41435672, 32'h3fb97b96} /* (8, 13, 6) {real, imag} */,
  {32'h40b18cee, 32'hc0a1d524} /* (8, 13, 5) {real, imag} */,
  {32'hc0cb0e2a, 32'h3fa4fce8} /* (8, 13, 4) {real, imag} */,
  {32'h41470a8a, 32'h40c60a50} /* (8, 13, 3) {real, imag} */,
  {32'h415f8476, 32'hc086bf90} /* (8, 13, 2) {real, imag} */,
  {32'hbfd60340, 32'h41df2a90} /* (8, 13, 1) {real, imag} */,
  {32'h4124106c, 32'h3fe7d78c} /* (8, 13, 0) {real, imag} */,
  {32'h40357610, 32'hc1256b63} /* (8, 12, 31) {real, imag} */,
  {32'h401d0cf0, 32'hc0b1f03c} /* (8, 12, 30) {real, imag} */,
  {32'h40fb81ee, 32'h40844b1c} /* (8, 12, 29) {real, imag} */,
  {32'hc0f1c692, 32'hc094ec5a} /* (8, 12, 28) {real, imag} */,
  {32'hc00cf69e, 32'hc1771a44} /* (8, 12, 27) {real, imag} */,
  {32'hc11fa9a6, 32'hc19922f0} /* (8, 12, 26) {real, imag} */,
  {32'h411bdbd0, 32'h414d104e} /* (8, 12, 25) {real, imag} */,
  {32'hbfd47254, 32'h40ac0f58} /* (8, 12, 24) {real, imag} */,
  {32'hc13740dd, 32'hc0d7cb75} /* (8, 12, 23) {real, imag} */,
  {32'h41a54578, 32'h41438cf4} /* (8, 12, 22) {real, imag} */,
  {32'h3f1eabb0, 32'h411b6490} /* (8, 12, 21) {real, imag} */,
  {32'hc1342018, 32'hc1ae2721} /* (8, 12, 20) {real, imag} */,
  {32'hc117baba, 32'h40e30d05} /* (8, 12, 19) {real, imag} */,
  {32'hc18f969b, 32'h40c33a74} /* (8, 12, 18) {real, imag} */,
  {32'hbe856ee0, 32'h409df81c} /* (8, 12, 17) {real, imag} */,
  {32'hc0411a54, 32'hbfa4a7fb} /* (8, 12, 16) {real, imag} */,
  {32'hbe8e81a0, 32'hc1370b26} /* (8, 12, 15) {real, imag} */,
  {32'hc032a3cf, 32'h4104ae1c} /* (8, 12, 14) {real, imag} */,
  {32'hc1a5fd20, 32'h3f2eaa56} /* (8, 12, 13) {real, imag} */,
  {32'h41667d72, 32'hc106a9d9} /* (8, 12, 12) {real, imag} */,
  {32'hc08b7635, 32'hc0a29e51} /* (8, 12, 11) {real, imag} */,
  {32'hc03f40d0, 32'h3ee8ac20} /* (8, 12, 10) {real, imag} */,
  {32'h4182d65b, 32'hc11e3488} /* (8, 12, 9) {real, imag} */,
  {32'hc06aa95c, 32'h41bcc3af} /* (8, 12, 8) {real, imag} */,
  {32'hc13c7917, 32'h401626de} /* (8, 12, 7) {real, imag} */,
  {32'h40ac6c5d, 32'hbfbea744} /* (8, 12, 6) {real, imag} */,
  {32'h41b31400, 32'h41498edf} /* (8, 12, 5) {real, imag} */,
  {32'hc0abb416, 32'hc03c0d68} /* (8, 12, 4) {real, imag} */,
  {32'h409690b5, 32'hc15008e3} /* (8, 12, 3) {real, imag} */,
  {32'hc0cf9ebc, 32'h41844609} /* (8, 12, 2) {real, imag} */,
  {32'h41164e44, 32'h40a767df} /* (8, 12, 1) {real, imag} */,
  {32'h40cdc9ca, 32'h41a4456d} /* (8, 12, 0) {real, imag} */,
  {32'h40fdfe98, 32'h4027f2ca} /* (8, 11, 31) {real, imag} */,
  {32'h407c0f6c, 32'h41603e2a} /* (8, 11, 30) {real, imag} */,
  {32'hc0249d82, 32'hc023a120} /* (8, 11, 29) {real, imag} */,
  {32'h40999a44, 32'h416a3174} /* (8, 11, 28) {real, imag} */,
  {32'h41a41030, 32'h4019b1ba} /* (8, 11, 27) {real, imag} */,
  {32'h405299e0, 32'hc1171ca4} /* (8, 11, 26) {real, imag} */,
  {32'hc09a6464, 32'hc06eb3aa} /* (8, 11, 25) {real, imag} */,
  {32'hc07316e6, 32'hc000e447} /* (8, 11, 24) {real, imag} */,
  {32'hc0962e51, 32'h3f9c200a} /* (8, 11, 23) {real, imag} */,
  {32'hc12809dd, 32'hc0080f88} /* (8, 11, 22) {real, imag} */,
  {32'h4111e5b4, 32'hc12629f5} /* (8, 11, 21) {real, imag} */,
  {32'h416e6cb2, 32'h41280ce9} /* (8, 11, 20) {real, imag} */,
  {32'h3fc1f4f6, 32'hc0f666f6} /* (8, 11, 19) {real, imag} */,
  {32'hbeae9c68, 32'hc1080698} /* (8, 11, 18) {real, imag} */,
  {32'h3ed31500, 32'h415b2730} /* (8, 11, 17) {real, imag} */,
  {32'h3f5f0d10, 32'hc0e1f965} /* (8, 11, 16) {real, imag} */,
  {32'h408c9fca, 32'hbf9e3f94} /* (8, 11, 15) {real, imag} */,
  {32'h40724476, 32'hc045c6de} /* (8, 11, 14) {real, imag} */,
  {32'hc21a57ec, 32'h40c217a2} /* (8, 11, 13) {real, imag} */,
  {32'hc13b9580, 32'hc0d529b4} /* (8, 11, 12) {real, imag} */,
  {32'h405aa7eb, 32'h40b61875} /* (8, 11, 11) {real, imag} */,
  {32'hc1ad1132, 32'h4209808d} /* (8, 11, 10) {real, imag} */,
  {32'h4153a870, 32'hbf6f63f0} /* (8, 11, 9) {real, imag} */,
  {32'hc1594768, 32'hc1823c90} /* (8, 11, 8) {real, imag} */,
  {32'hc0e5c5c7, 32'hc091e722} /* (8, 11, 7) {real, imag} */,
  {32'h406f1ea0, 32'h3fbae576} /* (8, 11, 6) {real, imag} */,
  {32'hc1d5675d, 32'hc051725d} /* (8, 11, 5) {real, imag} */,
  {32'h41405847, 32'hc0204283} /* (8, 11, 4) {real, imag} */,
  {32'hbfdb6708, 32'h4105d7ee} /* (8, 11, 3) {real, imag} */,
  {32'h41140654, 32'h41262ab4} /* (8, 11, 2) {real, imag} */,
  {32'hc06ffe40, 32'hc16dc1f0} /* (8, 11, 1) {real, imag} */,
  {32'hc1de58f0, 32'hc1f19ffb} /* (8, 11, 0) {real, imag} */,
  {32'h3e832b70, 32'hbfe17bc8} /* (8, 10, 31) {real, imag} */,
  {32'hc120172c, 32'hc00884f8} /* (8, 10, 30) {real, imag} */,
  {32'hbe35b3c0, 32'hc09983d6} /* (8, 10, 29) {real, imag} */,
  {32'h41a9b56d, 32'hbffb3d02} /* (8, 10, 28) {real, imag} */,
  {32'h4052d82c, 32'h40e9bf85} /* (8, 10, 27) {real, imag} */,
  {32'hc153bc4d, 32'h40cd4586} /* (8, 10, 26) {real, imag} */,
  {32'hc18ec2d2, 32'hc0372eea} /* (8, 10, 25) {real, imag} */,
  {32'hc0c067f1, 32'hc13b7f13} /* (8, 10, 24) {real, imag} */,
  {32'hc1686a9b, 32'hc0ee3314} /* (8, 10, 23) {real, imag} */,
  {32'hc0073572, 32'hc0ac138b} /* (8, 10, 22) {real, imag} */,
  {32'h412a4f8a, 32'h411e9dbc} /* (8, 10, 21) {real, imag} */,
  {32'h411d7941, 32'hbf3b224c} /* (8, 10, 20) {real, imag} */,
  {32'h41394fca, 32'h4105d9a4} /* (8, 10, 19) {real, imag} */,
  {32'h3f722020, 32'hc080fdc8} /* (8, 10, 18) {real, imag} */,
  {32'h4107b5ef, 32'hc05b90a8} /* (8, 10, 17) {real, imag} */,
  {32'hc0e9f8aa, 32'h4051bed6} /* (8, 10, 16) {real, imag} */,
  {32'h3fc7fd52, 32'h41069a98} /* (8, 10, 15) {real, imag} */,
  {32'hc0484b42, 32'hc05d3018} /* (8, 10, 14) {real, imag} */,
  {32'h40135819, 32'h41323515} /* (8, 10, 13) {real, imag} */,
  {32'h412e1097, 32'hc0973398} /* (8, 10, 12) {real, imag} */,
  {32'h3d240b00, 32'h40b6ad7c} /* (8, 10, 11) {real, imag} */,
  {32'h4093403a, 32'hc0f5245a} /* (8, 10, 10) {real, imag} */,
  {32'h41a562d9, 32'hc0cb6f1b} /* (8, 10, 9) {real, imag} */,
  {32'hbf7d9608, 32'h40ed07b5} /* (8, 10, 8) {real, imag} */,
  {32'h40cdfa1c, 32'hc115ff91} /* (8, 10, 7) {real, imag} */,
  {32'hc1a7dd91, 32'hbf2beaf8} /* (8, 10, 6) {real, imag} */,
  {32'hc14315e2, 32'hc0506771} /* (8, 10, 5) {real, imag} */,
  {32'h413f70de, 32'h410ac131} /* (8, 10, 4) {real, imag} */,
  {32'hc13b5051, 32'h3f6c78da} /* (8, 10, 3) {real, imag} */,
  {32'h414a5af5, 32'h40bfcc9a} /* (8, 10, 2) {real, imag} */,
  {32'hc0ad8c29, 32'hc04a7a20} /* (8, 10, 1) {real, imag} */,
  {32'hc0fa5f81, 32'h411d3b3a} /* (8, 10, 0) {real, imag} */,
  {32'hc1b75939, 32'h41aed1db} /* (8, 9, 31) {real, imag} */,
  {32'h41801be1, 32'hc1c82d02} /* (8, 9, 30) {real, imag} */,
  {32'h40c40757, 32'h3f237808} /* (8, 9, 29) {real, imag} */,
  {32'hc19a9344, 32'hbf5ea538} /* (8, 9, 28) {real, imag} */,
  {32'hc18ff435, 32'hc01502f0} /* (8, 9, 27) {real, imag} */,
  {32'hc0322c92, 32'hc1673680} /* (8, 9, 26) {real, imag} */,
  {32'hbf79a7f4, 32'hc19895d0} /* (8, 9, 25) {real, imag} */,
  {32'hc0a93a42, 32'h40de5bd6} /* (8, 9, 24) {real, imag} */,
  {32'hbf3d1fe0, 32'h40ffe028} /* (8, 9, 23) {real, imag} */,
  {32'h411cdd0c, 32'hc0e9511c} /* (8, 9, 22) {real, imag} */,
  {32'h40b222a0, 32'h41d4de4c} /* (8, 9, 21) {real, imag} */,
  {32'h416c6859, 32'h40b61877} /* (8, 9, 20) {real, imag} */,
  {32'hc0d363be, 32'hc106977a} /* (8, 9, 19) {real, imag} */,
  {32'hc0e51436, 32'h402c8e8e} /* (8, 9, 18) {real, imag} */,
  {32'hc01b7c33, 32'hc08e8632} /* (8, 9, 17) {real, imag} */,
  {32'h4002d384, 32'h40be27b1} /* (8, 9, 16) {real, imag} */,
  {32'hc0f2c9bc, 32'h415e0108} /* (8, 9, 15) {real, imag} */,
  {32'h3fbc5d70, 32'h4105b13e} /* (8, 9, 14) {real, imag} */,
  {32'h3faa1ac8, 32'hc1765ef1} /* (8, 9, 13) {real, imag} */,
  {32'h41a8f4ea, 32'hc149c5c7} /* (8, 9, 12) {real, imag} */,
  {32'h4075311c, 32'hbfc20a96} /* (8, 9, 11) {real, imag} */,
  {32'hc0c11e19, 32'h40e63bff} /* (8, 9, 10) {real, imag} */,
  {32'hc153f2af, 32'h418018ce} /* (8, 9, 9) {real, imag} */,
  {32'hc09b03f5, 32'hbf1a4628} /* (8, 9, 8) {real, imag} */,
  {32'hc0c90e47, 32'h411f85ba} /* (8, 9, 7) {real, imag} */,
  {32'hc1308120, 32'hc045997a} /* (8, 9, 6) {real, imag} */,
  {32'hc0227b2c, 32'hc1197c32} /* (8, 9, 5) {real, imag} */,
  {32'h4015ba23, 32'h409322b6} /* (8, 9, 4) {real, imag} */,
  {32'hbfefbaca, 32'hc0cfcd6b} /* (8, 9, 3) {real, imag} */,
  {32'hc057e46f, 32'hc183bd80} /* (8, 9, 2) {real, imag} */,
  {32'h40ae3e34, 32'h3f8722d4} /* (8, 9, 1) {real, imag} */,
  {32'hc1bf00d0, 32'hc1d687ce} /* (8, 9, 0) {real, imag} */,
  {32'hc22b588b, 32'hc1f37c8e} /* (8, 8, 31) {real, imag} */,
  {32'h41d9f388, 32'hc02f43d6} /* (8, 8, 30) {real, imag} */,
  {32'h408d2346, 32'h3fa8f49a} /* (8, 8, 29) {real, imag} */,
  {32'h41e01a48, 32'hbc9b8f80} /* (8, 8, 28) {real, imag} */,
  {32'h4175b960, 32'hc1036f92} /* (8, 8, 27) {real, imag} */,
  {32'h418e7085, 32'hc0a12d66} /* (8, 8, 26) {real, imag} */,
  {32'hc034541c, 32'h41554ef3} /* (8, 8, 25) {real, imag} */,
  {32'hbf43dca8, 32'hc1707c13} /* (8, 8, 24) {real, imag} */,
  {32'h404d317c, 32'hc0bdb690} /* (8, 8, 23) {real, imag} */,
  {32'hbf60ae0b, 32'hbfbfc020} /* (8, 8, 22) {real, imag} */,
  {32'h3fac2baa, 32'h403ae2c4} /* (8, 8, 21) {real, imag} */,
  {32'h4055a426, 32'h4170035b} /* (8, 8, 20) {real, imag} */,
  {32'hc0df9239, 32'hc05e8d58} /* (8, 8, 19) {real, imag} */,
  {32'hc0ffacf9, 32'hc13d1d44} /* (8, 8, 18) {real, imag} */,
  {32'h40c37693, 32'h4128a6b2} /* (8, 8, 17) {real, imag} */,
  {32'h40cba8de, 32'h408ad055} /* (8, 8, 16) {real, imag} */,
  {32'hbeb18a10, 32'h402e8d62} /* (8, 8, 15) {real, imag} */,
  {32'hc1573482, 32'h40e75785} /* (8, 8, 14) {real, imag} */,
  {32'h402d6963, 32'hc12cf958} /* (8, 8, 13) {real, imag} */,
  {32'h41200028, 32'hbea488c8} /* (8, 8, 12) {real, imag} */,
  {32'h40d910ca, 32'h3e59d600} /* (8, 8, 11) {real, imag} */,
  {32'h418f8dbb, 32'h410ea5bd} /* (8, 8, 10) {real, imag} */,
  {32'h3e1893e0, 32'h41391f5d} /* (8, 8, 9) {real, imag} */,
  {32'hc0c2fbc4, 32'hc14e4b69} /* (8, 8, 8) {real, imag} */,
  {32'hc152cfeb, 32'h41c0a1ed} /* (8, 8, 7) {real, imag} */,
  {32'hbfd327c0, 32'hc195483c} /* (8, 8, 6) {real, imag} */,
  {32'h411cd322, 32'h40201c7e} /* (8, 8, 5) {real, imag} */,
  {32'hc06fa31a, 32'hc194aa26} /* (8, 8, 4) {real, imag} */,
  {32'h401ebc3c, 32'h411e50d4} /* (8, 8, 3) {real, imag} */,
  {32'h41c4b48c, 32'hbded9780} /* (8, 8, 2) {real, imag} */,
  {32'hc1c71e19, 32'hc175166e} /* (8, 8, 1) {real, imag} */,
  {32'hc1936038, 32'h3f1c9980} /* (8, 8, 0) {real, imag} */,
  {32'hc0947a74, 32'hc0e6c954} /* (8, 7, 31) {real, imag} */,
  {32'h3f12f940, 32'hc160713a} /* (8, 7, 30) {real, imag} */,
  {32'h400bb6b6, 32'hc1172242} /* (8, 7, 29) {real, imag} */,
  {32'hc118ba23, 32'h4153e79f} /* (8, 7, 28) {real, imag} */,
  {32'hc08e45ce, 32'h3e74b720} /* (8, 7, 27) {real, imag} */,
  {32'h411c9b49, 32'hc0bfe0a8} /* (8, 7, 26) {real, imag} */,
  {32'hc1105f5e, 32'h40bd15d5} /* (8, 7, 25) {real, imag} */,
  {32'h405272c6, 32'hc0d4e389} /* (8, 7, 24) {real, imag} */,
  {32'hc161dde2, 32'h40598f37} /* (8, 7, 23) {real, imag} */,
  {32'hbf20a856, 32'h414ea660} /* (8, 7, 22) {real, imag} */,
  {32'hbff19858, 32'h409bf2a8} /* (8, 7, 21) {real, imag} */,
  {32'h4105e7e7, 32'h40531ec0} /* (8, 7, 20) {real, imag} */,
  {32'h4119e5c6, 32'hc079f117} /* (8, 7, 19) {real, imag} */,
  {32'h41422796, 32'hc1362cdc} /* (8, 7, 18) {real, imag} */,
  {32'h4080da92, 32'hc0c12dcd} /* (8, 7, 17) {real, imag} */,
  {32'h405ab75e, 32'hbe8c5a30} /* (8, 7, 16) {real, imag} */,
  {32'h40d78e06, 32'hc1494efe} /* (8, 7, 15) {real, imag} */,
  {32'h414f910f, 32'h40610a3a} /* (8, 7, 14) {real, imag} */,
  {32'hc173a30a, 32'h3fab1194} /* (8, 7, 13) {real, imag} */,
  {32'hc1496cbe, 32'hc0df5733} /* (8, 7, 12) {real, imag} */,
  {32'h418371a9, 32'h404c8b86} /* (8, 7, 11) {real, imag} */,
  {32'hc0204e30, 32'hbfb8f2b0} /* (8, 7, 10) {real, imag} */,
  {32'hc0e091b0, 32'h41714b59} /* (8, 7, 9) {real, imag} */,
  {32'h40e466f4, 32'h4136c616} /* (8, 7, 8) {real, imag} */,
  {32'h4111d480, 32'hc119ba82} /* (8, 7, 7) {real, imag} */,
  {32'hc114a574, 32'hc0c06b47} /* (8, 7, 6) {real, imag} */,
  {32'h410860d2, 32'h4092faa6} /* (8, 7, 5) {real, imag} */,
  {32'hc143ff04, 32'h3fa4ccc9} /* (8, 7, 4) {real, imag} */,
  {32'hc1f9ef90, 32'h41ccd28a} /* (8, 7, 3) {real, imag} */,
  {32'hbfba0994, 32'hc21b4ef0} /* (8, 7, 2) {real, imag} */,
  {32'h4147b797, 32'h41c725cf} /* (8, 7, 1) {real, imag} */,
  {32'h419f600c, 32'h410ba742} /* (8, 7, 0) {real, imag} */,
  {32'hc113337e, 32'hc11d0403} /* (8, 6, 31) {real, imag} */,
  {32'hbe223fc0, 32'h404a774a} /* (8, 6, 30) {real, imag} */,
  {32'h404391bc, 32'h40d19c6e} /* (8, 6, 29) {real, imag} */,
  {32'hc02b32e4, 32'hc0faf4b7} /* (8, 6, 28) {real, imag} */,
  {32'h41255606, 32'h41827fcf} /* (8, 6, 27) {real, imag} */,
  {32'hc1596dca, 32'h414e255c} /* (8, 6, 26) {real, imag} */,
  {32'h3e839ff8, 32'h4006ad42} /* (8, 6, 25) {real, imag} */,
  {32'h3eac5cd8, 32'hc0b22f40} /* (8, 6, 24) {real, imag} */,
  {32'h418d37be, 32'h4146f048} /* (8, 6, 23) {real, imag} */,
  {32'h416db58a, 32'hc07ae31e} /* (8, 6, 22) {real, imag} */,
  {32'h4138a24b, 32'hbf62e78c} /* (8, 6, 21) {real, imag} */,
  {32'hc19c9498, 32'hc1ba7193} /* (8, 6, 20) {real, imag} */,
  {32'hc08cda54, 32'h412d1013} /* (8, 6, 19) {real, imag} */,
  {32'h41014c70, 32'hc1281e2f} /* (8, 6, 18) {real, imag} */,
  {32'h4081d552, 32'hc102b2b7} /* (8, 6, 17) {real, imag} */,
  {32'hc0dfc13c, 32'hc046a443} /* (8, 6, 16) {real, imag} */,
  {32'h409cd784, 32'hc0f33dc2} /* (8, 6, 15) {real, imag} */,
  {32'h4103ab2e, 32'h402bbf04} /* (8, 6, 14) {real, imag} */,
  {32'h412c16ae, 32'hc081eea8} /* (8, 6, 13) {real, imag} */,
  {32'h41066f9f, 32'h4115083d} /* (8, 6, 12) {real, imag} */,
  {32'h41453715, 32'hc173b089} /* (8, 6, 11) {real, imag} */,
  {32'h416c69ea, 32'h4110c792} /* (8, 6, 10) {real, imag} */,
  {32'hc0fe0c32, 32'h3f62edb8} /* (8, 6, 9) {real, imag} */,
  {32'h40317a9a, 32'h40e7cab1} /* (8, 6, 8) {real, imag} */,
  {32'hc1078555, 32'h42132adc} /* (8, 6, 7) {real, imag} */,
  {32'h412525d6, 32'h41102f8f} /* (8, 6, 6) {real, imag} */,
  {32'h400b4c4c, 32'hc092a7a7} /* (8, 6, 5) {real, imag} */,
  {32'h41729525, 32'hc14f2690} /* (8, 6, 4) {real, imag} */,
  {32'h408c642c, 32'h40aa9c49} /* (8, 6, 3) {real, imag} */,
  {32'hc2026050, 32'hc163b8b4} /* (8, 6, 2) {real, imag} */,
  {32'hc141a9e0, 32'hc140adb2} /* (8, 6, 1) {real, imag} */,
  {32'hc128f784, 32'h416d50a2} /* (8, 6, 0) {real, imag} */,
  {32'hc2a45f32, 32'hc1268117} /* (8, 5, 31) {real, imag} */,
  {32'h42139c8f, 32'hc1cf5082} /* (8, 5, 30) {real, imag} */,
  {32'h41b96cb6, 32'h405ccd84} /* (8, 5, 29) {real, imag} */,
  {32'h3fec1680, 32'hc0b27da9} /* (8, 5, 28) {real, imag} */,
  {32'hc0af85c8, 32'hc0dc86c0} /* (8, 5, 27) {real, imag} */,
  {32'hc17fec05, 32'h41ecd200} /* (8, 5, 26) {real, imag} */,
  {32'h404812b8, 32'h41377a2e} /* (8, 5, 25) {real, imag} */,
  {32'h41675f10, 32'hc19b53a4} /* (8, 5, 24) {real, imag} */,
  {32'hbf59211c, 32'h412f0302} /* (8, 5, 23) {real, imag} */,
  {32'h41046867, 32'hbfdb52a8} /* (8, 5, 22) {real, imag} */,
  {32'h3f11f7f0, 32'hc1af835c} /* (8, 5, 21) {real, imag} */,
  {32'hc135eb5a, 32'hc14210f2} /* (8, 5, 20) {real, imag} */,
  {32'h41147cb8, 32'h40c2c4a4} /* (8, 5, 19) {real, imag} */,
  {32'hc0f480f6, 32'hc05d50da} /* (8, 5, 18) {real, imag} */,
  {32'hc0a1ecfa, 32'hc020f380} /* (8, 5, 17) {real, imag} */,
  {32'h410314b3, 32'h40263d22} /* (8, 5, 16) {real, imag} */,
  {32'h414ca738, 32'h3f8f37a4} /* (8, 5, 15) {real, imag} */,
  {32'hc12746a6, 32'h41b27688} /* (8, 5, 14) {real, imag} */,
  {32'hc104c9f6, 32'h406c48ec} /* (8, 5, 13) {real, imag} */,
  {32'h4121277a, 32'hc0d823c2} /* (8, 5, 12) {real, imag} */,
  {32'h411b0683, 32'hc1971048} /* (8, 5, 11) {real, imag} */,
  {32'h40e158e9, 32'h4002028c} /* (8, 5, 10) {real, imag} */,
  {32'hc04d9140, 32'h4117b90d} /* (8, 5, 9) {real, imag} */,
  {32'h41956503, 32'hc08601c4} /* (8, 5, 8) {real, imag} */,
  {32'hc1347a94, 32'hc11fbe62} /* (8, 5, 7) {real, imag} */,
  {32'hc050a0d8, 32'h4155a3bd} /* (8, 5, 6) {real, imag} */,
  {32'h4241590c, 32'h420f191d} /* (8, 5, 5) {real, imag} */,
  {32'hc199a4ea, 32'hc1110346} /* (8, 5, 4) {real, imag} */,
  {32'hc17f891e, 32'hbed0c570} /* (8, 5, 3) {real, imag} */,
  {32'h41c4c139, 32'h4235c15c} /* (8, 5, 2) {real, imag} */,
  {32'hc1e1dd3a, 32'hc2803406} /* (8, 5, 1) {real, imag} */,
  {32'hc285626f, 32'hc1af64cd} /* (8, 5, 0) {real, imag} */,
  {32'h41cd1bda, 32'h42c3a0d8} /* (8, 4, 31) {real, imag} */,
  {32'hc2ac3a41, 32'hc2a30b6d} /* (8, 4, 30) {real, imag} */,
  {32'hc1bd52fa, 32'hc0a1fec8} /* (8, 4, 29) {real, imag} */,
  {32'h41b762c1, 32'h4193291a} /* (8, 4, 28) {real, imag} */,
  {32'hc18e30f6, 32'hc175b074} /* (8, 4, 27) {real, imag} */,
  {32'hc102be28, 32'h4109bfce} /* (8, 4, 26) {real, imag} */,
  {32'h40f9daf2, 32'h40d571dc} /* (8, 4, 25) {real, imag} */,
  {32'hc1266fa4, 32'hc15f1371} /* (8, 4, 24) {real, imag} */,
  {32'h41b4e8f0, 32'hc083a134} /* (8, 4, 23) {real, imag} */,
  {32'h413c69c6, 32'hc1694c04} /* (8, 4, 22) {real, imag} */,
  {32'hbf85bf0c, 32'h41622b63} /* (8, 4, 21) {real, imag} */,
  {32'h4064a5ae, 32'h408acd0c} /* (8, 4, 20) {real, imag} */,
  {32'hc04f186e, 32'h40759e8d} /* (8, 4, 19) {real, imag} */,
  {32'h3f7887d8, 32'hc14984c5} /* (8, 4, 18) {real, imag} */,
  {32'hc1096498, 32'hbed20fe0} /* (8, 4, 17) {real, imag} */,
  {32'h41418759, 32'hbf6c4b78} /* (8, 4, 16) {real, imag} */,
  {32'hc0d7fe1a, 32'hc10b5554} /* (8, 4, 15) {real, imag} */,
  {32'h40d0ba30, 32'hc11b4534} /* (8, 4, 14) {real, imag} */,
  {32'hbe9c3290, 32'h41a7fdbe} /* (8, 4, 13) {real, imag} */,
  {32'h3fa32af4, 32'h405b2d12} /* (8, 4, 12) {real, imag} */,
  {32'h4194bde1, 32'h4072f5fa} /* (8, 4, 11) {real, imag} */,
  {32'hc119e39d, 32'h409558cb} /* (8, 4, 10) {real, imag} */,
  {32'hc0d0dfe5, 32'h4091c0a3} /* (8, 4, 9) {real, imag} */,
  {32'h4148bd09, 32'hc224d9bc} /* (8, 4, 8) {real, imag} */,
  {32'h4092b5da, 32'hbfd4d568} /* (8, 4, 7) {real, imag} */,
  {32'h41f62477, 32'hc064245c} /* (8, 4, 6) {real, imag} */,
  {32'hc073e91d, 32'hc21139ed} /* (8, 4, 5) {real, imag} */,
  {32'h41600eac, 32'h404f0ee8} /* (8, 4, 4) {real, imag} */,
  {32'hc23f514c, 32'h41ef7074} /* (8, 4, 3) {real, imag} */,
  {32'hc2d2d024, 32'hc28dc6d8} /* (8, 4, 2) {real, imag} */,
  {32'h431b5363, 32'h428fdba4} /* (8, 4, 1) {real, imag} */,
  {32'h425cba62, 32'h41cb1984} /* (8, 4, 0) {real, imag} */,
  {32'hc3093e46, 32'h423626fc} /* (8, 3, 31) {real, imag} */,
  {32'h42894744, 32'hc3190739} /* (8, 3, 30) {real, imag} */,
  {32'h4114dccb, 32'h420a6de0} /* (8, 3, 29) {real, imag} */,
  {32'h4206a215, 32'h40b00a0c} /* (8, 3, 28) {real, imag} */,
  {32'hc22c0982, 32'hc0c53252} /* (8, 3, 27) {real, imag} */,
  {32'hc1377f2f, 32'h3fb4a574} /* (8, 3, 26) {real, imag} */,
  {32'hc1c5f9d7, 32'h41b3ce37} /* (8, 3, 25) {real, imag} */,
  {32'hc1c19c86, 32'hc1dee8f4} /* (8, 3, 24) {real, imag} */,
  {32'h3ef3f120, 32'hc1120a8a} /* (8, 3, 23) {real, imag} */,
  {32'h41b014cf, 32'h4114608e} /* (8, 3, 22) {real, imag} */,
  {32'h3f9272ea, 32'h41107c32} /* (8, 3, 21) {real, imag} */,
  {32'h40b4b810, 32'h400f69e6} /* (8, 3, 20) {real, imag} */,
  {32'h414214fb, 32'h41875f48} /* (8, 3, 19) {real, imag} */,
  {32'hc0cbf336, 32'hc119a022} /* (8, 3, 18) {real, imag} */,
  {32'h41017329, 32'hbe050ff0} /* (8, 3, 17) {real, imag} */,
  {32'hc16f6542, 32'h412959d7} /* (8, 3, 16) {real, imag} */,
  {32'hc18d1aa0, 32'h405a01d8} /* (8, 3, 15) {real, imag} */,
  {32'hc072e101, 32'hc12a0b76} /* (8, 3, 14) {real, imag} */,
  {32'hc03ae50c, 32'hc0408295} /* (8, 3, 13) {real, imag} */,
  {32'h413e90cb, 32'hc0527004} /* (8, 3, 12) {real, imag} */,
  {32'h40cfac72, 32'hc06f0eaf} /* (8, 3, 11) {real, imag} */,
  {32'hc10ab030, 32'h3ee74d38} /* (8, 3, 10) {real, imag} */,
  {32'h3f175ec0, 32'h40ad7edd} /* (8, 3, 9) {real, imag} */,
  {32'h40539718, 32'h4157fcbc} /* (8, 3, 8) {real, imag} */,
  {32'hc1c471b5, 32'h40348a10} /* (8, 3, 7) {real, imag} */,
  {32'hc0e275de, 32'h4072ee5c} /* (8, 3, 6) {real, imag} */,
  {32'h4104af16, 32'h41d7e300} /* (8, 3, 5) {real, imag} */,
  {32'hc25a96f3, 32'h41c322c6} /* (8, 3, 4) {real, imag} */,
  {32'hc19fe610, 32'h41096a58} /* (8, 3, 3) {real, imag} */,
  {32'h41088d04, 32'hc2afbae0} /* (8, 3, 2) {real, imag} */,
  {32'h42e35e97, 32'h42cfbbd8} /* (8, 3, 1) {real, imag} */,
  {32'h418dfd16, 32'hc2084645} /* (8, 3, 0) {real, imag} */,
  {32'hc498727c, 32'hc1ffb2f2} /* (8, 2, 31) {real, imag} */,
  {32'h440a3d64, 32'hc319eda6} /* (8, 2, 30) {real, imag} */,
  {32'hc1fb0fdb, 32'h42920442} /* (8, 2, 29) {real, imag} */,
  {32'hc1ff7fdc, 32'h428ed330} /* (8, 2, 28) {real, imag} */,
  {32'h42a003a0, 32'hc21caf60} /* (8, 2, 27) {real, imag} */,
  {32'h41a6cd38, 32'hc13f15dd} /* (8, 2, 26) {real, imag} */,
  {32'h41b7d1e8, 32'h417e53be} /* (8, 2, 25) {real, imag} */,
  {32'h41958887, 32'h3d0cca00} /* (8, 2, 24) {real, imag} */,
  {32'hc10e917f, 32'hc01d929a} /* (8, 2, 23) {real, imag} */,
  {32'hc1152825, 32'hc06b0078} /* (8, 2, 22) {real, imag} */,
  {32'hc107f4f8, 32'hc0fc9800} /* (8, 2, 21) {real, imag} */,
  {32'h4178535d, 32'hc1cf1b82} /* (8, 2, 20) {real, imag} */,
  {32'h3f0e9734, 32'hc130bbed} /* (8, 2, 19) {real, imag} */,
  {32'hc11a609b, 32'hbea83950} /* (8, 2, 18) {real, imag} */,
  {32'h418739ba, 32'h411d214c} /* (8, 2, 17) {real, imag} */,
  {32'hc121e42e, 32'h411acf0c} /* (8, 2, 16) {real, imag} */,
  {32'hc148bf24, 32'h40d7b4b5} /* (8, 2, 15) {real, imag} */,
  {32'hc0fced45, 32'h41075247} /* (8, 2, 14) {real, imag} */,
  {32'h411e21f4, 32'hc0e13645} /* (8, 2, 13) {real, imag} */,
  {32'h4153a7cb, 32'hc131c74c} /* (8, 2, 12) {real, imag} */,
  {32'hbfda6a86, 32'h415848fc} /* (8, 2, 11) {real, imag} */,
  {32'hc0bbccc2, 32'hbf6216b0} /* (8, 2, 10) {real, imag} */,
  {32'h416c9750, 32'h40e19701} /* (8, 2, 9) {real, imag} */,
  {32'hc08f4426, 32'h40018f42} /* (8, 2, 8) {real, imag} */,
  {32'hc190a884, 32'hc2039adc} /* (8, 2, 7) {real, imag} */,
  {32'h3fe42078, 32'h40e0be35} /* (8, 2, 6) {real, imag} */,
  {32'h428c6076, 32'h41dbbdea} /* (8, 2, 5) {real, imag} */,
  {32'hc2d758c2, 32'hc1c3bede} /* (8, 2, 4) {real, imag} */,
  {32'hc1e50215, 32'h40602560} /* (8, 2, 3) {real, imag} */,
  {32'h43cce94e, 32'hc2ad8e00} /* (8, 2, 2) {real, imag} */,
  {32'hc4203dbc, 32'h43212c7c} /* (8, 2, 1) {real, imag} */,
  {32'hc41b20e7, 32'hc3158d32} /* (8, 2, 0) {real, imag} */,
  {32'h44c3e72d, 32'hc3c6ca94} /* (8, 1, 31) {real, imag} */,
  {32'hc3ab8065, 32'h42969374} /* (8, 1, 30) {real, imag} */,
  {32'hc100a106, 32'hc0fe2978} /* (8, 1, 29) {real, imag} */,
  {32'h428394cd, 32'h42a07ef2} /* (8, 1, 28) {real, imag} */,
  {32'hc2b5cc2c, 32'hc123a32d} /* (8, 1, 27) {real, imag} */,
  {32'hc19807b8, 32'h412ed425} /* (8, 1, 26) {real, imag} */,
  {32'h4195d823, 32'hc15cee22} /* (8, 1, 25) {real, imag} */,
  {32'hc211bc7d, 32'hbea24140} /* (8, 1, 24) {real, imag} */,
  {32'h40933ae0, 32'h415d209e} /* (8, 1, 23) {real, imag} */,
  {32'h400cc0b8, 32'h40dbd85f} /* (8, 1, 22) {real, imag} */,
  {32'hc22e581e, 32'h40c9eff2} /* (8, 1, 21) {real, imag} */,
  {32'h414e6234, 32'hc1a20ee9} /* (8, 1, 20) {real, imag} */,
  {32'hc03c7b21, 32'hc09ef37c} /* (8, 1, 19) {real, imag} */,
  {32'hc12a4c87, 32'h41989ca2} /* (8, 1, 18) {real, imag} */,
  {32'hc01f94a6, 32'h3f31bf3c} /* (8, 1, 17) {real, imag} */,
  {32'h409f1e63, 32'h3f77e51e} /* (8, 1, 16) {real, imag} */,
  {32'h4087c8b9, 32'h411b5098} /* (8, 1, 15) {real, imag} */,
  {32'h40e556b2, 32'hc18606e2} /* (8, 1, 14) {real, imag} */,
  {32'h40670ff6, 32'hbf8e4e50} /* (8, 1, 13) {real, imag} */,
  {32'h3fbe162c, 32'hc19ccdf0} /* (8, 1, 12) {real, imag} */,
  {32'hc1114d2c, 32'hc1aec71a} /* (8, 1, 11) {real, imag} */,
  {32'hc1bdb8a6, 32'hc0cda082} /* (8, 1, 10) {real, imag} */,
  {32'hc109eb2a, 32'hc18b9a8a} /* (8, 1, 9) {real, imag} */,
  {32'hc01f0128, 32'hc1e99d99} /* (8, 1, 8) {real, imag} */,
  {32'h412e5da6, 32'h4149af36} /* (8, 1, 7) {real, imag} */,
  {32'hc1d6180e, 32'hc069fab4} /* (8, 1, 6) {real, imag} */,
  {32'hc29f7400, 32'hc1a6fb00} /* (8, 1, 5) {real, imag} */,
  {32'h42699c56, 32'hc1835cb3} /* (8, 1, 4) {real, imag} */,
  {32'hc21060a1, 32'hc2435b96} /* (8, 1, 3) {real, imag} */,
  {32'hc40af8a8, 32'hc401b2e0} /* (8, 1, 2) {real, imag} */,
  {32'h450bb595, 32'h448a3849} /* (8, 1, 1) {real, imag} */,
  {32'h4504ce84, 32'h436653ae} /* (8, 1, 0) {real, imag} */,
  {32'h44a04da9, 32'hc4855672} /* (8, 0, 31) {real, imag} */,
  {32'hc32dcf1c, 32'h43a32011} /* (8, 0, 30) {real, imag} */,
  {32'hc106b557, 32'h409f5e94} /* (8, 0, 29) {real, imag} */,
  {32'hc0c079a0, 32'h41d89bdf} /* (8, 0, 28) {real, imag} */,
  {32'hc28e92c8, 32'h40aaefa2} /* (8, 0, 27) {real, imag} */,
  {32'h41fe832a, 32'hc16fa759} /* (8, 0, 26) {real, imag} */,
  {32'hc11fa627, 32'hc1956852} /* (8, 0, 25) {real, imag} */,
  {32'h41bdd5ec, 32'h41dfd780} /* (8, 0, 24) {real, imag} */,
  {32'h41018c46, 32'hbf8a9a0c} /* (8, 0, 23) {real, imag} */,
  {32'hbf95a502, 32'h41b61edd} /* (8, 0, 22) {real, imag} */,
  {32'hc1823ac5, 32'h4078373c} /* (8, 0, 21) {real, imag} */,
  {32'hc134a3e7, 32'hc1c47486} /* (8, 0, 20) {real, imag} */,
  {32'h41503e82, 32'hc06662b8} /* (8, 0, 19) {real, imag} */,
  {32'hc09536d3, 32'h40b0edf6} /* (8, 0, 18) {real, imag} */,
  {32'hc1149894, 32'h3deed660} /* (8, 0, 17) {real, imag} */,
  {32'hc1270673, 32'h00000000} /* (8, 0, 16) {real, imag} */,
  {32'hc1149894, 32'hbdeed660} /* (8, 0, 15) {real, imag} */,
  {32'hc09536d3, 32'hc0b0edf6} /* (8, 0, 14) {real, imag} */,
  {32'h41503e82, 32'h406662b8} /* (8, 0, 13) {real, imag} */,
  {32'hc134a3e7, 32'h41c47486} /* (8, 0, 12) {real, imag} */,
  {32'hc1823ac5, 32'hc078373c} /* (8, 0, 11) {real, imag} */,
  {32'hbf95a502, 32'hc1b61edd} /* (8, 0, 10) {real, imag} */,
  {32'h41018c46, 32'h3f8a9a0c} /* (8, 0, 9) {real, imag} */,
  {32'h41bdd5ec, 32'hc1dfd780} /* (8, 0, 8) {real, imag} */,
  {32'hc11fa627, 32'h41956852} /* (8, 0, 7) {real, imag} */,
  {32'h41fe832a, 32'h416fa759} /* (8, 0, 6) {real, imag} */,
  {32'hc28e92c8, 32'hc0aaefa2} /* (8, 0, 5) {real, imag} */,
  {32'hc0c079a0, 32'hc1d89bdf} /* (8, 0, 4) {real, imag} */,
  {32'hc106b557, 32'hc09f5e94} /* (8, 0, 3) {real, imag} */,
  {32'hc32dcf1c, 32'hc3a32011} /* (8, 0, 2) {real, imag} */,
  {32'h44a04da9, 32'h44855672} /* (8, 0, 1) {real, imag} */,
  {32'h4509bc66, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h44e46005, 32'hc45ac369} /* (7, 31, 31) {real, imag} */,
  {32'hc3e86dfe, 32'h43e6db87} /* (7, 31, 30) {real, imag} */,
  {32'hc233fe73, 32'h42bea9b8} /* (7, 31, 29) {real, imag} */,
  {32'h4245eefc, 32'h41582628} /* (7, 31, 28) {real, imag} */,
  {32'hc2947832, 32'h42051748} /* (7, 31, 27) {real, imag} */,
  {32'hc1a184f3, 32'h3fee1918} /* (7, 31, 26) {real, imag} */,
  {32'h41846d3d, 32'hc1aafaa4} /* (7, 31, 25) {real, imag} */,
  {32'hc165b8e3, 32'h422474f4} /* (7, 31, 24) {real, imag} */,
  {32'hc10ef8eb, 32'hbffe84c2} /* (7, 31, 23) {real, imag} */,
  {32'hc0a31a3c, 32'hc12874cf} /* (7, 31, 22) {real, imag} */,
  {32'hc18baf35, 32'h4173dd65} /* (7, 31, 21) {real, imag} */,
  {32'h3f9a5122, 32'h411f9a44} /* (7, 31, 20) {real, imag} */,
  {32'hc13eed78, 32'h412c31bb} /* (7, 31, 19) {real, imag} */,
  {32'hc11d4807, 32'hc04d7a80} /* (7, 31, 18) {real, imag} */,
  {32'hc058398b, 32'hc0f0c7a2} /* (7, 31, 17) {real, imag} */,
  {32'hbef30e68, 32'h41894ed0} /* (7, 31, 16) {real, imag} */,
  {32'hc0ec9447, 32'hbeab8dd8} /* (7, 31, 15) {real, imag} */,
  {32'h3f8eb8f4, 32'hc1a94be0} /* (7, 31, 14) {real, imag} */,
  {32'h4025fd46, 32'hc1039e28} /* (7, 31, 13) {real, imag} */,
  {32'h3f143e00, 32'hc08934b4} /* (7, 31, 12) {real, imag} */,
  {32'hc117b321, 32'hc1f4c342} /* (7, 31, 11) {real, imag} */,
  {32'h419bf955, 32'h4090a892} /* (7, 31, 10) {real, imag} */,
  {32'h40a3d984, 32'hc0f70729} /* (7, 31, 9) {real, imag} */,
  {32'hc1c5bb0f, 32'hc1c386b2} /* (7, 31, 8) {real, imag} */,
  {32'h41141749, 32'h40514667} /* (7, 31, 7) {real, imag} */,
  {32'hc198a781, 32'hc1e6c1b7} /* (7, 31, 6) {real, imag} */,
  {32'hc2bcfb34, 32'hbf4d7808} /* (7, 31, 5) {real, imag} */,
  {32'h4252bdee, 32'hc28425f4} /* (7, 31, 4) {real, imag} */,
  {32'h423125cc, 32'h421fd7f0} /* (7, 31, 3) {real, imag} */,
  {32'hc389f35d, 32'hc2181785} /* (7, 31, 2) {real, imag} */,
  {32'h44a4cfda, 32'h43a909f4} /* (7, 31, 1) {real, imag} */,
  {32'h44deaf4e, 32'hc3699daf} /* (7, 31, 0) {real, imag} */,
  {32'hc401a06e, 32'hc2c00cee} /* (7, 30, 31) {real, imag} */,
  {32'h43bfb028, 32'h4252eee3} /* (7, 30, 30) {real, imag} */,
  {32'hc1e510e5, 32'hc206f27a} /* (7, 30, 29) {real, imag} */,
  {32'hc2ed82c2, 32'h41a45c96} /* (7, 30, 28) {real, imag} */,
  {32'h425a86e0, 32'hc210dd2d} /* (7, 30, 27) {real, imag} */,
  {32'h4114d677, 32'hbf9d75c8} /* (7, 30, 26) {real, imag} */,
  {32'hc0d46ab6, 32'h41abb5e4} /* (7, 30, 25) {real, imag} */,
  {32'hc04a8438, 32'hc0e6ec32} /* (7, 30, 24) {real, imag} */,
  {32'h40fdfff3, 32'hc1ad5409} /* (7, 30, 23) {real, imag} */,
  {32'h411e3bfc, 32'hbe92d3a0} /* (7, 30, 22) {real, imag} */,
  {32'h417320d2, 32'hc1473896} /* (7, 30, 21) {real, imag} */,
  {32'hc1846e42, 32'hc12be0dc} /* (7, 30, 20) {real, imag} */,
  {32'hc18bbdb3, 32'h3f494fd0} /* (7, 30, 19) {real, imag} */,
  {32'h410ca669, 32'h41102aaf} /* (7, 30, 18) {real, imag} */,
  {32'h412490e8, 32'hc0d22017} /* (7, 30, 17) {real, imag} */,
  {32'hc05779f8, 32'hc074dd6a} /* (7, 30, 16) {real, imag} */,
  {32'hbda00920, 32'hbfb42c24} /* (7, 30, 15) {real, imag} */,
  {32'h4025f04c, 32'h40fa5f60} /* (7, 30, 14) {real, imag} */,
  {32'hc097bc02, 32'hbf0d77c0} /* (7, 30, 13) {real, imag} */,
  {32'h41813f15, 32'h418553c3} /* (7, 30, 12) {real, imag} */,
  {32'h41867f99, 32'h408ce1fb} /* (7, 30, 11) {real, imag} */,
  {32'h41ad37ac, 32'hc1b12e16} /* (7, 30, 10) {real, imag} */,
  {32'h40e886ca, 32'h40a44ae9} /* (7, 30, 9) {real, imag} */,
  {32'h41fd0b22, 32'hc10b4666} /* (7, 30, 8) {real, imag} */,
  {32'hc19e8dac, 32'hc06e44a0} /* (7, 30, 7) {real, imag} */,
  {32'h4197941f, 32'h413919e7} /* (7, 30, 6) {real, imag} */,
  {32'h4235edfc, 32'h42169f3e} /* (7, 30, 5) {real, imag} */,
  {32'hc0bc7818, 32'hc2250f79} /* (7, 30, 4) {real, imag} */,
  {32'hc241ec25, 32'hc249bce9} /* (7, 30, 3) {real, imag} */,
  {32'h43f44116, 32'h43049647} /* (7, 30, 2) {real, imag} */,
  {32'hc47c0336, 32'hc188d424} /* (7, 30, 1) {real, imag} */,
  {32'hc4020d36, 32'h4335fa66} /* (7, 30, 0) {real, imag} */,
  {32'h43043c7c, 32'hc3057b78} /* (7, 29, 31) {real, imag} */,
  {32'hc1a9105c, 32'h4261f7be} /* (7, 29, 30) {real, imag} */,
  {32'hc0a802b7, 32'h410ff03a} /* (7, 29, 29) {real, imag} */,
  {32'hc243bbb3, 32'hc1b62de3} /* (7, 29, 28) {real, imag} */,
  {32'h41fde1fa, 32'h409b275c} /* (7, 29, 27) {real, imag} */,
  {32'h4024ca54, 32'h412e0949} /* (7, 29, 26) {real, imag} */,
  {32'hc064a047, 32'hc09ebce2} /* (7, 29, 25) {real, imag} */,
  {32'hc09f597f, 32'hc12916c2} /* (7, 29, 24) {real, imag} */,
  {32'h40d684a1, 32'hc16f3847} /* (7, 29, 23) {real, imag} */,
  {32'hbfb8eaf2, 32'h3fd20ec0} /* (7, 29, 22) {real, imag} */,
  {32'hc0c37236, 32'h41a4e890} /* (7, 29, 21) {real, imag} */,
  {32'h3f5df110, 32'h41698afb} /* (7, 29, 20) {real, imag} */,
  {32'hc0c4cb0a, 32'h405c5322} /* (7, 29, 19) {real, imag} */,
  {32'h41704e0a, 32'hc11f7362} /* (7, 29, 18) {real, imag} */,
  {32'h404c3cc8, 32'hc08c597a} /* (7, 29, 17) {real, imag} */,
  {32'h3f9c0f3c, 32'h41320dcc} /* (7, 29, 16) {real, imag} */,
  {32'hc02ce640, 32'hbe52f7e0} /* (7, 29, 15) {real, imag} */,
  {32'h3ebaf8d0, 32'h40ff8842} /* (7, 29, 14) {real, imag} */,
  {32'h418b3650, 32'hc0be71e4} /* (7, 29, 13) {real, imag} */,
  {32'hc12c9c55, 32'h407810d4} /* (7, 29, 12) {real, imag} */,
  {32'h4053417b, 32'h418785b6} /* (7, 29, 11) {real, imag} */,
  {32'h3ead01e8, 32'hc05a4ed5} /* (7, 29, 10) {real, imag} */,
  {32'h3fd60968, 32'hbdcc3340} /* (7, 29, 9) {real, imag} */,
  {32'hc1b7a790, 32'h41b37252} /* (7, 29, 8) {real, imag} */,
  {32'hc1c0829c, 32'hc198d497} /* (7, 29, 7) {real, imag} */,
  {32'hc1b852fa, 32'h40355df0} /* (7, 29, 6) {real, imag} */,
  {32'hc058e7a2, 32'hc10c36d4} /* (7, 29, 5) {real, imag} */,
  {32'h42271c10, 32'hc1caaf40} /* (7, 29, 4) {real, imag} */,
  {32'hc16905a8, 32'h3f88cbd0} /* (7, 29, 3) {real, imag} */,
  {32'h4270769c, 32'h42eccdb2} /* (7, 29, 2) {real, imag} */,
  {32'hc30efc8b, 32'hc25d5adc} /* (7, 29, 1) {real, imag} */,
  {32'h41b2150d, 32'hc107d89d} /* (7, 29, 0) {real, imag} */,
  {32'h42f063b8, 32'hc2c57a32} /* (7, 28, 31) {real, imag} */,
  {32'hc2990dcb, 32'h42ab1fba} /* (7, 28, 30) {real, imag} */,
  {32'hc185c3a1, 32'h3faf91d4} /* (7, 28, 29) {real, imag} */,
  {32'h40ebe8f6, 32'hc22712dd} /* (7, 28, 28) {real, imag} */,
  {32'hbf5edd60, 32'h4211f9ac} /* (7, 28, 27) {real, imag} */,
  {32'h41030cb3, 32'hc12c2d98} /* (7, 28, 26) {real, imag} */,
  {32'hbfffc7d0, 32'hbf0f5dc0} /* (7, 28, 25) {real, imag} */,
  {32'hc0e6e362, 32'h41968b22} /* (7, 28, 24) {real, imag} */,
  {32'h41688ac6, 32'h41a9b961} /* (7, 28, 23) {real, imag} */,
  {32'h4067b9ff, 32'h3fa83df4} /* (7, 28, 22) {real, imag} */,
  {32'h40f46279, 32'h417abb78} /* (7, 28, 21) {real, imag} */,
  {32'hc0ec5af8, 32'hc0c475a4} /* (7, 28, 20) {real, imag} */,
  {32'h41676cc0, 32'hc06738e8} /* (7, 28, 19) {real, imag} */,
  {32'hc175f890, 32'h40c1ae46} /* (7, 28, 18) {real, imag} */,
  {32'hc1500cd0, 32'hc0ced7ab} /* (7, 28, 17) {real, imag} */,
  {32'h3eb2f91e, 32'hc0ce1870} /* (7, 28, 16) {real, imag} */,
  {32'h413ee65c, 32'hbe6689e0} /* (7, 28, 15) {real, imag} */,
  {32'hc10b6e3d, 32'h40d4d238} /* (7, 28, 14) {real, imag} */,
  {32'hc0064640, 32'hc158e026} /* (7, 28, 13) {real, imag} */,
  {32'hc09e878a, 32'hc1a416ee} /* (7, 28, 12) {real, imag} */,
  {32'h402bc3fe, 32'h41a60e9b} /* (7, 28, 11) {real, imag} */,
  {32'h415b850a, 32'h40807bca} /* (7, 28, 10) {real, imag} */,
  {32'hc120e940, 32'h4124124b} /* (7, 28, 9) {real, imag} */,
  {32'hbfefeb08, 32'h419b9cba} /* (7, 28, 8) {real, imag} */,
  {32'h40a68ac1, 32'hc0440a28} /* (7, 28, 7) {real, imag} */,
  {32'hc149cb68, 32'h404fe96c} /* (7, 28, 6) {real, imag} */,
  {32'hc0eb7eb1, 32'h405c04f6} /* (7, 28, 5) {real, imag} */,
  {32'h4213734a, 32'hc0eb6c8a} /* (7, 28, 4) {real, imag} */,
  {32'h41157314, 32'h4186ddf6} /* (7, 28, 3) {real, imag} */,
  {32'hc2a85c1c, 32'h4286f907} /* (7, 28, 2) {real, imag} */,
  {32'h41175e9a, 32'hc2acb87c} /* (7, 28, 1) {real, imag} */,
  {32'h426cdcee, 32'hc068c630} /* (7, 28, 0) {real, imag} */,
  {32'hc2245525, 32'h41c6695a} /* (7, 27, 31) {real, imag} */,
  {32'h422bcdc6, 32'hc215d816} /* (7, 27, 30) {real, imag} */,
  {32'hc02ea4b0, 32'hbe57ca00} /* (7, 27, 29) {real, imag} */,
  {32'h3f38c840, 32'hc03d9c08} /* (7, 27, 28) {real, imag} */,
  {32'h41b4209c, 32'hc1271331} /* (7, 27, 27) {real, imag} */,
  {32'h41a07657, 32'hc182c462} /* (7, 27, 26) {real, imag} */,
  {32'hc126cc80, 32'hc0ade43c} /* (7, 27, 25) {real, imag} */,
  {32'h40935f5c, 32'h412b7649} /* (7, 27, 24) {real, imag} */,
  {32'h40d1ea63, 32'hbf1bcab8} /* (7, 27, 23) {real, imag} */,
  {32'h40bd048e, 32'h41679b66} /* (7, 27, 22) {real, imag} */,
  {32'hc18e6e03, 32'h40edddd6} /* (7, 27, 21) {real, imag} */,
  {32'h401296a0, 32'h41317fe6} /* (7, 27, 20) {real, imag} */,
  {32'hbfbeb399, 32'h411f3793} /* (7, 27, 19) {real, imag} */,
  {32'hc1945932, 32'hc08eedc1} /* (7, 27, 18) {real, imag} */,
  {32'hc0ea741d, 32'h40718934} /* (7, 27, 17) {real, imag} */,
  {32'h40932f00, 32'h41258512} /* (7, 27, 16) {real, imag} */,
  {32'h40710008, 32'h3da36d90} /* (7, 27, 15) {real, imag} */,
  {32'hc0e3b8c2, 32'h4164fb40} /* (7, 27, 14) {real, imag} */,
  {32'h410f3b08, 32'h3fce455a} /* (7, 27, 13) {real, imag} */,
  {32'hc0691f84, 32'h408f2456} /* (7, 27, 12) {real, imag} */,
  {32'h411e0cba, 32'hc0e1ff8f} /* (7, 27, 11) {real, imag} */,
  {32'h40d3d02f, 32'hc0371ad8} /* (7, 27, 10) {real, imag} */,
  {32'hc0d3c55e, 32'h410d5f4a} /* (7, 27, 9) {real, imag} */,
  {32'h3de16da0, 32'h41434b04} /* (7, 27, 8) {real, imag} */,
  {32'hc16a7a8e, 32'hc0c30939} /* (7, 27, 7) {real, imag} */,
  {32'hc10ab28a, 32'hc08fe854} /* (7, 27, 6) {real, imag} */,
  {32'h4136d98f, 32'h412258a2} /* (7, 27, 5) {real, imag} */,
  {32'hc1422102, 32'hc07d4d28} /* (7, 27, 4) {real, imag} */,
  {32'hc07ba380, 32'h40b0f9c2} /* (7, 27, 3) {real, imag} */,
  {32'h424eb1ae, 32'h420b7256} /* (7, 27, 2) {real, imag} */,
  {32'hc2a473b8, 32'hc06037e4} /* (7, 27, 1) {real, imag} */,
  {32'hc291524c, 32'h41d14b9c} /* (7, 27, 0) {real, imag} */,
  {32'hc193b9d5, 32'hc0e9946b} /* (7, 26, 31) {real, imag} */,
  {32'hc1d113e2, 32'h40ec2cf0} /* (7, 26, 30) {real, imag} */,
  {32'hc12f9bba, 32'hc1d075a5} /* (7, 26, 29) {real, imag} */,
  {32'h4019aa8d, 32'hbfb934b0} /* (7, 26, 28) {real, imag} */,
  {32'hc02ecab3, 32'hc0308da5} /* (7, 26, 27) {real, imag} */,
  {32'hc0bccbb8, 32'h40094240} /* (7, 26, 26) {real, imag} */,
  {32'h41e93bd0, 32'hc1661d14} /* (7, 26, 25) {real, imag} */,
  {32'h415e53c4, 32'h40909405} /* (7, 26, 24) {real, imag} */,
  {32'hc154eb66, 32'h409182ce} /* (7, 26, 23) {real, imag} */,
  {32'h40255ca0, 32'h41280a7c} /* (7, 26, 22) {real, imag} */,
  {32'h4123c58f, 32'h411b1729} /* (7, 26, 21) {real, imag} */,
  {32'hc0ffb441, 32'hc16b2218} /* (7, 26, 20) {real, imag} */,
  {32'h40a3694b, 32'h40d5c90a} /* (7, 26, 19) {real, imag} */,
  {32'hc1035005, 32'hc120de34} /* (7, 26, 18) {real, imag} */,
  {32'hc0a7d23e, 32'h3e9f0050} /* (7, 26, 17) {real, imag} */,
  {32'hc13cde08, 32'h40c460b1} /* (7, 26, 16) {real, imag} */,
  {32'hc023ccdf, 32'hc09dfd7f} /* (7, 26, 15) {real, imag} */,
  {32'hc0b8ec60, 32'hc0402754} /* (7, 26, 14) {real, imag} */,
  {32'hc0b06ddb, 32'hc119f858} /* (7, 26, 13) {real, imag} */,
  {32'h3fa0ae34, 32'h40c22b18} /* (7, 26, 12) {real, imag} */,
  {32'hc0d2eb6b, 32'h4096b662} /* (7, 26, 11) {real, imag} */,
  {32'hc0920264, 32'hc068ad34} /* (7, 26, 10) {real, imag} */,
  {32'h419449ef, 32'h40c64a8b} /* (7, 26, 9) {real, imag} */,
  {32'h3fee5368, 32'h411bad3f} /* (7, 26, 8) {real, imag} */,
  {32'h4176317a, 32'hbf182130} /* (7, 26, 7) {real, imag} */,
  {32'hc0501ac8, 32'h3e0b0f80} /* (7, 26, 6) {real, imag} */,
  {32'h4195b2eb, 32'hc18ca3a8} /* (7, 26, 5) {real, imag} */,
  {32'hc0fac502, 32'hc15cfbeb} /* (7, 26, 4) {real, imag} */,
  {32'hc09780cf, 32'h4166be86} /* (7, 26, 3) {real, imag} */,
  {32'hc058836c, 32'h414c5e3d} /* (7, 26, 2) {real, imag} */,
  {32'h40d33625, 32'hc18933b2} /* (7, 26, 1) {real, imag} */,
  {32'hbff5e64c, 32'h413b646a} /* (7, 26, 0) {real, imag} */,
  {32'hc0dd6c84, 32'hc19536a7} /* (7, 25, 31) {real, imag} */,
  {32'hc097c106, 32'h42117784} /* (7, 25, 30) {real, imag} */,
  {32'hc158e1a7, 32'hc1cae47e} /* (7, 25, 29) {real, imag} */,
  {32'h40aeee4c, 32'hc1c2c4ed} /* (7, 25, 28) {real, imag} */,
  {32'h4216df1b, 32'h410c6c8e} /* (7, 25, 27) {real, imag} */,
  {32'h41a76907, 32'hc07b301c} /* (7, 25, 26) {real, imag} */,
  {32'hc103307d, 32'h41af7cd4} /* (7, 25, 25) {real, imag} */,
  {32'hc187e855, 32'h4121c52c} /* (7, 25, 24) {real, imag} */,
  {32'h415bee02, 32'hc1c8148e} /* (7, 25, 23) {real, imag} */,
  {32'h41bbe576, 32'hc156a8b7} /* (7, 25, 22) {real, imag} */,
  {32'hc1581164, 32'hbf211a40} /* (7, 25, 21) {real, imag} */,
  {32'hc0e66e14, 32'h418a44c0} /* (7, 25, 20) {real, imag} */,
  {32'h4092eede, 32'hc1551574} /* (7, 25, 19) {real, imag} */,
  {32'h405ed06a, 32'h40f7b616} /* (7, 25, 18) {real, imag} */,
  {32'hbe8aacd8, 32'h40a205ee} /* (7, 25, 17) {real, imag} */,
  {32'hc0b4ef65, 32'h40837ec5} /* (7, 25, 16) {real, imag} */,
  {32'hc0f390a4, 32'hc01b40ee} /* (7, 25, 15) {real, imag} */,
  {32'h406eb45a, 32'h401364be} /* (7, 25, 14) {real, imag} */,
  {32'hbfabb8d8, 32'hc0e7849d} /* (7, 25, 13) {real, imag} */,
  {32'hbfa041be, 32'hc0817d28} /* (7, 25, 12) {real, imag} */,
  {32'h4070ce72, 32'h4137e75b} /* (7, 25, 11) {real, imag} */,
  {32'hc0d01160, 32'hc02fb3ab} /* (7, 25, 10) {real, imag} */,
  {32'hc10e9fde, 32'h40be0516} /* (7, 25, 9) {real, imag} */,
  {32'h41194be8, 32'h41094afa} /* (7, 25, 8) {real, imag} */,
  {32'hc1187117, 32'hc1c7916c} /* (7, 25, 7) {real, imag} */,
  {32'hbfec870c, 32'hc171a2a0} /* (7, 25, 6) {real, imag} */,
  {32'h410b9255, 32'h40a89574} /* (7, 25, 5) {real, imag} */,
  {32'hc0177096, 32'hc0af4bf6} /* (7, 25, 4) {real, imag} */,
  {32'hc1c1cbe2, 32'hc082e6f2} /* (7, 25, 3) {real, imag} */,
  {32'h410b396a, 32'h408d12c4} /* (7, 25, 2) {real, imag} */,
  {32'hc08097ac, 32'h4103c292} /* (7, 25, 1) {real, imag} */,
  {32'h415c6cf6, 32'hc1080cec} /* (7, 25, 0) {real, imag} */,
  {32'hc185bea2, 32'h4208ba72} /* (7, 24, 31) {real, imag} */,
  {32'h41abc60a, 32'hc09a63d8} /* (7, 24, 30) {real, imag} */,
  {32'h40a71798, 32'hc0f9c8ad} /* (7, 24, 29) {real, imag} */,
  {32'hc1751275, 32'h418353c9} /* (7, 24, 28) {real, imag} */,
  {32'hc18a9c0a, 32'hc041f356} /* (7, 24, 27) {real, imag} */,
  {32'hc1839bc4, 32'hbfaab288} /* (7, 24, 26) {real, imag} */,
  {32'hc1562194, 32'hc0c2a799} /* (7, 24, 25) {real, imag} */,
  {32'hc082bea0, 32'hc1ed49e8} /* (7, 24, 24) {real, imag} */,
  {32'hc17c6ebc, 32'h413580c1} /* (7, 24, 23) {real, imag} */,
  {32'h40f224d9, 32'h40b27aeb} /* (7, 24, 22) {real, imag} */,
  {32'h406c51f4, 32'hc19448a2} /* (7, 24, 21) {real, imag} */,
  {32'hc013d438, 32'h4080b5a3} /* (7, 24, 20) {real, imag} */,
  {32'hc1a678ba, 32'hc0ab537b} /* (7, 24, 19) {real, imag} */,
  {32'h41abd7d9, 32'h411d457a} /* (7, 24, 18) {real, imag} */,
  {32'h408c8756, 32'h412fee88} /* (7, 24, 17) {real, imag} */,
  {32'hc10cce62, 32'hc08cbf28} /* (7, 24, 16) {real, imag} */,
  {32'hc185b17a, 32'hc111e174} /* (7, 24, 15) {real, imag} */,
  {32'h412e1656, 32'hc111e712} /* (7, 24, 14) {real, imag} */,
  {32'hc081fc1c, 32'hbf9fc260} /* (7, 24, 13) {real, imag} */,
  {32'hc0d0db5c, 32'hc18be5fb} /* (7, 24, 12) {real, imag} */,
  {32'hc0b3c6bd, 32'hc15468ce} /* (7, 24, 11) {real, imag} */,
  {32'h3f97da88, 32'hbf596878} /* (7, 24, 10) {real, imag} */,
  {32'h41000960, 32'h41733d78} /* (7, 24, 9) {real, imag} */,
  {32'h415a3f11, 32'h41b40aad} /* (7, 24, 8) {real, imag} */,
  {32'hc10ed724, 32'h415bc6aa} /* (7, 24, 7) {real, imag} */,
  {32'h412100f8, 32'h4143c935} /* (7, 24, 6) {real, imag} */,
  {32'h41fb1944, 32'h4159517a} /* (7, 24, 5) {real, imag} */,
  {32'h41569b50, 32'hc077efea} /* (7, 24, 4) {real, imag} */,
  {32'h4102b91c, 32'h410acfe4} /* (7, 24, 3) {real, imag} */,
  {32'h41e7772d, 32'hc18daf33} /* (7, 24, 2) {real, imag} */,
  {32'hc2445dc3, 32'h41b0f6f4} /* (7, 24, 1) {real, imag} */,
  {32'hc1d59ae1, 32'h419d5430} /* (7, 24, 0) {real, imag} */,
  {32'hc1a3e8b2, 32'hbfb53f94} /* (7, 23, 31) {real, imag} */,
  {32'hc17c6eb4, 32'h4090460c} /* (7, 23, 30) {real, imag} */,
  {32'hc010ddc5, 32'hc12a54ab} /* (7, 23, 29) {real, imag} */,
  {32'h4103b555, 32'hc0fd0e40} /* (7, 23, 28) {real, imag} */,
  {32'hc09c122e, 32'hc13099cb} /* (7, 23, 27) {real, imag} */,
  {32'hc1634717, 32'h40f38c0e} /* (7, 23, 26) {real, imag} */,
  {32'h3f81b375, 32'hc1809196} /* (7, 23, 25) {real, imag} */,
  {32'hc07344c6, 32'h40357eaa} /* (7, 23, 24) {real, imag} */,
  {32'hc125075c, 32'hc1add430} /* (7, 23, 23) {real, imag} */,
  {32'h40f1f827, 32'h40d0a882} /* (7, 23, 22) {real, imag} */,
  {32'h410f7d66, 32'hbf848a34} /* (7, 23, 21) {real, imag} */,
  {32'h4038f8d8, 32'hc0a62cc7} /* (7, 23, 20) {real, imag} */,
  {32'hc003aa64, 32'h41594fea} /* (7, 23, 19) {real, imag} */,
  {32'h4101c450, 32'hc01c057d} /* (7, 23, 18) {real, imag} */,
  {32'h40840bd2, 32'h41291a2e} /* (7, 23, 17) {real, imag} */,
  {32'h4059950a, 32'hc10b14f2} /* (7, 23, 16) {real, imag} */,
  {32'h407ef25a, 32'hc0f2c3b0} /* (7, 23, 15) {real, imag} */,
  {32'hc176a155, 32'h40ae0d62} /* (7, 23, 14) {real, imag} */,
  {32'h416d8db2, 32'hc137a2ad} /* (7, 23, 13) {real, imag} */,
  {32'h40118b70, 32'h4056a280} /* (7, 23, 12) {real, imag} */,
  {32'hbf43aa10, 32'h4115329b} /* (7, 23, 11) {real, imag} */,
  {32'h41a93f92, 32'h40ae5ddf} /* (7, 23, 10) {real, imag} */,
  {32'hc18d934e, 32'h4188890a} /* (7, 23, 9) {real, imag} */,
  {32'h40ba57d0, 32'h41576f5c} /* (7, 23, 8) {real, imag} */,
  {32'hc18c599b, 32'h40acb604} /* (7, 23, 7) {real, imag} */,
  {32'h3fe78818, 32'h40b594ca} /* (7, 23, 6) {real, imag} */,
  {32'hc168ea77, 32'hc0f0daf6} /* (7, 23, 5) {real, imag} */,
  {32'hbf818f2a, 32'hbebbfb90} /* (7, 23, 4) {real, imag} */,
  {32'hbf34d3a8, 32'h3f070108} /* (7, 23, 3) {real, imag} */,
  {32'h415f4c0a, 32'h41b3a7da} /* (7, 23, 2) {real, imag} */,
  {32'hc147f4f4, 32'hc1c8ff99} /* (7, 23, 1) {real, imag} */,
  {32'hc10cab70, 32'h40aa75bb} /* (7, 23, 0) {real, imag} */,
  {32'h418882a9, 32'h4095d1f6} /* (7, 22, 31) {real, imag} */,
  {32'h3f82fdbc, 32'h413cd440} /* (7, 22, 30) {real, imag} */,
  {32'hc0bbae5b, 32'hc1a5982e} /* (7, 22, 29) {real, imag} */,
  {32'hbfe87f66, 32'h3fccdc9c} /* (7, 22, 28) {real, imag} */,
  {32'h41a3294a, 32'h40add336} /* (7, 22, 27) {real, imag} */,
  {32'hc1251743, 32'hc1468402} /* (7, 22, 26) {real, imag} */,
  {32'hc0c4900e, 32'h4152e7ee} /* (7, 22, 25) {real, imag} */,
  {32'hc080ef45, 32'h405d1a5a} /* (7, 22, 24) {real, imag} */,
  {32'h40d9d1c7, 32'hc0be809b} /* (7, 22, 23) {real, imag} */,
  {32'hc14b8a6c, 32'hc06a8332} /* (7, 22, 22) {real, imag} */,
  {32'h40f8ab78, 32'h41a9c9e2} /* (7, 22, 21) {real, imag} */,
  {32'h41132994, 32'hc18c2d91} /* (7, 22, 20) {real, imag} */,
  {32'h4171a90e, 32'h40f572c3} /* (7, 22, 19) {real, imag} */,
  {32'hc14d89c3, 32'h41421b37} /* (7, 22, 18) {real, imag} */,
  {32'hbfc43ac6, 32'h40a5e844} /* (7, 22, 17) {real, imag} */,
  {32'hbe7c1ca0, 32'h40d8a611} /* (7, 22, 16) {real, imag} */,
  {32'hc1094e9a, 32'h40d07b9e} /* (7, 22, 15) {real, imag} */,
  {32'hc065f34c, 32'hbeebb9f0} /* (7, 22, 14) {real, imag} */,
  {32'h40f647c9, 32'hc18f47b8} /* (7, 22, 13) {real, imag} */,
  {32'h41c8129a, 32'hbf6d4e20} /* (7, 22, 12) {real, imag} */,
  {32'h41d6fd4b, 32'h3f1a2da0} /* (7, 22, 11) {real, imag} */,
  {32'hc1956590, 32'h4104fa9e} /* (7, 22, 10) {real, imag} */,
  {32'h40d1ca1c, 32'h40ea8bae} /* (7, 22, 9) {real, imag} */,
  {32'hc159c1e3, 32'hc081fc71} /* (7, 22, 8) {real, imag} */,
  {32'h406a54c2, 32'h417fd1dc} /* (7, 22, 7) {real, imag} */,
  {32'h41168c53, 32'h409623a9} /* (7, 22, 6) {real, imag} */,
  {32'h410a3e92, 32'h415a078d} /* (7, 22, 5) {real, imag} */,
  {32'h3f310efc, 32'hc185fc28} /* (7, 22, 4) {real, imag} */,
  {32'hc13719f2, 32'h4140d69b} /* (7, 22, 3) {real, imag} */,
  {32'hc14630ac, 32'hc0bd22a0} /* (7, 22, 2) {real, imag} */,
  {32'hbeb2af60, 32'hc0d42cf5} /* (7, 22, 1) {real, imag} */,
  {32'hc06b884c, 32'hc1d2b5c6} /* (7, 22, 0) {real, imag} */,
  {32'h3fcdb350, 32'h41d17db1} /* (7, 21, 31) {real, imag} */,
  {32'hc0969c6f, 32'hc1832e61} /* (7, 21, 30) {real, imag} */,
  {32'h416543e2, 32'h41b77cc1} /* (7, 21, 29) {real, imag} */,
  {32'h40cc5f40, 32'h41b2c1ce} /* (7, 21, 28) {real, imag} */,
  {32'hc03f3f74, 32'hc109e67c} /* (7, 21, 27) {real, imag} */,
  {32'h411bc99a, 32'hc1a789de} /* (7, 21, 26) {real, imag} */,
  {32'h411dbd94, 32'hc09d6376} /* (7, 21, 25) {real, imag} */,
  {32'hc018252c, 32'hc0902c8e} /* (7, 21, 24) {real, imag} */,
  {32'h414918f2, 32'h419376bf} /* (7, 21, 23) {real, imag} */,
  {32'hc18973e0, 32'hc19d56b6} /* (7, 21, 22) {real, imag} */,
  {32'hc075e3b8, 32'hc13a6fa0} /* (7, 21, 21) {real, imag} */,
  {32'h3f6f6e68, 32'h4149e075} /* (7, 21, 20) {real, imag} */,
  {32'hc00808e4, 32'h3f2baec8} /* (7, 21, 19) {real, imag} */,
  {32'hc144b906, 32'h415244d0} /* (7, 21, 18) {real, imag} */,
  {32'h4121e5d8, 32'hc0ccee7b} /* (7, 21, 17) {real, imag} */,
  {32'h411d38f0, 32'hc08d4c9e} /* (7, 21, 16) {real, imag} */,
  {32'hc0fa9f6b, 32'h40853ebd} /* (7, 21, 15) {real, imag} */,
  {32'h412b4a7f, 32'hc0b352f6} /* (7, 21, 14) {real, imag} */,
  {32'h40c7a9da, 32'h3f1864c8} /* (7, 21, 13) {real, imag} */,
  {32'h41c62406, 32'hbf589b24} /* (7, 21, 12) {real, imag} */,
  {32'h418962ff, 32'h411918f2} /* (7, 21, 11) {real, imag} */,
  {32'hc095bd6e, 32'h4105abdd} /* (7, 21, 10) {real, imag} */,
  {32'hc1d39410, 32'hc16c07e5} /* (7, 21, 9) {real, imag} */,
  {32'hc0eb2e5a, 32'hc161b4fe} /* (7, 21, 8) {real, imag} */,
  {32'hc1b5b176, 32'h4067affe} /* (7, 21, 7) {real, imag} */,
  {32'h410b401b, 32'hc0d0c105} /* (7, 21, 6) {real, imag} */,
  {32'h3fe61b48, 32'hc105c4f9} /* (7, 21, 5) {real, imag} */,
  {32'hc1328038, 32'h4118b778} /* (7, 21, 4) {real, imag} */,
  {32'h411bab4c, 32'hc13335a0} /* (7, 21, 3) {real, imag} */,
  {32'h41b2056c, 32'hbe26c680} /* (7, 21, 2) {real, imag} */,
  {32'h3f0e2b00, 32'h40e77718} /* (7, 21, 1) {real, imag} */,
  {32'hc122e90c, 32'h412458d1} /* (7, 21, 0) {real, imag} */,
  {32'h417bb391, 32'h3f7186dc} /* (7, 20, 31) {real, imag} */,
  {32'h3f82cfe8, 32'h4069a7a4} /* (7, 20, 30) {real, imag} */,
  {32'hc19545bc, 32'h40d505fb} /* (7, 20, 29) {real, imag} */,
  {32'h4190a7b4, 32'h4140f98f} /* (7, 20, 28) {real, imag} */,
  {32'hc1887442, 32'h400faf84} /* (7, 20, 27) {real, imag} */,
  {32'hc039d5a5, 32'hc162a084} /* (7, 20, 26) {real, imag} */,
  {32'h416141d8, 32'h40e3025e} /* (7, 20, 25) {real, imag} */,
  {32'h3dbfd940, 32'hc0da5c30} /* (7, 20, 24) {real, imag} */,
  {32'hc16444bc, 32'h401f49a0} /* (7, 20, 23) {real, imag} */,
  {32'h414b822c, 32'hc1aebbb2} /* (7, 20, 22) {real, imag} */,
  {32'hc0475460, 32'h408fcab2} /* (7, 20, 21) {real, imag} */,
  {32'h41599a99, 32'h3f27eb98} /* (7, 20, 20) {real, imag} */,
  {32'hc146d037, 32'hc12f92d9} /* (7, 20, 19) {real, imag} */,
  {32'h40a9b576, 32'hc15ad8ec} /* (7, 20, 18) {real, imag} */,
  {32'hc05e01bc, 32'hc0a53c40} /* (7, 20, 17) {real, imag} */,
  {32'h3efbdf68, 32'h414b2b0a} /* (7, 20, 16) {real, imag} */,
  {32'h4144dfd9, 32'hbf752dd8} /* (7, 20, 15) {real, imag} */,
  {32'hc0318f0a, 32'hbf524c74} /* (7, 20, 14) {real, imag} */,
  {32'hc1182b34, 32'h411fc0a0} /* (7, 20, 13) {real, imag} */,
  {32'h40d0f5a6, 32'hc0f179f9} /* (7, 20, 12) {real, imag} */,
  {32'hbff49c70, 32'h418925ac} /* (7, 20, 11) {real, imag} */,
  {32'hc1737009, 32'h3fd2ad0a} /* (7, 20, 10) {real, imag} */,
  {32'h404a60c8, 32'hc160a0d4} /* (7, 20, 9) {real, imag} */,
  {32'hc0e52549, 32'hbece9b38} /* (7, 20, 8) {real, imag} */,
  {32'h407383e4, 32'hbea5c390} /* (7, 20, 7) {real, imag} */,
  {32'h40d4237e, 32'hc16b17d3} /* (7, 20, 6) {real, imag} */,
  {32'hc032bab4, 32'h402ce1da} /* (7, 20, 5) {real, imag} */,
  {32'hc1480d48, 32'hc161a35a} /* (7, 20, 4) {real, imag} */,
  {32'h3f85e688, 32'hc0f5f75c} /* (7, 20, 3) {real, imag} */,
  {32'hc04d4a68, 32'h3e7120a0} /* (7, 20, 2) {real, imag} */,
  {32'h40bbbf3f, 32'h4038c002} /* (7, 20, 1) {real, imag} */,
  {32'h3f875290, 32'h3fce2638} /* (7, 20, 0) {real, imag} */,
  {32'h403d99d8, 32'h400d5caf} /* (7, 19, 31) {real, imag} */,
  {32'hc064611e, 32'h41852dee} /* (7, 19, 30) {real, imag} */,
  {32'hbf2401dc, 32'hc1853e70} /* (7, 19, 29) {real, imag} */,
  {32'hbfc43800, 32'hc0be6f38} /* (7, 19, 28) {real, imag} */,
  {32'h408277e3, 32'hbec9f240} /* (7, 19, 27) {real, imag} */,
  {32'hbf76df52, 32'hc00752b4} /* (7, 19, 26) {real, imag} */,
  {32'h40c38365, 32'hc0a18244} /* (7, 19, 25) {real, imag} */,
  {32'h3f294f20, 32'h41250654} /* (7, 19, 24) {real, imag} */,
  {32'hc0a8f11e, 32'hc128b7c8} /* (7, 19, 23) {real, imag} */,
  {32'hc1879be7, 32'hc072b803} /* (7, 19, 22) {real, imag} */,
  {32'h40874c6a, 32'hc17d1442} /* (7, 19, 21) {real, imag} */,
  {32'h4104509c, 32'hc196d098} /* (7, 19, 20) {real, imag} */,
  {32'h4146b91e, 32'h404ec295} /* (7, 19, 19) {real, imag} */,
  {32'hc17b6811, 32'hc0704fe4} /* (7, 19, 18) {real, imag} */,
  {32'h4109f7f2, 32'hc0b8d96e} /* (7, 19, 17) {real, imag} */,
  {32'h409a3d28, 32'h412e913f} /* (7, 19, 16) {real, imag} */,
  {32'h3fc7e5c8, 32'h40bcbe55} /* (7, 19, 15) {real, imag} */,
  {32'hc1a1e2a2, 32'h40faaa42} /* (7, 19, 14) {real, imag} */,
  {32'h419c4835, 32'hc1421c1e} /* (7, 19, 13) {real, imag} */,
  {32'hc15d9231, 32'h41234ee2} /* (7, 19, 12) {real, imag} */,
  {32'hc17f6fb7, 32'h3fd72648} /* (7, 19, 11) {real, imag} */,
  {32'hc0381c86, 32'h4020c01a} /* (7, 19, 10) {real, imag} */,
  {32'hc10b3242, 32'h3ea56240} /* (7, 19, 9) {real, imag} */,
  {32'hc107782a, 32'h41238236} /* (7, 19, 8) {real, imag} */,
  {32'h4158c5ef, 32'hbf8015f7} /* (7, 19, 7) {real, imag} */,
  {32'h413c0425, 32'h40dbd481} /* (7, 19, 6) {real, imag} */,
  {32'hbfd6da74, 32'h40e3a6a2} /* (7, 19, 5) {real, imag} */,
  {32'h3fd7359c, 32'hbfbb7c36} /* (7, 19, 4) {real, imag} */,
  {32'h409206f4, 32'hc15b394b} /* (7, 19, 3) {real, imag} */,
  {32'hc1397424, 32'hc0b7d039} /* (7, 19, 2) {real, imag} */,
  {32'h407bd264, 32'hc185c4a3} /* (7, 19, 1) {real, imag} */,
  {32'hc1fb397e, 32'hc111f938} /* (7, 19, 0) {real, imag} */,
  {32'h407510c3, 32'h410e3876} /* (7, 18, 31) {real, imag} */,
  {32'h40150098, 32'h3f87f502} /* (7, 18, 30) {real, imag} */,
  {32'h3f5042fc, 32'h3fb1ef7a} /* (7, 18, 29) {real, imag} */,
  {32'hc01eeefe, 32'hc0f26661} /* (7, 18, 28) {real, imag} */,
  {32'hc07bcb5c, 32'hc13d04bc} /* (7, 18, 27) {real, imag} */,
  {32'h408f65eb, 32'hc0f37ed1} /* (7, 18, 26) {real, imag} */,
  {32'hc10851d1, 32'hc0061c64} /* (7, 18, 25) {real, imag} */,
  {32'h405f5f28, 32'hc0c946fb} /* (7, 18, 24) {real, imag} */,
  {32'hc14112f2, 32'hc1549f0a} /* (7, 18, 23) {real, imag} */,
  {32'h40b7e22e, 32'h4193b553} /* (7, 18, 22) {real, imag} */,
  {32'hc02172fc, 32'h40a03442} /* (7, 18, 21) {real, imag} */,
  {32'h3e969d7c, 32'hc0da4ded} /* (7, 18, 20) {real, imag} */,
  {32'hc0d4050a, 32'h4106250e} /* (7, 18, 19) {real, imag} */,
  {32'hc136d7f9, 32'hc1384937} /* (7, 18, 18) {real, imag} */,
  {32'hc0fbaca8, 32'h3f7648d2} /* (7, 18, 17) {real, imag} */,
  {32'h3ea31ee0, 32'hc11d823d} /* (7, 18, 16) {real, imag} */,
  {32'h4097e3bf, 32'h4023a8a4} /* (7, 18, 15) {real, imag} */,
  {32'hc1de5060, 32'h412c2a5a} /* (7, 18, 14) {real, imag} */,
  {32'hc0d88c8a, 32'hc0075a36} /* (7, 18, 13) {real, imag} */,
  {32'h410de5f9, 32'h400b8bb8} /* (7, 18, 12) {real, imag} */,
  {32'h3fc86b98, 32'h4175521a} /* (7, 18, 11) {real, imag} */,
  {32'hbfefa308, 32'hc0720082} /* (7, 18, 10) {real, imag} */,
  {32'hc0a93415, 32'hc0f5f9e8} /* (7, 18, 9) {real, imag} */,
  {32'h40227ffb, 32'h40e6fb3c} /* (7, 18, 8) {real, imag} */,
  {32'hbfb82fa0, 32'h4129d277} /* (7, 18, 7) {real, imag} */,
  {32'h41249dcf, 32'h40c1649d} /* (7, 18, 6) {real, imag} */,
  {32'hc0abad20, 32'hc0d75517} /* (7, 18, 5) {real, imag} */,
  {32'hbf82c188, 32'hc0a25260} /* (7, 18, 4) {real, imag} */,
  {32'h40eceec2, 32'h412331b3} /* (7, 18, 3) {real, imag} */,
  {32'h3fa1eb46, 32'hc0142837} /* (7, 18, 2) {real, imag} */,
  {32'hc05579ac, 32'h41752167} /* (7, 18, 1) {real, imag} */,
  {32'h3f644210, 32'h3fc36878} /* (7, 18, 0) {real, imag} */,
  {32'hbf9a5630, 32'hc131a1ae} /* (7, 17, 31) {real, imag} */,
  {32'hc0ab5312, 32'hc09e506d} /* (7, 17, 30) {real, imag} */,
  {32'h4076ce39, 32'hc0946c30} /* (7, 17, 29) {real, imag} */,
  {32'hc0cf6fb6, 32'hc1799252} /* (7, 17, 28) {real, imag} */,
  {32'h417ac091, 32'hc02d2930} /* (7, 17, 27) {real, imag} */,
  {32'hbdd26ea0, 32'h3fc9347b} /* (7, 17, 26) {real, imag} */,
  {32'hc1930ff1, 32'hbd546600} /* (7, 17, 25) {real, imag} */,
  {32'h410c8707, 32'h4001977c} /* (7, 17, 24) {real, imag} */,
  {32'h410c45e0, 32'h41b4d70e} /* (7, 17, 23) {real, imag} */,
  {32'h41353b57, 32'hc15a02d3} /* (7, 17, 22) {real, imag} */,
  {32'h411ff032, 32'hbe9f1310} /* (7, 17, 21) {real, imag} */,
  {32'hc18c5bda, 32'h408f4022} /* (7, 17, 20) {real, imag} */,
  {32'h40b5191c, 32'hc0618967} /* (7, 17, 19) {real, imag} */,
  {32'h40c1c9ac, 32'hbf81b52c} /* (7, 17, 18) {real, imag} */,
  {32'h40a04870, 32'hc0f3cfaa} /* (7, 17, 17) {real, imag} */,
  {32'h3fa8c5e8, 32'h4026eae5} /* (7, 17, 16) {real, imag} */,
  {32'h3f7cc4a8, 32'h400f5cdf} /* (7, 17, 15) {real, imag} */,
  {32'hbfa5383c, 32'h3fa17690} /* (7, 17, 14) {real, imag} */,
  {32'hc11ae312, 32'hc06a00f9} /* (7, 17, 13) {real, imag} */,
  {32'h40ee959c, 32'hc1259852} /* (7, 17, 12) {real, imag} */,
  {32'hc1144dde, 32'hc0cab9a1} /* (7, 17, 11) {real, imag} */,
  {32'hbf60b400, 32'hc107b6c0} /* (7, 17, 10) {real, imag} */,
  {32'hc0ccc6c1, 32'h408b6d76} /* (7, 17, 9) {real, imag} */,
  {32'hbf09c1c4, 32'h41a4c34b} /* (7, 17, 8) {real, imag} */,
  {32'hbff8e47e, 32'hc15907a0} /* (7, 17, 7) {real, imag} */,
  {32'hbfd125e9, 32'hc13d0f10} /* (7, 17, 6) {real, imag} */,
  {32'h3fb60db2, 32'hc021e23e} /* (7, 17, 5) {real, imag} */,
  {32'h409abc20, 32'h40698cd2} /* (7, 17, 4) {real, imag} */,
  {32'h3e09d3b0, 32'h415e79de} /* (7, 17, 3) {real, imag} */,
  {32'h405f0dba, 32'hc077bbee} /* (7, 17, 2) {real, imag} */,
  {32'hc16603b6, 32'hc07fe5f6} /* (7, 17, 1) {real, imag} */,
  {32'h409455e5, 32'hc08b0b16} /* (7, 17, 0) {real, imag} */,
  {32'h4074e3b7, 32'hbfdf50e8} /* (7, 16, 31) {real, imag} */,
  {32'hbf8cdcd6, 32'h401c9011} /* (7, 16, 30) {real, imag} */,
  {32'h410040b6, 32'hc08d0173} /* (7, 16, 29) {real, imag} */,
  {32'hc03f8820, 32'h40a93748} /* (7, 16, 28) {real, imag} */,
  {32'hbf62850a, 32'h407f56ba} /* (7, 16, 27) {real, imag} */,
  {32'h402216bb, 32'h3e7253e0} /* (7, 16, 26) {real, imag} */,
  {32'h412b43b8, 32'hc0f28cc2} /* (7, 16, 25) {real, imag} */,
  {32'hc130e6d7, 32'h40aef458} /* (7, 16, 24) {real, imag} */,
  {32'h409c7e90, 32'h414e4b64} /* (7, 16, 23) {real, imag} */,
  {32'h401ea4d6, 32'hbfb01c84} /* (7, 16, 22) {real, imag} */,
  {32'h3f176c64, 32'hc1a02613} /* (7, 16, 21) {real, imag} */,
  {32'hc09eb12b, 32'h3fc1250c} /* (7, 16, 20) {real, imag} */,
  {32'h41440c76, 32'hbf1261ac} /* (7, 16, 19) {real, imag} */,
  {32'hbfaceb20, 32'hbdd5fec8} /* (7, 16, 18) {real, imag} */,
  {32'h408e6c82, 32'h40a435a2} /* (7, 16, 17) {real, imag} */,
  {32'h40b7514e, 32'h00000000} /* (7, 16, 16) {real, imag} */,
  {32'h408e6c82, 32'hc0a435a2} /* (7, 16, 15) {real, imag} */,
  {32'hbfaceb20, 32'h3dd5fec8} /* (7, 16, 14) {real, imag} */,
  {32'h41440c76, 32'h3f1261ac} /* (7, 16, 13) {real, imag} */,
  {32'hc09eb12b, 32'hbfc1250c} /* (7, 16, 12) {real, imag} */,
  {32'h3f176c64, 32'h41a02613} /* (7, 16, 11) {real, imag} */,
  {32'h401ea4d6, 32'h3fb01c84} /* (7, 16, 10) {real, imag} */,
  {32'h409c7e90, 32'hc14e4b64} /* (7, 16, 9) {real, imag} */,
  {32'hc130e6d7, 32'hc0aef458} /* (7, 16, 8) {real, imag} */,
  {32'h412b43b8, 32'h40f28cc2} /* (7, 16, 7) {real, imag} */,
  {32'h402216bb, 32'hbe7253e0} /* (7, 16, 6) {real, imag} */,
  {32'hbf62850a, 32'hc07f56ba} /* (7, 16, 5) {real, imag} */,
  {32'hc03f8820, 32'hc0a93748} /* (7, 16, 4) {real, imag} */,
  {32'h410040b6, 32'h408d0173} /* (7, 16, 3) {real, imag} */,
  {32'hbf8cdcd6, 32'hc01c9011} /* (7, 16, 2) {real, imag} */,
  {32'h4074e3b7, 32'h3fdf50e8} /* (7, 16, 1) {real, imag} */,
  {32'hc0e296d6, 32'h00000000} /* (7, 16, 0) {real, imag} */,
  {32'hc16603b6, 32'h407fe5f6} /* (7, 15, 31) {real, imag} */,
  {32'h405f0dba, 32'h4077bbee} /* (7, 15, 30) {real, imag} */,
  {32'h3e09d3b0, 32'hc15e79de} /* (7, 15, 29) {real, imag} */,
  {32'h409abc20, 32'hc0698cd2} /* (7, 15, 28) {real, imag} */,
  {32'h3fb60db2, 32'h4021e23e} /* (7, 15, 27) {real, imag} */,
  {32'hbfd125e9, 32'h413d0f10} /* (7, 15, 26) {real, imag} */,
  {32'hbff8e47e, 32'h415907a0} /* (7, 15, 25) {real, imag} */,
  {32'hbf09c1c4, 32'hc1a4c34b} /* (7, 15, 24) {real, imag} */,
  {32'hc0ccc6c1, 32'hc08b6d76} /* (7, 15, 23) {real, imag} */,
  {32'hbf60b400, 32'h4107b6c0} /* (7, 15, 22) {real, imag} */,
  {32'hc1144dde, 32'h40cab9a1} /* (7, 15, 21) {real, imag} */,
  {32'h40ee959c, 32'h41259852} /* (7, 15, 20) {real, imag} */,
  {32'hc11ae312, 32'h406a00f9} /* (7, 15, 19) {real, imag} */,
  {32'hbfa5383c, 32'hbfa17690} /* (7, 15, 18) {real, imag} */,
  {32'h3f7cc4a8, 32'hc00f5cdf} /* (7, 15, 17) {real, imag} */,
  {32'h3fa8c5e8, 32'hc026eae5} /* (7, 15, 16) {real, imag} */,
  {32'h40a04870, 32'h40f3cfaa} /* (7, 15, 15) {real, imag} */,
  {32'h40c1c9ac, 32'h3f81b52c} /* (7, 15, 14) {real, imag} */,
  {32'h40b5191c, 32'h40618967} /* (7, 15, 13) {real, imag} */,
  {32'hc18c5bda, 32'hc08f4022} /* (7, 15, 12) {real, imag} */,
  {32'h411ff032, 32'h3e9f1310} /* (7, 15, 11) {real, imag} */,
  {32'h41353b57, 32'h415a02d3} /* (7, 15, 10) {real, imag} */,
  {32'h410c45e0, 32'hc1b4d70e} /* (7, 15, 9) {real, imag} */,
  {32'h410c8707, 32'hc001977c} /* (7, 15, 8) {real, imag} */,
  {32'hc1930ff1, 32'h3d546600} /* (7, 15, 7) {real, imag} */,
  {32'hbdd26ea0, 32'hbfc9347b} /* (7, 15, 6) {real, imag} */,
  {32'h417ac091, 32'h402d2930} /* (7, 15, 5) {real, imag} */,
  {32'hc0cf6fb6, 32'h41799252} /* (7, 15, 4) {real, imag} */,
  {32'h4076ce39, 32'h40946c30} /* (7, 15, 3) {real, imag} */,
  {32'hc0ab5312, 32'h409e506d} /* (7, 15, 2) {real, imag} */,
  {32'hbf9a5630, 32'h4131a1ae} /* (7, 15, 1) {real, imag} */,
  {32'h409455e5, 32'h408b0b16} /* (7, 15, 0) {real, imag} */,
  {32'hc05579ac, 32'hc1752167} /* (7, 14, 31) {real, imag} */,
  {32'h3fa1eb46, 32'h40142837} /* (7, 14, 30) {real, imag} */,
  {32'h40eceec2, 32'hc12331b3} /* (7, 14, 29) {real, imag} */,
  {32'hbf82c188, 32'h40a25260} /* (7, 14, 28) {real, imag} */,
  {32'hc0abad20, 32'h40d75517} /* (7, 14, 27) {real, imag} */,
  {32'h41249dcf, 32'hc0c1649d} /* (7, 14, 26) {real, imag} */,
  {32'hbfb82fa0, 32'hc129d277} /* (7, 14, 25) {real, imag} */,
  {32'h40227ffb, 32'hc0e6fb3c} /* (7, 14, 24) {real, imag} */,
  {32'hc0a93415, 32'h40f5f9e8} /* (7, 14, 23) {real, imag} */,
  {32'hbfefa308, 32'h40720082} /* (7, 14, 22) {real, imag} */,
  {32'h3fc86b98, 32'hc175521a} /* (7, 14, 21) {real, imag} */,
  {32'h410de5f9, 32'hc00b8bb8} /* (7, 14, 20) {real, imag} */,
  {32'hc0d88c8a, 32'h40075a36} /* (7, 14, 19) {real, imag} */,
  {32'hc1de5060, 32'hc12c2a5a} /* (7, 14, 18) {real, imag} */,
  {32'h4097e3bf, 32'hc023a8a4} /* (7, 14, 17) {real, imag} */,
  {32'h3ea31ee0, 32'h411d823d} /* (7, 14, 16) {real, imag} */,
  {32'hc0fbaca8, 32'hbf7648d2} /* (7, 14, 15) {real, imag} */,
  {32'hc136d7f9, 32'h41384937} /* (7, 14, 14) {real, imag} */,
  {32'hc0d4050a, 32'hc106250e} /* (7, 14, 13) {real, imag} */,
  {32'h3e969d7c, 32'h40da4ded} /* (7, 14, 12) {real, imag} */,
  {32'hc02172fc, 32'hc0a03442} /* (7, 14, 11) {real, imag} */,
  {32'h40b7e22e, 32'hc193b553} /* (7, 14, 10) {real, imag} */,
  {32'hc14112f2, 32'h41549f0a} /* (7, 14, 9) {real, imag} */,
  {32'h405f5f28, 32'h40c946fb} /* (7, 14, 8) {real, imag} */,
  {32'hc10851d1, 32'h40061c64} /* (7, 14, 7) {real, imag} */,
  {32'h408f65eb, 32'h40f37ed1} /* (7, 14, 6) {real, imag} */,
  {32'hc07bcb5c, 32'h413d04bc} /* (7, 14, 5) {real, imag} */,
  {32'hc01eeefe, 32'h40f26661} /* (7, 14, 4) {real, imag} */,
  {32'h3f5042fc, 32'hbfb1ef7a} /* (7, 14, 3) {real, imag} */,
  {32'h40150098, 32'hbf87f502} /* (7, 14, 2) {real, imag} */,
  {32'h407510c3, 32'hc10e3876} /* (7, 14, 1) {real, imag} */,
  {32'h3f644210, 32'hbfc36878} /* (7, 14, 0) {real, imag} */,
  {32'h407bd264, 32'h4185c4a3} /* (7, 13, 31) {real, imag} */,
  {32'hc1397424, 32'h40b7d039} /* (7, 13, 30) {real, imag} */,
  {32'h409206f4, 32'h415b394b} /* (7, 13, 29) {real, imag} */,
  {32'h3fd7359c, 32'h3fbb7c36} /* (7, 13, 28) {real, imag} */,
  {32'hbfd6da74, 32'hc0e3a6a2} /* (7, 13, 27) {real, imag} */,
  {32'h413c0425, 32'hc0dbd481} /* (7, 13, 26) {real, imag} */,
  {32'h4158c5ef, 32'h3f8015f7} /* (7, 13, 25) {real, imag} */,
  {32'hc107782a, 32'hc1238236} /* (7, 13, 24) {real, imag} */,
  {32'hc10b3242, 32'hbea56240} /* (7, 13, 23) {real, imag} */,
  {32'hc0381c86, 32'hc020c01a} /* (7, 13, 22) {real, imag} */,
  {32'hc17f6fb7, 32'hbfd72648} /* (7, 13, 21) {real, imag} */,
  {32'hc15d9231, 32'hc1234ee2} /* (7, 13, 20) {real, imag} */,
  {32'h419c4835, 32'h41421c1e} /* (7, 13, 19) {real, imag} */,
  {32'hc1a1e2a2, 32'hc0faaa42} /* (7, 13, 18) {real, imag} */,
  {32'h3fc7e5c8, 32'hc0bcbe55} /* (7, 13, 17) {real, imag} */,
  {32'h409a3d28, 32'hc12e913f} /* (7, 13, 16) {real, imag} */,
  {32'h4109f7f2, 32'h40b8d96e} /* (7, 13, 15) {real, imag} */,
  {32'hc17b6811, 32'h40704fe4} /* (7, 13, 14) {real, imag} */,
  {32'h4146b91e, 32'hc04ec295} /* (7, 13, 13) {real, imag} */,
  {32'h4104509c, 32'h4196d098} /* (7, 13, 12) {real, imag} */,
  {32'h40874c6a, 32'h417d1442} /* (7, 13, 11) {real, imag} */,
  {32'hc1879be7, 32'h4072b803} /* (7, 13, 10) {real, imag} */,
  {32'hc0a8f11e, 32'h4128b7c8} /* (7, 13, 9) {real, imag} */,
  {32'h3f294f20, 32'hc1250654} /* (7, 13, 8) {real, imag} */,
  {32'h40c38365, 32'h40a18244} /* (7, 13, 7) {real, imag} */,
  {32'hbf76df52, 32'h400752b4} /* (7, 13, 6) {real, imag} */,
  {32'h408277e3, 32'h3ec9f240} /* (7, 13, 5) {real, imag} */,
  {32'hbfc43800, 32'h40be6f38} /* (7, 13, 4) {real, imag} */,
  {32'hbf2401dc, 32'h41853e70} /* (7, 13, 3) {real, imag} */,
  {32'hc064611e, 32'hc1852dee} /* (7, 13, 2) {real, imag} */,
  {32'h403d99d8, 32'hc00d5caf} /* (7, 13, 1) {real, imag} */,
  {32'hc1fb397e, 32'h4111f938} /* (7, 13, 0) {real, imag} */,
  {32'h40bbbf3f, 32'hc038c002} /* (7, 12, 31) {real, imag} */,
  {32'hc04d4a68, 32'hbe7120a0} /* (7, 12, 30) {real, imag} */,
  {32'h3f85e688, 32'h40f5f75c} /* (7, 12, 29) {real, imag} */,
  {32'hc1480d48, 32'h4161a35a} /* (7, 12, 28) {real, imag} */,
  {32'hc032bab4, 32'hc02ce1da} /* (7, 12, 27) {real, imag} */,
  {32'h40d4237e, 32'h416b17d3} /* (7, 12, 26) {real, imag} */,
  {32'h407383e4, 32'h3ea5c390} /* (7, 12, 25) {real, imag} */,
  {32'hc0e52549, 32'h3ece9b38} /* (7, 12, 24) {real, imag} */,
  {32'h404a60c8, 32'h4160a0d4} /* (7, 12, 23) {real, imag} */,
  {32'hc1737009, 32'hbfd2ad0a} /* (7, 12, 22) {real, imag} */,
  {32'hbff49c70, 32'hc18925ac} /* (7, 12, 21) {real, imag} */,
  {32'h40d0f5a6, 32'h40f179f9} /* (7, 12, 20) {real, imag} */,
  {32'hc1182b34, 32'hc11fc0a0} /* (7, 12, 19) {real, imag} */,
  {32'hc0318f0a, 32'h3f524c74} /* (7, 12, 18) {real, imag} */,
  {32'h4144dfd9, 32'h3f752dd8} /* (7, 12, 17) {real, imag} */,
  {32'h3efbdf68, 32'hc14b2b0a} /* (7, 12, 16) {real, imag} */,
  {32'hc05e01bc, 32'h40a53c40} /* (7, 12, 15) {real, imag} */,
  {32'h40a9b576, 32'h415ad8ec} /* (7, 12, 14) {real, imag} */,
  {32'hc146d037, 32'h412f92d9} /* (7, 12, 13) {real, imag} */,
  {32'h41599a99, 32'hbf27eb98} /* (7, 12, 12) {real, imag} */,
  {32'hc0475460, 32'hc08fcab2} /* (7, 12, 11) {real, imag} */,
  {32'h414b822c, 32'h41aebbb2} /* (7, 12, 10) {real, imag} */,
  {32'hc16444bc, 32'hc01f49a0} /* (7, 12, 9) {real, imag} */,
  {32'h3dbfd940, 32'h40da5c30} /* (7, 12, 8) {real, imag} */,
  {32'h416141d8, 32'hc0e3025e} /* (7, 12, 7) {real, imag} */,
  {32'hc039d5a5, 32'h4162a084} /* (7, 12, 6) {real, imag} */,
  {32'hc1887442, 32'hc00faf84} /* (7, 12, 5) {real, imag} */,
  {32'h4190a7b4, 32'hc140f98f} /* (7, 12, 4) {real, imag} */,
  {32'hc19545bc, 32'hc0d505fb} /* (7, 12, 3) {real, imag} */,
  {32'h3f82cfe8, 32'hc069a7a4} /* (7, 12, 2) {real, imag} */,
  {32'h417bb391, 32'hbf7186dc} /* (7, 12, 1) {real, imag} */,
  {32'h3f875290, 32'hbfce2638} /* (7, 12, 0) {real, imag} */,
  {32'h3f0e2b00, 32'hc0e77718} /* (7, 11, 31) {real, imag} */,
  {32'h41b2056c, 32'h3e26c680} /* (7, 11, 30) {real, imag} */,
  {32'h411bab4c, 32'h413335a0} /* (7, 11, 29) {real, imag} */,
  {32'hc1328038, 32'hc118b778} /* (7, 11, 28) {real, imag} */,
  {32'h3fe61b48, 32'h4105c4f9} /* (7, 11, 27) {real, imag} */,
  {32'h410b401b, 32'h40d0c105} /* (7, 11, 26) {real, imag} */,
  {32'hc1b5b176, 32'hc067affe} /* (7, 11, 25) {real, imag} */,
  {32'hc0eb2e5a, 32'h4161b4fe} /* (7, 11, 24) {real, imag} */,
  {32'hc1d39410, 32'h416c07e5} /* (7, 11, 23) {real, imag} */,
  {32'hc095bd6e, 32'hc105abdd} /* (7, 11, 22) {real, imag} */,
  {32'h418962ff, 32'hc11918f2} /* (7, 11, 21) {real, imag} */,
  {32'h41c62406, 32'h3f589b24} /* (7, 11, 20) {real, imag} */,
  {32'h40c7a9da, 32'hbf1864c8} /* (7, 11, 19) {real, imag} */,
  {32'h412b4a7f, 32'h40b352f6} /* (7, 11, 18) {real, imag} */,
  {32'hc0fa9f6b, 32'hc0853ebd} /* (7, 11, 17) {real, imag} */,
  {32'h411d38f0, 32'h408d4c9e} /* (7, 11, 16) {real, imag} */,
  {32'h4121e5d8, 32'h40ccee7b} /* (7, 11, 15) {real, imag} */,
  {32'hc144b906, 32'hc15244d0} /* (7, 11, 14) {real, imag} */,
  {32'hc00808e4, 32'hbf2baec8} /* (7, 11, 13) {real, imag} */,
  {32'h3f6f6e68, 32'hc149e075} /* (7, 11, 12) {real, imag} */,
  {32'hc075e3b8, 32'h413a6fa0} /* (7, 11, 11) {real, imag} */,
  {32'hc18973e0, 32'h419d56b6} /* (7, 11, 10) {real, imag} */,
  {32'h414918f2, 32'hc19376bf} /* (7, 11, 9) {real, imag} */,
  {32'hc018252c, 32'h40902c8e} /* (7, 11, 8) {real, imag} */,
  {32'h411dbd94, 32'h409d6376} /* (7, 11, 7) {real, imag} */,
  {32'h411bc99a, 32'h41a789de} /* (7, 11, 6) {real, imag} */,
  {32'hc03f3f74, 32'h4109e67c} /* (7, 11, 5) {real, imag} */,
  {32'h40cc5f40, 32'hc1b2c1ce} /* (7, 11, 4) {real, imag} */,
  {32'h416543e2, 32'hc1b77cc1} /* (7, 11, 3) {real, imag} */,
  {32'hc0969c6f, 32'h41832e61} /* (7, 11, 2) {real, imag} */,
  {32'h3fcdb350, 32'hc1d17db1} /* (7, 11, 1) {real, imag} */,
  {32'hc122e90c, 32'hc12458d1} /* (7, 11, 0) {real, imag} */,
  {32'hbeb2af60, 32'h40d42cf5} /* (7, 10, 31) {real, imag} */,
  {32'hc14630ac, 32'h40bd22a0} /* (7, 10, 30) {real, imag} */,
  {32'hc13719f2, 32'hc140d69b} /* (7, 10, 29) {real, imag} */,
  {32'h3f310efc, 32'h4185fc28} /* (7, 10, 28) {real, imag} */,
  {32'h410a3e92, 32'hc15a078d} /* (7, 10, 27) {real, imag} */,
  {32'h41168c53, 32'hc09623a9} /* (7, 10, 26) {real, imag} */,
  {32'h406a54c2, 32'hc17fd1dc} /* (7, 10, 25) {real, imag} */,
  {32'hc159c1e3, 32'h4081fc71} /* (7, 10, 24) {real, imag} */,
  {32'h40d1ca1c, 32'hc0ea8bae} /* (7, 10, 23) {real, imag} */,
  {32'hc1956590, 32'hc104fa9e} /* (7, 10, 22) {real, imag} */,
  {32'h41d6fd4b, 32'hbf1a2da0} /* (7, 10, 21) {real, imag} */,
  {32'h41c8129a, 32'h3f6d4e20} /* (7, 10, 20) {real, imag} */,
  {32'h40f647c9, 32'h418f47b8} /* (7, 10, 19) {real, imag} */,
  {32'hc065f34c, 32'h3eebb9f0} /* (7, 10, 18) {real, imag} */,
  {32'hc1094e9a, 32'hc0d07b9e} /* (7, 10, 17) {real, imag} */,
  {32'hbe7c1ca0, 32'hc0d8a611} /* (7, 10, 16) {real, imag} */,
  {32'hbfc43ac6, 32'hc0a5e844} /* (7, 10, 15) {real, imag} */,
  {32'hc14d89c3, 32'hc1421b37} /* (7, 10, 14) {real, imag} */,
  {32'h4171a90e, 32'hc0f572c3} /* (7, 10, 13) {real, imag} */,
  {32'h41132994, 32'h418c2d91} /* (7, 10, 12) {real, imag} */,
  {32'h40f8ab78, 32'hc1a9c9e2} /* (7, 10, 11) {real, imag} */,
  {32'hc14b8a6c, 32'h406a8332} /* (7, 10, 10) {real, imag} */,
  {32'h40d9d1c7, 32'h40be809b} /* (7, 10, 9) {real, imag} */,
  {32'hc080ef45, 32'hc05d1a5a} /* (7, 10, 8) {real, imag} */,
  {32'hc0c4900e, 32'hc152e7ee} /* (7, 10, 7) {real, imag} */,
  {32'hc1251743, 32'h41468402} /* (7, 10, 6) {real, imag} */,
  {32'h41a3294a, 32'hc0add336} /* (7, 10, 5) {real, imag} */,
  {32'hbfe87f66, 32'hbfccdc9c} /* (7, 10, 4) {real, imag} */,
  {32'hc0bbae5b, 32'h41a5982e} /* (7, 10, 3) {real, imag} */,
  {32'h3f82fdbc, 32'hc13cd440} /* (7, 10, 2) {real, imag} */,
  {32'h418882a9, 32'hc095d1f6} /* (7, 10, 1) {real, imag} */,
  {32'hc06b884c, 32'h41d2b5c6} /* (7, 10, 0) {real, imag} */,
  {32'hc147f4f4, 32'h41c8ff99} /* (7, 9, 31) {real, imag} */,
  {32'h415f4c0a, 32'hc1b3a7da} /* (7, 9, 30) {real, imag} */,
  {32'hbf34d3a8, 32'hbf070108} /* (7, 9, 29) {real, imag} */,
  {32'hbf818f2a, 32'h3ebbfb90} /* (7, 9, 28) {real, imag} */,
  {32'hc168ea77, 32'h40f0daf6} /* (7, 9, 27) {real, imag} */,
  {32'h3fe78818, 32'hc0b594ca} /* (7, 9, 26) {real, imag} */,
  {32'hc18c599b, 32'hc0acb604} /* (7, 9, 25) {real, imag} */,
  {32'h40ba57d0, 32'hc1576f5c} /* (7, 9, 24) {real, imag} */,
  {32'hc18d934e, 32'hc188890a} /* (7, 9, 23) {real, imag} */,
  {32'h41a93f92, 32'hc0ae5ddf} /* (7, 9, 22) {real, imag} */,
  {32'hbf43aa10, 32'hc115329b} /* (7, 9, 21) {real, imag} */,
  {32'h40118b70, 32'hc056a280} /* (7, 9, 20) {real, imag} */,
  {32'h416d8db2, 32'h4137a2ad} /* (7, 9, 19) {real, imag} */,
  {32'hc176a155, 32'hc0ae0d62} /* (7, 9, 18) {real, imag} */,
  {32'h407ef25a, 32'h40f2c3b0} /* (7, 9, 17) {real, imag} */,
  {32'h4059950a, 32'h410b14f2} /* (7, 9, 16) {real, imag} */,
  {32'h40840bd2, 32'hc1291a2e} /* (7, 9, 15) {real, imag} */,
  {32'h4101c450, 32'h401c057d} /* (7, 9, 14) {real, imag} */,
  {32'hc003aa64, 32'hc1594fea} /* (7, 9, 13) {real, imag} */,
  {32'h4038f8d8, 32'h40a62cc7} /* (7, 9, 12) {real, imag} */,
  {32'h410f7d66, 32'h3f848a34} /* (7, 9, 11) {real, imag} */,
  {32'h40f1f827, 32'hc0d0a882} /* (7, 9, 10) {real, imag} */,
  {32'hc125075c, 32'h41add430} /* (7, 9, 9) {real, imag} */,
  {32'hc07344c6, 32'hc0357eaa} /* (7, 9, 8) {real, imag} */,
  {32'h3f81b375, 32'h41809196} /* (7, 9, 7) {real, imag} */,
  {32'hc1634717, 32'hc0f38c0e} /* (7, 9, 6) {real, imag} */,
  {32'hc09c122e, 32'h413099cb} /* (7, 9, 5) {real, imag} */,
  {32'h4103b555, 32'h40fd0e40} /* (7, 9, 4) {real, imag} */,
  {32'hc010ddc5, 32'h412a54ab} /* (7, 9, 3) {real, imag} */,
  {32'hc17c6eb4, 32'hc090460c} /* (7, 9, 2) {real, imag} */,
  {32'hc1a3e8b2, 32'h3fb53f94} /* (7, 9, 1) {real, imag} */,
  {32'hc10cab70, 32'hc0aa75bb} /* (7, 9, 0) {real, imag} */,
  {32'hc2445dc3, 32'hc1b0f6f4} /* (7, 8, 31) {real, imag} */,
  {32'h41e7772d, 32'h418daf33} /* (7, 8, 30) {real, imag} */,
  {32'h4102b91c, 32'hc10acfe4} /* (7, 8, 29) {real, imag} */,
  {32'h41569b50, 32'h4077efea} /* (7, 8, 28) {real, imag} */,
  {32'h41fb1944, 32'hc159517a} /* (7, 8, 27) {real, imag} */,
  {32'h412100f8, 32'hc143c935} /* (7, 8, 26) {real, imag} */,
  {32'hc10ed724, 32'hc15bc6aa} /* (7, 8, 25) {real, imag} */,
  {32'h415a3f11, 32'hc1b40aad} /* (7, 8, 24) {real, imag} */,
  {32'h41000960, 32'hc1733d78} /* (7, 8, 23) {real, imag} */,
  {32'h3f97da88, 32'h3f596878} /* (7, 8, 22) {real, imag} */,
  {32'hc0b3c6bd, 32'h415468ce} /* (7, 8, 21) {real, imag} */,
  {32'hc0d0db5c, 32'h418be5fb} /* (7, 8, 20) {real, imag} */,
  {32'hc081fc1c, 32'h3f9fc260} /* (7, 8, 19) {real, imag} */,
  {32'h412e1656, 32'h4111e712} /* (7, 8, 18) {real, imag} */,
  {32'hc185b17a, 32'h4111e174} /* (7, 8, 17) {real, imag} */,
  {32'hc10cce62, 32'h408cbf28} /* (7, 8, 16) {real, imag} */,
  {32'h408c8756, 32'hc12fee88} /* (7, 8, 15) {real, imag} */,
  {32'h41abd7d9, 32'hc11d457a} /* (7, 8, 14) {real, imag} */,
  {32'hc1a678ba, 32'h40ab537b} /* (7, 8, 13) {real, imag} */,
  {32'hc013d438, 32'hc080b5a3} /* (7, 8, 12) {real, imag} */,
  {32'h406c51f4, 32'h419448a2} /* (7, 8, 11) {real, imag} */,
  {32'h40f224d9, 32'hc0b27aeb} /* (7, 8, 10) {real, imag} */,
  {32'hc17c6ebc, 32'hc13580c1} /* (7, 8, 9) {real, imag} */,
  {32'hc082bea0, 32'h41ed49e8} /* (7, 8, 8) {real, imag} */,
  {32'hc1562194, 32'h40c2a799} /* (7, 8, 7) {real, imag} */,
  {32'hc1839bc4, 32'h3faab288} /* (7, 8, 6) {real, imag} */,
  {32'hc18a9c0a, 32'h4041f356} /* (7, 8, 5) {real, imag} */,
  {32'hc1751275, 32'hc18353c9} /* (7, 8, 4) {real, imag} */,
  {32'h40a71798, 32'h40f9c8ad} /* (7, 8, 3) {real, imag} */,
  {32'h41abc60a, 32'h409a63d8} /* (7, 8, 2) {real, imag} */,
  {32'hc185bea2, 32'hc208ba72} /* (7, 8, 1) {real, imag} */,
  {32'hc1d59ae1, 32'hc19d5430} /* (7, 8, 0) {real, imag} */,
  {32'hc08097ac, 32'hc103c292} /* (7, 7, 31) {real, imag} */,
  {32'h410b396a, 32'hc08d12c4} /* (7, 7, 30) {real, imag} */,
  {32'hc1c1cbe2, 32'h4082e6f2} /* (7, 7, 29) {real, imag} */,
  {32'hc0177096, 32'h40af4bf6} /* (7, 7, 28) {real, imag} */,
  {32'h410b9255, 32'hc0a89574} /* (7, 7, 27) {real, imag} */,
  {32'hbfec870c, 32'h4171a2a0} /* (7, 7, 26) {real, imag} */,
  {32'hc1187117, 32'h41c7916c} /* (7, 7, 25) {real, imag} */,
  {32'h41194be8, 32'hc1094afa} /* (7, 7, 24) {real, imag} */,
  {32'hc10e9fde, 32'hc0be0516} /* (7, 7, 23) {real, imag} */,
  {32'hc0d01160, 32'h402fb3ab} /* (7, 7, 22) {real, imag} */,
  {32'h4070ce72, 32'hc137e75b} /* (7, 7, 21) {real, imag} */,
  {32'hbfa041be, 32'h40817d28} /* (7, 7, 20) {real, imag} */,
  {32'hbfabb8d8, 32'h40e7849d} /* (7, 7, 19) {real, imag} */,
  {32'h406eb45a, 32'hc01364be} /* (7, 7, 18) {real, imag} */,
  {32'hc0f390a4, 32'h401b40ee} /* (7, 7, 17) {real, imag} */,
  {32'hc0b4ef65, 32'hc0837ec5} /* (7, 7, 16) {real, imag} */,
  {32'hbe8aacd8, 32'hc0a205ee} /* (7, 7, 15) {real, imag} */,
  {32'h405ed06a, 32'hc0f7b616} /* (7, 7, 14) {real, imag} */,
  {32'h4092eede, 32'h41551574} /* (7, 7, 13) {real, imag} */,
  {32'hc0e66e14, 32'hc18a44c0} /* (7, 7, 12) {real, imag} */,
  {32'hc1581164, 32'h3f211a40} /* (7, 7, 11) {real, imag} */,
  {32'h41bbe576, 32'h4156a8b7} /* (7, 7, 10) {real, imag} */,
  {32'h415bee02, 32'h41c8148e} /* (7, 7, 9) {real, imag} */,
  {32'hc187e855, 32'hc121c52c} /* (7, 7, 8) {real, imag} */,
  {32'hc103307d, 32'hc1af7cd4} /* (7, 7, 7) {real, imag} */,
  {32'h41a76907, 32'h407b301c} /* (7, 7, 6) {real, imag} */,
  {32'h4216df1b, 32'hc10c6c8e} /* (7, 7, 5) {real, imag} */,
  {32'h40aeee4c, 32'h41c2c4ed} /* (7, 7, 4) {real, imag} */,
  {32'hc158e1a7, 32'h41cae47e} /* (7, 7, 3) {real, imag} */,
  {32'hc097c106, 32'hc2117784} /* (7, 7, 2) {real, imag} */,
  {32'hc0dd6c84, 32'h419536a7} /* (7, 7, 1) {real, imag} */,
  {32'h415c6cf6, 32'h41080cec} /* (7, 7, 0) {real, imag} */,
  {32'h40d33625, 32'h418933b2} /* (7, 6, 31) {real, imag} */,
  {32'hc058836c, 32'hc14c5e3d} /* (7, 6, 30) {real, imag} */,
  {32'hc09780cf, 32'hc166be86} /* (7, 6, 29) {real, imag} */,
  {32'hc0fac502, 32'h415cfbeb} /* (7, 6, 28) {real, imag} */,
  {32'h4195b2eb, 32'h418ca3a8} /* (7, 6, 27) {real, imag} */,
  {32'hc0501ac8, 32'hbe0b0f80} /* (7, 6, 26) {real, imag} */,
  {32'h4176317a, 32'h3f182130} /* (7, 6, 25) {real, imag} */,
  {32'h3fee5368, 32'hc11bad3f} /* (7, 6, 24) {real, imag} */,
  {32'h419449ef, 32'hc0c64a8b} /* (7, 6, 23) {real, imag} */,
  {32'hc0920264, 32'h4068ad34} /* (7, 6, 22) {real, imag} */,
  {32'hc0d2eb6b, 32'hc096b662} /* (7, 6, 21) {real, imag} */,
  {32'h3fa0ae34, 32'hc0c22b18} /* (7, 6, 20) {real, imag} */,
  {32'hc0b06ddb, 32'h4119f858} /* (7, 6, 19) {real, imag} */,
  {32'hc0b8ec60, 32'h40402754} /* (7, 6, 18) {real, imag} */,
  {32'hc023ccdf, 32'h409dfd7f} /* (7, 6, 17) {real, imag} */,
  {32'hc13cde08, 32'hc0c460b1} /* (7, 6, 16) {real, imag} */,
  {32'hc0a7d23e, 32'hbe9f0050} /* (7, 6, 15) {real, imag} */,
  {32'hc1035005, 32'h4120de34} /* (7, 6, 14) {real, imag} */,
  {32'h40a3694b, 32'hc0d5c90a} /* (7, 6, 13) {real, imag} */,
  {32'hc0ffb441, 32'h416b2218} /* (7, 6, 12) {real, imag} */,
  {32'h4123c58f, 32'hc11b1729} /* (7, 6, 11) {real, imag} */,
  {32'h40255ca0, 32'hc1280a7c} /* (7, 6, 10) {real, imag} */,
  {32'hc154eb66, 32'hc09182ce} /* (7, 6, 9) {real, imag} */,
  {32'h415e53c4, 32'hc0909405} /* (7, 6, 8) {real, imag} */,
  {32'h41e93bd0, 32'h41661d14} /* (7, 6, 7) {real, imag} */,
  {32'hc0bccbb8, 32'hc0094240} /* (7, 6, 6) {real, imag} */,
  {32'hc02ecab3, 32'h40308da5} /* (7, 6, 5) {real, imag} */,
  {32'h4019aa8d, 32'h3fb934b0} /* (7, 6, 4) {real, imag} */,
  {32'hc12f9bba, 32'h41d075a5} /* (7, 6, 3) {real, imag} */,
  {32'hc1d113e2, 32'hc0ec2cf0} /* (7, 6, 2) {real, imag} */,
  {32'hc193b9d5, 32'h40e9946b} /* (7, 6, 1) {real, imag} */,
  {32'hbff5e64c, 32'hc13b646a} /* (7, 6, 0) {real, imag} */,
  {32'hc2a473b8, 32'h406037e4} /* (7, 5, 31) {real, imag} */,
  {32'h424eb1ae, 32'hc20b7256} /* (7, 5, 30) {real, imag} */,
  {32'hc07ba380, 32'hc0b0f9c2} /* (7, 5, 29) {real, imag} */,
  {32'hc1422102, 32'h407d4d28} /* (7, 5, 28) {real, imag} */,
  {32'h4136d98f, 32'hc12258a2} /* (7, 5, 27) {real, imag} */,
  {32'hc10ab28a, 32'h408fe854} /* (7, 5, 26) {real, imag} */,
  {32'hc16a7a8e, 32'h40c30939} /* (7, 5, 25) {real, imag} */,
  {32'h3de16da0, 32'hc1434b04} /* (7, 5, 24) {real, imag} */,
  {32'hc0d3c55e, 32'hc10d5f4a} /* (7, 5, 23) {real, imag} */,
  {32'h40d3d02f, 32'h40371ad8} /* (7, 5, 22) {real, imag} */,
  {32'h411e0cba, 32'h40e1ff8f} /* (7, 5, 21) {real, imag} */,
  {32'hc0691f84, 32'hc08f2456} /* (7, 5, 20) {real, imag} */,
  {32'h410f3b08, 32'hbfce455a} /* (7, 5, 19) {real, imag} */,
  {32'hc0e3b8c2, 32'hc164fb40} /* (7, 5, 18) {real, imag} */,
  {32'h40710008, 32'hbda36d90} /* (7, 5, 17) {real, imag} */,
  {32'h40932f00, 32'hc1258512} /* (7, 5, 16) {real, imag} */,
  {32'hc0ea741d, 32'hc0718934} /* (7, 5, 15) {real, imag} */,
  {32'hc1945932, 32'h408eedc1} /* (7, 5, 14) {real, imag} */,
  {32'hbfbeb399, 32'hc11f3793} /* (7, 5, 13) {real, imag} */,
  {32'h401296a0, 32'hc1317fe6} /* (7, 5, 12) {real, imag} */,
  {32'hc18e6e03, 32'hc0edddd6} /* (7, 5, 11) {real, imag} */,
  {32'h40bd048e, 32'hc1679b66} /* (7, 5, 10) {real, imag} */,
  {32'h40d1ea63, 32'h3f1bcab8} /* (7, 5, 9) {real, imag} */,
  {32'h40935f5c, 32'hc12b7649} /* (7, 5, 8) {real, imag} */,
  {32'hc126cc80, 32'h40ade43c} /* (7, 5, 7) {real, imag} */,
  {32'h41a07657, 32'h4182c462} /* (7, 5, 6) {real, imag} */,
  {32'h41b4209c, 32'h41271331} /* (7, 5, 5) {real, imag} */,
  {32'h3f38c840, 32'h403d9c08} /* (7, 5, 4) {real, imag} */,
  {32'hc02ea4b0, 32'h3e57ca00} /* (7, 5, 3) {real, imag} */,
  {32'h422bcdc6, 32'h4215d816} /* (7, 5, 2) {real, imag} */,
  {32'hc2245525, 32'hc1c6695a} /* (7, 5, 1) {real, imag} */,
  {32'hc291524c, 32'hc1d14b9c} /* (7, 5, 0) {real, imag} */,
  {32'h41175e9a, 32'h42acb87c} /* (7, 4, 31) {real, imag} */,
  {32'hc2a85c1c, 32'hc286f907} /* (7, 4, 30) {real, imag} */,
  {32'h41157314, 32'hc186ddf6} /* (7, 4, 29) {real, imag} */,
  {32'h4213734a, 32'h40eb6c8a} /* (7, 4, 28) {real, imag} */,
  {32'hc0eb7eb1, 32'hc05c04f6} /* (7, 4, 27) {real, imag} */,
  {32'hc149cb68, 32'hc04fe96c} /* (7, 4, 26) {real, imag} */,
  {32'h40a68ac1, 32'h40440a28} /* (7, 4, 25) {real, imag} */,
  {32'hbfefeb08, 32'hc19b9cba} /* (7, 4, 24) {real, imag} */,
  {32'hc120e940, 32'hc124124b} /* (7, 4, 23) {real, imag} */,
  {32'h415b850a, 32'hc0807bca} /* (7, 4, 22) {real, imag} */,
  {32'h402bc3fe, 32'hc1a60e9b} /* (7, 4, 21) {real, imag} */,
  {32'hc09e878a, 32'h41a416ee} /* (7, 4, 20) {real, imag} */,
  {32'hc0064640, 32'h4158e026} /* (7, 4, 19) {real, imag} */,
  {32'hc10b6e3d, 32'hc0d4d238} /* (7, 4, 18) {real, imag} */,
  {32'h413ee65c, 32'h3e6689e0} /* (7, 4, 17) {real, imag} */,
  {32'h3eb2f91e, 32'h40ce1870} /* (7, 4, 16) {real, imag} */,
  {32'hc1500cd0, 32'h40ced7ab} /* (7, 4, 15) {real, imag} */,
  {32'hc175f890, 32'hc0c1ae46} /* (7, 4, 14) {real, imag} */,
  {32'h41676cc0, 32'h406738e8} /* (7, 4, 13) {real, imag} */,
  {32'hc0ec5af8, 32'h40c475a4} /* (7, 4, 12) {real, imag} */,
  {32'h40f46279, 32'hc17abb78} /* (7, 4, 11) {real, imag} */,
  {32'h4067b9ff, 32'hbfa83df4} /* (7, 4, 10) {real, imag} */,
  {32'h41688ac6, 32'hc1a9b961} /* (7, 4, 9) {real, imag} */,
  {32'hc0e6e362, 32'hc1968b22} /* (7, 4, 8) {real, imag} */,
  {32'hbfffc7d0, 32'h3f0f5dc0} /* (7, 4, 7) {real, imag} */,
  {32'h41030cb3, 32'h412c2d98} /* (7, 4, 6) {real, imag} */,
  {32'hbf5edd60, 32'hc211f9ac} /* (7, 4, 5) {real, imag} */,
  {32'h40ebe8f6, 32'h422712dd} /* (7, 4, 4) {real, imag} */,
  {32'hc185c3a1, 32'hbfaf91d4} /* (7, 4, 3) {real, imag} */,
  {32'hc2990dcb, 32'hc2ab1fba} /* (7, 4, 2) {real, imag} */,
  {32'h42f063b8, 32'h42c57a32} /* (7, 4, 1) {real, imag} */,
  {32'h426cdcee, 32'h4068c630} /* (7, 4, 0) {real, imag} */,
  {32'hc30efc8b, 32'h425d5adc} /* (7, 3, 31) {real, imag} */,
  {32'h4270769c, 32'hc2eccdb2} /* (7, 3, 30) {real, imag} */,
  {32'hc16905a8, 32'hbf88cbd0} /* (7, 3, 29) {real, imag} */,
  {32'h42271c10, 32'h41caaf40} /* (7, 3, 28) {real, imag} */,
  {32'hc058e7a2, 32'h410c36d4} /* (7, 3, 27) {real, imag} */,
  {32'hc1b852fa, 32'hc0355df0} /* (7, 3, 26) {real, imag} */,
  {32'hc1c0829c, 32'h4198d497} /* (7, 3, 25) {real, imag} */,
  {32'hc1b7a790, 32'hc1b37252} /* (7, 3, 24) {real, imag} */,
  {32'h3fd60968, 32'h3dcc3340} /* (7, 3, 23) {real, imag} */,
  {32'h3ead01e8, 32'h405a4ed5} /* (7, 3, 22) {real, imag} */,
  {32'h4053417b, 32'hc18785b6} /* (7, 3, 21) {real, imag} */,
  {32'hc12c9c55, 32'hc07810d4} /* (7, 3, 20) {real, imag} */,
  {32'h418b3650, 32'h40be71e4} /* (7, 3, 19) {real, imag} */,
  {32'h3ebaf8d0, 32'hc0ff8842} /* (7, 3, 18) {real, imag} */,
  {32'hc02ce640, 32'h3e52f7e0} /* (7, 3, 17) {real, imag} */,
  {32'h3f9c0f3c, 32'hc1320dcc} /* (7, 3, 16) {real, imag} */,
  {32'h404c3cc8, 32'h408c597a} /* (7, 3, 15) {real, imag} */,
  {32'h41704e0a, 32'h411f7362} /* (7, 3, 14) {real, imag} */,
  {32'hc0c4cb0a, 32'hc05c5322} /* (7, 3, 13) {real, imag} */,
  {32'h3f5df110, 32'hc1698afb} /* (7, 3, 12) {real, imag} */,
  {32'hc0c37236, 32'hc1a4e890} /* (7, 3, 11) {real, imag} */,
  {32'hbfb8eaf2, 32'hbfd20ec0} /* (7, 3, 10) {real, imag} */,
  {32'h40d684a1, 32'h416f3847} /* (7, 3, 9) {real, imag} */,
  {32'hc09f597f, 32'h412916c2} /* (7, 3, 8) {real, imag} */,
  {32'hc064a047, 32'h409ebce2} /* (7, 3, 7) {real, imag} */,
  {32'h4024ca54, 32'hc12e0949} /* (7, 3, 6) {real, imag} */,
  {32'h41fde1fa, 32'hc09b275c} /* (7, 3, 5) {real, imag} */,
  {32'hc243bbb3, 32'h41b62de3} /* (7, 3, 4) {real, imag} */,
  {32'hc0a802b7, 32'hc10ff03a} /* (7, 3, 3) {real, imag} */,
  {32'hc1a9105c, 32'hc261f7be} /* (7, 3, 2) {real, imag} */,
  {32'h43043c7c, 32'h43057b78} /* (7, 3, 1) {real, imag} */,
  {32'h41b2150d, 32'h4107d89d} /* (7, 3, 0) {real, imag} */,
  {32'hc47c0336, 32'h4188d424} /* (7, 2, 31) {real, imag} */,
  {32'h43f44116, 32'hc3049647} /* (7, 2, 30) {real, imag} */,
  {32'hc241ec25, 32'h4249bce9} /* (7, 2, 29) {real, imag} */,
  {32'hc0bc7818, 32'h42250f79} /* (7, 2, 28) {real, imag} */,
  {32'h4235edfc, 32'hc2169f3e} /* (7, 2, 27) {real, imag} */,
  {32'h4197941f, 32'hc13919e7} /* (7, 2, 26) {real, imag} */,
  {32'hc19e8dac, 32'h406e44a0} /* (7, 2, 25) {real, imag} */,
  {32'h41fd0b22, 32'h410b4666} /* (7, 2, 24) {real, imag} */,
  {32'h40e886ca, 32'hc0a44ae9} /* (7, 2, 23) {real, imag} */,
  {32'h41ad37ac, 32'h41b12e16} /* (7, 2, 22) {real, imag} */,
  {32'h41867f99, 32'hc08ce1fb} /* (7, 2, 21) {real, imag} */,
  {32'h41813f15, 32'hc18553c3} /* (7, 2, 20) {real, imag} */,
  {32'hc097bc02, 32'h3f0d77c0} /* (7, 2, 19) {real, imag} */,
  {32'h4025f04c, 32'hc0fa5f60} /* (7, 2, 18) {real, imag} */,
  {32'hbda00920, 32'h3fb42c24} /* (7, 2, 17) {real, imag} */,
  {32'hc05779f8, 32'h4074dd6a} /* (7, 2, 16) {real, imag} */,
  {32'h412490e8, 32'h40d22017} /* (7, 2, 15) {real, imag} */,
  {32'h410ca669, 32'hc1102aaf} /* (7, 2, 14) {real, imag} */,
  {32'hc18bbdb3, 32'hbf494fd0} /* (7, 2, 13) {real, imag} */,
  {32'hc1846e42, 32'h412be0dc} /* (7, 2, 12) {real, imag} */,
  {32'h417320d2, 32'h41473896} /* (7, 2, 11) {real, imag} */,
  {32'h411e3bfc, 32'h3e92d3a0} /* (7, 2, 10) {real, imag} */,
  {32'h40fdfff3, 32'h41ad5409} /* (7, 2, 9) {real, imag} */,
  {32'hc04a8438, 32'h40e6ec32} /* (7, 2, 8) {real, imag} */,
  {32'hc0d46ab6, 32'hc1abb5e4} /* (7, 2, 7) {real, imag} */,
  {32'h4114d677, 32'h3f9d75c8} /* (7, 2, 6) {real, imag} */,
  {32'h425a86e0, 32'h4210dd2d} /* (7, 2, 5) {real, imag} */,
  {32'hc2ed82c2, 32'hc1a45c96} /* (7, 2, 4) {real, imag} */,
  {32'hc1e510e5, 32'h4206f27a} /* (7, 2, 3) {real, imag} */,
  {32'h43bfb028, 32'hc252eee3} /* (7, 2, 2) {real, imag} */,
  {32'hc401a06e, 32'h42c00cee} /* (7, 2, 1) {real, imag} */,
  {32'hc4020d36, 32'hc335fa66} /* (7, 2, 0) {real, imag} */,
  {32'h44a4cfda, 32'hc3a909f4} /* (7, 1, 31) {real, imag} */,
  {32'hc389f35d, 32'h42181785} /* (7, 1, 30) {real, imag} */,
  {32'h423125cc, 32'hc21fd7f0} /* (7, 1, 29) {real, imag} */,
  {32'h4252bdee, 32'h428425f4} /* (7, 1, 28) {real, imag} */,
  {32'hc2bcfb34, 32'h3f4d7808} /* (7, 1, 27) {real, imag} */,
  {32'hc198a781, 32'h41e6c1b7} /* (7, 1, 26) {real, imag} */,
  {32'h41141749, 32'hc0514667} /* (7, 1, 25) {real, imag} */,
  {32'hc1c5bb0f, 32'h41c386b2} /* (7, 1, 24) {real, imag} */,
  {32'h40a3d984, 32'h40f70729} /* (7, 1, 23) {real, imag} */,
  {32'h419bf955, 32'hc090a892} /* (7, 1, 22) {real, imag} */,
  {32'hc117b321, 32'h41f4c342} /* (7, 1, 21) {real, imag} */,
  {32'h3f143e00, 32'h408934b4} /* (7, 1, 20) {real, imag} */,
  {32'h4025fd46, 32'h41039e28} /* (7, 1, 19) {real, imag} */,
  {32'h3f8eb8f4, 32'h41a94be0} /* (7, 1, 18) {real, imag} */,
  {32'hc0ec9447, 32'h3eab8dd8} /* (7, 1, 17) {real, imag} */,
  {32'hbef30e68, 32'hc1894ed0} /* (7, 1, 16) {real, imag} */,
  {32'hc058398b, 32'h40f0c7a2} /* (7, 1, 15) {real, imag} */,
  {32'hc11d4807, 32'h404d7a80} /* (7, 1, 14) {real, imag} */,
  {32'hc13eed78, 32'hc12c31bb} /* (7, 1, 13) {real, imag} */,
  {32'h3f9a5122, 32'hc11f9a44} /* (7, 1, 12) {real, imag} */,
  {32'hc18baf35, 32'hc173dd65} /* (7, 1, 11) {real, imag} */,
  {32'hc0a31a3c, 32'h412874cf} /* (7, 1, 10) {real, imag} */,
  {32'hc10ef8eb, 32'h3ffe84c2} /* (7, 1, 9) {real, imag} */,
  {32'hc165b8e3, 32'hc22474f4} /* (7, 1, 8) {real, imag} */,
  {32'h41846d3d, 32'h41aafaa4} /* (7, 1, 7) {real, imag} */,
  {32'hc1a184f3, 32'hbfee1918} /* (7, 1, 6) {real, imag} */,
  {32'hc2947832, 32'hc2051748} /* (7, 1, 5) {real, imag} */,
  {32'h4245eefc, 32'hc1582628} /* (7, 1, 4) {real, imag} */,
  {32'hc233fe73, 32'hc2bea9b8} /* (7, 1, 3) {real, imag} */,
  {32'hc3e86dfe, 32'hc3e6db87} /* (7, 1, 2) {real, imag} */,
  {32'h44e46005, 32'h445ac369} /* (7, 1, 1) {real, imag} */,
  {32'h44deaf4e, 32'h43699daf} /* (7, 1, 0) {real, imag} */,
  {32'h44846afa, 32'hc45b6a80} /* (7, 0, 31) {real, imag} */,
  {32'hc2ceac6a, 32'h438336f2} /* (7, 0, 30) {real, imag} */,
  {32'hc08e4fcc, 32'hc1b3fe6b} /* (7, 0, 29) {real, imag} */,
  {32'h41635448, 32'h407d0fa0} /* (7, 0, 28) {real, imag} */,
  {32'hc27f0831, 32'h41d16c1a} /* (7, 0, 27) {real, imag} */,
  {32'h403f935e, 32'h41430877} /* (7, 0, 26) {real, imag} */,
  {32'h416f6a72, 32'hc23195fa} /* (7, 0, 25) {real, imag} */,
  {32'hc18874d8, 32'h3ff60830} /* (7, 0, 24) {real, imag} */,
  {32'h412b376c, 32'hc05520a8} /* (7, 0, 23) {real, imag} */,
  {32'hc15145dc, 32'h4040b683} /* (7, 0, 22) {real, imag} */,
  {32'hc12f2eea, 32'h412b4290} /* (7, 0, 21) {real, imag} */,
  {32'h3fc057d8, 32'hc199f9a7} /* (7, 0, 20) {real, imag} */,
  {32'h40245ecc, 32'hbf147a5c} /* (7, 0, 19) {real, imag} */,
  {32'h40b6ba40, 32'h4181ca2b} /* (7, 0, 18) {real, imag} */,
  {32'h408432d0, 32'hc0d29cc9} /* (7, 0, 17) {real, imag} */,
  {32'hc0a07d94, 32'h00000000} /* (7, 0, 16) {real, imag} */,
  {32'h408432d0, 32'h40d29cc9} /* (7, 0, 15) {real, imag} */,
  {32'h40b6ba40, 32'hc181ca2b} /* (7, 0, 14) {real, imag} */,
  {32'h40245ecc, 32'h3f147a5c} /* (7, 0, 13) {real, imag} */,
  {32'h3fc057d8, 32'h4199f9a7} /* (7, 0, 12) {real, imag} */,
  {32'hc12f2eea, 32'hc12b4290} /* (7, 0, 11) {real, imag} */,
  {32'hc15145dc, 32'hc040b683} /* (7, 0, 10) {real, imag} */,
  {32'h412b376c, 32'h405520a8} /* (7, 0, 9) {real, imag} */,
  {32'hc18874d8, 32'hbff60830} /* (7, 0, 8) {real, imag} */,
  {32'h416f6a72, 32'h423195fa} /* (7, 0, 7) {real, imag} */,
  {32'h403f935e, 32'hc1430877} /* (7, 0, 6) {real, imag} */,
  {32'hc27f0831, 32'hc1d16c1a} /* (7, 0, 5) {real, imag} */,
  {32'h41635448, 32'hc07d0fa0} /* (7, 0, 4) {real, imag} */,
  {32'hc08e4fcc, 32'h41b3fe6b} /* (7, 0, 3) {real, imag} */,
  {32'hc2ceac6a, 32'hc38336f2} /* (7, 0, 2) {real, imag} */,
  {32'h44846afa, 32'h445b6a80} /* (7, 0, 1) {real, imag} */,
  {32'h44f18902, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h449cbd4a, 32'hc4081355} /* (6, 31, 31) {real, imag} */,
  {32'hc3a4e64a, 32'h439b9bf8} /* (6, 31, 30) {real, imag} */,
  {32'hc1a575ee, 32'h4287893d} /* (6, 31, 29) {real, imag} */,
  {32'h424182cd, 32'h41d536de} /* (6, 31, 28) {real, imag} */,
  {32'hc2702b8e, 32'h4118e236} /* (6, 31, 27) {real, imag} */,
  {32'hc1751b62, 32'h3f9dba94} /* (6, 31, 26) {real, imag} */,
  {32'h41c30ac0, 32'hc0e26ffa} /* (6, 31, 25) {real, imag} */,
  {32'hc124d526, 32'h4206c0c2} /* (6, 31, 24) {real, imag} */,
  {32'h412e01e9, 32'h3e0a9480} /* (6, 31, 23) {real, imag} */,
  {32'hc11af5bc, 32'h400c86b1} /* (6, 31, 22) {real, imag} */,
  {32'hc19db160, 32'h41be8369} /* (6, 31, 21) {real, imag} */,
  {32'hc010ba32, 32'hbfc8daac} /* (6, 31, 20) {real, imag} */,
  {32'h3eafa580, 32'hbfbad3db} /* (6, 31, 19) {real, imag} */,
  {32'h410d0e80, 32'h41807478} /* (6, 31, 18) {real, imag} */,
  {32'hc1213968, 32'hc025f118} /* (6, 31, 17) {real, imag} */,
  {32'hc0eb0cce, 32'hc05e0e18} /* (6, 31, 16) {real, imag} */,
  {32'h404b5712, 32'hc0678f7a} /* (6, 31, 15) {real, imag} */,
  {32'hc1769b04, 32'hc0855a8b} /* (6, 31, 14) {real, imag} */,
  {32'h401c0e6e, 32'h41026814} /* (6, 31, 13) {real, imag} */,
  {32'h416bc1d6, 32'hc0bde156} /* (6, 31, 12) {real, imag} */,
  {32'hc1ab8a8c, 32'hc200b772} /* (6, 31, 11) {real, imag} */,
  {32'h412f1eac, 32'h40f3cda2} /* (6, 31, 10) {real, imag} */,
  {32'h3fc92f8c, 32'h4164a539} /* (6, 31, 9) {real, imag} */,
  {32'hc1af5090, 32'hc0abc1d1} /* (6, 31, 8) {real, imag} */,
  {32'hc1893dee, 32'h3fb26728} /* (6, 31, 7) {real, imag} */,
  {32'h41417d26, 32'hc05fc2fa} /* (6, 31, 6) {real, imag} */,
  {32'hc2b74f0c, 32'h41628e0a} /* (6, 31, 5) {real, imag} */,
  {32'h423ed70e, 32'hc24619ab} /* (6, 31, 4) {real, imag} */,
  {32'h42849d73, 32'h4185217f} /* (6, 31, 3) {real, imag} */,
  {32'hc3393089, 32'h3eb45180} /* (6, 31, 2) {real, imag} */,
  {32'h445e82cb, 32'h437286c0} /* (6, 31, 1) {real, imag} */,
  {32'h449fd30a, 32'hc36b3175} /* (6, 31, 0) {real, imag} */,
  {32'hc39ecffa, 32'hc2a7fa80} /* (6, 30, 31) {real, imag} */,
  {32'h43587e37, 32'h3fc528c0} /* (6, 30, 30) {real, imag} */,
  {32'hc1667c55, 32'hc2203d1e} /* (6, 30, 29) {real, imag} */,
  {32'hc2ae24a7, 32'h4022a7b0} /* (6, 30, 28) {real, imag} */,
  {32'h42340b32, 32'hc116e888} /* (6, 30, 27) {real, imag} */,
  {32'h40a8c640, 32'hc1894c50} /* (6, 30, 26) {real, imag} */,
  {32'hc096b2b2, 32'h41831a6c} /* (6, 30, 25) {real, imag} */,
  {32'h41d86070, 32'hc09d26fc} /* (6, 30, 24) {real, imag} */,
  {32'h41430072, 32'hc172c842} /* (6, 30, 23) {real, imag} */,
  {32'h40c7f755, 32'h3fd7fb10} /* (6, 30, 22) {real, imag} */,
  {32'h412e24dc, 32'hc1bdc8dc} /* (6, 30, 21) {real, imag} */,
  {32'hc13c19f0, 32'h40315e10} /* (6, 30, 20) {real, imag} */,
  {32'h40181f1e, 32'h3f7fed15} /* (6, 30, 19) {real, imag} */,
  {32'h40b8db14, 32'hc035f704} /* (6, 30, 18) {real, imag} */,
  {32'h403f3712, 32'h4106dd8c} /* (6, 30, 17) {real, imag} */,
  {32'hbe16e840, 32'h3f6291a8} /* (6, 30, 16) {real, imag} */,
  {32'hc050d590, 32'hc0568cb6} /* (6, 30, 15) {real, imag} */,
  {32'hc1367104, 32'h4148d701} /* (6, 30, 14) {real, imag} */,
  {32'h40f990fa, 32'hc11849d3} /* (6, 30, 13) {real, imag} */,
  {32'h3fc4a074, 32'hc14a98a3} /* (6, 30, 12) {real, imag} */,
  {32'h40458a1d, 32'h4183d576} /* (6, 30, 11) {real, imag} */,
  {32'h3eb2a800, 32'h40128536} /* (6, 30, 10) {real, imag} */,
  {32'hc178c1be, 32'hbf7957e0} /* (6, 30, 9) {real, imag} */,
  {32'h422d6493, 32'hc1287c6b} /* (6, 30, 8) {real, imag} */,
  {32'hc04aef3c, 32'h4116ee08} /* (6, 30, 7) {real, imag} */,
  {32'h4101b47c, 32'hbf855b60} /* (6, 30, 6) {real, imag} */,
  {32'h41b08e0d, 32'h41fc1d8b} /* (6, 30, 5) {real, imag} */,
  {32'h41094bd4, 32'hc1f6120d} /* (6, 30, 4) {real, imag} */,
  {32'hc2488758, 32'hc21287ec} /* (6, 30, 3) {real, imag} */,
  {32'h43b07012, 32'h42ac400d} /* (6, 30, 2) {real, imag} */,
  {32'hc41ffd87, 32'h3fc49930} /* (6, 30, 1) {real, imag} */,
  {32'hc3aed24a, 32'h43125213} /* (6, 30, 0) {real, imag} */,
  {32'h42b45df8, 32'hc2ed5064} /* (6, 29, 31) {real, imag} */,
  {32'h40bc4c3c, 32'h413546da} /* (6, 29, 30) {real, imag} */,
  {32'hc1cc68e0, 32'h413cb546} /* (6, 29, 29) {real, imag} */,
  {32'hc1d1e1ba, 32'hc10b9f11} /* (6, 29, 28) {real, imag} */,
  {32'h41f5f994, 32'h41d49451} /* (6, 29, 27) {real, imag} */,
  {32'h402fb600, 32'h420e3130} /* (6, 29, 26) {real, imag} */,
  {32'hc1218e82, 32'hc01f6da6} /* (6, 29, 25) {real, imag} */,
  {32'hc17bed88, 32'h41999556} /* (6, 29, 24) {real, imag} */,
  {32'h41948835, 32'hbfa958d0} /* (6, 29, 23) {real, imag} */,
  {32'hc1950e76, 32'hc0cfa509} /* (6, 29, 22) {real, imag} */,
  {32'h417ea02c, 32'hbf4fda6c} /* (6, 29, 21) {real, imag} */,
  {32'hc039026c, 32'h416a9420} /* (6, 29, 20) {real, imag} */,
  {32'h4006d394, 32'h4127f34b} /* (6, 29, 19) {real, imag} */,
  {32'h41cbcf8a, 32'hc0bae89a} /* (6, 29, 18) {real, imag} */,
  {32'hc151dd8e, 32'hc10c2277} /* (6, 29, 17) {real, imag} */,
  {32'hbf4ab9f4, 32'hbfe4e2ca} /* (6, 29, 16) {real, imag} */,
  {32'h41311e3c, 32'hc0c84078} /* (6, 29, 15) {real, imag} */,
  {32'hbfa6261c, 32'h409f8920} /* (6, 29, 14) {real, imag} */,
  {32'h41a3faa6, 32'hc1390170} /* (6, 29, 13) {real, imag} */,
  {32'hc035145c, 32'hc125aad0} /* (6, 29, 12) {real, imag} */,
  {32'hc11cd648, 32'hc173e68d} /* (6, 29, 11) {real, imag} */,
  {32'h3ed07750, 32'h409d62cf} /* (6, 29, 10) {real, imag} */,
  {32'h410eb618, 32'h4024a6cc} /* (6, 29, 9) {real, imag} */,
  {32'h410637ef, 32'h41b2ed8c} /* (6, 29, 8) {real, imag} */,
  {32'hbf6be0a0, 32'h4115739a} /* (6, 29, 7) {real, imag} */,
  {32'hc2112008, 32'hc0e65e23} /* (6, 29, 6) {real, imag} */,
  {32'h409591c0, 32'h40bfc9e7} /* (6, 29, 5) {real, imag} */,
  {32'h41ce4a34, 32'hc1d4a4a1} /* (6, 29, 4) {real, imag} */,
  {32'h40d75f26, 32'h3ea30910} /* (6, 29, 3) {real, imag} */,
  {32'h419eac7a, 32'h42fcaf3a} /* (6, 29, 2) {real, imag} */,
  {32'hc2bb06ef, 32'hc1f5c638} /* (6, 29, 1) {real, imag} */,
  {32'h41c5c137, 32'hc281562d} /* (6, 29, 0) {real, imag} */,
  {32'h42694d46, 32'hc2922f85} /* (6, 28, 31) {real, imag} */,
  {32'hc25b88d7, 32'h42463d81} /* (6, 28, 30) {real, imag} */,
  {32'hc10cc302, 32'hc0abf7cc} /* (6, 28, 29) {real, imag} */,
  {32'h410935ba, 32'hc19139ee} /* (6, 28, 28) {real, imag} */,
  {32'hc18b23d4, 32'h415f882c} /* (6, 28, 27) {real, imag} */,
  {32'hc17ad5f8, 32'hc1f05d98} /* (6, 28, 26) {real, imag} */,
  {32'h403eec46, 32'hc0032086} /* (6, 28, 25) {real, imag} */,
  {32'hc1ba7c42, 32'hc13384fd} /* (6, 28, 24) {real, imag} */,
  {32'h41700d3c, 32'h41513acf} /* (6, 28, 23) {real, imag} */,
  {32'hc1201d00, 32'hc004a154} /* (6, 28, 22) {real, imag} */,
  {32'h3fbfa660, 32'h40782686} /* (6, 28, 21) {real, imag} */,
  {32'hbf115ad0, 32'hc1c27f36} /* (6, 28, 20) {real, imag} */,
  {32'h415482d6, 32'h41945c59} /* (6, 28, 19) {real, imag} */,
  {32'h3f636570, 32'h41594274} /* (6, 28, 18) {real, imag} */,
  {32'hc0c0b34d, 32'hc119a613} /* (6, 28, 17) {real, imag} */,
  {32'hc03ba422, 32'hc0c78412} /* (6, 28, 16) {real, imag} */,
  {32'h40ed938a, 32'h405d3a06} /* (6, 28, 15) {real, imag} */,
  {32'h415c3030, 32'h41433461} /* (6, 28, 14) {real, imag} */,
  {32'hbff049ac, 32'h406f67c2} /* (6, 28, 13) {real, imag} */,
  {32'h4176841e, 32'h3ef1e348} /* (6, 28, 12) {real, imag} */,
  {32'h4124f472, 32'hbffdfa78} /* (6, 28, 11) {real, imag} */,
  {32'hc19a3ab7, 32'h3fc14a5a} /* (6, 28, 10) {real, imag} */,
  {32'hc0f96c39, 32'h4089e54c} /* (6, 28, 9) {real, imag} */,
  {32'hc1a270ce, 32'h40e9add8} /* (6, 28, 8) {real, imag} */,
  {32'hc0325355, 32'hc104d2ef} /* (6, 28, 7) {real, imag} */,
  {32'h400a21b4, 32'h419ae96e} /* (6, 28, 6) {real, imag} */,
  {32'h3ff00f0a, 32'hc1444c9e} /* (6, 28, 5) {real, imag} */,
  {32'h4139a3ff, 32'h415341c9} /* (6, 28, 4) {real, imag} */,
  {32'h410e828e, 32'hc14496fe} /* (6, 28, 3) {real, imag} */,
  {32'hc236af96, 32'h425036cd} /* (6, 28, 2) {real, imag} */,
  {32'h41171e0e, 32'hc25e02ae} /* (6, 28, 1) {real, imag} */,
  {32'h423ff7ff, 32'h40e215a8} /* (6, 28, 0) {real, imag} */,
  {32'hc188b77c, 32'h42501214} /* (6, 27, 31) {real, imag} */,
  {32'h41eb0e63, 32'hc21b3060} /* (6, 27, 30) {real, imag} */,
  {32'hbdcec240, 32'hc14ff8c1} /* (6, 27, 29) {real, imag} */,
  {32'hc0b7f7a2, 32'h412bd8e5} /* (6, 27, 28) {real, imag} */,
  {32'h40033d94, 32'hc0f27dc0} /* (6, 27, 27) {real, imag} */,
  {32'h414310f8, 32'hc10564d2} /* (6, 27, 26) {real, imag} */,
  {32'hc10bff0d, 32'h4079e8f8} /* (6, 27, 25) {real, imag} */,
  {32'h40563eac, 32'h414bdfd9} /* (6, 27, 24) {real, imag} */,
  {32'hc118c2e6, 32'h41091009} /* (6, 27, 23) {real, imag} */,
  {32'hc0a42274, 32'hc11dfa80} /* (6, 27, 22) {real, imag} */,
  {32'h4130dca6, 32'hc137c138} /* (6, 27, 21) {real, imag} */,
  {32'hc0efae90, 32'h41be7872} /* (6, 27, 20) {real, imag} */,
  {32'h40d7544c, 32'hc12b5fde} /* (6, 27, 19) {real, imag} */,
  {32'h3f96ab78, 32'hc00f2bf4} /* (6, 27, 18) {real, imag} */,
  {32'h3fc9d02c, 32'h3c8529c0} /* (6, 27, 17) {real, imag} */,
  {32'h3da6b440, 32'h40dd36f9} /* (6, 27, 16) {real, imag} */,
  {32'hc0f662e1, 32'hbf8164ac} /* (6, 27, 15) {real, imag} */,
  {32'hbd875d60, 32'h3ff046f4} /* (6, 27, 14) {real, imag} */,
  {32'hc0626f96, 32'h413253e6} /* (6, 27, 13) {real, imag} */,
  {32'h41241177, 32'h41580c18} /* (6, 27, 12) {real, imag} */,
  {32'h40eea60b, 32'h41da0ec7} /* (6, 27, 11) {real, imag} */,
  {32'hc1762ffc, 32'hc1bef540} /* (6, 27, 10) {real, imag} */,
  {32'h400ebfca, 32'h408d85e3} /* (6, 27, 9) {real, imag} */,
  {32'hc0f04bf9, 32'hc0fa7c4f} /* (6, 27, 8) {real, imag} */,
  {32'hc09b52d6, 32'hc0cb9210} /* (6, 27, 7) {real, imag} */,
  {32'h40a3f8b1, 32'h3ffb6f42} /* (6, 27, 6) {real, imag} */,
  {32'h42040590, 32'hc1545966} /* (6, 27, 5) {real, imag} */,
  {32'hc21219f4, 32'h40adb710} /* (6, 27, 4) {real, imag} */,
  {32'hc19598a2, 32'hc0625794} /* (6, 27, 3) {real, imag} */,
  {32'h42461b96, 32'hc1a59a98} /* (6, 27, 2) {real, imag} */,
  {32'hc26929f8, 32'hc23528e2} /* (6, 27, 1) {real, imag} */,
  {32'hc25de6d8, 32'h41e02773} /* (6, 27, 0) {real, imag} */,
  {32'hc1f25449, 32'hc1ba5230} /* (6, 26, 31) {real, imag} */,
  {32'hc2323dbd, 32'hc1387a7e} /* (6, 26, 30) {real, imag} */,
  {32'hc1ba26b1, 32'h419fc4f8} /* (6, 26, 29) {real, imag} */,
  {32'h411b2dc6, 32'hc09521bc} /* (6, 26, 28) {real, imag} */,
  {32'hc0f52a8c, 32'hc15241eb} /* (6, 26, 27) {real, imag} */,
  {32'hbcf91200, 32'hc129fe2c} /* (6, 26, 26) {real, imag} */,
  {32'h41c354a0, 32'h41422846} /* (6, 26, 25) {real, imag} */,
  {32'h3f46d490, 32'hc1015a9a} /* (6, 26, 24) {real, imag} */,
  {32'h404cd7a8, 32'hc1c2697a} /* (6, 26, 23) {real, imag} */,
  {32'h40c7178b, 32'hc0d809a2} /* (6, 26, 22) {real, imag} */,
  {32'h4155870c, 32'h3f219fd0} /* (6, 26, 21) {real, imag} */,
  {32'hc089dd10, 32'h40849a1f} /* (6, 26, 20) {real, imag} */,
  {32'hc078291c, 32'h40ecdc0a} /* (6, 26, 19) {real, imag} */,
  {32'hbfa7852a, 32'h4071f654} /* (6, 26, 18) {real, imag} */,
  {32'h3ca36900, 32'hc109df2c} /* (6, 26, 17) {real, imag} */,
  {32'hbfb2243c, 32'hc00431d0} /* (6, 26, 16) {real, imag} */,
  {32'hc1a2b1f6, 32'h41707c04} /* (6, 26, 15) {real, imag} */,
  {32'h408ed292, 32'hc1261958} /* (6, 26, 14) {real, imag} */,
  {32'hc105bcb2, 32'h41ac5708} /* (6, 26, 13) {real, imag} */,
  {32'h3f8cbbc6, 32'hc0287c12} /* (6, 26, 12) {real, imag} */,
  {32'hc15e5b16, 32'h4108b3ef} /* (6, 26, 11) {real, imag} */,
  {32'h4093aefc, 32'hc04c3652} /* (6, 26, 10) {real, imag} */,
  {32'hc00b0936, 32'h418a3c23} /* (6, 26, 9) {real, imag} */,
  {32'hbf821c32, 32'h3fa00d60} /* (6, 26, 8) {real, imag} */,
  {32'h410cc555, 32'hc1858720} /* (6, 26, 7) {real, imag} */,
  {32'h41853e5a, 32'h4122980e} /* (6, 26, 6) {real, imag} */,
  {32'hbfb6bffc, 32'hc0f7c3e6} /* (6, 26, 5) {real, imag} */,
  {32'h40f47737, 32'h40f202ba} /* (6, 26, 4) {real, imag} */,
  {32'hc118f380, 32'hc05ae2c4} /* (6, 26, 3) {real, imag} */,
  {32'hc15a9cf6, 32'h419195f0} /* (6, 26, 2) {real, imag} */,
  {32'h4147d0d2, 32'hc1bdc1ec} /* (6, 26, 1) {real, imag} */,
  {32'h3f76d520, 32'h41b91890} /* (6, 26, 0) {real, imag} */,
  {32'hc0a5e802, 32'hc1aa930f} /* (6, 25, 31) {real, imag} */,
  {32'h40ae506c, 32'h41a5af8c} /* (6, 25, 30) {real, imag} */,
  {32'h3fb921c8, 32'hc128c78a} /* (6, 25, 29) {real, imag} */,
  {32'h41996716, 32'hc15f5b22} /* (6, 25, 28) {real, imag} */,
  {32'h41530722, 32'h4075e6c2} /* (6, 25, 27) {real, imag} */,
  {32'h41c3ecb4, 32'hc0b2e572} /* (6, 25, 26) {real, imag} */,
  {32'hbfac60c8, 32'hc0b31cb9} /* (6, 25, 25) {real, imag} */,
  {32'hc07de2d2, 32'hc0f0d761} /* (6, 25, 24) {real, imag} */,
  {32'h41980028, 32'hbfea490c} /* (6, 25, 23) {real, imag} */,
  {32'h3f627ac0, 32'h409385b9} /* (6, 25, 22) {real, imag} */,
  {32'hc096216c, 32'h4065748e} /* (6, 25, 21) {real, imag} */,
  {32'hbf411de0, 32'h4087f729} /* (6, 25, 20) {real, imag} */,
  {32'h410b6d3c, 32'hc00215d1} /* (6, 25, 19) {real, imag} */,
  {32'h41048564, 32'h3fd62005} /* (6, 25, 18) {real, imag} */,
  {32'hc14cd932, 32'hc0d119ce} /* (6, 25, 17) {real, imag} */,
  {32'hc1772f22, 32'h400f89d1} /* (6, 25, 16) {real, imag} */,
  {32'hbf14f88a, 32'h40d173dc} /* (6, 25, 15) {real, imag} */,
  {32'h40034462, 32'h418c8496} /* (6, 25, 14) {real, imag} */,
  {32'hc168c74a, 32'hc13da0e6} /* (6, 25, 13) {real, imag} */,
  {32'hc083e732, 32'h412979fe} /* (6, 25, 12) {real, imag} */,
  {32'h40feebc2, 32'hbfe92808} /* (6, 25, 11) {real, imag} */,
  {32'hc0e106c7, 32'hc1ccfa39} /* (6, 25, 10) {real, imag} */,
  {32'hc15c88d2, 32'hc0644d00} /* (6, 25, 9) {real, imag} */,
  {32'h40aa2e4a, 32'h3fcc0168} /* (6, 25, 8) {real, imag} */,
  {32'h4129dc72, 32'h41ae2f00} /* (6, 25, 7) {real, imag} */,
  {32'hc1a23f48, 32'h3ef113c0} /* (6, 25, 6) {real, imag} */,
  {32'hc003be64, 32'hc192afb1} /* (6, 25, 5) {real, imag} */,
  {32'hc1d6b4e8, 32'h4081b000} /* (6, 25, 4) {real, imag} */,
  {32'hc17274f6, 32'hc16590e5} /* (6, 25, 3) {real, imag} */,
  {32'hc01232a4, 32'hc17ade4b} /* (6, 25, 2) {real, imag} */,
  {32'h4188278e, 32'hc19b5262} /* (6, 25, 1) {real, imag} */,
  {32'h40ff5802, 32'h40708bed} /* (6, 25, 0) {real, imag} */,
  {32'hc1e94d0c, 32'h41c80658} /* (6, 24, 31) {real, imag} */,
  {32'h41edbb79, 32'hc124b57d} /* (6, 24, 30) {real, imag} */,
  {32'h3fd28dc0, 32'hc0d77852} /* (6, 24, 29) {real, imag} */,
  {32'hc1568347, 32'h417c68f3} /* (6, 24, 28) {real, imag} */,
  {32'hc1870efe, 32'hc0c3ea96} /* (6, 24, 27) {real, imag} */,
  {32'hc1c2933c, 32'hc0361ffd} /* (6, 24, 26) {real, imag} */,
  {32'h409c97c8, 32'hc043b98c} /* (6, 24, 25) {real, imag} */,
  {32'hc00591a4, 32'hc18a90ec} /* (6, 24, 24) {real, imag} */,
  {32'hc1828819, 32'hc188bd20} /* (6, 24, 23) {real, imag} */,
  {32'hc0aef400, 32'h3d9cf000} /* (6, 24, 22) {real, imag} */,
  {32'h411a4d44, 32'hc0f0dc23} /* (6, 24, 21) {real, imag} */,
  {32'h3f38a91e, 32'hc13eaca8} /* (6, 24, 20) {real, imag} */,
  {32'h40a9b190, 32'h3fb7515a} /* (6, 24, 19) {real, imag} */,
  {32'h4095d88f, 32'h41324ddb} /* (6, 24, 18) {real, imag} */,
  {32'h412793e2, 32'hc11f2b87} /* (6, 24, 17) {real, imag} */,
  {32'h40ecc261, 32'hc10837df} /* (6, 24, 16) {real, imag} */,
  {32'hc0ff0707, 32'hbe9366a0} /* (6, 24, 15) {real, imag} */,
  {32'hc00644c8, 32'h4030405b} /* (6, 24, 14) {real, imag} */,
  {32'h40a3beff, 32'hc07827ee} /* (6, 24, 13) {real, imag} */,
  {32'hc104844e, 32'h4048abd2} /* (6, 24, 12) {real, imag} */,
  {32'h4152de4a, 32'hc0b76523} /* (6, 24, 11) {real, imag} */,
  {32'hc07d1440, 32'hc0da7b1a} /* (6, 24, 10) {real, imag} */,
  {32'h41137530, 32'hc00adae6} /* (6, 24, 9) {real, imag} */,
  {32'h4132582e, 32'h411dcacc} /* (6, 24, 8) {real, imag} */,
  {32'hbe4be340, 32'h41363465} /* (6, 24, 7) {real, imag} */,
  {32'h3fd7a6c8, 32'h408c094a} /* (6, 24, 6) {real, imag} */,
  {32'h41b9e2a0, 32'h416b7a88} /* (6, 24, 5) {real, imag} */,
  {32'hc1ac51df, 32'hc191b442} /* (6, 24, 4) {real, imag} */,
  {32'h4150e104, 32'hc1ac9af2} /* (6, 24, 3) {real, imag} */,
  {32'h4199af10, 32'hc070a2e7} /* (6, 24, 2) {real, imag} */,
  {32'hc1f0afaa, 32'h41a2f0a1} /* (6, 24, 1) {real, imag} */,
  {32'hc1f2cf56, 32'h4207d76e} /* (6, 24, 0) {real, imag} */,
  {32'h3f4e5bf4, 32'hc09c9553} /* (6, 23, 31) {real, imag} */,
  {32'hc077f940, 32'h419459c4} /* (6, 23, 30) {real, imag} */,
  {32'h41dc493b, 32'hc108a96e} /* (6, 23, 29) {real, imag} */,
  {32'hc09a39c2, 32'h41881570} /* (6, 23, 28) {real, imag} */,
  {32'h41408947, 32'h3f75cf70} /* (6, 23, 27) {real, imag} */,
  {32'h410a79d8, 32'hc0d0e5e9} /* (6, 23, 26) {real, imag} */,
  {32'h4180addf, 32'h3fba01c8} /* (6, 23, 25) {real, imag} */,
  {32'h40d4b958, 32'hbf9a0578} /* (6, 23, 24) {real, imag} */,
  {32'h410a5192, 32'hc1909d0d} /* (6, 23, 23) {real, imag} */,
  {32'hc0239f27, 32'h42335d9a} /* (6, 23, 22) {real, imag} */,
  {32'hc0b52fd7, 32'h3fc31454} /* (6, 23, 21) {real, imag} */,
  {32'hbf4b9760, 32'hc10be03e} /* (6, 23, 20) {real, imag} */,
  {32'hbeee6230, 32'hc0e2c92f} /* (6, 23, 19) {real, imag} */,
  {32'hbfa013cc, 32'hbf953b81} /* (6, 23, 18) {real, imag} */,
  {32'hc1671edd, 32'hc0da9202} /* (6, 23, 17) {real, imag} */,
  {32'hbfe1fe60, 32'hc06d0371} /* (6, 23, 16) {real, imag} */,
  {32'hc0a7da75, 32'hc180523f} /* (6, 23, 15) {real, imag} */,
  {32'h410fcd0c, 32'h3f7701e0} /* (6, 23, 14) {real, imag} */,
  {32'hc1eed2e7, 32'hc1852710} /* (6, 23, 13) {real, imag} */,
  {32'h4166138f, 32'hc1cecede} /* (6, 23, 12) {real, imag} */,
  {32'h40646ef2, 32'h414b4c3a} /* (6, 23, 11) {real, imag} */,
  {32'hc091229d, 32'h411b054f} /* (6, 23, 10) {real, imag} */,
  {32'h3fe528c9, 32'hc04538a4} /* (6, 23, 9) {real, imag} */,
  {32'hc085a6f4, 32'hc16e75a0} /* (6, 23, 8) {real, imag} */,
  {32'hbf402e40, 32'hc1156fd3} /* (6, 23, 7) {real, imag} */,
  {32'hc05b1b77, 32'h417a202d} /* (6, 23, 6) {real, imag} */,
  {32'hbfc946c6, 32'hc0f8137a} /* (6, 23, 5) {real, imag} */,
  {32'hc053a2d6, 32'hc18db652} /* (6, 23, 4) {real, imag} */,
  {32'hc14487f8, 32'h41668f96} /* (6, 23, 3) {real, imag} */,
  {32'h3e63eb40, 32'hc0deb6b6} /* (6, 23, 2) {real, imag} */,
  {32'hc0291446, 32'hc1d60dc0} /* (6, 23, 1) {real, imag} */,
  {32'hc1410ec0, 32'hc192713c} /* (6, 23, 0) {real, imag} */,
  {32'h418ff111, 32'h40d1efee} /* (6, 22, 31) {real, imag} */,
  {32'hc15515e8, 32'h41cd9bfa} /* (6, 22, 30) {real, imag} */,
  {32'hc180027c, 32'hc0307a14} /* (6, 22, 29) {real, imag} */,
  {32'hbf956669, 32'hc08e48ca} /* (6, 22, 28) {real, imag} */,
  {32'h40cab31c, 32'h4115d26b} /* (6, 22, 27) {real, imag} */,
  {32'h3f05f5f0, 32'hc13e755f} /* (6, 22, 26) {real, imag} */,
  {32'h4158df24, 32'hc0b0fc8a} /* (6, 22, 25) {real, imag} */,
  {32'h4131462a, 32'h417306be} /* (6, 22, 24) {real, imag} */,
  {32'hc17c7dad, 32'h41acf84a} /* (6, 22, 23) {real, imag} */,
  {32'hc1ad4f58, 32'hc1c63174} /* (6, 22, 22) {real, imag} */,
  {32'h417500b2, 32'h41333171} /* (6, 22, 21) {real, imag} */,
  {32'hc09ec6ba, 32'hc0e1c4a4} /* (6, 22, 20) {real, imag} */,
  {32'hc18d9cce, 32'hc10925aa} /* (6, 22, 19) {real, imag} */,
  {32'h4126951e, 32'hc1a780e8} /* (6, 22, 18) {real, imag} */,
  {32'hbff339b6, 32'hc0d49d4b} /* (6, 22, 17) {real, imag} */,
  {32'hc0c44769, 32'h40f00cda} /* (6, 22, 16) {real, imag} */,
  {32'h4111f71c, 32'hbcd57e40} /* (6, 22, 15) {real, imag} */,
  {32'hc0fdd2f2, 32'hbf3bf0f0} /* (6, 22, 14) {real, imag} */,
  {32'hc1039fa8, 32'hc0a24a5a} /* (6, 22, 13) {real, imag} */,
  {32'hc082e346, 32'h40ae9ec9} /* (6, 22, 12) {real, imag} */,
  {32'hc0c24b6a, 32'h414adcae} /* (6, 22, 11) {real, imag} */,
  {32'h3feeeaf8, 32'hc1b229a6} /* (6, 22, 10) {real, imag} */,
  {32'h4049d454, 32'h3fc5b920} /* (6, 22, 9) {real, imag} */,
  {32'h40ccce45, 32'h41572acc} /* (6, 22, 8) {real, imag} */,
  {32'h400ca2ac, 32'hc055916a} /* (6, 22, 7) {real, imag} */,
  {32'h4167e346, 32'h41731b00} /* (6, 22, 6) {real, imag} */,
  {32'h3fc65e04, 32'hbfb74894} /* (6, 22, 5) {real, imag} */,
  {32'h414bc55e, 32'hbe8f17b4} /* (6, 22, 4) {real, imag} */,
  {32'hc0af7e17, 32'h41a69520} /* (6, 22, 3) {real, imag} */,
  {32'hc0e45c46, 32'h41f184d0} /* (6, 22, 2) {real, imag} */,
  {32'hc19044d4, 32'hc0e5fece} /* (6, 22, 1) {real, imag} */,
  {32'hc12071da, 32'hc206e6e9} /* (6, 22, 0) {real, imag} */,
  {32'hbfb7f768, 32'h41edb7e6} /* (6, 21, 31) {real, imag} */,
  {32'hc059996d, 32'hc1dbeb42} /* (6, 21, 30) {real, imag} */,
  {32'hc0ff92cc, 32'hc13646dc} /* (6, 21, 29) {real, imag} */,
  {32'hc11fdb73, 32'hc19a6a70} /* (6, 21, 28) {real, imag} */,
  {32'h40d2859e, 32'h3f147108} /* (6, 21, 27) {real, imag} */,
  {32'hc091a11d, 32'h410557e7} /* (6, 21, 26) {real, imag} */,
  {32'hc148d70a, 32'h411404d3} /* (6, 21, 25) {real, imag} */,
  {32'hc0b5955e, 32'hc15e14a7} /* (6, 21, 24) {real, imag} */,
  {32'hbf97ae9e, 32'h4197bedd} /* (6, 21, 23) {real, imag} */,
  {32'hc09024b4, 32'h4183142c} /* (6, 21, 22) {real, imag} */,
  {32'hc11b0f5c, 32'hbed76300} /* (6, 21, 21) {real, imag} */,
  {32'h41882813, 32'hc0267abe} /* (6, 21, 20) {real, imag} */,
  {32'h40cfae3a, 32'hc152e5a7} /* (6, 21, 19) {real, imag} */,
  {32'hc0a2462e, 32'hc039feb3} /* (6, 21, 18) {real, imag} */,
  {32'hbc99d200, 32'hc1545cfa} /* (6, 21, 17) {real, imag} */,
  {32'hc0244595, 32'hbf8ce07c} /* (6, 21, 16) {real, imag} */,
  {32'hc0c458a1, 32'h3f39c6b0} /* (6, 21, 15) {real, imag} */,
  {32'hc087e2a4, 32'h4019176c} /* (6, 21, 14) {real, imag} */,
  {32'h41233bdf, 32'h41ad7946} /* (6, 21, 13) {real, imag} */,
  {32'hc0be7283, 32'hc045ff8a} /* (6, 21, 12) {real, imag} */,
  {32'hc10fefee, 32'hc1afe4c0} /* (6, 21, 11) {real, imag} */,
  {32'hc0f38ee1, 32'hc14b77a8} /* (6, 21, 10) {real, imag} */,
  {32'h4140c697, 32'hc0d0aa52} /* (6, 21, 9) {real, imag} */,
  {32'h4148ac3c, 32'hc08fe6e7} /* (6, 21, 8) {real, imag} */,
  {32'h411fa7ec, 32'h412b5800} /* (6, 21, 7) {real, imag} */,
  {32'h411140fd, 32'h41148570} /* (6, 21, 6) {real, imag} */,
  {32'hc06da93c, 32'hc033c00e} /* (6, 21, 5) {real, imag} */,
  {32'hc032f47c, 32'h40ae7080} /* (6, 21, 4) {real, imag} */,
  {32'hc036736e, 32'hc048e4e8} /* (6, 21, 3) {real, imag} */,
  {32'h40a4a528, 32'hc0eb88ba} /* (6, 21, 2) {real, imag} */,
  {32'hc134a1f9, 32'h419a9502} /* (6, 21, 1) {real, imag} */,
  {32'h4147da22, 32'h4121e9e4} /* (6, 21, 0) {real, imag} */,
  {32'hc0ced62d, 32'h415aa48c} /* (6, 20, 31) {real, imag} */,
  {32'hbf8fc158, 32'hc09d2c56} /* (6, 20, 30) {real, imag} */,
  {32'hc183f567, 32'hc02882c2} /* (6, 20, 29) {real, imag} */,
  {32'h40ff155f, 32'hc031dc27} /* (6, 20, 28) {real, imag} */,
  {32'h3f0d16a8, 32'hc0a30e64} /* (6, 20, 27) {real, imag} */,
  {32'hc0abe016, 32'hc0ec3316} /* (6, 20, 26) {real, imag} */,
  {32'h414a39c4, 32'h40188ce8} /* (6, 20, 25) {real, imag} */,
  {32'h40d67a64, 32'hc16d9831} /* (6, 20, 24) {real, imag} */,
  {32'h410747b1, 32'hc12769fc} /* (6, 20, 23) {real, imag} */,
  {32'hc17ec0df, 32'hbf8e52d4} /* (6, 20, 22) {real, imag} */,
  {32'hc0dcd7bf, 32'hbf2734b8} /* (6, 20, 21) {real, imag} */,
  {32'h40155a42, 32'h41743535} /* (6, 20, 20) {real, imag} */,
  {32'h40da52e5, 32'h414b18c0} /* (6, 20, 19) {real, imag} */,
  {32'hc1397bd8, 32'hbf92bcd6} /* (6, 20, 18) {real, imag} */,
  {32'h408d8432, 32'hc18a4295} /* (6, 20, 17) {real, imag} */,
  {32'hbf8ddca4, 32'hc0d7546a} /* (6, 20, 16) {real, imag} */,
  {32'h4119cc85, 32'h40f3e896} /* (6, 20, 15) {real, imag} */,
  {32'h40994d21, 32'h3ff5cf3a} /* (6, 20, 14) {real, imag} */,
  {32'h40c1eb62, 32'hc1516cb2} /* (6, 20, 13) {real, imag} */,
  {32'hbfe5cd34, 32'h41653052} /* (6, 20, 12) {real, imag} */,
  {32'h41344244, 32'hc0a11ca6} /* (6, 20, 11) {real, imag} */,
  {32'h40a94351, 32'hc08f4ea8} /* (6, 20, 10) {real, imag} */,
  {32'h40b121b8, 32'h40dc1c5f} /* (6, 20, 9) {real, imag} */,
  {32'hc0f84860, 32'h4090cdfb} /* (6, 20, 8) {real, imag} */,
  {32'hc15f9120, 32'hc1169f67} /* (6, 20, 7) {real, imag} */,
  {32'h40c481cd, 32'hc10256d8} /* (6, 20, 6) {real, imag} */,
  {32'h412be18c, 32'hbfafa3a8} /* (6, 20, 5) {real, imag} */,
  {32'h40bae797, 32'h412b363d} /* (6, 20, 4) {real, imag} */,
  {32'hbddb9980, 32'h3fa447c0} /* (6, 20, 3) {real, imag} */,
  {32'hc055bb68, 32'h4095d054} /* (6, 20, 2) {real, imag} */,
  {32'h41165b8e, 32'h4112a665} /* (6, 20, 1) {real, imag} */,
  {32'hc0b82c6d, 32'hc12ff3fb} /* (6, 20, 0) {real, imag} */,
  {32'h410dbce0, 32'hc1636ef1} /* (6, 19, 31) {real, imag} */,
  {32'h40ee07ef, 32'h415b1e67} /* (6, 19, 30) {real, imag} */,
  {32'hbed7e720, 32'h3f8de098} /* (6, 19, 29) {real, imag} */,
  {32'hbe9da860, 32'hc0c62b30} /* (6, 19, 28) {real, imag} */,
  {32'h40eb2508, 32'h3e4e38c0} /* (6, 19, 27) {real, imag} */,
  {32'h4185fd17, 32'h40965e2c} /* (6, 19, 26) {real, imag} */,
  {32'hc125e8ff, 32'hc1073b4c} /* (6, 19, 25) {real, imag} */,
  {32'h40f53082, 32'hc16f2f3c} /* (6, 19, 24) {real, imag} */,
  {32'hc1891b2a, 32'h401233cc} /* (6, 19, 23) {real, imag} */,
  {32'hc08332c3, 32'h40b2fdd0} /* (6, 19, 22) {real, imag} */,
  {32'hc0031afc, 32'hc11b34a4} /* (6, 19, 21) {real, imag} */,
  {32'h40cfd7c7, 32'h403f0d94} /* (6, 19, 20) {real, imag} */,
  {32'hc155dff2, 32'hc1254b22} /* (6, 19, 19) {real, imag} */,
  {32'h403f30cc, 32'hc00aa9ac} /* (6, 19, 18) {real, imag} */,
  {32'hc032cf15, 32'h415acb83} /* (6, 19, 17) {real, imag} */,
  {32'h3fc23c69, 32'hc08b07aa} /* (6, 19, 16) {real, imag} */,
  {32'h404a2956, 32'hbdf4d020} /* (6, 19, 15) {real, imag} */,
  {32'hc090d9d0, 32'hc0b59d22} /* (6, 19, 14) {real, imag} */,
  {32'h40db5c0c, 32'h415388e0} /* (6, 19, 13) {real, imag} */,
  {32'hc1600398, 32'h409adec6} /* (6, 19, 12) {real, imag} */,
  {32'hc0945755, 32'hc0b824ad} /* (6, 19, 11) {real, imag} */,
  {32'h412f4f85, 32'h41147e7c} /* (6, 19, 10) {real, imag} */,
  {32'h404007ec, 32'h4103fdcd} /* (6, 19, 9) {real, imag} */,
  {32'h3ff4bdd2, 32'hc0c4d71c} /* (6, 19, 8) {real, imag} */,
  {32'h412cc9fc, 32'hc01f30b1} /* (6, 19, 7) {real, imag} */,
  {32'hbf271a80, 32'hbde47d20} /* (6, 19, 6) {real, imag} */,
  {32'hc1683e9e, 32'h3fe0d5c8} /* (6, 19, 5) {real, imag} */,
  {32'hc01f39d6, 32'h40960674} /* (6, 19, 4) {real, imag} */,
  {32'h410a05fc, 32'hc0d77f42} /* (6, 19, 3) {real, imag} */,
  {32'hc0d5c405, 32'hbd676e00} /* (6, 19, 2) {real, imag} */,
  {32'hbfc8976c, 32'h41924165} /* (6, 19, 1) {real, imag} */,
  {32'h40ba8ad4, 32'hc1770261} /* (6, 19, 0) {real, imag} */,
  {32'hc102f185, 32'h3ec0a250} /* (6, 18, 31) {real, imag} */,
  {32'h414ac3cd, 32'hc0a5643b} /* (6, 18, 30) {real, imag} */,
  {32'h410e9177, 32'hc006d5e0} /* (6, 18, 29) {real, imag} */,
  {32'hc11108cd, 32'h3f9482fe} /* (6, 18, 28) {real, imag} */,
  {32'hbf8f22ca, 32'hc152e9de} /* (6, 18, 27) {real, imag} */,
  {32'hc07251f1, 32'hc15c36ab} /* (6, 18, 26) {real, imag} */,
  {32'hc122c903, 32'hc106e040} /* (6, 18, 25) {real, imag} */,
  {32'hc1041503, 32'h3ea78f8c} /* (6, 18, 24) {real, imag} */,
  {32'h409bb96e, 32'h40430c34} /* (6, 18, 23) {real, imag} */,
  {32'h41725a54, 32'hc0a3eecb} /* (6, 18, 22) {real, imag} */,
  {32'hc1f1a9d2, 32'hbc459c00} /* (6, 18, 21) {real, imag} */,
  {32'hbf8fee60, 32'hbfad7970} /* (6, 18, 20) {real, imag} */,
  {32'h40d4d026, 32'h40a1ca1a} /* (6, 18, 19) {real, imag} */,
  {32'h40721caa, 32'hc104c775} /* (6, 18, 18) {real, imag} */,
  {32'h41124ea5, 32'hc10982cb} /* (6, 18, 17) {real, imag} */,
  {32'hc0eba45d, 32'hc066018d} /* (6, 18, 16) {real, imag} */,
  {32'hc1075ab4, 32'hc0c83d84} /* (6, 18, 15) {real, imag} */,
  {32'h412f5613, 32'h40fa4688} /* (6, 18, 14) {real, imag} */,
  {32'hc0c4d74e, 32'h4135534a} /* (6, 18, 13) {real, imag} */,
  {32'h40a5dc33, 32'hc1b35d1c} /* (6, 18, 12) {real, imag} */,
  {32'h4101cbd8, 32'h3eff4a1c} /* (6, 18, 11) {real, imag} */,
  {32'hc1934589, 32'h416066d4} /* (6, 18, 10) {real, imag} */,
  {32'hc1237c36, 32'h415ae775} /* (6, 18, 9) {real, imag} */,
  {32'hc15e746a, 32'h41a4235c} /* (6, 18, 8) {real, imag} */,
  {32'hc1678cb6, 32'h3f98e298} /* (6, 18, 7) {real, imag} */,
  {32'hbdb19e80, 32'hc093b5b0} /* (6, 18, 6) {real, imag} */,
  {32'h4007038a, 32'hc0d5fa26} /* (6, 18, 5) {real, imag} */,
  {32'h3fae7a76, 32'hc1030567} /* (6, 18, 4) {real, imag} */,
  {32'h40898c6c, 32'hc153724e} /* (6, 18, 3) {real, imag} */,
  {32'hc0a6fa77, 32'hc10f1400} /* (6, 18, 2) {real, imag} */,
  {32'h4145b862, 32'h41e842cb} /* (6, 18, 1) {real, imag} */,
  {32'hbfd4305a, 32'h40b3f654} /* (6, 18, 0) {real, imag} */,
  {32'h419afcd5, 32'hc0587615} /* (6, 17, 31) {real, imag} */,
  {32'hbe73d8ac, 32'h4103ae97} /* (6, 17, 30) {real, imag} */,
  {32'hbf828770, 32'hc09f5162} /* (6, 17, 29) {real, imag} */,
  {32'hc053b349, 32'h4134afaa} /* (6, 17, 28) {real, imag} */,
  {32'hc0a32944, 32'hc0f6c924} /* (6, 17, 27) {real, imag} */,
  {32'h3f8e4ec7, 32'h409f85e6} /* (6, 17, 26) {real, imag} */,
  {32'h3fd2125a, 32'hc0e89ea9} /* (6, 17, 25) {real, imag} */,
  {32'h407092c6, 32'hbffb747f} /* (6, 17, 24) {real, imag} */,
  {32'hc0e0568a, 32'hc05488be} /* (6, 17, 23) {real, imag} */,
  {32'h408bcedd, 32'h40c5db8e} /* (6, 17, 22) {real, imag} */,
  {32'h3ea01520, 32'hc08c7cb5} /* (6, 17, 21) {real, imag} */,
  {32'h41dbac1c, 32'hc0bf0a02} /* (6, 17, 20) {real, imag} */,
  {32'hbfce231a, 32'h3f6105f4} /* (6, 17, 19) {real, imag} */,
  {32'hc0bd0bb8, 32'hbd4e8880} /* (6, 17, 18) {real, imag} */,
  {32'h404c515f, 32'hc00277d0} /* (6, 17, 17) {real, imag} */,
  {32'h400f7799, 32'hc0e72008} /* (6, 17, 16) {real, imag} */,
  {32'hc073b8c2, 32'h40938784} /* (6, 17, 15) {real, imag} */,
  {32'h402b3009, 32'h414146c8} /* (6, 17, 14) {real, imag} */,
  {32'h40fb13e4, 32'hbf647030} /* (6, 17, 13) {real, imag} */,
  {32'hc08f6dd6, 32'h40cbf2c2} /* (6, 17, 12) {real, imag} */,
  {32'hc12fa412, 32'h3ec4f178} /* (6, 17, 11) {real, imag} */,
  {32'hc121d247, 32'hc00cf674} /* (6, 17, 10) {real, imag} */,
  {32'hc109a6a4, 32'hc163382c} /* (6, 17, 9) {real, imag} */,
  {32'hc1001617, 32'hc003cee5} /* (6, 17, 8) {real, imag} */,
  {32'hc141223e, 32'h41334b8d} /* (6, 17, 7) {real, imag} */,
  {32'hbecce680, 32'hc057daca} /* (6, 17, 6) {real, imag} */,
  {32'hc0ae1419, 32'hc09b375b} /* (6, 17, 5) {real, imag} */,
  {32'hc0c64bdc, 32'hc0dec928} /* (6, 17, 4) {real, imag} */,
  {32'h41100784, 32'h4051e196} /* (6, 17, 3) {real, imag} */,
  {32'h3fd9a640, 32'hc03aa65e} /* (6, 17, 2) {real, imag} */,
  {32'hc04c4072, 32'hc0fea9b8} /* (6, 17, 1) {real, imag} */,
  {32'h40bc5de9, 32'hc185407f} /* (6, 17, 0) {real, imag} */,
  {32'h410eb71d, 32'h410e33a8} /* (6, 16, 31) {real, imag} */,
  {32'hc097d354, 32'h406395a8} /* (6, 16, 30) {real, imag} */,
  {32'hc0790023, 32'h401a2dfe} /* (6, 16, 29) {real, imag} */,
  {32'hc1317221, 32'h40929320} /* (6, 16, 28) {real, imag} */,
  {32'hc12c5cc6, 32'h4097071e} /* (6, 16, 27) {real, imag} */,
  {32'h40bc0cbc, 32'h3f824932} /* (6, 16, 26) {real, imag} */,
  {32'h4105dc86, 32'h40b67cea} /* (6, 16, 25) {real, imag} */,
  {32'h3e981170, 32'h4184b9bd} /* (6, 16, 24) {real, imag} */,
  {32'hc0d38b17, 32'hc1118f54} /* (6, 16, 23) {real, imag} */,
  {32'h4101e50c, 32'hc0f14794} /* (6, 16, 22) {real, imag} */,
  {32'hbefaad38, 32'h41069a4b} /* (6, 16, 21) {real, imag} */,
  {32'h4098b88b, 32'h409505bc} /* (6, 16, 20) {real, imag} */,
  {32'h40dc9502, 32'hc100211a} /* (6, 16, 19) {real, imag} */,
  {32'h4153fafc, 32'hc12a6044} /* (6, 16, 18) {real, imag} */,
  {32'hc03d87f6, 32'h415e7e4a} /* (6, 16, 17) {real, imag} */,
  {32'hc103e90f, 32'h00000000} /* (6, 16, 16) {real, imag} */,
  {32'hc03d87f6, 32'hc15e7e4a} /* (6, 16, 15) {real, imag} */,
  {32'h4153fafc, 32'h412a6044} /* (6, 16, 14) {real, imag} */,
  {32'h40dc9502, 32'h4100211a} /* (6, 16, 13) {real, imag} */,
  {32'h4098b88b, 32'hc09505bc} /* (6, 16, 12) {real, imag} */,
  {32'hbefaad38, 32'hc1069a4b} /* (6, 16, 11) {real, imag} */,
  {32'h4101e50c, 32'h40f14794} /* (6, 16, 10) {real, imag} */,
  {32'hc0d38b17, 32'h41118f54} /* (6, 16, 9) {real, imag} */,
  {32'h3e981170, 32'hc184b9bd} /* (6, 16, 8) {real, imag} */,
  {32'h4105dc86, 32'hc0b67cea} /* (6, 16, 7) {real, imag} */,
  {32'h40bc0cbc, 32'hbf824932} /* (6, 16, 6) {real, imag} */,
  {32'hc12c5cc6, 32'hc097071e} /* (6, 16, 5) {real, imag} */,
  {32'hc1317221, 32'hc0929320} /* (6, 16, 4) {real, imag} */,
  {32'hc0790023, 32'hc01a2dfe} /* (6, 16, 3) {real, imag} */,
  {32'hc097d354, 32'hc06395a8} /* (6, 16, 2) {real, imag} */,
  {32'h410eb71d, 32'hc10e33a8} /* (6, 16, 1) {real, imag} */,
  {32'h413e759d, 32'h00000000} /* (6, 16, 0) {real, imag} */,
  {32'hc04c4072, 32'h40fea9b8} /* (6, 15, 31) {real, imag} */,
  {32'h3fd9a640, 32'h403aa65e} /* (6, 15, 30) {real, imag} */,
  {32'h41100784, 32'hc051e196} /* (6, 15, 29) {real, imag} */,
  {32'hc0c64bdc, 32'h40dec928} /* (6, 15, 28) {real, imag} */,
  {32'hc0ae1419, 32'h409b375b} /* (6, 15, 27) {real, imag} */,
  {32'hbecce680, 32'h4057daca} /* (6, 15, 26) {real, imag} */,
  {32'hc141223e, 32'hc1334b8d} /* (6, 15, 25) {real, imag} */,
  {32'hc1001617, 32'h4003cee5} /* (6, 15, 24) {real, imag} */,
  {32'hc109a6a4, 32'h4163382c} /* (6, 15, 23) {real, imag} */,
  {32'hc121d247, 32'h400cf674} /* (6, 15, 22) {real, imag} */,
  {32'hc12fa412, 32'hbec4f178} /* (6, 15, 21) {real, imag} */,
  {32'hc08f6dd6, 32'hc0cbf2c2} /* (6, 15, 20) {real, imag} */,
  {32'h40fb13e4, 32'h3f647030} /* (6, 15, 19) {real, imag} */,
  {32'h402b3009, 32'hc14146c8} /* (6, 15, 18) {real, imag} */,
  {32'hc073b8c2, 32'hc0938784} /* (6, 15, 17) {real, imag} */,
  {32'h400f7799, 32'h40e72008} /* (6, 15, 16) {real, imag} */,
  {32'h404c515f, 32'h400277d0} /* (6, 15, 15) {real, imag} */,
  {32'hc0bd0bb8, 32'h3d4e8880} /* (6, 15, 14) {real, imag} */,
  {32'hbfce231a, 32'hbf6105f4} /* (6, 15, 13) {real, imag} */,
  {32'h41dbac1c, 32'h40bf0a02} /* (6, 15, 12) {real, imag} */,
  {32'h3ea01520, 32'h408c7cb5} /* (6, 15, 11) {real, imag} */,
  {32'h408bcedd, 32'hc0c5db8e} /* (6, 15, 10) {real, imag} */,
  {32'hc0e0568a, 32'h405488be} /* (6, 15, 9) {real, imag} */,
  {32'h407092c6, 32'h3ffb747f} /* (6, 15, 8) {real, imag} */,
  {32'h3fd2125a, 32'h40e89ea9} /* (6, 15, 7) {real, imag} */,
  {32'h3f8e4ec7, 32'hc09f85e6} /* (6, 15, 6) {real, imag} */,
  {32'hc0a32944, 32'h40f6c924} /* (6, 15, 5) {real, imag} */,
  {32'hc053b349, 32'hc134afaa} /* (6, 15, 4) {real, imag} */,
  {32'hbf828770, 32'h409f5162} /* (6, 15, 3) {real, imag} */,
  {32'hbe73d8ac, 32'hc103ae97} /* (6, 15, 2) {real, imag} */,
  {32'h419afcd5, 32'h40587615} /* (6, 15, 1) {real, imag} */,
  {32'h40bc5de9, 32'h4185407f} /* (6, 15, 0) {real, imag} */,
  {32'h4145b862, 32'hc1e842cb} /* (6, 14, 31) {real, imag} */,
  {32'hc0a6fa77, 32'h410f1400} /* (6, 14, 30) {real, imag} */,
  {32'h40898c6c, 32'h4153724e} /* (6, 14, 29) {real, imag} */,
  {32'h3fae7a76, 32'h41030567} /* (6, 14, 28) {real, imag} */,
  {32'h4007038a, 32'h40d5fa26} /* (6, 14, 27) {real, imag} */,
  {32'hbdb19e80, 32'h4093b5b0} /* (6, 14, 26) {real, imag} */,
  {32'hc1678cb6, 32'hbf98e298} /* (6, 14, 25) {real, imag} */,
  {32'hc15e746a, 32'hc1a4235c} /* (6, 14, 24) {real, imag} */,
  {32'hc1237c36, 32'hc15ae775} /* (6, 14, 23) {real, imag} */,
  {32'hc1934589, 32'hc16066d4} /* (6, 14, 22) {real, imag} */,
  {32'h4101cbd8, 32'hbeff4a1c} /* (6, 14, 21) {real, imag} */,
  {32'h40a5dc33, 32'h41b35d1c} /* (6, 14, 20) {real, imag} */,
  {32'hc0c4d74e, 32'hc135534a} /* (6, 14, 19) {real, imag} */,
  {32'h412f5613, 32'hc0fa4688} /* (6, 14, 18) {real, imag} */,
  {32'hc1075ab4, 32'h40c83d84} /* (6, 14, 17) {real, imag} */,
  {32'hc0eba45d, 32'h4066018d} /* (6, 14, 16) {real, imag} */,
  {32'h41124ea5, 32'h410982cb} /* (6, 14, 15) {real, imag} */,
  {32'h40721caa, 32'h4104c775} /* (6, 14, 14) {real, imag} */,
  {32'h40d4d026, 32'hc0a1ca1a} /* (6, 14, 13) {real, imag} */,
  {32'hbf8fee60, 32'h3fad7970} /* (6, 14, 12) {real, imag} */,
  {32'hc1f1a9d2, 32'h3c459c00} /* (6, 14, 11) {real, imag} */,
  {32'h41725a54, 32'h40a3eecb} /* (6, 14, 10) {real, imag} */,
  {32'h409bb96e, 32'hc0430c34} /* (6, 14, 9) {real, imag} */,
  {32'hc1041503, 32'hbea78f8c} /* (6, 14, 8) {real, imag} */,
  {32'hc122c903, 32'h4106e040} /* (6, 14, 7) {real, imag} */,
  {32'hc07251f1, 32'h415c36ab} /* (6, 14, 6) {real, imag} */,
  {32'hbf8f22ca, 32'h4152e9de} /* (6, 14, 5) {real, imag} */,
  {32'hc11108cd, 32'hbf9482fe} /* (6, 14, 4) {real, imag} */,
  {32'h410e9177, 32'h4006d5e0} /* (6, 14, 3) {real, imag} */,
  {32'h414ac3cd, 32'h40a5643b} /* (6, 14, 2) {real, imag} */,
  {32'hc102f185, 32'hbec0a250} /* (6, 14, 1) {real, imag} */,
  {32'hbfd4305a, 32'hc0b3f654} /* (6, 14, 0) {real, imag} */,
  {32'hbfc8976c, 32'hc1924165} /* (6, 13, 31) {real, imag} */,
  {32'hc0d5c405, 32'h3d676e00} /* (6, 13, 30) {real, imag} */,
  {32'h410a05fc, 32'h40d77f42} /* (6, 13, 29) {real, imag} */,
  {32'hc01f39d6, 32'hc0960674} /* (6, 13, 28) {real, imag} */,
  {32'hc1683e9e, 32'hbfe0d5c8} /* (6, 13, 27) {real, imag} */,
  {32'hbf271a80, 32'h3de47d20} /* (6, 13, 26) {real, imag} */,
  {32'h412cc9fc, 32'h401f30b1} /* (6, 13, 25) {real, imag} */,
  {32'h3ff4bdd2, 32'h40c4d71c} /* (6, 13, 24) {real, imag} */,
  {32'h404007ec, 32'hc103fdcd} /* (6, 13, 23) {real, imag} */,
  {32'h412f4f85, 32'hc1147e7c} /* (6, 13, 22) {real, imag} */,
  {32'hc0945755, 32'h40b824ad} /* (6, 13, 21) {real, imag} */,
  {32'hc1600398, 32'hc09adec6} /* (6, 13, 20) {real, imag} */,
  {32'h40db5c0c, 32'hc15388e0} /* (6, 13, 19) {real, imag} */,
  {32'hc090d9d0, 32'h40b59d22} /* (6, 13, 18) {real, imag} */,
  {32'h404a2956, 32'h3df4d020} /* (6, 13, 17) {real, imag} */,
  {32'h3fc23c69, 32'h408b07aa} /* (6, 13, 16) {real, imag} */,
  {32'hc032cf15, 32'hc15acb83} /* (6, 13, 15) {real, imag} */,
  {32'h403f30cc, 32'h400aa9ac} /* (6, 13, 14) {real, imag} */,
  {32'hc155dff2, 32'h41254b22} /* (6, 13, 13) {real, imag} */,
  {32'h40cfd7c7, 32'hc03f0d94} /* (6, 13, 12) {real, imag} */,
  {32'hc0031afc, 32'h411b34a4} /* (6, 13, 11) {real, imag} */,
  {32'hc08332c3, 32'hc0b2fdd0} /* (6, 13, 10) {real, imag} */,
  {32'hc1891b2a, 32'hc01233cc} /* (6, 13, 9) {real, imag} */,
  {32'h40f53082, 32'h416f2f3c} /* (6, 13, 8) {real, imag} */,
  {32'hc125e8ff, 32'h41073b4c} /* (6, 13, 7) {real, imag} */,
  {32'h4185fd17, 32'hc0965e2c} /* (6, 13, 6) {real, imag} */,
  {32'h40eb2508, 32'hbe4e38c0} /* (6, 13, 5) {real, imag} */,
  {32'hbe9da860, 32'h40c62b30} /* (6, 13, 4) {real, imag} */,
  {32'hbed7e720, 32'hbf8de098} /* (6, 13, 3) {real, imag} */,
  {32'h40ee07ef, 32'hc15b1e67} /* (6, 13, 2) {real, imag} */,
  {32'h410dbce0, 32'h41636ef1} /* (6, 13, 1) {real, imag} */,
  {32'h40ba8ad4, 32'h41770261} /* (6, 13, 0) {real, imag} */,
  {32'h41165b8e, 32'hc112a665} /* (6, 12, 31) {real, imag} */,
  {32'hc055bb68, 32'hc095d054} /* (6, 12, 30) {real, imag} */,
  {32'hbddb9980, 32'hbfa447c0} /* (6, 12, 29) {real, imag} */,
  {32'h40bae797, 32'hc12b363d} /* (6, 12, 28) {real, imag} */,
  {32'h412be18c, 32'h3fafa3a8} /* (6, 12, 27) {real, imag} */,
  {32'h40c481cd, 32'h410256d8} /* (6, 12, 26) {real, imag} */,
  {32'hc15f9120, 32'h41169f67} /* (6, 12, 25) {real, imag} */,
  {32'hc0f84860, 32'hc090cdfb} /* (6, 12, 24) {real, imag} */,
  {32'h40b121b8, 32'hc0dc1c5f} /* (6, 12, 23) {real, imag} */,
  {32'h40a94351, 32'h408f4ea8} /* (6, 12, 22) {real, imag} */,
  {32'h41344244, 32'h40a11ca6} /* (6, 12, 21) {real, imag} */,
  {32'hbfe5cd34, 32'hc1653052} /* (6, 12, 20) {real, imag} */,
  {32'h40c1eb62, 32'h41516cb2} /* (6, 12, 19) {real, imag} */,
  {32'h40994d21, 32'hbff5cf3a} /* (6, 12, 18) {real, imag} */,
  {32'h4119cc85, 32'hc0f3e896} /* (6, 12, 17) {real, imag} */,
  {32'hbf8ddca4, 32'h40d7546a} /* (6, 12, 16) {real, imag} */,
  {32'h408d8432, 32'h418a4295} /* (6, 12, 15) {real, imag} */,
  {32'hc1397bd8, 32'h3f92bcd6} /* (6, 12, 14) {real, imag} */,
  {32'h40da52e5, 32'hc14b18c0} /* (6, 12, 13) {real, imag} */,
  {32'h40155a42, 32'hc1743535} /* (6, 12, 12) {real, imag} */,
  {32'hc0dcd7bf, 32'h3f2734b8} /* (6, 12, 11) {real, imag} */,
  {32'hc17ec0df, 32'h3f8e52d4} /* (6, 12, 10) {real, imag} */,
  {32'h410747b1, 32'h412769fc} /* (6, 12, 9) {real, imag} */,
  {32'h40d67a64, 32'h416d9831} /* (6, 12, 8) {real, imag} */,
  {32'h414a39c4, 32'hc0188ce8} /* (6, 12, 7) {real, imag} */,
  {32'hc0abe016, 32'h40ec3316} /* (6, 12, 6) {real, imag} */,
  {32'h3f0d16a8, 32'h40a30e64} /* (6, 12, 5) {real, imag} */,
  {32'h40ff155f, 32'h4031dc27} /* (6, 12, 4) {real, imag} */,
  {32'hc183f567, 32'h402882c2} /* (6, 12, 3) {real, imag} */,
  {32'hbf8fc158, 32'h409d2c56} /* (6, 12, 2) {real, imag} */,
  {32'hc0ced62d, 32'hc15aa48c} /* (6, 12, 1) {real, imag} */,
  {32'hc0b82c6d, 32'h412ff3fb} /* (6, 12, 0) {real, imag} */,
  {32'hc134a1f9, 32'hc19a9502} /* (6, 11, 31) {real, imag} */,
  {32'h40a4a528, 32'h40eb88ba} /* (6, 11, 30) {real, imag} */,
  {32'hc036736e, 32'h4048e4e8} /* (6, 11, 29) {real, imag} */,
  {32'hc032f47c, 32'hc0ae7080} /* (6, 11, 28) {real, imag} */,
  {32'hc06da93c, 32'h4033c00e} /* (6, 11, 27) {real, imag} */,
  {32'h411140fd, 32'hc1148570} /* (6, 11, 26) {real, imag} */,
  {32'h411fa7ec, 32'hc12b5800} /* (6, 11, 25) {real, imag} */,
  {32'h4148ac3c, 32'h408fe6e7} /* (6, 11, 24) {real, imag} */,
  {32'h4140c697, 32'h40d0aa52} /* (6, 11, 23) {real, imag} */,
  {32'hc0f38ee1, 32'h414b77a8} /* (6, 11, 22) {real, imag} */,
  {32'hc10fefee, 32'h41afe4c0} /* (6, 11, 21) {real, imag} */,
  {32'hc0be7283, 32'h4045ff8a} /* (6, 11, 20) {real, imag} */,
  {32'h41233bdf, 32'hc1ad7946} /* (6, 11, 19) {real, imag} */,
  {32'hc087e2a4, 32'hc019176c} /* (6, 11, 18) {real, imag} */,
  {32'hc0c458a1, 32'hbf39c6b0} /* (6, 11, 17) {real, imag} */,
  {32'hc0244595, 32'h3f8ce07c} /* (6, 11, 16) {real, imag} */,
  {32'hbc99d200, 32'h41545cfa} /* (6, 11, 15) {real, imag} */,
  {32'hc0a2462e, 32'h4039feb3} /* (6, 11, 14) {real, imag} */,
  {32'h40cfae3a, 32'h4152e5a7} /* (6, 11, 13) {real, imag} */,
  {32'h41882813, 32'h40267abe} /* (6, 11, 12) {real, imag} */,
  {32'hc11b0f5c, 32'h3ed76300} /* (6, 11, 11) {real, imag} */,
  {32'hc09024b4, 32'hc183142c} /* (6, 11, 10) {real, imag} */,
  {32'hbf97ae9e, 32'hc197bedd} /* (6, 11, 9) {real, imag} */,
  {32'hc0b5955e, 32'h415e14a7} /* (6, 11, 8) {real, imag} */,
  {32'hc148d70a, 32'hc11404d3} /* (6, 11, 7) {real, imag} */,
  {32'hc091a11d, 32'hc10557e7} /* (6, 11, 6) {real, imag} */,
  {32'h40d2859e, 32'hbf147108} /* (6, 11, 5) {real, imag} */,
  {32'hc11fdb73, 32'h419a6a70} /* (6, 11, 4) {real, imag} */,
  {32'hc0ff92cc, 32'h413646dc} /* (6, 11, 3) {real, imag} */,
  {32'hc059996d, 32'h41dbeb42} /* (6, 11, 2) {real, imag} */,
  {32'hbfb7f768, 32'hc1edb7e6} /* (6, 11, 1) {real, imag} */,
  {32'h4147da22, 32'hc121e9e4} /* (6, 11, 0) {real, imag} */,
  {32'hc19044d4, 32'h40e5fece} /* (6, 10, 31) {real, imag} */,
  {32'hc0e45c46, 32'hc1f184d0} /* (6, 10, 30) {real, imag} */,
  {32'hc0af7e17, 32'hc1a69520} /* (6, 10, 29) {real, imag} */,
  {32'h414bc55e, 32'h3e8f17b4} /* (6, 10, 28) {real, imag} */,
  {32'h3fc65e04, 32'h3fb74894} /* (6, 10, 27) {real, imag} */,
  {32'h4167e346, 32'hc1731b00} /* (6, 10, 26) {real, imag} */,
  {32'h400ca2ac, 32'h4055916a} /* (6, 10, 25) {real, imag} */,
  {32'h40ccce45, 32'hc1572acc} /* (6, 10, 24) {real, imag} */,
  {32'h4049d454, 32'hbfc5b920} /* (6, 10, 23) {real, imag} */,
  {32'h3feeeaf8, 32'h41b229a6} /* (6, 10, 22) {real, imag} */,
  {32'hc0c24b6a, 32'hc14adcae} /* (6, 10, 21) {real, imag} */,
  {32'hc082e346, 32'hc0ae9ec9} /* (6, 10, 20) {real, imag} */,
  {32'hc1039fa8, 32'h40a24a5a} /* (6, 10, 19) {real, imag} */,
  {32'hc0fdd2f2, 32'h3f3bf0f0} /* (6, 10, 18) {real, imag} */,
  {32'h4111f71c, 32'h3cd57e40} /* (6, 10, 17) {real, imag} */,
  {32'hc0c44769, 32'hc0f00cda} /* (6, 10, 16) {real, imag} */,
  {32'hbff339b6, 32'h40d49d4b} /* (6, 10, 15) {real, imag} */,
  {32'h4126951e, 32'h41a780e8} /* (6, 10, 14) {real, imag} */,
  {32'hc18d9cce, 32'h410925aa} /* (6, 10, 13) {real, imag} */,
  {32'hc09ec6ba, 32'h40e1c4a4} /* (6, 10, 12) {real, imag} */,
  {32'h417500b2, 32'hc1333171} /* (6, 10, 11) {real, imag} */,
  {32'hc1ad4f58, 32'h41c63174} /* (6, 10, 10) {real, imag} */,
  {32'hc17c7dad, 32'hc1acf84a} /* (6, 10, 9) {real, imag} */,
  {32'h4131462a, 32'hc17306be} /* (6, 10, 8) {real, imag} */,
  {32'h4158df24, 32'h40b0fc8a} /* (6, 10, 7) {real, imag} */,
  {32'h3f05f5f0, 32'h413e755f} /* (6, 10, 6) {real, imag} */,
  {32'h40cab31c, 32'hc115d26b} /* (6, 10, 5) {real, imag} */,
  {32'hbf956669, 32'h408e48ca} /* (6, 10, 4) {real, imag} */,
  {32'hc180027c, 32'h40307a14} /* (6, 10, 3) {real, imag} */,
  {32'hc15515e8, 32'hc1cd9bfa} /* (6, 10, 2) {real, imag} */,
  {32'h418ff111, 32'hc0d1efee} /* (6, 10, 1) {real, imag} */,
  {32'hc12071da, 32'h4206e6e9} /* (6, 10, 0) {real, imag} */,
  {32'hc0291446, 32'h41d60dc0} /* (6, 9, 31) {real, imag} */,
  {32'h3e63eb40, 32'h40deb6b6} /* (6, 9, 30) {real, imag} */,
  {32'hc14487f8, 32'hc1668f96} /* (6, 9, 29) {real, imag} */,
  {32'hc053a2d6, 32'h418db652} /* (6, 9, 28) {real, imag} */,
  {32'hbfc946c6, 32'h40f8137a} /* (6, 9, 27) {real, imag} */,
  {32'hc05b1b77, 32'hc17a202d} /* (6, 9, 26) {real, imag} */,
  {32'hbf402e40, 32'h41156fd3} /* (6, 9, 25) {real, imag} */,
  {32'hc085a6f4, 32'h416e75a0} /* (6, 9, 24) {real, imag} */,
  {32'h3fe528c9, 32'h404538a4} /* (6, 9, 23) {real, imag} */,
  {32'hc091229d, 32'hc11b054f} /* (6, 9, 22) {real, imag} */,
  {32'h40646ef2, 32'hc14b4c3a} /* (6, 9, 21) {real, imag} */,
  {32'h4166138f, 32'h41cecede} /* (6, 9, 20) {real, imag} */,
  {32'hc1eed2e7, 32'h41852710} /* (6, 9, 19) {real, imag} */,
  {32'h410fcd0c, 32'hbf7701e0} /* (6, 9, 18) {real, imag} */,
  {32'hc0a7da75, 32'h4180523f} /* (6, 9, 17) {real, imag} */,
  {32'hbfe1fe60, 32'h406d0371} /* (6, 9, 16) {real, imag} */,
  {32'hc1671edd, 32'h40da9202} /* (6, 9, 15) {real, imag} */,
  {32'hbfa013cc, 32'h3f953b81} /* (6, 9, 14) {real, imag} */,
  {32'hbeee6230, 32'h40e2c92f} /* (6, 9, 13) {real, imag} */,
  {32'hbf4b9760, 32'h410be03e} /* (6, 9, 12) {real, imag} */,
  {32'hc0b52fd7, 32'hbfc31454} /* (6, 9, 11) {real, imag} */,
  {32'hc0239f27, 32'hc2335d9a} /* (6, 9, 10) {real, imag} */,
  {32'h410a5192, 32'h41909d0d} /* (6, 9, 9) {real, imag} */,
  {32'h40d4b958, 32'h3f9a0578} /* (6, 9, 8) {real, imag} */,
  {32'h4180addf, 32'hbfba01c8} /* (6, 9, 7) {real, imag} */,
  {32'h410a79d8, 32'h40d0e5e9} /* (6, 9, 6) {real, imag} */,
  {32'h41408947, 32'hbf75cf70} /* (6, 9, 5) {real, imag} */,
  {32'hc09a39c2, 32'hc1881570} /* (6, 9, 4) {real, imag} */,
  {32'h41dc493b, 32'h4108a96e} /* (6, 9, 3) {real, imag} */,
  {32'hc077f940, 32'hc19459c4} /* (6, 9, 2) {real, imag} */,
  {32'h3f4e5bf4, 32'h409c9553} /* (6, 9, 1) {real, imag} */,
  {32'hc1410ec0, 32'h4192713c} /* (6, 9, 0) {real, imag} */,
  {32'hc1f0afaa, 32'hc1a2f0a1} /* (6, 8, 31) {real, imag} */,
  {32'h4199af10, 32'h4070a2e7} /* (6, 8, 30) {real, imag} */,
  {32'h4150e104, 32'h41ac9af2} /* (6, 8, 29) {real, imag} */,
  {32'hc1ac51df, 32'h4191b442} /* (6, 8, 28) {real, imag} */,
  {32'h41b9e2a0, 32'hc16b7a88} /* (6, 8, 27) {real, imag} */,
  {32'h3fd7a6c8, 32'hc08c094a} /* (6, 8, 26) {real, imag} */,
  {32'hbe4be340, 32'hc1363465} /* (6, 8, 25) {real, imag} */,
  {32'h4132582e, 32'hc11dcacc} /* (6, 8, 24) {real, imag} */,
  {32'h41137530, 32'h400adae6} /* (6, 8, 23) {real, imag} */,
  {32'hc07d1440, 32'h40da7b1a} /* (6, 8, 22) {real, imag} */,
  {32'h4152de4a, 32'h40b76523} /* (6, 8, 21) {real, imag} */,
  {32'hc104844e, 32'hc048abd2} /* (6, 8, 20) {real, imag} */,
  {32'h40a3beff, 32'h407827ee} /* (6, 8, 19) {real, imag} */,
  {32'hc00644c8, 32'hc030405b} /* (6, 8, 18) {real, imag} */,
  {32'hc0ff0707, 32'h3e9366a0} /* (6, 8, 17) {real, imag} */,
  {32'h40ecc261, 32'h410837df} /* (6, 8, 16) {real, imag} */,
  {32'h412793e2, 32'h411f2b87} /* (6, 8, 15) {real, imag} */,
  {32'h4095d88f, 32'hc1324ddb} /* (6, 8, 14) {real, imag} */,
  {32'h40a9b190, 32'hbfb7515a} /* (6, 8, 13) {real, imag} */,
  {32'h3f38a91e, 32'h413eaca8} /* (6, 8, 12) {real, imag} */,
  {32'h411a4d44, 32'h40f0dc23} /* (6, 8, 11) {real, imag} */,
  {32'hc0aef400, 32'hbd9cf000} /* (6, 8, 10) {real, imag} */,
  {32'hc1828819, 32'h4188bd20} /* (6, 8, 9) {real, imag} */,
  {32'hc00591a4, 32'h418a90ec} /* (6, 8, 8) {real, imag} */,
  {32'h409c97c8, 32'h4043b98c} /* (6, 8, 7) {real, imag} */,
  {32'hc1c2933c, 32'h40361ffd} /* (6, 8, 6) {real, imag} */,
  {32'hc1870efe, 32'h40c3ea96} /* (6, 8, 5) {real, imag} */,
  {32'hc1568347, 32'hc17c68f3} /* (6, 8, 4) {real, imag} */,
  {32'h3fd28dc0, 32'h40d77852} /* (6, 8, 3) {real, imag} */,
  {32'h41edbb79, 32'h4124b57d} /* (6, 8, 2) {real, imag} */,
  {32'hc1e94d0c, 32'hc1c80658} /* (6, 8, 1) {real, imag} */,
  {32'hc1f2cf56, 32'hc207d76e} /* (6, 8, 0) {real, imag} */,
  {32'h4188278e, 32'h419b5262} /* (6, 7, 31) {real, imag} */,
  {32'hc01232a4, 32'h417ade4b} /* (6, 7, 30) {real, imag} */,
  {32'hc17274f6, 32'h416590e5} /* (6, 7, 29) {real, imag} */,
  {32'hc1d6b4e8, 32'hc081b000} /* (6, 7, 28) {real, imag} */,
  {32'hc003be64, 32'h4192afb1} /* (6, 7, 27) {real, imag} */,
  {32'hc1a23f48, 32'hbef113c0} /* (6, 7, 26) {real, imag} */,
  {32'h4129dc72, 32'hc1ae2f00} /* (6, 7, 25) {real, imag} */,
  {32'h40aa2e4a, 32'hbfcc0168} /* (6, 7, 24) {real, imag} */,
  {32'hc15c88d2, 32'h40644d00} /* (6, 7, 23) {real, imag} */,
  {32'hc0e106c7, 32'h41ccfa39} /* (6, 7, 22) {real, imag} */,
  {32'h40feebc2, 32'h3fe92808} /* (6, 7, 21) {real, imag} */,
  {32'hc083e732, 32'hc12979fe} /* (6, 7, 20) {real, imag} */,
  {32'hc168c74a, 32'h413da0e6} /* (6, 7, 19) {real, imag} */,
  {32'h40034462, 32'hc18c8496} /* (6, 7, 18) {real, imag} */,
  {32'hbf14f88a, 32'hc0d173dc} /* (6, 7, 17) {real, imag} */,
  {32'hc1772f22, 32'hc00f89d1} /* (6, 7, 16) {real, imag} */,
  {32'hc14cd932, 32'h40d119ce} /* (6, 7, 15) {real, imag} */,
  {32'h41048564, 32'hbfd62005} /* (6, 7, 14) {real, imag} */,
  {32'h410b6d3c, 32'h400215d1} /* (6, 7, 13) {real, imag} */,
  {32'hbf411de0, 32'hc087f729} /* (6, 7, 12) {real, imag} */,
  {32'hc096216c, 32'hc065748e} /* (6, 7, 11) {real, imag} */,
  {32'h3f627ac0, 32'hc09385b9} /* (6, 7, 10) {real, imag} */,
  {32'h41980028, 32'h3fea490c} /* (6, 7, 9) {real, imag} */,
  {32'hc07de2d2, 32'h40f0d761} /* (6, 7, 8) {real, imag} */,
  {32'hbfac60c8, 32'h40b31cb9} /* (6, 7, 7) {real, imag} */,
  {32'h41c3ecb4, 32'h40b2e572} /* (6, 7, 6) {real, imag} */,
  {32'h41530722, 32'hc075e6c2} /* (6, 7, 5) {real, imag} */,
  {32'h41996716, 32'h415f5b22} /* (6, 7, 4) {real, imag} */,
  {32'h3fb921c8, 32'h4128c78a} /* (6, 7, 3) {real, imag} */,
  {32'h40ae506c, 32'hc1a5af8c} /* (6, 7, 2) {real, imag} */,
  {32'hc0a5e802, 32'h41aa930f} /* (6, 7, 1) {real, imag} */,
  {32'h40ff5802, 32'hc0708bed} /* (6, 7, 0) {real, imag} */,
  {32'h4147d0d2, 32'h41bdc1ec} /* (6, 6, 31) {real, imag} */,
  {32'hc15a9cf6, 32'hc19195f0} /* (6, 6, 30) {real, imag} */,
  {32'hc118f380, 32'h405ae2c4} /* (6, 6, 29) {real, imag} */,
  {32'h40f47737, 32'hc0f202ba} /* (6, 6, 28) {real, imag} */,
  {32'hbfb6bffc, 32'h40f7c3e6} /* (6, 6, 27) {real, imag} */,
  {32'h41853e5a, 32'hc122980e} /* (6, 6, 26) {real, imag} */,
  {32'h410cc555, 32'h41858720} /* (6, 6, 25) {real, imag} */,
  {32'hbf821c32, 32'hbfa00d60} /* (6, 6, 24) {real, imag} */,
  {32'hc00b0936, 32'hc18a3c23} /* (6, 6, 23) {real, imag} */,
  {32'h4093aefc, 32'h404c3652} /* (6, 6, 22) {real, imag} */,
  {32'hc15e5b16, 32'hc108b3ef} /* (6, 6, 21) {real, imag} */,
  {32'h3f8cbbc6, 32'h40287c12} /* (6, 6, 20) {real, imag} */,
  {32'hc105bcb2, 32'hc1ac5708} /* (6, 6, 19) {real, imag} */,
  {32'h408ed292, 32'h41261958} /* (6, 6, 18) {real, imag} */,
  {32'hc1a2b1f6, 32'hc1707c04} /* (6, 6, 17) {real, imag} */,
  {32'hbfb2243c, 32'h400431d0} /* (6, 6, 16) {real, imag} */,
  {32'h3ca36900, 32'h4109df2c} /* (6, 6, 15) {real, imag} */,
  {32'hbfa7852a, 32'hc071f654} /* (6, 6, 14) {real, imag} */,
  {32'hc078291c, 32'hc0ecdc0a} /* (6, 6, 13) {real, imag} */,
  {32'hc089dd10, 32'hc0849a1f} /* (6, 6, 12) {real, imag} */,
  {32'h4155870c, 32'hbf219fd0} /* (6, 6, 11) {real, imag} */,
  {32'h40c7178b, 32'h40d809a2} /* (6, 6, 10) {real, imag} */,
  {32'h404cd7a8, 32'h41c2697a} /* (6, 6, 9) {real, imag} */,
  {32'h3f46d490, 32'h41015a9a} /* (6, 6, 8) {real, imag} */,
  {32'h41c354a0, 32'hc1422846} /* (6, 6, 7) {real, imag} */,
  {32'hbcf91200, 32'h4129fe2c} /* (6, 6, 6) {real, imag} */,
  {32'hc0f52a8c, 32'h415241eb} /* (6, 6, 5) {real, imag} */,
  {32'h411b2dc6, 32'h409521bc} /* (6, 6, 4) {real, imag} */,
  {32'hc1ba26b1, 32'hc19fc4f8} /* (6, 6, 3) {real, imag} */,
  {32'hc2323dbd, 32'h41387a7e} /* (6, 6, 2) {real, imag} */,
  {32'hc1f25449, 32'h41ba5230} /* (6, 6, 1) {real, imag} */,
  {32'h3f76d520, 32'hc1b91890} /* (6, 6, 0) {real, imag} */,
  {32'hc26929f8, 32'h423528e2} /* (6, 5, 31) {real, imag} */,
  {32'h42461b96, 32'h41a59a98} /* (6, 5, 30) {real, imag} */,
  {32'hc19598a2, 32'h40625794} /* (6, 5, 29) {real, imag} */,
  {32'hc21219f4, 32'hc0adb710} /* (6, 5, 28) {real, imag} */,
  {32'h42040590, 32'h41545966} /* (6, 5, 27) {real, imag} */,
  {32'h40a3f8b1, 32'hbffb6f42} /* (6, 5, 26) {real, imag} */,
  {32'hc09b52d6, 32'h40cb9210} /* (6, 5, 25) {real, imag} */,
  {32'hc0f04bf9, 32'h40fa7c4f} /* (6, 5, 24) {real, imag} */,
  {32'h400ebfca, 32'hc08d85e3} /* (6, 5, 23) {real, imag} */,
  {32'hc1762ffc, 32'h41bef540} /* (6, 5, 22) {real, imag} */,
  {32'h40eea60b, 32'hc1da0ec7} /* (6, 5, 21) {real, imag} */,
  {32'h41241177, 32'hc1580c18} /* (6, 5, 20) {real, imag} */,
  {32'hc0626f96, 32'hc13253e6} /* (6, 5, 19) {real, imag} */,
  {32'hbd875d60, 32'hbff046f4} /* (6, 5, 18) {real, imag} */,
  {32'hc0f662e1, 32'h3f8164ac} /* (6, 5, 17) {real, imag} */,
  {32'h3da6b440, 32'hc0dd36f9} /* (6, 5, 16) {real, imag} */,
  {32'h3fc9d02c, 32'hbc8529c0} /* (6, 5, 15) {real, imag} */,
  {32'h3f96ab78, 32'h400f2bf4} /* (6, 5, 14) {real, imag} */,
  {32'h40d7544c, 32'h412b5fde} /* (6, 5, 13) {real, imag} */,
  {32'hc0efae90, 32'hc1be7872} /* (6, 5, 12) {real, imag} */,
  {32'h4130dca6, 32'h4137c138} /* (6, 5, 11) {real, imag} */,
  {32'hc0a42274, 32'h411dfa80} /* (6, 5, 10) {real, imag} */,
  {32'hc118c2e6, 32'hc1091009} /* (6, 5, 9) {real, imag} */,
  {32'h40563eac, 32'hc14bdfd9} /* (6, 5, 8) {real, imag} */,
  {32'hc10bff0d, 32'hc079e8f8} /* (6, 5, 7) {real, imag} */,
  {32'h414310f8, 32'h410564d2} /* (6, 5, 6) {real, imag} */,
  {32'h40033d94, 32'h40f27dc0} /* (6, 5, 5) {real, imag} */,
  {32'hc0b7f7a2, 32'hc12bd8e5} /* (6, 5, 4) {real, imag} */,
  {32'hbdcec240, 32'h414ff8c1} /* (6, 5, 3) {real, imag} */,
  {32'h41eb0e63, 32'h421b3060} /* (6, 5, 2) {real, imag} */,
  {32'hc188b77c, 32'hc2501214} /* (6, 5, 1) {real, imag} */,
  {32'hc25de6d8, 32'hc1e02773} /* (6, 5, 0) {real, imag} */,
  {32'h41171e0e, 32'h425e02ae} /* (6, 4, 31) {real, imag} */,
  {32'hc236af96, 32'hc25036cd} /* (6, 4, 30) {real, imag} */,
  {32'h410e828e, 32'h414496fe} /* (6, 4, 29) {real, imag} */,
  {32'h4139a3ff, 32'hc15341c9} /* (6, 4, 28) {real, imag} */,
  {32'h3ff00f0a, 32'h41444c9e} /* (6, 4, 27) {real, imag} */,
  {32'h400a21b4, 32'hc19ae96e} /* (6, 4, 26) {real, imag} */,
  {32'hc0325355, 32'h4104d2ef} /* (6, 4, 25) {real, imag} */,
  {32'hc1a270ce, 32'hc0e9add8} /* (6, 4, 24) {real, imag} */,
  {32'hc0f96c39, 32'hc089e54c} /* (6, 4, 23) {real, imag} */,
  {32'hc19a3ab7, 32'hbfc14a5a} /* (6, 4, 22) {real, imag} */,
  {32'h4124f472, 32'h3ffdfa78} /* (6, 4, 21) {real, imag} */,
  {32'h4176841e, 32'hbef1e348} /* (6, 4, 20) {real, imag} */,
  {32'hbff049ac, 32'hc06f67c2} /* (6, 4, 19) {real, imag} */,
  {32'h415c3030, 32'hc1433461} /* (6, 4, 18) {real, imag} */,
  {32'h40ed938a, 32'hc05d3a06} /* (6, 4, 17) {real, imag} */,
  {32'hc03ba422, 32'h40c78412} /* (6, 4, 16) {real, imag} */,
  {32'hc0c0b34d, 32'h4119a613} /* (6, 4, 15) {real, imag} */,
  {32'h3f636570, 32'hc1594274} /* (6, 4, 14) {real, imag} */,
  {32'h415482d6, 32'hc1945c59} /* (6, 4, 13) {real, imag} */,
  {32'hbf115ad0, 32'h41c27f36} /* (6, 4, 12) {real, imag} */,
  {32'h3fbfa660, 32'hc0782686} /* (6, 4, 11) {real, imag} */,
  {32'hc1201d00, 32'h4004a154} /* (6, 4, 10) {real, imag} */,
  {32'h41700d3c, 32'hc1513acf} /* (6, 4, 9) {real, imag} */,
  {32'hc1ba7c42, 32'h413384fd} /* (6, 4, 8) {real, imag} */,
  {32'h403eec46, 32'h40032086} /* (6, 4, 7) {real, imag} */,
  {32'hc17ad5f8, 32'h41f05d98} /* (6, 4, 6) {real, imag} */,
  {32'hc18b23d4, 32'hc15f882c} /* (6, 4, 5) {real, imag} */,
  {32'h410935ba, 32'h419139ee} /* (6, 4, 4) {real, imag} */,
  {32'hc10cc302, 32'h40abf7cc} /* (6, 4, 3) {real, imag} */,
  {32'hc25b88d7, 32'hc2463d81} /* (6, 4, 2) {real, imag} */,
  {32'h42694d46, 32'h42922f85} /* (6, 4, 1) {real, imag} */,
  {32'h423ff7ff, 32'hc0e215a8} /* (6, 4, 0) {real, imag} */,
  {32'hc2bb06ef, 32'h41f5c638} /* (6, 3, 31) {real, imag} */,
  {32'h419eac7a, 32'hc2fcaf3a} /* (6, 3, 30) {real, imag} */,
  {32'h40d75f26, 32'hbea30910} /* (6, 3, 29) {real, imag} */,
  {32'h41ce4a34, 32'h41d4a4a1} /* (6, 3, 28) {real, imag} */,
  {32'h409591c0, 32'hc0bfc9e7} /* (6, 3, 27) {real, imag} */,
  {32'hc2112008, 32'h40e65e23} /* (6, 3, 26) {real, imag} */,
  {32'hbf6be0a0, 32'hc115739a} /* (6, 3, 25) {real, imag} */,
  {32'h410637ef, 32'hc1b2ed8c} /* (6, 3, 24) {real, imag} */,
  {32'h410eb618, 32'hc024a6cc} /* (6, 3, 23) {real, imag} */,
  {32'h3ed07750, 32'hc09d62cf} /* (6, 3, 22) {real, imag} */,
  {32'hc11cd648, 32'h4173e68d} /* (6, 3, 21) {real, imag} */,
  {32'hc035145c, 32'h4125aad0} /* (6, 3, 20) {real, imag} */,
  {32'h41a3faa6, 32'h41390170} /* (6, 3, 19) {real, imag} */,
  {32'hbfa6261c, 32'hc09f8920} /* (6, 3, 18) {real, imag} */,
  {32'h41311e3c, 32'h40c84078} /* (6, 3, 17) {real, imag} */,
  {32'hbf4ab9f4, 32'h3fe4e2ca} /* (6, 3, 16) {real, imag} */,
  {32'hc151dd8e, 32'h410c2277} /* (6, 3, 15) {real, imag} */,
  {32'h41cbcf8a, 32'h40bae89a} /* (6, 3, 14) {real, imag} */,
  {32'h4006d394, 32'hc127f34b} /* (6, 3, 13) {real, imag} */,
  {32'hc039026c, 32'hc16a9420} /* (6, 3, 12) {real, imag} */,
  {32'h417ea02c, 32'h3f4fda6c} /* (6, 3, 11) {real, imag} */,
  {32'hc1950e76, 32'h40cfa509} /* (6, 3, 10) {real, imag} */,
  {32'h41948835, 32'h3fa958d0} /* (6, 3, 9) {real, imag} */,
  {32'hc17bed88, 32'hc1999556} /* (6, 3, 8) {real, imag} */,
  {32'hc1218e82, 32'h401f6da6} /* (6, 3, 7) {real, imag} */,
  {32'h402fb600, 32'hc20e3130} /* (6, 3, 6) {real, imag} */,
  {32'h41f5f994, 32'hc1d49451} /* (6, 3, 5) {real, imag} */,
  {32'hc1d1e1ba, 32'h410b9f11} /* (6, 3, 4) {real, imag} */,
  {32'hc1cc68e0, 32'hc13cb546} /* (6, 3, 3) {real, imag} */,
  {32'h40bc4c3c, 32'hc13546da} /* (6, 3, 2) {real, imag} */,
  {32'h42b45df8, 32'h42ed5064} /* (6, 3, 1) {real, imag} */,
  {32'h41c5c137, 32'h4281562d} /* (6, 3, 0) {real, imag} */,
  {32'hc41ffd87, 32'hbfc49930} /* (6, 2, 31) {real, imag} */,
  {32'h43b07012, 32'hc2ac400d} /* (6, 2, 30) {real, imag} */,
  {32'hc2488758, 32'h421287ec} /* (6, 2, 29) {real, imag} */,
  {32'h41094bd4, 32'h41f6120d} /* (6, 2, 28) {real, imag} */,
  {32'h41b08e0d, 32'hc1fc1d8b} /* (6, 2, 27) {real, imag} */,
  {32'h4101b47c, 32'h3f855b60} /* (6, 2, 26) {real, imag} */,
  {32'hc04aef3c, 32'hc116ee08} /* (6, 2, 25) {real, imag} */,
  {32'h422d6493, 32'h41287c6b} /* (6, 2, 24) {real, imag} */,
  {32'hc178c1be, 32'h3f7957e0} /* (6, 2, 23) {real, imag} */,
  {32'h3eb2a800, 32'hc0128536} /* (6, 2, 22) {real, imag} */,
  {32'h40458a1d, 32'hc183d576} /* (6, 2, 21) {real, imag} */,
  {32'h3fc4a074, 32'h414a98a3} /* (6, 2, 20) {real, imag} */,
  {32'h40f990fa, 32'h411849d3} /* (6, 2, 19) {real, imag} */,
  {32'hc1367104, 32'hc148d701} /* (6, 2, 18) {real, imag} */,
  {32'hc050d590, 32'h40568cb6} /* (6, 2, 17) {real, imag} */,
  {32'hbe16e840, 32'hbf6291a8} /* (6, 2, 16) {real, imag} */,
  {32'h403f3712, 32'hc106dd8c} /* (6, 2, 15) {real, imag} */,
  {32'h40b8db14, 32'h4035f704} /* (6, 2, 14) {real, imag} */,
  {32'h40181f1e, 32'hbf7fed15} /* (6, 2, 13) {real, imag} */,
  {32'hc13c19f0, 32'hc0315e10} /* (6, 2, 12) {real, imag} */,
  {32'h412e24dc, 32'h41bdc8dc} /* (6, 2, 11) {real, imag} */,
  {32'h40c7f755, 32'hbfd7fb10} /* (6, 2, 10) {real, imag} */,
  {32'h41430072, 32'h4172c842} /* (6, 2, 9) {real, imag} */,
  {32'h41d86070, 32'h409d26fc} /* (6, 2, 8) {real, imag} */,
  {32'hc096b2b2, 32'hc1831a6c} /* (6, 2, 7) {real, imag} */,
  {32'h40a8c640, 32'h41894c50} /* (6, 2, 6) {real, imag} */,
  {32'h42340b32, 32'h4116e888} /* (6, 2, 5) {real, imag} */,
  {32'hc2ae24a7, 32'hc022a7b0} /* (6, 2, 4) {real, imag} */,
  {32'hc1667c55, 32'h42203d1e} /* (6, 2, 3) {real, imag} */,
  {32'h43587e37, 32'hbfc528c0} /* (6, 2, 2) {real, imag} */,
  {32'hc39ecffa, 32'h42a7fa80} /* (6, 2, 1) {real, imag} */,
  {32'hc3aed24a, 32'hc3125213} /* (6, 2, 0) {real, imag} */,
  {32'h445e82cb, 32'hc37286c0} /* (6, 1, 31) {real, imag} */,
  {32'hc3393089, 32'hbeb45180} /* (6, 1, 30) {real, imag} */,
  {32'h42849d73, 32'hc185217f} /* (6, 1, 29) {real, imag} */,
  {32'h423ed70e, 32'h424619ab} /* (6, 1, 28) {real, imag} */,
  {32'hc2b74f0c, 32'hc1628e0a} /* (6, 1, 27) {real, imag} */,
  {32'h41417d26, 32'h405fc2fa} /* (6, 1, 26) {real, imag} */,
  {32'hc1893dee, 32'hbfb26728} /* (6, 1, 25) {real, imag} */,
  {32'hc1af5090, 32'h40abc1d1} /* (6, 1, 24) {real, imag} */,
  {32'h3fc92f8c, 32'hc164a539} /* (6, 1, 23) {real, imag} */,
  {32'h412f1eac, 32'hc0f3cda2} /* (6, 1, 22) {real, imag} */,
  {32'hc1ab8a8c, 32'h4200b772} /* (6, 1, 21) {real, imag} */,
  {32'h416bc1d6, 32'h40bde156} /* (6, 1, 20) {real, imag} */,
  {32'h401c0e6e, 32'hc1026814} /* (6, 1, 19) {real, imag} */,
  {32'hc1769b04, 32'h40855a8b} /* (6, 1, 18) {real, imag} */,
  {32'h404b5712, 32'h40678f7a} /* (6, 1, 17) {real, imag} */,
  {32'hc0eb0cce, 32'h405e0e18} /* (6, 1, 16) {real, imag} */,
  {32'hc1213968, 32'h4025f118} /* (6, 1, 15) {real, imag} */,
  {32'h410d0e80, 32'hc1807478} /* (6, 1, 14) {real, imag} */,
  {32'h3eafa580, 32'h3fbad3db} /* (6, 1, 13) {real, imag} */,
  {32'hc010ba32, 32'h3fc8daac} /* (6, 1, 12) {real, imag} */,
  {32'hc19db160, 32'hc1be8369} /* (6, 1, 11) {real, imag} */,
  {32'hc11af5bc, 32'hc00c86b1} /* (6, 1, 10) {real, imag} */,
  {32'h412e01e9, 32'hbe0a9480} /* (6, 1, 9) {real, imag} */,
  {32'hc124d526, 32'hc206c0c2} /* (6, 1, 8) {real, imag} */,
  {32'h41c30ac0, 32'h40e26ffa} /* (6, 1, 7) {real, imag} */,
  {32'hc1751b62, 32'hbf9dba94} /* (6, 1, 6) {real, imag} */,
  {32'hc2702b8e, 32'hc118e236} /* (6, 1, 5) {real, imag} */,
  {32'h424182cd, 32'hc1d536de} /* (6, 1, 4) {real, imag} */,
  {32'hc1a575ee, 32'hc287893d} /* (6, 1, 3) {real, imag} */,
  {32'hc3a4e64a, 32'hc39b9bf8} /* (6, 1, 2) {real, imag} */,
  {32'h449cbd4a, 32'h44081355} /* (6, 1, 1) {real, imag} */,
  {32'h449fd30a, 32'h436b3175} /* (6, 1, 0) {real, imag} */,
  {32'h4434b0b3, 32'hc41ddcf1} /* (6, 0, 31) {real, imag} */,
  {32'hc2279c50, 32'h4327e5d8} /* (6, 0, 30) {real, imag} */,
  {32'h4192fde1, 32'hc22c198c} /* (6, 0, 29) {real, imag} */,
  {32'h40206320, 32'hc22aa057} /* (6, 0, 28) {real, imag} */,
  {32'hc21de18c, 32'h418d89e8} /* (6, 0, 27) {real, imag} */,
  {32'h41d0e4d7, 32'h40d7dbc4} /* (6, 0, 26) {real, imag} */,
  {32'h41c8a551, 32'hc21805d5} /* (6, 0, 25) {real, imag} */,
  {32'hc0aad428, 32'h410bf166} /* (6, 0, 24) {real, imag} */,
  {32'hc19e1595, 32'h409ada58} /* (6, 0, 23) {real, imag} */,
  {32'hc06a688c, 32'hc0f98d73} /* (6, 0, 22) {real, imag} */,
  {32'hc1809f9b, 32'h419a9d37} /* (6, 0, 21) {real, imag} */,
  {32'h41042066, 32'hc0d45dd4} /* (6, 0, 20) {real, imag} */,
  {32'h41347180, 32'h417acb18} /* (6, 0, 19) {real, imag} */,
  {32'hc0cc7530, 32'h41684676} /* (6, 0, 18) {real, imag} */,
  {32'hc0184504, 32'h3f7d14f2} /* (6, 0, 17) {real, imag} */,
  {32'h4136c008, 32'h00000000} /* (6, 0, 16) {real, imag} */,
  {32'hc0184504, 32'hbf7d14f2} /* (6, 0, 15) {real, imag} */,
  {32'hc0cc7530, 32'hc1684676} /* (6, 0, 14) {real, imag} */,
  {32'h41347180, 32'hc17acb18} /* (6, 0, 13) {real, imag} */,
  {32'h41042066, 32'h40d45dd4} /* (6, 0, 12) {real, imag} */,
  {32'hc1809f9b, 32'hc19a9d37} /* (6, 0, 11) {real, imag} */,
  {32'hc06a688c, 32'h40f98d73} /* (6, 0, 10) {real, imag} */,
  {32'hc19e1595, 32'hc09ada58} /* (6, 0, 9) {real, imag} */,
  {32'hc0aad428, 32'hc10bf166} /* (6, 0, 8) {real, imag} */,
  {32'h41c8a551, 32'h421805d5} /* (6, 0, 7) {real, imag} */,
  {32'h41d0e4d7, 32'hc0d7dbc4} /* (6, 0, 6) {real, imag} */,
  {32'hc21de18c, 32'hc18d89e8} /* (6, 0, 5) {real, imag} */,
  {32'h40206320, 32'h422aa057} /* (6, 0, 4) {real, imag} */,
  {32'h4192fde1, 32'h422c198c} /* (6, 0, 3) {real, imag} */,
  {32'hc2279c50, 32'hc327e5d8} /* (6, 0, 2) {real, imag} */,
  {32'h4434b0b3, 32'h441ddcf1} /* (6, 0, 1) {real, imag} */,
  {32'h44c34370, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'h43bdb712, 32'hc26e91b4} /* (5, 31, 31) {real, imag} */,
  {32'hc0d733e0, 32'h4160f640} /* (5, 31, 30) {real, imag} */,
  {32'hc10d3652, 32'h425c2658} /* (5, 31, 29) {real, imag} */,
  {32'h41cad6a5, 32'h420f0810} /* (5, 31, 28) {real, imag} */,
  {32'hc12e5fb8, 32'hc1b8a617} /* (5, 31, 27) {real, imag} */,
  {32'hc1aee3e4, 32'h414e317d} /* (5, 31, 26) {real, imag} */,
  {32'hc0a5dcbc, 32'hc1858868} /* (5, 31, 25) {real, imag} */,
  {32'h41da4d77, 32'hc0e83474} /* (5, 31, 24) {real, imag} */,
  {32'hc189c200, 32'hc15b87cb} /* (5, 31, 23) {real, imag} */,
  {32'hc10c54b5, 32'h41238f9a} /* (5, 31, 22) {real, imag} */,
  {32'h41592f8f, 32'h4142139a} /* (5, 31, 21) {real, imag} */,
  {32'h40ce8303, 32'h401a8872} /* (5, 31, 20) {real, imag} */,
  {32'h4123cbba, 32'hc0974527} /* (5, 31, 19) {real, imag} */,
  {32'h41177e17, 32'h4129c5c3} /* (5, 31, 18) {real, imag} */,
  {32'h408d8ff3, 32'hc0af6c15} /* (5, 31, 17) {real, imag} */,
  {32'h40004ef8, 32'h40b29433} /* (5, 31, 16) {real, imag} */,
  {32'h40476a4a, 32'h3eda9ad0} /* (5, 31, 15) {real, imag} */,
  {32'hc08f312c, 32'h4130c575} /* (5, 31, 14) {real, imag} */,
  {32'h4003e909, 32'h410817c7} /* (5, 31, 13) {real, imag} */,
  {32'h40b23de7, 32'h4140ed13} /* (5, 31, 12) {real, imag} */,
  {32'hc10faa5a, 32'hbdddf380} /* (5, 31, 11) {real, imag} */,
  {32'hc072237e, 32'h403cf99a} /* (5, 31, 10) {real, imag} */,
  {32'h4158dd67, 32'h410f8268} /* (5, 31, 9) {real, imag} */,
  {32'h40748864, 32'h41145451} /* (5, 31, 8) {real, imag} */,
  {32'hc22bb13e, 32'h406b6a01} /* (5, 31, 7) {real, imag} */,
  {32'h41162453, 32'h413b854e} /* (5, 31, 6) {real, imag} */,
  {32'h418af44c, 32'hc15f17a4} /* (5, 31, 5) {real, imag} */,
  {32'h40abdf6e, 32'h41bf581d} /* (5, 31, 4) {real, imag} */,
  {32'h42671a97, 32'h41616697} /* (5, 31, 3) {real, imag} */,
  {32'h41b6ace0, 32'h3fa8e240} /* (5, 31, 2) {real, imag} */,
  {32'h4364b078, 32'h42d6416a} /* (5, 31, 1) {real, imag} */,
  {32'h440da16e, 32'hc31b2d54} /* (5, 31, 0) {real, imag} */,
  {32'h41b7f910, 32'hc21e8910} /* (5, 30, 31) {real, imag} */,
  {32'hc26434ce, 32'hc2a33f10} /* (5, 30, 30) {real, imag} */,
  {32'hbf0c5e20, 32'hc0d3845a} /* (5, 30, 29) {real, imag} */,
  {32'h40e9d564, 32'hc1b7755f} /* (5, 30, 28) {real, imag} */,
  {32'h41d7b7b1, 32'h420572b9} /* (5, 30, 27) {real, imag} */,
  {32'h40643a27, 32'hc18aa4ce} /* (5, 30, 26) {real, imag} */,
  {32'hc08e2d9e, 32'h415ad9da} /* (5, 30, 25) {real, imag} */,
  {32'h3fbc7780, 32'h40781028} /* (5, 30, 24) {real, imag} */,
  {32'h408d99a5, 32'hc1f2d973} /* (5, 30, 23) {real, imag} */,
  {32'hc13ba530, 32'hc0a734c4} /* (5, 30, 22) {real, imag} */,
  {32'hc0850fc0, 32'h4105ed4b} /* (5, 30, 21) {real, imag} */,
  {32'h3f893194, 32'h4072a765} /* (5, 30, 20) {real, imag} */,
  {32'hbf7721f6, 32'hbc96c400} /* (5, 30, 19) {real, imag} */,
  {32'h3c983500, 32'h40fa9fd2} /* (5, 30, 18) {real, imag} */,
  {32'hc0e9b948, 32'hc0baa6bc} /* (5, 30, 17) {real, imag} */,
  {32'h40ad36a2, 32'h4077a9c0} /* (5, 30, 16) {real, imag} */,
  {32'h40c89513, 32'h40e6a7aa} /* (5, 30, 15) {real, imag} */,
  {32'hbfc4fca8, 32'h4063166a} /* (5, 30, 14) {real, imag} */,
  {32'hc08a04a7, 32'h416593ee} /* (5, 30, 13) {real, imag} */,
  {32'h415c5e12, 32'hc03bf454} /* (5, 30, 12) {real, imag} */,
  {32'hc0bca46b, 32'hc10931f6} /* (5, 30, 11) {real, imag} */,
  {32'h40322634, 32'h40dd055c} /* (5, 30, 10) {real, imag} */,
  {32'hbf922184, 32'h403564d5} /* (5, 30, 9) {real, imag} */,
  {32'h410a1216, 32'hc217f9fd} /* (5, 30, 8) {real, imag} */,
  {32'h415844fa, 32'h4119bcf4} /* (5, 30, 7) {real, imag} */,
  {32'hc1ddc0ea, 32'hc1a79de6} /* (5, 30, 6) {real, imag} */,
  {32'hc1fbb23d, 32'hc09478f8} /* (5, 30, 5) {real, imag} */,
  {32'h4148cbb6, 32'h41a03f07} /* (5, 30, 4) {real, imag} */,
  {32'h3ee8f2a0, 32'hc1caec4b} /* (5, 30, 3) {real, imag} */,
  {32'h41cc8e18, 32'h4120cfc0} /* (5, 30, 2) {real, imag} */,
  {32'hc133b740, 32'hbfa13220} /* (5, 30, 1) {real, imag} */,
  {32'hc294f34e, 32'h426141c1} /* (5, 30, 0) {real, imag} */,
  {32'h414dc5ec, 32'hc2472d42} /* (5, 29, 31) {real, imag} */,
  {32'h420ccf79, 32'hc28f49d4} /* (5, 29, 30) {real, imag} */,
  {32'hc11be700, 32'hc1304cda} /* (5, 29, 29) {real, imag} */,
  {32'h4119a51e, 32'hc0f2991e} /* (5, 29, 28) {real, imag} */,
  {32'hc139ce16, 32'h412959d8} /* (5, 29, 27) {real, imag} */,
  {32'h3f9133d8, 32'h4189c1ca} /* (5, 29, 26) {real, imag} */,
  {32'hc124e860, 32'h41d88e82} /* (5, 29, 25) {real, imag} */,
  {32'hc0675284, 32'hc168f030} /* (5, 29, 24) {real, imag} */,
  {32'h3ea04300, 32'h40cade51} /* (5, 29, 23) {real, imag} */,
  {32'h40b8ed07, 32'h41035e4b} /* (5, 29, 22) {real, imag} */,
  {32'hc164a6f0, 32'h4184311a} /* (5, 29, 21) {real, imag} */,
  {32'hc0caedd3, 32'h4063fdbc} /* (5, 29, 20) {real, imag} */,
  {32'h4145e166, 32'hc08737b9} /* (5, 29, 19) {real, imag} */,
  {32'h40f27b56, 32'h413bdd81} /* (5, 29, 18) {real, imag} */,
  {32'h413e8ced, 32'h40502368} /* (5, 29, 17) {real, imag} */,
  {32'hc0e3e7d6, 32'h402f8c2e} /* (5, 29, 16) {real, imag} */,
  {32'hc00b5172, 32'hc09722b0} /* (5, 29, 15) {real, imag} */,
  {32'hc04af1af, 32'h40322665} /* (5, 29, 14) {real, imag} */,
  {32'h3fc381a2, 32'hc132229f} /* (5, 29, 13) {real, imag} */,
  {32'h41c25ffc, 32'h3ea4ff00} /* (5, 29, 12) {real, imag} */,
  {32'hc0646820, 32'hc107ea03} /* (5, 29, 11) {real, imag} */,
  {32'hc03ab9b4, 32'h40fd48bf} /* (5, 29, 10) {real, imag} */,
  {32'h417f16f8, 32'h4066b7cc} /* (5, 29, 9) {real, imag} */,
  {32'h41b2f2b8, 32'h4080b4a0} /* (5, 29, 8) {real, imag} */,
  {32'hc148c62a, 32'hc18575b2} /* (5, 29, 7) {real, imag} */,
  {32'hc1d6869f, 32'h40b1d670} /* (5, 29, 6) {real, imag} */,
  {32'hc12280e9, 32'h41a9ae8a} /* (5, 29, 5) {real, imag} */,
  {32'hc147d1a5, 32'hc0685338} /* (5, 29, 4) {real, imag} */,
  {32'h4000ca96, 32'hc165ae72} /* (5, 29, 3) {real, imag} */,
  {32'hc128df48, 32'h42272ee2} /* (5, 29, 2) {real, imag} */,
  {32'h40e66eb8, 32'h42321549} /* (5, 29, 1) {real, imag} */,
  {32'h4180fbc1, 32'hc2502bfb} /* (5, 29, 0) {real, imag} */,
  {32'hc29bb8b4, 32'hc17eec40} /* (5, 28, 31) {real, imag} */,
  {32'h41c95216, 32'h414f0d84} /* (5, 28, 30) {real, imag} */,
  {32'hc1c0fcdb, 32'hc1d55504} /* (5, 28, 29) {real, imag} */,
  {32'h41ac6584, 32'h4057dc70} /* (5, 28, 28) {real, imag} */,
  {32'h412869ff, 32'hc078d2e8} /* (5, 28, 27) {real, imag} */,
  {32'hbff564a8, 32'hc00440a2} /* (5, 28, 26) {real, imag} */,
  {32'hc1a154e8, 32'h401cf48c} /* (5, 28, 25) {real, imag} */,
  {32'h40c286f5, 32'hc15bdea7} /* (5, 28, 24) {real, imag} */,
  {32'hc186559a, 32'h402b3a16} /* (5, 28, 23) {real, imag} */,
  {32'h40b4f5f8, 32'h41c12023} /* (5, 28, 22) {real, imag} */,
  {32'h416c92c8, 32'hc138d52b} /* (5, 28, 21) {real, imag} */,
  {32'hc0f7a766, 32'hc15d9f64} /* (5, 28, 20) {real, imag} */,
  {32'hc17fb710, 32'h40b45d8e} /* (5, 28, 19) {real, imag} */,
  {32'h411636c0, 32'hc17555e4} /* (5, 28, 18) {real, imag} */,
  {32'hbf922ef4, 32'h4005d776} /* (5, 28, 17) {real, imag} */,
  {32'hc0b5a500, 32'hc0c0947a} /* (5, 28, 16) {real, imag} */,
  {32'h40d093aa, 32'hc00f0679} /* (5, 28, 15) {real, imag} */,
  {32'hc1459a7d, 32'hc0ec0dc0} /* (5, 28, 14) {real, imag} */,
  {32'hc10757a0, 32'hc0da7be6} /* (5, 28, 13) {real, imag} */,
  {32'h411c0740, 32'hc1b0f3f4} /* (5, 28, 12) {real, imag} */,
  {32'h411d3956, 32'h4141769a} /* (5, 28, 11) {real, imag} */,
  {32'h40fc4804, 32'hc0613fb9} /* (5, 28, 10) {real, imag} */,
  {32'h409053ae, 32'hc028cc36} /* (5, 28, 9) {real, imag} */,
  {32'h418513a0, 32'h413f80f6} /* (5, 28, 8) {real, imag} */,
  {32'h40833a1c, 32'hc18ca0ee} /* (5, 28, 7) {real, imag} */,
  {32'hc1b3df08, 32'h4123a6f8} /* (5, 28, 6) {real, imag} */,
  {32'h4123e4e8, 32'h41b9a4fa} /* (5, 28, 5) {real, imag} */,
  {32'h404aacb2, 32'hc1838016} /* (5, 28, 4) {real, imag} */,
  {32'h4063e05d, 32'hbed388e0} /* (5, 28, 3) {real, imag} */,
  {32'h40963ce8, 32'hc1cfc354} /* (5, 28, 2) {real, imag} */,
  {32'hc1bdc213, 32'h41da51e3} /* (5, 28, 1) {real, imag} */,
  {32'h416cc939, 32'h419148c0} /* (5, 28, 0) {real, imag} */,
  {32'h41b0f85b, 32'hc0c2a416} /* (5, 27, 31) {real, imag} */,
  {32'hc0335e44, 32'hc1a8c87a} /* (5, 27, 30) {real, imag} */,
  {32'h41921aa2, 32'hc015bdc8} /* (5, 27, 29) {real, imag} */,
  {32'hc1ac5ab0, 32'hc0f5a5a7} /* (5, 27, 28) {real, imag} */,
  {32'hc1a5ea98, 32'hc0b13d60} /* (5, 27, 27) {real, imag} */,
  {32'h4119459e, 32'h40f6ff96} /* (5, 27, 26) {real, imag} */,
  {32'hc1100a19, 32'h409db134} /* (5, 27, 25) {real, imag} */,
  {32'h408314cb, 32'hbf304f04} /* (5, 27, 24) {real, imag} */,
  {32'hc13c02c4, 32'hc06bb5b2} /* (5, 27, 23) {real, imag} */,
  {32'h400bf216, 32'hc18b22d7} /* (5, 27, 22) {real, imag} */,
  {32'h4129aed5, 32'h40e43aae} /* (5, 27, 21) {real, imag} */,
  {32'h4065d141, 32'hbf852890} /* (5, 27, 20) {real, imag} */,
  {32'h4143b0f5, 32'hc172e301} /* (5, 27, 19) {real, imag} */,
  {32'h4110f440, 32'hbfa79ab0} /* (5, 27, 18) {real, imag} */,
  {32'hc0c37a24, 32'hbf4e99d0} /* (5, 27, 17) {real, imag} */,
  {32'h403c5b44, 32'hc00bc834} /* (5, 27, 16) {real, imag} */,
  {32'hbf723f26, 32'h40d8b7c0} /* (5, 27, 15) {real, imag} */,
  {32'hc129bb6a, 32'hbfdc5dd0} /* (5, 27, 14) {real, imag} */,
  {32'hc197544b, 32'hc124f7b0} /* (5, 27, 13) {real, imag} */,
  {32'hc0f9b317, 32'h41242bfc} /* (5, 27, 12) {real, imag} */,
  {32'hc0951511, 32'h41350d00} /* (5, 27, 11) {real, imag} */,
  {32'hc1894323, 32'h41a47f57} /* (5, 27, 10) {real, imag} */,
  {32'hc0e48fd3, 32'hc171ab4c} /* (5, 27, 9) {real, imag} */,
  {32'hc206198c, 32'hc0f13ff4} /* (5, 27, 8) {real, imag} */,
  {32'h408c633e, 32'hc0b357cb} /* (5, 27, 7) {real, imag} */,
  {32'h41043aba, 32'hc19c612a} /* (5, 27, 6) {real, imag} */,
  {32'hc18e1474, 32'hc18cc338} /* (5, 27, 5) {real, imag} */,
  {32'hc1255a2d, 32'h409cb3a8} /* (5, 27, 4) {real, imag} */,
  {32'hc1aa7356, 32'h418ffdd3} /* (5, 27, 3) {real, imag} */,
  {32'hc117236a, 32'h4116ccb4} /* (5, 27, 2) {real, imag} */,
  {32'h41d3eb6e, 32'hc24bbef5} /* (5, 27, 1) {real, imag} */,
  {32'h414555c0, 32'hc13d4a1d} /* (5, 27, 0) {real, imag} */,
  {32'hc0c7c574, 32'hc111f4fc} /* (5, 26, 31) {real, imag} */,
  {32'hc1a7baa6, 32'h41147dc7} /* (5, 26, 30) {real, imag} */,
  {32'hc190c6c7, 32'h41d18a6a} /* (5, 26, 29) {real, imag} */,
  {32'hc076ee08, 32'hc0edf240} /* (5, 26, 28) {real, imag} */,
  {32'hc082b7ec, 32'hc133b206} /* (5, 26, 27) {real, imag} */,
  {32'hc1665fb4, 32'hc15859f0} /* (5, 26, 26) {real, imag} */,
  {32'h41b0b280, 32'hc14b180e} /* (5, 26, 25) {real, imag} */,
  {32'hc16656ca, 32'h411d9254} /* (5, 26, 24) {real, imag} */,
  {32'h403e11b5, 32'h415b7dc6} /* (5, 26, 23) {real, imag} */,
  {32'h4171ac8c, 32'hc0335291} /* (5, 26, 22) {real, imag} */,
  {32'hc0b4b2c8, 32'hc1ca9f41} /* (5, 26, 21) {real, imag} */,
  {32'h41776cf8, 32'h411fda51} /* (5, 26, 20) {real, imag} */,
  {32'hbf6ebc44, 32'hc02115cc} /* (5, 26, 19) {real, imag} */,
  {32'h411e5949, 32'hc110a921} /* (5, 26, 18) {real, imag} */,
  {32'hc0b5093c, 32'h3f1d8fb0} /* (5, 26, 17) {real, imag} */,
  {32'h411d9664, 32'h409e84f9} /* (5, 26, 16) {real, imag} */,
  {32'hc141dec0, 32'h40e73c00} /* (5, 26, 15) {real, imag} */,
  {32'h40da7398, 32'hc0b755c4} /* (5, 26, 14) {real, imag} */,
  {32'h41041f64, 32'hc0ec22ca} /* (5, 26, 13) {real, imag} */,
  {32'hc0b51ba0, 32'h40038da6} /* (5, 26, 12) {real, imag} */,
  {32'hc1128324, 32'h3f922710} /* (5, 26, 11) {real, imag} */,
  {32'hc0c10445, 32'hc11a4a3e} /* (5, 26, 10) {real, imag} */,
  {32'hc1320f12, 32'hc003fec0} /* (5, 26, 9) {real, imag} */,
  {32'hc09a1248, 32'h410a33c2} /* (5, 26, 8) {real, imag} */,
  {32'h3fbe8ef0, 32'hc1bf54c4} /* (5, 26, 7) {real, imag} */,
  {32'hc0d43026, 32'h41228410} /* (5, 26, 6) {real, imag} */,
  {32'h411fd09a, 32'hc11117ca} /* (5, 26, 5) {real, imag} */,
  {32'h40a46f0c, 32'hc048b702} /* (5, 26, 4) {real, imag} */,
  {32'h4159d75c, 32'h407818f2} /* (5, 26, 3) {real, imag} */,
  {32'hc1513f72, 32'h40ddfb50} /* (5, 26, 2) {real, imag} */,
  {32'h41198fc4, 32'hc18085d1} /* (5, 26, 1) {real, imag} */,
  {32'h41dfb55f, 32'hc019fc88} /* (5, 26, 0) {real, imag} */,
  {32'hc0c04a2c, 32'h40c12c74} /* (5, 25, 31) {real, imag} */,
  {32'hc036ac94, 32'hc1a84746} /* (5, 25, 30) {real, imag} */,
  {32'hc15cdeb8, 32'h410c5c02} /* (5, 25, 29) {real, imag} */,
  {32'h409e4d49, 32'hc07467e9} /* (5, 25, 28) {real, imag} */,
  {32'h40f39498, 32'hc1d53d65} /* (5, 25, 27) {real, imag} */,
  {32'h41719e32, 32'hc10074f6} /* (5, 25, 26) {real, imag} */,
  {32'hbce74b00, 32'h40c71e1a} /* (5, 25, 25) {real, imag} */,
  {32'h40eecada, 32'h410f0c44} /* (5, 25, 24) {real, imag} */,
  {32'h41393cf0, 32'hc0a35dd0} /* (5, 25, 23) {real, imag} */,
  {32'h4161f372, 32'hc1a52934} /* (5, 25, 22) {real, imag} */,
  {32'hc0691222, 32'hbf765400} /* (5, 25, 21) {real, imag} */,
  {32'hc05b13d8, 32'h4046b91b} /* (5, 25, 20) {real, imag} */,
  {32'hc157c307, 32'hc0a89e3a} /* (5, 25, 19) {real, imag} */,
  {32'hc1920707, 32'h40d3b173} /* (5, 25, 18) {real, imag} */,
  {32'hc108002e, 32'hc12a0ed7} /* (5, 25, 17) {real, imag} */,
  {32'hbc0ca000, 32'h40f862e6} /* (5, 25, 16) {real, imag} */,
  {32'h40e1d406, 32'hbfcc68ca} /* (5, 25, 15) {real, imag} */,
  {32'h40c6bf23, 32'hc06a803c} /* (5, 25, 14) {real, imag} */,
  {32'hc155d0e7, 32'hbf7dc1bc} /* (5, 25, 13) {real, imag} */,
  {32'h41a3d00a, 32'h41357b93} /* (5, 25, 12) {real, imag} */,
  {32'h40b31f54, 32'hc1a4a22c} /* (5, 25, 11) {real, imag} */,
  {32'h418c4dce, 32'hbe14a840} /* (5, 25, 10) {real, imag} */,
  {32'hc13261c1, 32'hc127cffe} /* (5, 25, 9) {real, imag} */,
  {32'hc1320a57, 32'hbf0d35c0} /* (5, 25, 8) {real, imag} */,
  {32'h41588aaa, 32'h411614e8} /* (5, 25, 7) {real, imag} */,
  {32'hbf1f5088, 32'h3fee2380} /* (5, 25, 6) {real, imag} */,
  {32'hc194175a, 32'h4032148b} /* (5, 25, 5) {real, imag} */,
  {32'hc1b87f12, 32'h41a9df0d} /* (5, 25, 4) {real, imag} */,
  {32'hc0e8f533, 32'h408af9b9} /* (5, 25, 3) {real, imag} */,
  {32'hc17d8e0f, 32'h411ecef2} /* (5, 25, 2) {real, imag} */,
  {32'h3fc581c8, 32'hc070a808} /* (5, 25, 1) {real, imag} */,
  {32'hc1cd6622, 32'h413f51a2} /* (5, 25, 0) {real, imag} */,
  {32'hc1112e80, 32'h40f53e30} /* (5, 24, 31) {real, imag} */,
  {32'h40f13ecb, 32'h40ef1504} /* (5, 24, 30) {real, imag} */,
  {32'hc0b44206, 32'h409a4529} /* (5, 24, 29) {real, imag} */,
  {32'h40e6258a, 32'h404b7efa} /* (5, 24, 28) {real, imag} */,
  {32'hc1b5eea0, 32'hc1409eed} /* (5, 24, 27) {real, imag} */,
  {32'h4156a992, 32'h40034150} /* (5, 24, 26) {real, imag} */,
  {32'h3e9451a0, 32'h41c57def} /* (5, 24, 25) {real, imag} */,
  {32'h41a2d6f9, 32'h419d4ef0} /* (5, 24, 24) {real, imag} */,
  {32'h414b9567, 32'hc1ea13d1} /* (5, 24, 23) {real, imag} */,
  {32'h40a29406, 32'h3f96a530} /* (5, 24, 22) {real, imag} */,
  {32'hc0806a5d, 32'h406a46d8} /* (5, 24, 21) {real, imag} */,
  {32'hc06032ec, 32'h41176986} /* (5, 24, 20) {real, imag} */,
  {32'h4108043d, 32'h40145a0c} /* (5, 24, 19) {real, imag} */,
  {32'hc1a46d56, 32'h3f438f70} /* (5, 24, 18) {real, imag} */,
  {32'h408404e8, 32'hc15579f0} /* (5, 24, 17) {real, imag} */,
  {32'h3fd50078, 32'hbd959f00} /* (5, 24, 16) {real, imag} */,
  {32'hbfa28ffe, 32'h40ff0ae5} /* (5, 24, 15) {real, imag} */,
  {32'h40818228, 32'hc108c96f} /* (5, 24, 14) {real, imag} */,
  {32'hc02a7c90, 32'h3f0f4f8c} /* (5, 24, 13) {real, imag} */,
  {32'hc07d75ec, 32'h41aae442} /* (5, 24, 12) {real, imag} */,
  {32'hc10895d0, 32'h3fb520fc} /* (5, 24, 11) {real, imag} */,
  {32'hc13b29f2, 32'hc0083ea6} /* (5, 24, 10) {real, imag} */,
  {32'h406ed3b4, 32'h41c9870d} /* (5, 24, 9) {real, imag} */,
  {32'hc1219344, 32'hc10adec8} /* (5, 24, 8) {real, imag} */,
  {32'h41197b30, 32'hc17cb568} /* (5, 24, 7) {real, imag} */,
  {32'h414d5601, 32'hc13262ae} /* (5, 24, 6) {real, imag} */,
  {32'hbf470b30, 32'h40ae78c8} /* (5, 24, 5) {real, imag} */,
  {32'hc17708f6, 32'h3f1ab9f8} /* (5, 24, 4) {real, imag} */,
  {32'h421cdcc2, 32'hc1bae395} /* (5, 24, 3) {real, imag} */,
  {32'hc184ca1b, 32'hc0fc7f3c} /* (5, 24, 2) {real, imag} */,
  {32'h41c8c834, 32'hc0378f20} /* (5, 24, 1) {real, imag} */,
  {32'h41808bc4, 32'h3d7da380} /* (5, 24, 0) {real, imag} */,
  {32'hbe620460, 32'h4042bd24} /* (5, 23, 31) {real, imag} */,
  {32'h4050b726, 32'h41cf311e} /* (5, 23, 30) {real, imag} */,
  {32'h412b8df4, 32'hc185d461} /* (5, 23, 29) {real, imag} */,
  {32'hbfff1fc9, 32'h4186e5ad} /* (5, 23, 28) {real, imag} */,
  {32'hc06f98d2, 32'hbfb3b218} /* (5, 23, 27) {real, imag} */,
  {32'hc0fd489a, 32'hc03b11f4} /* (5, 23, 26) {real, imag} */,
  {32'h4139749e, 32'h40a621b5} /* (5, 23, 25) {real, imag} */,
  {32'h417d1c13, 32'hc060c50e} /* (5, 23, 24) {real, imag} */,
  {32'h40a09265, 32'h3edebbe0} /* (5, 23, 23) {real, imag} */,
  {32'hbf45e3f0, 32'hc0d6f1f7} /* (5, 23, 22) {real, imag} */,
  {32'hbf840fa8, 32'hc0135475} /* (5, 23, 21) {real, imag} */,
  {32'hbfe4dd5a, 32'h3f47e6b4} /* (5, 23, 20) {real, imag} */,
  {32'h41569261, 32'hc12596f1} /* (5, 23, 19) {real, imag} */,
  {32'hc026930c, 32'h40042717} /* (5, 23, 18) {real, imag} */,
  {32'hc1515fac, 32'hc01f29bd} /* (5, 23, 17) {real, imag} */,
  {32'h4134b578, 32'hbfbbcba4} /* (5, 23, 16) {real, imag} */,
  {32'hc13a543b, 32'hc1782337} /* (5, 23, 15) {real, imag} */,
  {32'hc08a96b0, 32'hbf413bb0} /* (5, 23, 14) {real, imag} */,
  {32'hc008a902, 32'hc07f1d1e} /* (5, 23, 13) {real, imag} */,
  {32'hc11d05cb, 32'hc1ac9d6f} /* (5, 23, 12) {real, imag} */,
  {32'h40f5fd1e, 32'h41cb0d00} /* (5, 23, 11) {real, imag} */,
  {32'h4160129a, 32'hc1b03b75} /* (5, 23, 10) {real, imag} */,
  {32'hc11510a3, 32'hc120a68c} /* (5, 23, 9) {real, imag} */,
  {32'h41200395, 32'h4195590e} /* (5, 23, 8) {real, imag} */,
  {32'h4103f7d9, 32'h3f8a971e} /* (5, 23, 7) {real, imag} */,
  {32'h410ca1db, 32'hc0cbe539} /* (5, 23, 6) {real, imag} */,
  {32'h4121adaa, 32'hc046052e} /* (5, 23, 5) {real, imag} */,
  {32'hbf0d0ef0, 32'hc00a337b} /* (5, 23, 4) {real, imag} */,
  {32'hc0cf04b8, 32'hc05a12e7} /* (5, 23, 3) {real, imag} */,
  {32'h416caea1, 32'hc03b0e50} /* (5, 23, 2) {real, imag} */,
  {32'h3efe92c0, 32'h414ba3d6} /* (5, 23, 1) {real, imag} */,
  {32'hc1cb01aa, 32'hc0e99c2b} /* (5, 23, 0) {real, imag} */,
  {32'hc08dabc1, 32'hc0574f13} /* (5, 22, 31) {real, imag} */,
  {32'hbfbfcfc0, 32'h3e2808c0} /* (5, 22, 30) {real, imag} */,
  {32'hc0c0d714, 32'h4167400a} /* (5, 22, 29) {real, imag} */,
  {32'h40f6b8ec, 32'h41512cfb} /* (5, 22, 28) {real, imag} */,
  {32'hc114e008, 32'hbfd3c355} /* (5, 22, 27) {real, imag} */,
  {32'hc0b8f7ae, 32'hc0d4b468} /* (5, 22, 26) {real, imag} */,
  {32'h417a40ef, 32'hc1e912dc} /* (5, 22, 25) {real, imag} */,
  {32'h4120c52b, 32'h4035ad86} /* (5, 22, 24) {real, imag} */,
  {32'hc1358b81, 32'hc0d1b6d8} /* (5, 22, 23) {real, imag} */,
  {32'hc0f3928f, 32'hc0ab51c0} /* (5, 22, 22) {real, imag} */,
  {32'hc1271ce0, 32'hc0fcc2e8} /* (5, 22, 21) {real, imag} */,
  {32'hc0a9ffeb, 32'h41830938} /* (5, 22, 20) {real, imag} */,
  {32'h410bdff8, 32'h3f864b18} /* (5, 22, 19) {real, imag} */,
  {32'hc05f35bf, 32'h412103e9} /* (5, 22, 18) {real, imag} */,
  {32'h4175f945, 32'hc0010e84} /* (5, 22, 17) {real, imag} */,
  {32'h4073b228, 32'h416704f8} /* (5, 22, 16) {real, imag} */,
  {32'h40cc5d40, 32'h4076f8e0} /* (5, 22, 15) {real, imag} */,
  {32'h4149bc5b, 32'h3f77b5a0} /* (5, 22, 14) {real, imag} */,
  {32'h41324e00, 32'h4115c321} /* (5, 22, 13) {real, imag} */,
  {32'hc085de3c, 32'hbf8b5d20} /* (5, 22, 12) {real, imag} */,
  {32'hc1737412, 32'h417363c6} /* (5, 22, 11) {real, imag} */,
  {32'h412216bb, 32'hbfae9bd0} /* (5, 22, 10) {real, imag} */,
  {32'h3e02ad60, 32'hc04b63d0} /* (5, 22, 9) {real, imag} */,
  {32'hc17940ab, 32'h40493e24} /* (5, 22, 8) {real, imag} */,
  {32'h41763b46, 32'hbf6d8c98} /* (5, 22, 7) {real, imag} */,
  {32'hbfea1660, 32'hc1c0d422} /* (5, 22, 6) {real, imag} */,
  {32'h41a45438, 32'hc1535840} /* (5, 22, 5) {real, imag} */,
  {32'hc0e65807, 32'h41734f98} /* (5, 22, 4) {real, imag} */,
  {32'hc188572e, 32'h3f0c3ef0} /* (5, 22, 3) {real, imag} */,
  {32'hc00228fa, 32'h414f340e} /* (5, 22, 2) {real, imag} */,
  {32'h3e485d00, 32'h41a04356} /* (5, 22, 1) {real, imag} */,
  {32'hc0181a96, 32'h407a0e62} /* (5, 22, 0) {real, imag} */,
  {32'h3f73e850, 32'h4052a51c} /* (5, 21, 31) {real, imag} */,
  {32'h407263ba, 32'h4065f150} /* (5, 21, 30) {real, imag} */,
  {32'h41385ce4, 32'h414e1650} /* (5, 21, 29) {real, imag} */,
  {32'h40715e5c, 32'hc0a5fda6} /* (5, 21, 28) {real, imag} */,
  {32'hc06b6e30, 32'hbe203940} /* (5, 21, 27) {real, imag} */,
  {32'hc19d2e01, 32'hc144937d} /* (5, 21, 26) {real, imag} */,
  {32'hc18ab3bc, 32'hc0b726a1} /* (5, 21, 25) {real, imag} */,
  {32'h41113596, 32'h4199388d} /* (5, 21, 24) {real, imag} */,
  {32'h41193f90, 32'hc0fcb2aa} /* (5, 21, 23) {real, imag} */,
  {32'hc1c19235, 32'h414e4880} /* (5, 21, 22) {real, imag} */,
  {32'h420669de, 32'h41091faf} /* (5, 21, 21) {real, imag} */,
  {32'hbf18dfa8, 32'h40db7208} /* (5, 21, 20) {real, imag} */,
  {32'hbfafb4f0, 32'hbfd1925c} /* (5, 21, 19) {real, imag} */,
  {32'h40f92761, 32'h3fbb1e6e} /* (5, 21, 18) {real, imag} */,
  {32'hc128055f, 32'h4141d208} /* (5, 21, 17) {real, imag} */,
  {32'h40c1cf64, 32'hc1780adc} /* (5, 21, 16) {real, imag} */,
  {32'h404dca04, 32'h41170c31} /* (5, 21, 15) {real, imag} */,
  {32'h3fafe550, 32'hc0c281dc} /* (5, 21, 14) {real, imag} */,
  {32'h41055f9e, 32'hc1b682dc} /* (5, 21, 13) {real, imag} */,
  {32'h3f89294c, 32'hc1568298} /* (5, 21, 12) {real, imag} */,
  {32'hc1a391b8, 32'hc0b6cba8} /* (5, 21, 11) {real, imag} */,
  {32'h401ea37f, 32'h41be2b62} /* (5, 21, 10) {real, imag} */,
  {32'h410ddaa7, 32'h3e00a580} /* (5, 21, 9) {real, imag} */,
  {32'h3fb649ec, 32'hbed250f4} /* (5, 21, 8) {real, imag} */,
  {32'hc0af601e, 32'hc0dae229} /* (5, 21, 7) {real, imag} */,
  {32'h3fba3cbe, 32'h403b1007} /* (5, 21, 6) {real, imag} */,
  {32'h3fb5225d, 32'hc0f07d85} /* (5, 21, 5) {real, imag} */,
  {32'h412660cc, 32'hc113e792} /* (5, 21, 4) {real, imag} */,
  {32'hc13d9c4a, 32'hc08808ea} /* (5, 21, 3) {real, imag} */,
  {32'h4103f4c8, 32'hc100b28b} /* (5, 21, 2) {real, imag} */,
  {32'h410452f9, 32'hbfb4856c} /* (5, 21, 1) {real, imag} */,
  {32'h41428fa2, 32'hc082283a} /* (5, 21, 0) {real, imag} */,
  {32'hc0bc0c8a, 32'hc18dc2fd} /* (5, 20, 31) {real, imag} */,
  {32'hbfae3164, 32'hc04bf450} /* (5, 20, 30) {real, imag} */,
  {32'h40a4241b, 32'h40f3a5c4} /* (5, 20, 29) {real, imag} */,
  {32'hc150da8d, 32'hc05081b4} /* (5, 20, 28) {real, imag} */,
  {32'h41223ef4, 32'h40376ea4} /* (5, 20, 27) {real, imag} */,
  {32'hc084ab83, 32'h40b7d11e} /* (5, 20, 26) {real, imag} */,
  {32'hc09055fc, 32'hc1236c39} /* (5, 20, 25) {real, imag} */,
  {32'hc18c6683, 32'h3f82331a} /* (5, 20, 24) {real, imag} */,
  {32'h41a1872b, 32'h41357864} /* (5, 20, 23) {real, imag} */,
  {32'hc131f893, 32'h417d427d} /* (5, 20, 22) {real, imag} */,
  {32'hc146574e, 32'hc0b10006} /* (5, 20, 21) {real, imag} */,
  {32'hc05093c2, 32'hc03c14c6} /* (5, 20, 20) {real, imag} */,
  {32'hc0e25e4f, 32'h3da2cae0} /* (5, 20, 19) {real, imag} */,
  {32'h40b48476, 32'h41fb357e} /* (5, 20, 18) {real, imag} */,
  {32'h415c9a3b, 32'h40c01e7c} /* (5, 20, 17) {real, imag} */,
  {32'hbe202378, 32'hbf8ee302} /* (5, 20, 16) {real, imag} */,
  {32'hc0969107, 32'hc0babffc} /* (5, 20, 15) {real, imag} */,
  {32'hc1a6a305, 32'h410552b2} /* (5, 20, 14) {real, imag} */,
  {32'h402180c9, 32'h3f25d5e8} /* (5, 20, 13) {real, imag} */,
  {32'h4180e988, 32'hc1316ad8} /* (5, 20, 12) {real, imag} */,
  {32'h4006d1f0, 32'h3f1fd600} /* (5, 20, 11) {real, imag} */,
  {32'h4007c3dc, 32'hbf9b2e48} /* (5, 20, 10) {real, imag} */,
  {32'h40504df8, 32'hbe065ec0} /* (5, 20, 9) {real, imag} */,
  {32'h4063e5ac, 32'h40ea61aa} /* (5, 20, 8) {real, imag} */,
  {32'h41943038, 32'h4129a46f} /* (5, 20, 7) {real, imag} */,
  {32'hc17a2a50, 32'h416f3b9b} /* (5, 20, 6) {real, imag} */,
  {32'h40a9bbd0, 32'hc10f5b2e} /* (5, 20, 5) {real, imag} */,
  {32'h40440aae, 32'h4103d723} /* (5, 20, 4) {real, imag} */,
  {32'h4130e622, 32'h40a69f62} /* (5, 20, 3) {real, imag} */,
  {32'hc13a82db, 32'hc0501010} /* (5, 20, 2) {real, imag} */,
  {32'h41010ec2, 32'hc055e8ff} /* (5, 20, 1) {real, imag} */,
  {32'hc036b83b, 32'h408de54f} /* (5, 20, 0) {real, imag} */,
  {32'h4139855c, 32'hc079b093} /* (5, 19, 31) {real, imag} */,
  {32'h4198f6e2, 32'h404a2038} /* (5, 19, 30) {real, imag} */,
  {32'hbf478968, 32'hc095b681} /* (5, 19, 29) {real, imag} */,
  {32'hc02865aa, 32'h4045e060} /* (5, 19, 28) {real, imag} */,
  {32'hbfd42d0c, 32'hc0237863} /* (5, 19, 27) {real, imag} */,
  {32'h40fd2ebd, 32'hbf31f160} /* (5, 19, 26) {real, imag} */,
  {32'hc201b858, 32'h40c288e3} /* (5, 19, 25) {real, imag} */,
  {32'hc08e4869, 32'hc0931f24} /* (5, 19, 24) {real, imag} */,
  {32'hc10deca8, 32'h41b73d28} /* (5, 19, 23) {real, imag} */,
  {32'hc0f8ace0, 32'hc005cb6f} /* (5, 19, 22) {real, imag} */,
  {32'h408a3995, 32'hc0572415} /* (5, 19, 21) {real, imag} */,
  {32'h3f81dcf0, 32'hc0e8e627} /* (5, 19, 20) {real, imag} */,
  {32'h419b2ba8, 32'h3e8d2b00} /* (5, 19, 19) {real, imag} */,
  {32'hc108b50a, 32'hc0ae82b3} /* (5, 19, 18) {real, imag} */,
  {32'hbebfba30, 32'hbd0361c0} /* (5, 19, 17) {real, imag} */,
  {32'hc187f109, 32'hc0ba3a99} /* (5, 19, 16) {real, imag} */,
  {32'hc1900920, 32'hc027b89e} /* (5, 19, 15) {real, imag} */,
  {32'h3faa9c4c, 32'hc13164bf} /* (5, 19, 14) {real, imag} */,
  {32'hc100feaf, 32'h41152e21} /* (5, 19, 13) {real, imag} */,
  {32'h418084d0, 32'h40c51996} /* (5, 19, 12) {real, imag} */,
  {32'h40fc8d94, 32'h41607f4a} /* (5, 19, 11) {real, imag} */,
  {32'h4133c7ad, 32'hc15ab884} /* (5, 19, 10) {real, imag} */,
  {32'hc199aeab, 32'h410a5c4e} /* (5, 19, 9) {real, imag} */,
  {32'h40f316e3, 32'h40ebebea} /* (5, 19, 8) {real, imag} */,
  {32'hbfa9b7ac, 32'h416d1c26} /* (5, 19, 7) {real, imag} */,
  {32'hc100aafb, 32'h406afedf} /* (5, 19, 6) {real, imag} */,
  {32'hc0ebf916, 32'hbfae7a75} /* (5, 19, 5) {real, imag} */,
  {32'hc0b553f5, 32'hc0f02624} /* (5, 19, 4) {real, imag} */,
  {32'hc0a5f7a8, 32'h3ffeb500} /* (5, 19, 3) {real, imag} */,
  {32'h414febe8, 32'hc143690e} /* (5, 19, 2) {real, imag} */,
  {32'hc14c137a, 32'h40a495e0} /* (5, 19, 1) {real, imag} */,
  {32'hc06f7c10, 32'h410885ee} /* (5, 19, 0) {real, imag} */,
  {32'hc0c5f160, 32'hbf60ee68} /* (5, 18, 31) {real, imag} */,
  {32'h414ac6fb, 32'h4009f858} /* (5, 18, 30) {real, imag} */,
  {32'hc1027a36, 32'h40baa91e} /* (5, 18, 29) {real, imag} */,
  {32'hc18953d5, 32'hc0aca796} /* (5, 18, 28) {real, imag} */,
  {32'h40b3dbc6, 32'hc12b6ecb} /* (5, 18, 27) {real, imag} */,
  {32'h3fb4f0e2, 32'hc1225b9a} /* (5, 18, 26) {real, imag} */,
  {32'hbf827480, 32'hc119c425} /* (5, 18, 25) {real, imag} */,
  {32'h41756960, 32'h41392c5e} /* (5, 18, 24) {real, imag} */,
  {32'h40626e82, 32'hc075728e} /* (5, 18, 23) {real, imag} */,
  {32'hc10ff64f, 32'hc10ee591} /* (5, 18, 22) {real, imag} */,
  {32'h411322d0, 32'h405f69ed} /* (5, 18, 21) {real, imag} */,
  {32'hc0b07fd2, 32'hc0d718bc} /* (5, 18, 20) {real, imag} */,
  {32'h415cf6aa, 32'h405e1e5b} /* (5, 18, 19) {real, imag} */,
  {32'hc055a78c, 32'h3fa6bde0} /* (5, 18, 18) {real, imag} */,
  {32'h411d2856, 32'hbef92c80} /* (5, 18, 17) {real, imag} */,
  {32'h3fd97eb6, 32'h40e931e8} /* (5, 18, 16) {real, imag} */,
  {32'hc10e125b, 32'hc02242f0} /* (5, 18, 15) {real, imag} */,
  {32'h3f9f72a0, 32'hbf84ba49} /* (5, 18, 14) {real, imag} */,
  {32'h40942203, 32'h408c05ea} /* (5, 18, 13) {real, imag} */,
  {32'hc1c014d6, 32'h418917a9} /* (5, 18, 12) {real, imag} */,
  {32'h415794c4, 32'h411a96ee} /* (5, 18, 11) {real, imag} */,
  {32'h4078a6e0, 32'h405893e8} /* (5, 18, 10) {real, imag} */,
  {32'h40931115, 32'h3e675f60} /* (5, 18, 9) {real, imag} */,
  {32'hc12ab1bd, 32'h4004f46e} /* (5, 18, 8) {real, imag} */,
  {32'hc0bba65c, 32'h4139c137} /* (5, 18, 7) {real, imag} */,
  {32'hc0ab839e, 32'hc1c37dd4} /* (5, 18, 6) {real, imag} */,
  {32'hbf3f6192, 32'hc0dd055b} /* (5, 18, 5) {real, imag} */,
  {32'hbfd7b380, 32'h3f80d494} /* (5, 18, 4) {real, imag} */,
  {32'h3fe12bb2, 32'hc0b4571c} /* (5, 18, 3) {real, imag} */,
  {32'hbe75afc0, 32'h4133d49e} /* (5, 18, 2) {real, imag} */,
  {32'hc069ea98, 32'hbfbb6d14} /* (5, 18, 1) {real, imag} */,
  {32'h40f8027d, 32'hc0789667} /* (5, 18, 0) {real, imag} */,
  {32'h40e0fedc, 32'hc04fbb1a} /* (5, 17, 31) {real, imag} */,
  {32'hbfa09aec, 32'hc03b95c4} /* (5, 17, 30) {real, imag} */,
  {32'h40a740f3, 32'h40f2522c} /* (5, 17, 29) {real, imag} */,
  {32'h3ddcd830, 32'h407ec538} /* (5, 17, 28) {real, imag} */,
  {32'hc0f5fa7e, 32'h400d809e} /* (5, 17, 27) {real, imag} */,
  {32'h3faccb6a, 32'h411a91b3} /* (5, 17, 26) {real, imag} */,
  {32'hc0e359f1, 32'hc05a3ab8} /* (5, 17, 25) {real, imag} */,
  {32'hc100b9b4, 32'h400c1a7f} /* (5, 17, 24) {real, imag} */,
  {32'hc16afb42, 32'hbfc01b70} /* (5, 17, 23) {real, imag} */,
  {32'h3f69b578, 32'h4087e303} /* (5, 17, 22) {real, imag} */,
  {32'hc16e822e, 32'hc028a9a0} /* (5, 17, 21) {real, imag} */,
  {32'h40fe2638, 32'hbf71a7bc} /* (5, 17, 20) {real, imag} */,
  {32'hc1300d40, 32'hc1365ca3} /* (5, 17, 19) {real, imag} */,
  {32'h40cff076, 32'h40210e90} /* (5, 17, 18) {real, imag} */,
  {32'hc09de6c6, 32'hbeecb940} /* (5, 17, 17) {real, imag} */,
  {32'h415395fc, 32'h40817a56} /* (5, 17, 16) {real, imag} */,
  {32'h3dde14e0, 32'hc120a528} /* (5, 17, 15) {real, imag} */,
  {32'hc03c3826, 32'h409e534a} /* (5, 17, 14) {real, imag} */,
  {32'hc0590254, 32'h414c16ee} /* (5, 17, 13) {real, imag} */,
  {32'hc113ce23, 32'hc1a05cec} /* (5, 17, 12) {real, imag} */,
  {32'h4139af98, 32'hc0dd49a3} /* (5, 17, 11) {real, imag} */,
  {32'hbff6f309, 32'h40bf0b98} /* (5, 17, 10) {real, imag} */,
  {32'hc0c0ded7, 32'h4133d3ce} /* (5, 17, 9) {real, imag} */,
  {32'hc0035b20, 32'hc02f2b16} /* (5, 17, 8) {real, imag} */,
  {32'hc09a46af, 32'hbedd8c3c} /* (5, 17, 7) {real, imag} */,
  {32'h40a624ff, 32'h412f5ee6} /* (5, 17, 6) {real, imag} */,
  {32'hc0e6afe8, 32'hbf24b638} /* (5, 17, 5) {real, imag} */,
  {32'h40d5378b, 32'hc12122ec} /* (5, 17, 4) {real, imag} */,
  {32'h40352118, 32'hc093a120} /* (5, 17, 3) {real, imag} */,
  {32'h40417a50, 32'hc0362afa} /* (5, 17, 2) {real, imag} */,
  {32'hc0969fa5, 32'h41c6d50c} /* (5, 17, 1) {real, imag} */,
  {32'h40aa6297, 32'h412828a1} /* (5, 17, 0) {real, imag} */,
  {32'h40341599, 32'hbea07780} /* (5, 16, 31) {real, imag} */,
  {32'h3f00112c, 32'h40972c8e} /* (5, 16, 30) {real, imag} */,
  {32'h409829ee, 32'h40a5ef6e} /* (5, 16, 29) {real, imag} */,
  {32'hc0fa71f0, 32'h3ef3ffa0} /* (5, 16, 28) {real, imag} */,
  {32'h4071b6f1, 32'hc1181466} /* (5, 16, 27) {real, imag} */,
  {32'hc144b57c, 32'h403ee64f} /* (5, 16, 26) {real, imag} */,
  {32'hc019108e, 32'hbff67f28} /* (5, 16, 25) {real, imag} */,
  {32'hc06375d6, 32'hbeb95448} /* (5, 16, 24) {real, imag} */,
  {32'hbf323e72, 32'hc0e505a2} /* (5, 16, 23) {real, imag} */,
  {32'hc0d2b9ea, 32'h3fd02c79} /* (5, 16, 22) {real, imag} */,
  {32'h40d79aea, 32'h4102946c} /* (5, 16, 21) {real, imag} */,
  {32'h41238c95, 32'hbff29e50} /* (5, 16, 20) {real, imag} */,
  {32'h411bc8a7, 32'h4169cb23} /* (5, 16, 19) {real, imag} */,
  {32'hc084d942, 32'hbfe67c24} /* (5, 16, 18) {real, imag} */,
  {32'h3da96dc0, 32'hc0bd5427} /* (5, 16, 17) {real, imag} */,
  {32'hc0562ad7, 32'h00000000} /* (5, 16, 16) {real, imag} */,
  {32'h3da96dc0, 32'h40bd5427} /* (5, 16, 15) {real, imag} */,
  {32'hc084d942, 32'h3fe67c24} /* (5, 16, 14) {real, imag} */,
  {32'h411bc8a7, 32'hc169cb23} /* (5, 16, 13) {real, imag} */,
  {32'h41238c95, 32'h3ff29e50} /* (5, 16, 12) {real, imag} */,
  {32'h40d79aea, 32'hc102946c} /* (5, 16, 11) {real, imag} */,
  {32'hc0d2b9ea, 32'hbfd02c79} /* (5, 16, 10) {real, imag} */,
  {32'hbf323e72, 32'h40e505a2} /* (5, 16, 9) {real, imag} */,
  {32'hc06375d6, 32'h3eb95448} /* (5, 16, 8) {real, imag} */,
  {32'hc019108e, 32'h3ff67f28} /* (5, 16, 7) {real, imag} */,
  {32'hc144b57c, 32'hc03ee64f} /* (5, 16, 6) {real, imag} */,
  {32'h4071b6f1, 32'h41181466} /* (5, 16, 5) {real, imag} */,
  {32'hc0fa71f0, 32'hbef3ffa0} /* (5, 16, 4) {real, imag} */,
  {32'h409829ee, 32'hc0a5ef6e} /* (5, 16, 3) {real, imag} */,
  {32'h3f00112c, 32'hc0972c8e} /* (5, 16, 2) {real, imag} */,
  {32'h40341599, 32'h3ea07780} /* (5, 16, 1) {real, imag} */,
  {32'h4148d2a7, 32'h00000000} /* (5, 16, 0) {real, imag} */,
  {32'hc0969fa5, 32'hc1c6d50c} /* (5, 15, 31) {real, imag} */,
  {32'h40417a50, 32'h40362afa} /* (5, 15, 30) {real, imag} */,
  {32'h40352118, 32'h4093a120} /* (5, 15, 29) {real, imag} */,
  {32'h40d5378b, 32'h412122ec} /* (5, 15, 28) {real, imag} */,
  {32'hc0e6afe8, 32'h3f24b638} /* (5, 15, 27) {real, imag} */,
  {32'h40a624ff, 32'hc12f5ee6} /* (5, 15, 26) {real, imag} */,
  {32'hc09a46af, 32'h3edd8c3c} /* (5, 15, 25) {real, imag} */,
  {32'hc0035b20, 32'h402f2b16} /* (5, 15, 24) {real, imag} */,
  {32'hc0c0ded7, 32'hc133d3ce} /* (5, 15, 23) {real, imag} */,
  {32'hbff6f309, 32'hc0bf0b98} /* (5, 15, 22) {real, imag} */,
  {32'h4139af98, 32'h40dd49a3} /* (5, 15, 21) {real, imag} */,
  {32'hc113ce23, 32'h41a05cec} /* (5, 15, 20) {real, imag} */,
  {32'hc0590254, 32'hc14c16ee} /* (5, 15, 19) {real, imag} */,
  {32'hc03c3826, 32'hc09e534a} /* (5, 15, 18) {real, imag} */,
  {32'h3dde14e0, 32'h4120a528} /* (5, 15, 17) {real, imag} */,
  {32'h415395fc, 32'hc0817a56} /* (5, 15, 16) {real, imag} */,
  {32'hc09de6c6, 32'h3eecb940} /* (5, 15, 15) {real, imag} */,
  {32'h40cff076, 32'hc0210e90} /* (5, 15, 14) {real, imag} */,
  {32'hc1300d40, 32'h41365ca3} /* (5, 15, 13) {real, imag} */,
  {32'h40fe2638, 32'h3f71a7bc} /* (5, 15, 12) {real, imag} */,
  {32'hc16e822e, 32'h4028a9a0} /* (5, 15, 11) {real, imag} */,
  {32'h3f69b578, 32'hc087e303} /* (5, 15, 10) {real, imag} */,
  {32'hc16afb42, 32'h3fc01b70} /* (5, 15, 9) {real, imag} */,
  {32'hc100b9b4, 32'hc00c1a7f} /* (5, 15, 8) {real, imag} */,
  {32'hc0e359f1, 32'h405a3ab8} /* (5, 15, 7) {real, imag} */,
  {32'h3faccb6a, 32'hc11a91b3} /* (5, 15, 6) {real, imag} */,
  {32'hc0f5fa7e, 32'hc00d809e} /* (5, 15, 5) {real, imag} */,
  {32'h3ddcd830, 32'hc07ec538} /* (5, 15, 4) {real, imag} */,
  {32'h40a740f3, 32'hc0f2522c} /* (5, 15, 3) {real, imag} */,
  {32'hbfa09aec, 32'h403b95c4} /* (5, 15, 2) {real, imag} */,
  {32'h40e0fedc, 32'h404fbb1a} /* (5, 15, 1) {real, imag} */,
  {32'h40aa6297, 32'hc12828a1} /* (5, 15, 0) {real, imag} */,
  {32'hc069ea98, 32'h3fbb6d14} /* (5, 14, 31) {real, imag} */,
  {32'hbe75afc0, 32'hc133d49e} /* (5, 14, 30) {real, imag} */,
  {32'h3fe12bb2, 32'h40b4571c} /* (5, 14, 29) {real, imag} */,
  {32'hbfd7b380, 32'hbf80d494} /* (5, 14, 28) {real, imag} */,
  {32'hbf3f6192, 32'h40dd055b} /* (5, 14, 27) {real, imag} */,
  {32'hc0ab839e, 32'h41c37dd4} /* (5, 14, 26) {real, imag} */,
  {32'hc0bba65c, 32'hc139c137} /* (5, 14, 25) {real, imag} */,
  {32'hc12ab1bd, 32'hc004f46e} /* (5, 14, 24) {real, imag} */,
  {32'h40931115, 32'hbe675f60} /* (5, 14, 23) {real, imag} */,
  {32'h4078a6e0, 32'hc05893e8} /* (5, 14, 22) {real, imag} */,
  {32'h415794c4, 32'hc11a96ee} /* (5, 14, 21) {real, imag} */,
  {32'hc1c014d6, 32'hc18917a9} /* (5, 14, 20) {real, imag} */,
  {32'h40942203, 32'hc08c05ea} /* (5, 14, 19) {real, imag} */,
  {32'h3f9f72a0, 32'h3f84ba49} /* (5, 14, 18) {real, imag} */,
  {32'hc10e125b, 32'h402242f0} /* (5, 14, 17) {real, imag} */,
  {32'h3fd97eb6, 32'hc0e931e8} /* (5, 14, 16) {real, imag} */,
  {32'h411d2856, 32'h3ef92c80} /* (5, 14, 15) {real, imag} */,
  {32'hc055a78c, 32'hbfa6bde0} /* (5, 14, 14) {real, imag} */,
  {32'h415cf6aa, 32'hc05e1e5b} /* (5, 14, 13) {real, imag} */,
  {32'hc0b07fd2, 32'h40d718bc} /* (5, 14, 12) {real, imag} */,
  {32'h411322d0, 32'hc05f69ed} /* (5, 14, 11) {real, imag} */,
  {32'hc10ff64f, 32'h410ee591} /* (5, 14, 10) {real, imag} */,
  {32'h40626e82, 32'h4075728e} /* (5, 14, 9) {real, imag} */,
  {32'h41756960, 32'hc1392c5e} /* (5, 14, 8) {real, imag} */,
  {32'hbf827480, 32'h4119c425} /* (5, 14, 7) {real, imag} */,
  {32'h3fb4f0e2, 32'h41225b9a} /* (5, 14, 6) {real, imag} */,
  {32'h40b3dbc6, 32'h412b6ecb} /* (5, 14, 5) {real, imag} */,
  {32'hc18953d5, 32'h40aca796} /* (5, 14, 4) {real, imag} */,
  {32'hc1027a36, 32'hc0baa91e} /* (5, 14, 3) {real, imag} */,
  {32'h414ac6fb, 32'hc009f858} /* (5, 14, 2) {real, imag} */,
  {32'hc0c5f160, 32'h3f60ee68} /* (5, 14, 1) {real, imag} */,
  {32'h40f8027d, 32'h40789667} /* (5, 14, 0) {real, imag} */,
  {32'hc14c137a, 32'hc0a495e0} /* (5, 13, 31) {real, imag} */,
  {32'h414febe8, 32'h4143690e} /* (5, 13, 30) {real, imag} */,
  {32'hc0a5f7a8, 32'hbffeb500} /* (5, 13, 29) {real, imag} */,
  {32'hc0b553f5, 32'h40f02624} /* (5, 13, 28) {real, imag} */,
  {32'hc0ebf916, 32'h3fae7a75} /* (5, 13, 27) {real, imag} */,
  {32'hc100aafb, 32'hc06afedf} /* (5, 13, 26) {real, imag} */,
  {32'hbfa9b7ac, 32'hc16d1c26} /* (5, 13, 25) {real, imag} */,
  {32'h40f316e3, 32'hc0ebebea} /* (5, 13, 24) {real, imag} */,
  {32'hc199aeab, 32'hc10a5c4e} /* (5, 13, 23) {real, imag} */,
  {32'h4133c7ad, 32'h415ab884} /* (5, 13, 22) {real, imag} */,
  {32'h40fc8d94, 32'hc1607f4a} /* (5, 13, 21) {real, imag} */,
  {32'h418084d0, 32'hc0c51996} /* (5, 13, 20) {real, imag} */,
  {32'hc100feaf, 32'hc1152e21} /* (5, 13, 19) {real, imag} */,
  {32'h3faa9c4c, 32'h413164bf} /* (5, 13, 18) {real, imag} */,
  {32'hc1900920, 32'h4027b89e} /* (5, 13, 17) {real, imag} */,
  {32'hc187f109, 32'h40ba3a99} /* (5, 13, 16) {real, imag} */,
  {32'hbebfba30, 32'h3d0361c0} /* (5, 13, 15) {real, imag} */,
  {32'hc108b50a, 32'h40ae82b3} /* (5, 13, 14) {real, imag} */,
  {32'h419b2ba8, 32'hbe8d2b00} /* (5, 13, 13) {real, imag} */,
  {32'h3f81dcf0, 32'h40e8e627} /* (5, 13, 12) {real, imag} */,
  {32'h408a3995, 32'h40572415} /* (5, 13, 11) {real, imag} */,
  {32'hc0f8ace0, 32'h4005cb6f} /* (5, 13, 10) {real, imag} */,
  {32'hc10deca8, 32'hc1b73d28} /* (5, 13, 9) {real, imag} */,
  {32'hc08e4869, 32'h40931f24} /* (5, 13, 8) {real, imag} */,
  {32'hc201b858, 32'hc0c288e3} /* (5, 13, 7) {real, imag} */,
  {32'h40fd2ebd, 32'h3f31f160} /* (5, 13, 6) {real, imag} */,
  {32'hbfd42d0c, 32'h40237863} /* (5, 13, 5) {real, imag} */,
  {32'hc02865aa, 32'hc045e060} /* (5, 13, 4) {real, imag} */,
  {32'hbf478968, 32'h4095b681} /* (5, 13, 3) {real, imag} */,
  {32'h4198f6e2, 32'hc04a2038} /* (5, 13, 2) {real, imag} */,
  {32'h4139855c, 32'h4079b093} /* (5, 13, 1) {real, imag} */,
  {32'hc06f7c10, 32'hc10885ee} /* (5, 13, 0) {real, imag} */,
  {32'h41010ec2, 32'h4055e8ff} /* (5, 12, 31) {real, imag} */,
  {32'hc13a82db, 32'h40501010} /* (5, 12, 30) {real, imag} */,
  {32'h4130e622, 32'hc0a69f62} /* (5, 12, 29) {real, imag} */,
  {32'h40440aae, 32'hc103d723} /* (5, 12, 28) {real, imag} */,
  {32'h40a9bbd0, 32'h410f5b2e} /* (5, 12, 27) {real, imag} */,
  {32'hc17a2a50, 32'hc16f3b9b} /* (5, 12, 26) {real, imag} */,
  {32'h41943038, 32'hc129a46f} /* (5, 12, 25) {real, imag} */,
  {32'h4063e5ac, 32'hc0ea61aa} /* (5, 12, 24) {real, imag} */,
  {32'h40504df8, 32'h3e065ec0} /* (5, 12, 23) {real, imag} */,
  {32'h4007c3dc, 32'h3f9b2e48} /* (5, 12, 22) {real, imag} */,
  {32'h4006d1f0, 32'hbf1fd600} /* (5, 12, 21) {real, imag} */,
  {32'h4180e988, 32'h41316ad8} /* (5, 12, 20) {real, imag} */,
  {32'h402180c9, 32'hbf25d5e8} /* (5, 12, 19) {real, imag} */,
  {32'hc1a6a305, 32'hc10552b2} /* (5, 12, 18) {real, imag} */,
  {32'hc0969107, 32'h40babffc} /* (5, 12, 17) {real, imag} */,
  {32'hbe202378, 32'h3f8ee302} /* (5, 12, 16) {real, imag} */,
  {32'h415c9a3b, 32'hc0c01e7c} /* (5, 12, 15) {real, imag} */,
  {32'h40b48476, 32'hc1fb357e} /* (5, 12, 14) {real, imag} */,
  {32'hc0e25e4f, 32'hbda2cae0} /* (5, 12, 13) {real, imag} */,
  {32'hc05093c2, 32'h403c14c6} /* (5, 12, 12) {real, imag} */,
  {32'hc146574e, 32'h40b10006} /* (5, 12, 11) {real, imag} */,
  {32'hc131f893, 32'hc17d427d} /* (5, 12, 10) {real, imag} */,
  {32'h41a1872b, 32'hc1357864} /* (5, 12, 9) {real, imag} */,
  {32'hc18c6683, 32'hbf82331a} /* (5, 12, 8) {real, imag} */,
  {32'hc09055fc, 32'h41236c39} /* (5, 12, 7) {real, imag} */,
  {32'hc084ab83, 32'hc0b7d11e} /* (5, 12, 6) {real, imag} */,
  {32'h41223ef4, 32'hc0376ea4} /* (5, 12, 5) {real, imag} */,
  {32'hc150da8d, 32'h405081b4} /* (5, 12, 4) {real, imag} */,
  {32'h40a4241b, 32'hc0f3a5c4} /* (5, 12, 3) {real, imag} */,
  {32'hbfae3164, 32'h404bf450} /* (5, 12, 2) {real, imag} */,
  {32'hc0bc0c8a, 32'h418dc2fd} /* (5, 12, 1) {real, imag} */,
  {32'hc036b83b, 32'hc08de54f} /* (5, 12, 0) {real, imag} */,
  {32'h410452f9, 32'h3fb4856c} /* (5, 11, 31) {real, imag} */,
  {32'h4103f4c8, 32'h4100b28b} /* (5, 11, 30) {real, imag} */,
  {32'hc13d9c4a, 32'h408808ea} /* (5, 11, 29) {real, imag} */,
  {32'h412660cc, 32'h4113e792} /* (5, 11, 28) {real, imag} */,
  {32'h3fb5225d, 32'h40f07d85} /* (5, 11, 27) {real, imag} */,
  {32'h3fba3cbe, 32'hc03b1007} /* (5, 11, 26) {real, imag} */,
  {32'hc0af601e, 32'h40dae229} /* (5, 11, 25) {real, imag} */,
  {32'h3fb649ec, 32'h3ed250f4} /* (5, 11, 24) {real, imag} */,
  {32'h410ddaa7, 32'hbe00a580} /* (5, 11, 23) {real, imag} */,
  {32'h401ea37f, 32'hc1be2b62} /* (5, 11, 22) {real, imag} */,
  {32'hc1a391b8, 32'h40b6cba8} /* (5, 11, 21) {real, imag} */,
  {32'h3f89294c, 32'h41568298} /* (5, 11, 20) {real, imag} */,
  {32'h41055f9e, 32'h41b682dc} /* (5, 11, 19) {real, imag} */,
  {32'h3fafe550, 32'h40c281dc} /* (5, 11, 18) {real, imag} */,
  {32'h404dca04, 32'hc1170c31} /* (5, 11, 17) {real, imag} */,
  {32'h40c1cf64, 32'h41780adc} /* (5, 11, 16) {real, imag} */,
  {32'hc128055f, 32'hc141d208} /* (5, 11, 15) {real, imag} */,
  {32'h40f92761, 32'hbfbb1e6e} /* (5, 11, 14) {real, imag} */,
  {32'hbfafb4f0, 32'h3fd1925c} /* (5, 11, 13) {real, imag} */,
  {32'hbf18dfa8, 32'hc0db7208} /* (5, 11, 12) {real, imag} */,
  {32'h420669de, 32'hc1091faf} /* (5, 11, 11) {real, imag} */,
  {32'hc1c19235, 32'hc14e4880} /* (5, 11, 10) {real, imag} */,
  {32'h41193f90, 32'h40fcb2aa} /* (5, 11, 9) {real, imag} */,
  {32'h41113596, 32'hc199388d} /* (5, 11, 8) {real, imag} */,
  {32'hc18ab3bc, 32'h40b726a1} /* (5, 11, 7) {real, imag} */,
  {32'hc19d2e01, 32'h4144937d} /* (5, 11, 6) {real, imag} */,
  {32'hc06b6e30, 32'h3e203940} /* (5, 11, 5) {real, imag} */,
  {32'h40715e5c, 32'h40a5fda6} /* (5, 11, 4) {real, imag} */,
  {32'h41385ce4, 32'hc14e1650} /* (5, 11, 3) {real, imag} */,
  {32'h407263ba, 32'hc065f150} /* (5, 11, 2) {real, imag} */,
  {32'h3f73e850, 32'hc052a51c} /* (5, 11, 1) {real, imag} */,
  {32'h41428fa2, 32'h4082283a} /* (5, 11, 0) {real, imag} */,
  {32'h3e485d00, 32'hc1a04356} /* (5, 10, 31) {real, imag} */,
  {32'hc00228fa, 32'hc14f340e} /* (5, 10, 30) {real, imag} */,
  {32'hc188572e, 32'hbf0c3ef0} /* (5, 10, 29) {real, imag} */,
  {32'hc0e65807, 32'hc1734f98} /* (5, 10, 28) {real, imag} */,
  {32'h41a45438, 32'h41535840} /* (5, 10, 27) {real, imag} */,
  {32'hbfea1660, 32'h41c0d422} /* (5, 10, 26) {real, imag} */,
  {32'h41763b46, 32'h3f6d8c98} /* (5, 10, 25) {real, imag} */,
  {32'hc17940ab, 32'hc0493e24} /* (5, 10, 24) {real, imag} */,
  {32'h3e02ad60, 32'h404b63d0} /* (5, 10, 23) {real, imag} */,
  {32'h412216bb, 32'h3fae9bd0} /* (5, 10, 22) {real, imag} */,
  {32'hc1737412, 32'hc17363c6} /* (5, 10, 21) {real, imag} */,
  {32'hc085de3c, 32'h3f8b5d20} /* (5, 10, 20) {real, imag} */,
  {32'h41324e00, 32'hc115c321} /* (5, 10, 19) {real, imag} */,
  {32'h4149bc5b, 32'hbf77b5a0} /* (5, 10, 18) {real, imag} */,
  {32'h40cc5d40, 32'hc076f8e0} /* (5, 10, 17) {real, imag} */,
  {32'h4073b228, 32'hc16704f8} /* (5, 10, 16) {real, imag} */,
  {32'h4175f945, 32'h40010e84} /* (5, 10, 15) {real, imag} */,
  {32'hc05f35bf, 32'hc12103e9} /* (5, 10, 14) {real, imag} */,
  {32'h410bdff8, 32'hbf864b18} /* (5, 10, 13) {real, imag} */,
  {32'hc0a9ffeb, 32'hc1830938} /* (5, 10, 12) {real, imag} */,
  {32'hc1271ce0, 32'h40fcc2e8} /* (5, 10, 11) {real, imag} */,
  {32'hc0f3928f, 32'h40ab51c0} /* (5, 10, 10) {real, imag} */,
  {32'hc1358b81, 32'h40d1b6d8} /* (5, 10, 9) {real, imag} */,
  {32'h4120c52b, 32'hc035ad86} /* (5, 10, 8) {real, imag} */,
  {32'h417a40ef, 32'h41e912dc} /* (5, 10, 7) {real, imag} */,
  {32'hc0b8f7ae, 32'h40d4b468} /* (5, 10, 6) {real, imag} */,
  {32'hc114e008, 32'h3fd3c355} /* (5, 10, 5) {real, imag} */,
  {32'h40f6b8ec, 32'hc1512cfb} /* (5, 10, 4) {real, imag} */,
  {32'hc0c0d714, 32'hc167400a} /* (5, 10, 3) {real, imag} */,
  {32'hbfbfcfc0, 32'hbe2808c0} /* (5, 10, 2) {real, imag} */,
  {32'hc08dabc1, 32'h40574f13} /* (5, 10, 1) {real, imag} */,
  {32'hc0181a96, 32'hc07a0e62} /* (5, 10, 0) {real, imag} */,
  {32'h3efe92c0, 32'hc14ba3d6} /* (5, 9, 31) {real, imag} */,
  {32'h416caea1, 32'h403b0e50} /* (5, 9, 30) {real, imag} */,
  {32'hc0cf04b8, 32'h405a12e7} /* (5, 9, 29) {real, imag} */,
  {32'hbf0d0ef0, 32'h400a337b} /* (5, 9, 28) {real, imag} */,
  {32'h4121adaa, 32'h4046052e} /* (5, 9, 27) {real, imag} */,
  {32'h410ca1db, 32'h40cbe539} /* (5, 9, 26) {real, imag} */,
  {32'h4103f7d9, 32'hbf8a971e} /* (5, 9, 25) {real, imag} */,
  {32'h41200395, 32'hc195590e} /* (5, 9, 24) {real, imag} */,
  {32'hc11510a3, 32'h4120a68c} /* (5, 9, 23) {real, imag} */,
  {32'h4160129a, 32'h41b03b75} /* (5, 9, 22) {real, imag} */,
  {32'h40f5fd1e, 32'hc1cb0d00} /* (5, 9, 21) {real, imag} */,
  {32'hc11d05cb, 32'h41ac9d6f} /* (5, 9, 20) {real, imag} */,
  {32'hc008a902, 32'h407f1d1e} /* (5, 9, 19) {real, imag} */,
  {32'hc08a96b0, 32'h3f413bb0} /* (5, 9, 18) {real, imag} */,
  {32'hc13a543b, 32'h41782337} /* (5, 9, 17) {real, imag} */,
  {32'h4134b578, 32'h3fbbcba4} /* (5, 9, 16) {real, imag} */,
  {32'hc1515fac, 32'h401f29bd} /* (5, 9, 15) {real, imag} */,
  {32'hc026930c, 32'hc0042717} /* (5, 9, 14) {real, imag} */,
  {32'h41569261, 32'h412596f1} /* (5, 9, 13) {real, imag} */,
  {32'hbfe4dd5a, 32'hbf47e6b4} /* (5, 9, 12) {real, imag} */,
  {32'hbf840fa8, 32'h40135475} /* (5, 9, 11) {real, imag} */,
  {32'hbf45e3f0, 32'h40d6f1f7} /* (5, 9, 10) {real, imag} */,
  {32'h40a09265, 32'hbedebbe0} /* (5, 9, 9) {real, imag} */,
  {32'h417d1c13, 32'h4060c50e} /* (5, 9, 8) {real, imag} */,
  {32'h4139749e, 32'hc0a621b5} /* (5, 9, 7) {real, imag} */,
  {32'hc0fd489a, 32'h403b11f4} /* (5, 9, 6) {real, imag} */,
  {32'hc06f98d2, 32'h3fb3b218} /* (5, 9, 5) {real, imag} */,
  {32'hbfff1fc9, 32'hc186e5ad} /* (5, 9, 4) {real, imag} */,
  {32'h412b8df4, 32'h4185d461} /* (5, 9, 3) {real, imag} */,
  {32'h4050b726, 32'hc1cf311e} /* (5, 9, 2) {real, imag} */,
  {32'hbe620460, 32'hc042bd24} /* (5, 9, 1) {real, imag} */,
  {32'hc1cb01aa, 32'h40e99c2b} /* (5, 9, 0) {real, imag} */,
  {32'h41c8c834, 32'h40378f20} /* (5, 8, 31) {real, imag} */,
  {32'hc184ca1b, 32'h40fc7f3c} /* (5, 8, 30) {real, imag} */,
  {32'h421cdcc2, 32'h41bae395} /* (5, 8, 29) {real, imag} */,
  {32'hc17708f6, 32'hbf1ab9f8} /* (5, 8, 28) {real, imag} */,
  {32'hbf470b30, 32'hc0ae78c8} /* (5, 8, 27) {real, imag} */,
  {32'h414d5601, 32'h413262ae} /* (5, 8, 26) {real, imag} */,
  {32'h41197b30, 32'h417cb568} /* (5, 8, 25) {real, imag} */,
  {32'hc1219344, 32'h410adec8} /* (5, 8, 24) {real, imag} */,
  {32'h406ed3b4, 32'hc1c9870d} /* (5, 8, 23) {real, imag} */,
  {32'hc13b29f2, 32'h40083ea6} /* (5, 8, 22) {real, imag} */,
  {32'hc10895d0, 32'hbfb520fc} /* (5, 8, 21) {real, imag} */,
  {32'hc07d75ec, 32'hc1aae442} /* (5, 8, 20) {real, imag} */,
  {32'hc02a7c90, 32'hbf0f4f8c} /* (5, 8, 19) {real, imag} */,
  {32'h40818228, 32'h4108c96f} /* (5, 8, 18) {real, imag} */,
  {32'hbfa28ffe, 32'hc0ff0ae5} /* (5, 8, 17) {real, imag} */,
  {32'h3fd50078, 32'h3d959f00} /* (5, 8, 16) {real, imag} */,
  {32'h408404e8, 32'h415579f0} /* (5, 8, 15) {real, imag} */,
  {32'hc1a46d56, 32'hbf438f70} /* (5, 8, 14) {real, imag} */,
  {32'h4108043d, 32'hc0145a0c} /* (5, 8, 13) {real, imag} */,
  {32'hc06032ec, 32'hc1176986} /* (5, 8, 12) {real, imag} */,
  {32'hc0806a5d, 32'hc06a46d8} /* (5, 8, 11) {real, imag} */,
  {32'h40a29406, 32'hbf96a530} /* (5, 8, 10) {real, imag} */,
  {32'h414b9567, 32'h41ea13d1} /* (5, 8, 9) {real, imag} */,
  {32'h41a2d6f9, 32'hc19d4ef0} /* (5, 8, 8) {real, imag} */,
  {32'h3e9451a0, 32'hc1c57def} /* (5, 8, 7) {real, imag} */,
  {32'h4156a992, 32'hc0034150} /* (5, 8, 6) {real, imag} */,
  {32'hc1b5eea0, 32'h41409eed} /* (5, 8, 5) {real, imag} */,
  {32'h40e6258a, 32'hc04b7efa} /* (5, 8, 4) {real, imag} */,
  {32'hc0b44206, 32'hc09a4529} /* (5, 8, 3) {real, imag} */,
  {32'h40f13ecb, 32'hc0ef1504} /* (5, 8, 2) {real, imag} */,
  {32'hc1112e80, 32'hc0f53e30} /* (5, 8, 1) {real, imag} */,
  {32'h41808bc4, 32'hbd7da380} /* (5, 8, 0) {real, imag} */,
  {32'h3fc581c8, 32'h4070a808} /* (5, 7, 31) {real, imag} */,
  {32'hc17d8e0f, 32'hc11ecef2} /* (5, 7, 30) {real, imag} */,
  {32'hc0e8f533, 32'hc08af9b9} /* (5, 7, 29) {real, imag} */,
  {32'hc1b87f12, 32'hc1a9df0d} /* (5, 7, 28) {real, imag} */,
  {32'hc194175a, 32'hc032148b} /* (5, 7, 27) {real, imag} */,
  {32'hbf1f5088, 32'hbfee2380} /* (5, 7, 26) {real, imag} */,
  {32'h41588aaa, 32'hc11614e8} /* (5, 7, 25) {real, imag} */,
  {32'hc1320a57, 32'h3f0d35c0} /* (5, 7, 24) {real, imag} */,
  {32'hc13261c1, 32'h4127cffe} /* (5, 7, 23) {real, imag} */,
  {32'h418c4dce, 32'h3e14a840} /* (5, 7, 22) {real, imag} */,
  {32'h40b31f54, 32'h41a4a22c} /* (5, 7, 21) {real, imag} */,
  {32'h41a3d00a, 32'hc1357b93} /* (5, 7, 20) {real, imag} */,
  {32'hc155d0e7, 32'h3f7dc1bc} /* (5, 7, 19) {real, imag} */,
  {32'h40c6bf23, 32'h406a803c} /* (5, 7, 18) {real, imag} */,
  {32'h40e1d406, 32'h3fcc68ca} /* (5, 7, 17) {real, imag} */,
  {32'hbc0ca000, 32'hc0f862e6} /* (5, 7, 16) {real, imag} */,
  {32'hc108002e, 32'h412a0ed7} /* (5, 7, 15) {real, imag} */,
  {32'hc1920707, 32'hc0d3b173} /* (5, 7, 14) {real, imag} */,
  {32'hc157c307, 32'h40a89e3a} /* (5, 7, 13) {real, imag} */,
  {32'hc05b13d8, 32'hc046b91b} /* (5, 7, 12) {real, imag} */,
  {32'hc0691222, 32'h3f765400} /* (5, 7, 11) {real, imag} */,
  {32'h4161f372, 32'h41a52934} /* (5, 7, 10) {real, imag} */,
  {32'h41393cf0, 32'h40a35dd0} /* (5, 7, 9) {real, imag} */,
  {32'h40eecada, 32'hc10f0c44} /* (5, 7, 8) {real, imag} */,
  {32'hbce74b00, 32'hc0c71e1a} /* (5, 7, 7) {real, imag} */,
  {32'h41719e32, 32'h410074f6} /* (5, 7, 6) {real, imag} */,
  {32'h40f39498, 32'h41d53d65} /* (5, 7, 5) {real, imag} */,
  {32'h409e4d49, 32'h407467e9} /* (5, 7, 4) {real, imag} */,
  {32'hc15cdeb8, 32'hc10c5c02} /* (5, 7, 3) {real, imag} */,
  {32'hc036ac94, 32'h41a84746} /* (5, 7, 2) {real, imag} */,
  {32'hc0c04a2c, 32'hc0c12c74} /* (5, 7, 1) {real, imag} */,
  {32'hc1cd6622, 32'hc13f51a2} /* (5, 7, 0) {real, imag} */,
  {32'h41198fc4, 32'h418085d1} /* (5, 6, 31) {real, imag} */,
  {32'hc1513f72, 32'hc0ddfb50} /* (5, 6, 30) {real, imag} */,
  {32'h4159d75c, 32'hc07818f2} /* (5, 6, 29) {real, imag} */,
  {32'h40a46f0c, 32'h4048b702} /* (5, 6, 28) {real, imag} */,
  {32'h411fd09a, 32'h411117ca} /* (5, 6, 27) {real, imag} */,
  {32'hc0d43026, 32'hc1228410} /* (5, 6, 26) {real, imag} */,
  {32'h3fbe8ef0, 32'h41bf54c4} /* (5, 6, 25) {real, imag} */,
  {32'hc09a1248, 32'hc10a33c2} /* (5, 6, 24) {real, imag} */,
  {32'hc1320f12, 32'h4003fec0} /* (5, 6, 23) {real, imag} */,
  {32'hc0c10445, 32'h411a4a3e} /* (5, 6, 22) {real, imag} */,
  {32'hc1128324, 32'hbf922710} /* (5, 6, 21) {real, imag} */,
  {32'hc0b51ba0, 32'hc0038da6} /* (5, 6, 20) {real, imag} */,
  {32'h41041f64, 32'h40ec22ca} /* (5, 6, 19) {real, imag} */,
  {32'h40da7398, 32'h40b755c4} /* (5, 6, 18) {real, imag} */,
  {32'hc141dec0, 32'hc0e73c00} /* (5, 6, 17) {real, imag} */,
  {32'h411d9664, 32'hc09e84f9} /* (5, 6, 16) {real, imag} */,
  {32'hc0b5093c, 32'hbf1d8fb0} /* (5, 6, 15) {real, imag} */,
  {32'h411e5949, 32'h4110a921} /* (5, 6, 14) {real, imag} */,
  {32'hbf6ebc44, 32'h402115cc} /* (5, 6, 13) {real, imag} */,
  {32'h41776cf8, 32'hc11fda51} /* (5, 6, 12) {real, imag} */,
  {32'hc0b4b2c8, 32'h41ca9f41} /* (5, 6, 11) {real, imag} */,
  {32'h4171ac8c, 32'h40335291} /* (5, 6, 10) {real, imag} */,
  {32'h403e11b5, 32'hc15b7dc6} /* (5, 6, 9) {real, imag} */,
  {32'hc16656ca, 32'hc11d9254} /* (5, 6, 8) {real, imag} */,
  {32'h41b0b280, 32'h414b180e} /* (5, 6, 7) {real, imag} */,
  {32'hc1665fb4, 32'h415859f0} /* (5, 6, 6) {real, imag} */,
  {32'hc082b7ec, 32'h4133b206} /* (5, 6, 5) {real, imag} */,
  {32'hc076ee08, 32'h40edf240} /* (5, 6, 4) {real, imag} */,
  {32'hc190c6c7, 32'hc1d18a6a} /* (5, 6, 3) {real, imag} */,
  {32'hc1a7baa6, 32'hc1147dc7} /* (5, 6, 2) {real, imag} */,
  {32'hc0c7c574, 32'h4111f4fc} /* (5, 6, 1) {real, imag} */,
  {32'h41dfb55f, 32'h4019fc88} /* (5, 6, 0) {real, imag} */,
  {32'h41d3eb6e, 32'h424bbef5} /* (5, 5, 31) {real, imag} */,
  {32'hc117236a, 32'hc116ccb4} /* (5, 5, 30) {real, imag} */,
  {32'hc1aa7356, 32'hc18ffdd3} /* (5, 5, 29) {real, imag} */,
  {32'hc1255a2d, 32'hc09cb3a8} /* (5, 5, 28) {real, imag} */,
  {32'hc18e1474, 32'h418cc338} /* (5, 5, 27) {real, imag} */,
  {32'h41043aba, 32'h419c612a} /* (5, 5, 26) {real, imag} */,
  {32'h408c633e, 32'h40b357cb} /* (5, 5, 25) {real, imag} */,
  {32'hc206198c, 32'h40f13ff4} /* (5, 5, 24) {real, imag} */,
  {32'hc0e48fd3, 32'h4171ab4c} /* (5, 5, 23) {real, imag} */,
  {32'hc1894323, 32'hc1a47f57} /* (5, 5, 22) {real, imag} */,
  {32'hc0951511, 32'hc1350d00} /* (5, 5, 21) {real, imag} */,
  {32'hc0f9b317, 32'hc1242bfc} /* (5, 5, 20) {real, imag} */,
  {32'hc197544b, 32'h4124f7b0} /* (5, 5, 19) {real, imag} */,
  {32'hc129bb6a, 32'h3fdc5dd0} /* (5, 5, 18) {real, imag} */,
  {32'hbf723f26, 32'hc0d8b7c0} /* (5, 5, 17) {real, imag} */,
  {32'h403c5b44, 32'h400bc834} /* (5, 5, 16) {real, imag} */,
  {32'hc0c37a24, 32'h3f4e99d0} /* (5, 5, 15) {real, imag} */,
  {32'h4110f440, 32'h3fa79ab0} /* (5, 5, 14) {real, imag} */,
  {32'h4143b0f5, 32'h4172e301} /* (5, 5, 13) {real, imag} */,
  {32'h4065d141, 32'h3f852890} /* (5, 5, 12) {real, imag} */,
  {32'h4129aed5, 32'hc0e43aae} /* (5, 5, 11) {real, imag} */,
  {32'h400bf216, 32'h418b22d7} /* (5, 5, 10) {real, imag} */,
  {32'hc13c02c4, 32'h406bb5b2} /* (5, 5, 9) {real, imag} */,
  {32'h408314cb, 32'h3f304f04} /* (5, 5, 8) {real, imag} */,
  {32'hc1100a19, 32'hc09db134} /* (5, 5, 7) {real, imag} */,
  {32'h4119459e, 32'hc0f6ff96} /* (5, 5, 6) {real, imag} */,
  {32'hc1a5ea98, 32'h40b13d60} /* (5, 5, 5) {real, imag} */,
  {32'hc1ac5ab0, 32'h40f5a5a7} /* (5, 5, 4) {real, imag} */,
  {32'h41921aa2, 32'h4015bdc8} /* (5, 5, 3) {real, imag} */,
  {32'hc0335e44, 32'h41a8c87a} /* (5, 5, 2) {real, imag} */,
  {32'h41b0f85b, 32'h40c2a416} /* (5, 5, 1) {real, imag} */,
  {32'h414555c0, 32'h413d4a1d} /* (5, 5, 0) {real, imag} */,
  {32'hc1bdc213, 32'hc1da51e3} /* (5, 4, 31) {real, imag} */,
  {32'h40963ce8, 32'h41cfc354} /* (5, 4, 30) {real, imag} */,
  {32'h4063e05d, 32'h3ed388e0} /* (5, 4, 29) {real, imag} */,
  {32'h404aacb2, 32'h41838016} /* (5, 4, 28) {real, imag} */,
  {32'h4123e4e8, 32'hc1b9a4fa} /* (5, 4, 27) {real, imag} */,
  {32'hc1b3df08, 32'hc123a6f8} /* (5, 4, 26) {real, imag} */,
  {32'h40833a1c, 32'h418ca0ee} /* (5, 4, 25) {real, imag} */,
  {32'h418513a0, 32'hc13f80f6} /* (5, 4, 24) {real, imag} */,
  {32'h409053ae, 32'h4028cc36} /* (5, 4, 23) {real, imag} */,
  {32'h40fc4804, 32'h40613fb9} /* (5, 4, 22) {real, imag} */,
  {32'h411d3956, 32'hc141769a} /* (5, 4, 21) {real, imag} */,
  {32'h411c0740, 32'h41b0f3f4} /* (5, 4, 20) {real, imag} */,
  {32'hc10757a0, 32'h40da7be6} /* (5, 4, 19) {real, imag} */,
  {32'hc1459a7d, 32'h40ec0dc0} /* (5, 4, 18) {real, imag} */,
  {32'h40d093aa, 32'h400f0679} /* (5, 4, 17) {real, imag} */,
  {32'hc0b5a500, 32'h40c0947a} /* (5, 4, 16) {real, imag} */,
  {32'hbf922ef4, 32'hc005d776} /* (5, 4, 15) {real, imag} */,
  {32'h411636c0, 32'h417555e4} /* (5, 4, 14) {real, imag} */,
  {32'hc17fb710, 32'hc0b45d8e} /* (5, 4, 13) {real, imag} */,
  {32'hc0f7a766, 32'h415d9f64} /* (5, 4, 12) {real, imag} */,
  {32'h416c92c8, 32'h4138d52b} /* (5, 4, 11) {real, imag} */,
  {32'h40b4f5f8, 32'hc1c12023} /* (5, 4, 10) {real, imag} */,
  {32'hc186559a, 32'hc02b3a16} /* (5, 4, 9) {real, imag} */,
  {32'h40c286f5, 32'h415bdea7} /* (5, 4, 8) {real, imag} */,
  {32'hc1a154e8, 32'hc01cf48c} /* (5, 4, 7) {real, imag} */,
  {32'hbff564a8, 32'h400440a2} /* (5, 4, 6) {real, imag} */,
  {32'h412869ff, 32'h4078d2e8} /* (5, 4, 5) {real, imag} */,
  {32'h41ac6584, 32'hc057dc70} /* (5, 4, 4) {real, imag} */,
  {32'hc1c0fcdb, 32'h41d55504} /* (5, 4, 3) {real, imag} */,
  {32'h41c95216, 32'hc14f0d84} /* (5, 4, 2) {real, imag} */,
  {32'hc29bb8b4, 32'h417eec40} /* (5, 4, 1) {real, imag} */,
  {32'h416cc939, 32'hc19148c0} /* (5, 4, 0) {real, imag} */,
  {32'h40e66eb8, 32'hc2321549} /* (5, 3, 31) {real, imag} */,
  {32'hc128df48, 32'hc2272ee2} /* (5, 3, 30) {real, imag} */,
  {32'h4000ca96, 32'h4165ae72} /* (5, 3, 29) {real, imag} */,
  {32'hc147d1a5, 32'h40685338} /* (5, 3, 28) {real, imag} */,
  {32'hc12280e9, 32'hc1a9ae8a} /* (5, 3, 27) {real, imag} */,
  {32'hc1d6869f, 32'hc0b1d670} /* (5, 3, 26) {real, imag} */,
  {32'hc148c62a, 32'h418575b2} /* (5, 3, 25) {real, imag} */,
  {32'h41b2f2b8, 32'hc080b4a0} /* (5, 3, 24) {real, imag} */,
  {32'h417f16f8, 32'hc066b7cc} /* (5, 3, 23) {real, imag} */,
  {32'hc03ab9b4, 32'hc0fd48bf} /* (5, 3, 22) {real, imag} */,
  {32'hc0646820, 32'h4107ea03} /* (5, 3, 21) {real, imag} */,
  {32'h41c25ffc, 32'hbea4ff00} /* (5, 3, 20) {real, imag} */,
  {32'h3fc381a2, 32'h4132229f} /* (5, 3, 19) {real, imag} */,
  {32'hc04af1af, 32'hc0322665} /* (5, 3, 18) {real, imag} */,
  {32'hc00b5172, 32'h409722b0} /* (5, 3, 17) {real, imag} */,
  {32'hc0e3e7d6, 32'hc02f8c2e} /* (5, 3, 16) {real, imag} */,
  {32'h413e8ced, 32'hc0502368} /* (5, 3, 15) {real, imag} */,
  {32'h40f27b56, 32'hc13bdd81} /* (5, 3, 14) {real, imag} */,
  {32'h4145e166, 32'h408737b9} /* (5, 3, 13) {real, imag} */,
  {32'hc0caedd3, 32'hc063fdbc} /* (5, 3, 12) {real, imag} */,
  {32'hc164a6f0, 32'hc184311a} /* (5, 3, 11) {real, imag} */,
  {32'h40b8ed07, 32'hc1035e4b} /* (5, 3, 10) {real, imag} */,
  {32'h3ea04300, 32'hc0cade51} /* (5, 3, 9) {real, imag} */,
  {32'hc0675284, 32'h4168f030} /* (5, 3, 8) {real, imag} */,
  {32'hc124e860, 32'hc1d88e82} /* (5, 3, 7) {real, imag} */,
  {32'h3f9133d8, 32'hc189c1ca} /* (5, 3, 6) {real, imag} */,
  {32'hc139ce16, 32'hc12959d8} /* (5, 3, 5) {real, imag} */,
  {32'h4119a51e, 32'h40f2991e} /* (5, 3, 4) {real, imag} */,
  {32'hc11be700, 32'h41304cda} /* (5, 3, 3) {real, imag} */,
  {32'h420ccf79, 32'h428f49d4} /* (5, 3, 2) {real, imag} */,
  {32'h414dc5ec, 32'h42472d42} /* (5, 3, 1) {real, imag} */,
  {32'h4180fbc1, 32'h42502bfb} /* (5, 3, 0) {real, imag} */,
  {32'hc133b740, 32'h3fa13220} /* (5, 2, 31) {real, imag} */,
  {32'h41cc8e18, 32'hc120cfc0} /* (5, 2, 30) {real, imag} */,
  {32'h3ee8f2a0, 32'h41caec4b} /* (5, 2, 29) {real, imag} */,
  {32'h4148cbb6, 32'hc1a03f07} /* (5, 2, 28) {real, imag} */,
  {32'hc1fbb23d, 32'h409478f8} /* (5, 2, 27) {real, imag} */,
  {32'hc1ddc0ea, 32'h41a79de6} /* (5, 2, 26) {real, imag} */,
  {32'h415844fa, 32'hc119bcf4} /* (5, 2, 25) {real, imag} */,
  {32'h410a1216, 32'h4217f9fd} /* (5, 2, 24) {real, imag} */,
  {32'hbf922184, 32'hc03564d5} /* (5, 2, 23) {real, imag} */,
  {32'h40322634, 32'hc0dd055c} /* (5, 2, 22) {real, imag} */,
  {32'hc0bca46b, 32'h410931f6} /* (5, 2, 21) {real, imag} */,
  {32'h415c5e12, 32'h403bf454} /* (5, 2, 20) {real, imag} */,
  {32'hc08a04a7, 32'hc16593ee} /* (5, 2, 19) {real, imag} */,
  {32'hbfc4fca8, 32'hc063166a} /* (5, 2, 18) {real, imag} */,
  {32'h40c89513, 32'hc0e6a7aa} /* (5, 2, 17) {real, imag} */,
  {32'h40ad36a2, 32'hc077a9c0} /* (5, 2, 16) {real, imag} */,
  {32'hc0e9b948, 32'h40baa6bc} /* (5, 2, 15) {real, imag} */,
  {32'h3c983500, 32'hc0fa9fd2} /* (5, 2, 14) {real, imag} */,
  {32'hbf7721f6, 32'h3c96c400} /* (5, 2, 13) {real, imag} */,
  {32'h3f893194, 32'hc072a765} /* (5, 2, 12) {real, imag} */,
  {32'hc0850fc0, 32'hc105ed4b} /* (5, 2, 11) {real, imag} */,
  {32'hc13ba530, 32'h40a734c4} /* (5, 2, 10) {real, imag} */,
  {32'h408d99a5, 32'h41f2d973} /* (5, 2, 9) {real, imag} */,
  {32'h3fbc7780, 32'hc0781028} /* (5, 2, 8) {real, imag} */,
  {32'hc08e2d9e, 32'hc15ad9da} /* (5, 2, 7) {real, imag} */,
  {32'h40643a27, 32'h418aa4ce} /* (5, 2, 6) {real, imag} */,
  {32'h41d7b7b1, 32'hc20572b9} /* (5, 2, 5) {real, imag} */,
  {32'h40e9d564, 32'h41b7755f} /* (5, 2, 4) {real, imag} */,
  {32'hbf0c5e20, 32'h40d3845a} /* (5, 2, 3) {real, imag} */,
  {32'hc26434ce, 32'h42a33f10} /* (5, 2, 2) {real, imag} */,
  {32'h41b7f910, 32'h421e8910} /* (5, 2, 1) {real, imag} */,
  {32'hc294f34e, 32'hc26141c1} /* (5, 2, 0) {real, imag} */,
  {32'h4364b078, 32'hc2d6416a} /* (5, 1, 31) {real, imag} */,
  {32'h41b6ace0, 32'hbfa8e240} /* (5, 1, 30) {real, imag} */,
  {32'h42671a97, 32'hc1616697} /* (5, 1, 29) {real, imag} */,
  {32'h40abdf6e, 32'hc1bf581d} /* (5, 1, 28) {real, imag} */,
  {32'h418af44c, 32'h415f17a4} /* (5, 1, 27) {real, imag} */,
  {32'h41162453, 32'hc13b854e} /* (5, 1, 26) {real, imag} */,
  {32'hc22bb13e, 32'hc06b6a01} /* (5, 1, 25) {real, imag} */,
  {32'h40748864, 32'hc1145451} /* (5, 1, 24) {real, imag} */,
  {32'h4158dd67, 32'hc10f8268} /* (5, 1, 23) {real, imag} */,
  {32'hc072237e, 32'hc03cf99a} /* (5, 1, 22) {real, imag} */,
  {32'hc10faa5a, 32'h3dddf380} /* (5, 1, 21) {real, imag} */,
  {32'h40b23de7, 32'hc140ed13} /* (5, 1, 20) {real, imag} */,
  {32'h4003e909, 32'hc10817c7} /* (5, 1, 19) {real, imag} */,
  {32'hc08f312c, 32'hc130c575} /* (5, 1, 18) {real, imag} */,
  {32'h40476a4a, 32'hbeda9ad0} /* (5, 1, 17) {real, imag} */,
  {32'h40004ef8, 32'hc0b29433} /* (5, 1, 16) {real, imag} */,
  {32'h408d8ff3, 32'h40af6c15} /* (5, 1, 15) {real, imag} */,
  {32'h41177e17, 32'hc129c5c3} /* (5, 1, 14) {real, imag} */,
  {32'h4123cbba, 32'h40974527} /* (5, 1, 13) {real, imag} */,
  {32'h40ce8303, 32'hc01a8872} /* (5, 1, 12) {real, imag} */,
  {32'h41592f8f, 32'hc142139a} /* (5, 1, 11) {real, imag} */,
  {32'hc10c54b5, 32'hc1238f9a} /* (5, 1, 10) {real, imag} */,
  {32'hc189c200, 32'h415b87cb} /* (5, 1, 9) {real, imag} */,
  {32'h41da4d77, 32'h40e83474} /* (5, 1, 8) {real, imag} */,
  {32'hc0a5dcbc, 32'h41858868} /* (5, 1, 7) {real, imag} */,
  {32'hc1aee3e4, 32'hc14e317d} /* (5, 1, 6) {real, imag} */,
  {32'hc12e5fb8, 32'h41b8a617} /* (5, 1, 5) {real, imag} */,
  {32'h41cad6a5, 32'hc20f0810} /* (5, 1, 4) {real, imag} */,
  {32'hc10d3652, 32'hc25c2658} /* (5, 1, 3) {real, imag} */,
  {32'hc0d733e0, 32'hc160f640} /* (5, 1, 2) {real, imag} */,
  {32'h43bdb712, 32'h426e91b4} /* (5, 1, 1) {real, imag} */,
  {32'h440da16e, 32'h431b2d54} /* (5, 1, 0) {real, imag} */,
  {32'h438356ac, 32'hc3793bbd} /* (5, 0, 31) {real, imag} */,
  {32'h41c3ad50, 32'h423c8958} /* (5, 0, 30) {real, imag} */,
  {32'h42add7ae, 32'hc271b01a} /* (5, 0, 29) {real, imag} */,
  {32'hc0b71328, 32'hc207e979} /* (5, 0, 28) {real, imag} */,
  {32'hc09187dc, 32'h41467ab6} /* (5, 0, 27) {real, imag} */,
  {32'h421dceac, 32'h40a16244} /* (5, 0, 26) {real, imag} */,
  {32'h3ffa7ad0, 32'h411f5024} /* (5, 0, 25) {real, imag} */,
  {32'h3e2b5990, 32'hc1d52410} /* (5, 0, 24) {real, imag} */,
  {32'hbfb75518, 32'h41e67ff8} /* (5, 0, 23) {real, imag} */,
  {32'hc19fab31, 32'h418ff853} /* (5, 0, 22) {real, imag} */,
  {32'hc1381530, 32'h408008e0} /* (5, 0, 21) {real, imag} */,
  {32'hc1a2b0b6, 32'h3e8047b0} /* (5, 0, 20) {real, imag} */,
  {32'hc0bf891d, 32'h41084f85} /* (5, 0, 19) {real, imag} */,
  {32'hbf553c18, 32'h4127789c} /* (5, 0, 18) {real, imag} */,
  {32'hc12fc400, 32'h40b80350} /* (5, 0, 17) {real, imag} */,
  {32'hc1396b34, 32'h00000000} /* (5, 0, 16) {real, imag} */,
  {32'hc12fc400, 32'hc0b80350} /* (5, 0, 15) {real, imag} */,
  {32'hbf553c18, 32'hc127789c} /* (5, 0, 14) {real, imag} */,
  {32'hc0bf891d, 32'hc1084f85} /* (5, 0, 13) {real, imag} */,
  {32'hc1a2b0b6, 32'hbe8047b0} /* (5, 0, 12) {real, imag} */,
  {32'hc1381530, 32'hc08008e0} /* (5, 0, 11) {real, imag} */,
  {32'hc19fab31, 32'hc18ff853} /* (5, 0, 10) {real, imag} */,
  {32'hbfb75518, 32'hc1e67ff8} /* (5, 0, 9) {real, imag} */,
  {32'h3e2b5990, 32'h41d52410} /* (5, 0, 8) {real, imag} */,
  {32'h3ffa7ad0, 32'hc11f5024} /* (5, 0, 7) {real, imag} */,
  {32'h421dceac, 32'hc0a16244} /* (5, 0, 6) {real, imag} */,
  {32'hc09187dc, 32'hc1467ab6} /* (5, 0, 5) {real, imag} */,
  {32'hc0b71328, 32'h4207e979} /* (5, 0, 4) {real, imag} */,
  {32'h42add7ae, 32'h4271b01a} /* (5, 0, 3) {real, imag} */,
  {32'h41c3ad50, 32'hc23c8958} /* (5, 0, 2) {real, imag} */,
  {32'h438356ac, 32'h43793bbd} /* (5, 0, 1) {real, imag} */,
  {32'h4476a686, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hc3bb4b8d, 32'h43ad18d3} /* (4, 31, 31) {real, imag} */,
  {32'h436356ee, 32'hc33bd49a} /* (4, 31, 30) {real, imag} */,
  {32'h414bffd6, 32'h424b2118} /* (4, 31, 29) {real, imag} */,
  {32'h409f04c4, 32'h4223ec2c} /* (4, 31, 28) {real, imag} */,
  {32'h4278e9ef, 32'hc1d3ca10} /* (4, 31, 27) {real, imag} */,
  {32'hc1b11f6b, 32'h41cbc0dd} /* (4, 31, 26) {real, imag} */,
  {32'hc16b9284, 32'h40351bf0} /* (4, 31, 25) {real, imag} */,
  {32'h3f874130, 32'hc2164f38} /* (4, 31, 24) {real, imag} */,
  {32'hc1aba055, 32'hc185b886} /* (4, 31, 23) {real, imag} */,
  {32'h4100b80e, 32'hc071e4ad} /* (4, 31, 22) {real, imag} */,
  {32'hc0bbadc9, 32'hc18922e1} /* (4, 31, 21) {real, imag} */,
  {32'hc06e09ec, 32'h40ad394b} /* (4, 31, 20) {real, imag} */,
  {32'h40b73c2e, 32'h405aeacf} /* (4, 31, 19) {real, imag} */,
  {32'hc1c63230, 32'hc191c066} /* (4, 31, 18) {real, imag} */,
  {32'h4139a562, 32'hc01c5e2a} /* (4, 31, 17) {real, imag} */,
  {32'hc1563d96, 32'h4107be28} /* (4, 31, 16) {real, imag} */,
  {32'h411b17d8, 32'hc127b11e} /* (4, 31, 15) {real, imag} */,
  {32'h4096341b, 32'h418e4304} /* (4, 31, 14) {real, imag} */,
  {32'h40b40592, 32'h40c212ce} /* (4, 31, 13) {real, imag} */,
  {32'h40614bda, 32'hc05941ec} /* (4, 31, 12) {real, imag} */,
  {32'h41bf87c2, 32'h410fe028} /* (4, 31, 11) {real, imag} */,
  {32'hc0ad9324, 32'h418bf683} /* (4, 31, 10) {real, imag} */,
  {32'hc088855e, 32'hc01f0d88} /* (4, 31, 9) {real, imag} */,
  {32'h41bacac0, 32'h414b082a} /* (4, 31, 8) {real, imag} */,
  {32'hc1c1b6c6, 32'h407e6a5a} /* (4, 31, 7) {real, imag} */,
  {32'h4176b5ca, 32'h418101b6} /* (4, 31, 6) {real, imag} */,
  {32'h42cb796e, 32'hc0a90a2e} /* (4, 31, 5) {real, imag} */,
  {32'hc25eee70, 32'h428f469a} /* (4, 31, 4) {real, imag} */,
  {32'h42482ec2, 32'h4220f71e} /* (4, 31, 3) {real, imag} */,
  {32'h43268dc8, 32'hc1fc72eb} /* (4, 31, 2) {real, imag} */,
  {32'hc3931668, 32'hc19a93d0} /* (4, 31, 1) {real, imag} */,
  {32'hc1a2e928, 32'hc25fb30c} /* (4, 31, 0) {real, imag} */,
  {32'h4389ad3f, 32'hbfe65600} /* (4, 30, 31) {real, imag} */,
  {32'hc3631e4d, 32'hc2f92c8a} /* (4, 30, 30) {real, imag} */,
  {32'hc17a7a2c, 32'hc114b956} /* (4, 30, 29) {real, imag} */,
  {32'h42b5abc9, 32'hc0a026fe} /* (4, 30, 28) {real, imag} */,
  {32'hc1a71aba, 32'h42713038} /* (4, 30, 27) {real, imag} */,
  {32'h4138a4d6, 32'hc18b1eda} /* (4, 30, 26) {real, imag} */,
  {32'h41b1302c, 32'h40e13a6d} /* (4, 30, 25) {real, imag} */,
  {32'hc1f238c7, 32'h4146e651} /* (4, 30, 24) {real, imag} */,
  {32'h40bc9e98, 32'hc09f63ce} /* (4, 30, 23) {real, imag} */,
  {32'h410ce546, 32'hc1ad22cf} /* (4, 30, 22) {real, imag} */,
  {32'hc11bf068, 32'h412c79e1} /* (4, 30, 21) {real, imag} */,
  {32'h41347e97, 32'hc11c15f8} /* (4, 30, 20) {real, imag} */,
  {32'hc0bd1688, 32'h408bf04b} /* (4, 30, 19) {real, imag} */,
  {32'hc098bb90, 32'h419c22a7} /* (4, 30, 18) {real, imag} */,
  {32'h409adc31, 32'hc13aa487} /* (4, 30, 17) {real, imag} */,
  {32'h40e6aef0, 32'h40d2a889} /* (4, 30, 16) {real, imag} */,
  {32'hbfa36e56, 32'h418d98d2} /* (4, 30, 15) {real, imag} */,
  {32'h409776e0, 32'hc0690e34} /* (4, 30, 14) {real, imag} */,
  {32'hc0667f96, 32'h410bb15a} /* (4, 30, 13) {real, imag} */,
  {32'h412518f8, 32'h40616509} /* (4, 30, 12) {real, imag} */,
  {32'hc1276fd4, 32'hc1a028fa} /* (4, 30, 11) {real, imag} */,
  {32'h3f00fd80, 32'hc124ad02} /* (4, 30, 10) {real, imag} */,
  {32'hc122c4dc, 32'hc0a27409} /* (4, 30, 9) {real, imag} */,
  {32'hc121c3ec, 32'hc27ee26a} /* (4, 30, 8) {real, imag} */,
  {32'h410819cc, 32'h420ac40f} /* (4, 30, 7) {real, imag} */,
  {32'hc1d336de, 32'hc1ff7bee} /* (4, 30, 6) {real, imag} */,
  {32'hc2477ed0, 32'hc1a7ce8e} /* (4, 30, 5) {real, imag} */,
  {32'h411b3a96, 32'h428ba956} /* (4, 30, 4) {real, imag} */,
  {32'h3f76fe20, 32'hc1f4cdb0} /* (4, 30, 3) {real, imag} */,
  {32'hc36d9e45, 32'hc24bfea8} /* (4, 30, 2) {real, imag} */,
  {32'h43eccb8f, 32'hc1e09371} /* (4, 30, 1) {real, imag} */,
  {32'h432f23e6, 32'hc10f84c4} /* (4, 30, 0) {real, imag} */,
  {32'hc2978967, 32'hc12990d8} /* (4, 29, 31) {real, imag} */,
  {32'h415b17d7, 32'hc2e13b1e} /* (4, 29, 30) {real, imag} */,
  {32'hc10f8a99, 32'h418e8801} /* (4, 29, 29) {real, imag} */,
  {32'h41d50140, 32'h41be00e3} /* (4, 29, 28) {real, imag} */,
  {32'hc1daba0f, 32'h411c7bec} /* (4, 29, 27) {real, imag} */,
  {32'h3e685580, 32'h4126a326} /* (4, 29, 26) {real, imag} */,
  {32'hc091466c, 32'h41f8531c} /* (4, 29, 25) {real, imag} */,
  {32'h3f552ca8, 32'hc1670325} /* (4, 29, 24) {real, imag} */,
  {32'hc0aa23b5, 32'h4052ad2c} /* (4, 29, 23) {real, imag} */,
  {32'h3f945574, 32'h408afe0c} /* (4, 29, 22) {real, imag} */,
  {32'hc1704451, 32'h4084d772} /* (4, 29, 21) {real, imag} */,
  {32'h411e4222, 32'h411d30db} /* (4, 29, 20) {real, imag} */,
  {32'h411d5c2e, 32'hc04cbda8} /* (4, 29, 19) {real, imag} */,
  {32'hbfb58f34, 32'hc152fef7} /* (4, 29, 18) {real, imag} */,
  {32'h4096a47c, 32'hbe8ec6a8} /* (4, 29, 17) {real, imag} */,
  {32'h411a36fe, 32'h4128093b} /* (4, 29, 16) {real, imag} */,
  {32'h411d0c24, 32'hc037d1b9} /* (4, 29, 15) {real, imag} */,
  {32'hc196f64a, 32'h40631ac6} /* (4, 29, 14) {real, imag} */,
  {32'hc0f9d999, 32'h40d17123} /* (4, 29, 13) {real, imag} */,
  {32'h3fcae430, 32'h3e49e8f4} /* (4, 29, 12) {real, imag} */,
  {32'hc1273458, 32'h40fa333c} /* (4, 29, 11) {real, imag} */,
  {32'h41301c06, 32'h417bac9d} /* (4, 29, 10) {real, imag} */,
  {32'hc0a0fa2c, 32'h41979d86} /* (4, 29, 9) {real, imag} */,
  {32'h4078f89e, 32'hc1b2c1a8} /* (4, 29, 8) {real, imag} */,
  {32'hc0f9a733, 32'hc151590e} /* (4, 29, 7) {real, imag} */,
  {32'hc0fd5344, 32'h416bf55c} /* (4, 29, 6) {real, imag} */,
  {32'h42017646, 32'h41c49091} /* (4, 29, 5) {real, imag} */,
  {32'hc1cb52c6, 32'h4138f8bd} /* (4, 29, 4) {real, imag} */,
  {32'hbef56a00, 32'hc10f23ed} /* (4, 29, 3) {real, imag} */,
  {32'hc23ae113, 32'hc20d1e00} /* (4, 29, 2) {real, imag} */,
  {32'h42a89fe7, 32'h42597180} /* (4, 29, 1) {real, imag} */,
  {32'h4153a6a1, 32'hc1ccb1aa} /* (4, 29, 0) {real, imag} */,
  {32'hc318991c, 32'h424626ac} /* (4, 28, 31) {real, imag} */,
  {32'h42b21df1, 32'hc24393a6} /* (4, 28, 30) {real, imag} */,
  {32'hc19e1673, 32'hc1e59480} /* (4, 28, 29) {real, imag} */,
  {32'h41b820bc, 32'h41875424} /* (4, 28, 28) {real, imag} */,
  {32'h41a74907, 32'h40bdd40c} /* (4, 28, 27) {real, imag} */,
  {32'h405ecf00, 32'h412c1a5e} /* (4, 28, 26) {real, imag} */,
  {32'hc1a56632, 32'hc0d1664a} /* (4, 28, 25) {real, imag} */,
  {32'h40348c1a, 32'hc10dd106} /* (4, 28, 24) {real, imag} */,
  {32'hbefef2d0, 32'hc156adb8} /* (4, 28, 23) {real, imag} */,
  {32'h4144f75c, 32'h4159ae4a} /* (4, 28, 22) {real, imag} */,
  {32'hbedfd01c, 32'h4128f18f} /* (4, 28, 21) {real, imag} */,
  {32'hbf28b274, 32'h3eeca9c0} /* (4, 28, 20) {real, imag} */,
  {32'hc08385e5, 32'h401add16} /* (4, 28, 19) {real, imag} */,
  {32'hc0479f21, 32'hc1515276} /* (4, 28, 18) {real, imag} */,
  {32'hc0fb58e8, 32'h3fa74958} /* (4, 28, 17) {real, imag} */,
  {32'hc0cf493b, 32'h40fd1e16} /* (4, 28, 16) {real, imag} */,
  {32'hc03e688e, 32'hc13b3a58} /* (4, 28, 15) {real, imag} */,
  {32'h3d8bd940, 32'hc0d4eab6} /* (4, 28, 14) {real, imag} */,
  {32'h40d7c127, 32'h40aafcbc} /* (4, 28, 13) {real, imag} */,
  {32'hc091bdc4, 32'hc089679a} /* (4, 28, 12) {real, imag} */,
  {32'h41f2c0ca, 32'h40fdac7d} /* (4, 28, 11) {real, imag} */,
  {32'h412dcdbb, 32'h4057924f} /* (4, 28, 10) {real, imag} */,
  {32'h3fa460c8, 32'hc07ec0db} /* (4, 28, 9) {real, imag} */,
  {32'h4116f687, 32'h3eb75778} /* (4, 28, 8) {real, imag} */,
  {32'h4113b0b0, 32'hbe09ec20} /* (4, 28, 7) {real, imag} */,
  {32'hc223cb80, 32'h41398b2c} /* (4, 28, 6) {real, imag} */,
  {32'h3faa71c2, 32'h416c7ef0} /* (4, 28, 5) {real, imag} */,
  {32'hc18fc2ba, 32'hc0f3c6e3} /* (4, 28, 4) {real, imag} */,
  {32'hc0c83d1a, 32'hc0f2d4fc} /* (4, 28, 3) {real, imag} */,
  {32'h42291cb5, 32'hc2b9daec} /* (4, 28, 2) {real, imag} */,
  {32'hc2223b39, 32'h42a4f48e} /* (4, 28, 1) {real, imag} */,
  {32'hc237cfd6, 32'h41204cc8} /* (4, 28, 0) {real, imag} */,
  {32'h42a47c5e, 32'hc2217a40} /* (4, 27, 31) {real, imag} */,
  {32'h40f9080c, 32'hc1c62afb} /* (4, 27, 30) {real, imag} */,
  {32'h41a8b277, 32'hc0641184} /* (4, 27, 29) {real, imag} */,
  {32'h418ac180, 32'h40f32361} /* (4, 27, 28) {real, imag} */,
  {32'hc1cd0fde, 32'h41f5e207} /* (4, 27, 27) {real, imag} */,
  {32'hc12a11f4, 32'h415aaea5} /* (4, 27, 26) {real, imag} */,
  {32'hbf94a736, 32'hc09b60f2} /* (4, 27, 25) {real, imag} */,
  {32'h404c4244, 32'h4048e5ae} /* (4, 27, 24) {real, imag} */,
  {32'hbed7a1f0, 32'hbfb3ff90} /* (4, 27, 23) {real, imag} */,
  {32'h40dbab23, 32'hc18dbbd8} /* (4, 27, 22) {real, imag} */,
  {32'hc055cc9e, 32'h41d22e0e} /* (4, 27, 21) {real, imag} */,
  {32'hc0984681, 32'hc04bee1c} /* (4, 27, 20) {real, imag} */,
  {32'hc050a042, 32'h412a4d8f} /* (4, 27, 19) {real, imag} */,
  {32'h412a229e, 32'h40df34f4} /* (4, 27, 18) {real, imag} */,
  {32'h40e91b94, 32'h40a48f20} /* (4, 27, 17) {real, imag} */,
  {32'hc007ff72, 32'hc1024680} /* (4, 27, 16) {real, imag} */,
  {32'hc0e1e64c, 32'hc0f4062e} /* (4, 27, 15) {real, imag} */,
  {32'h412fd40e, 32'hc0e0cafe} /* (4, 27, 14) {real, imag} */,
  {32'hc13a10a6, 32'hbfa54dc0} /* (4, 27, 13) {real, imag} */,
  {32'hc0ede98c, 32'hc08eaf0e} /* (4, 27, 12) {real, imag} */,
  {32'hc10a65c0, 32'hc1e962b4} /* (4, 27, 11) {real, imag} */,
  {32'hc0076fa0, 32'hbf15ce48} /* (4, 27, 10) {real, imag} */,
  {32'h40b5de95, 32'h41610bf2} /* (4, 27, 9) {real, imag} */,
  {32'hc10a68f8, 32'h3fcbb67e} /* (4, 27, 8) {real, imag} */,
  {32'h41c45c7e, 32'hc127cbc8} /* (4, 27, 7) {real, imag} */,
  {32'hc11a5dea, 32'hc1295625} /* (4, 27, 6) {real, imag} */,
  {32'hc1a819a3, 32'h40999575} /* (4, 27, 5) {real, imag} */,
  {32'h41ba9428, 32'h41af9882} /* (4, 27, 4) {real, imag} */,
  {32'hc03b7eaa, 32'h413b7e25} /* (4, 27, 3) {real, imag} */,
  {32'hc22feab3, 32'h414d9c0a} /* (4, 27, 2) {real, imag} */,
  {32'h425a6421, 32'hc1b24c80} /* (4, 27, 1) {real, imag} */,
  {32'h42a3bf55, 32'h40b2cd1c} /* (4, 27, 0) {real, imag} */,
  {32'h4188b211, 32'hc144fc49} /* (4, 26, 31) {real, imag} */,
  {32'hc1ae8ad9, 32'h40891fca} /* (4, 26, 30) {real, imag} */,
  {32'hc134a0be, 32'hc0c159b7} /* (4, 26, 29) {real, imag} */,
  {32'hc0b9af60, 32'h411a5db0} /* (4, 26, 28) {real, imag} */,
  {32'hc09d9fa9, 32'hc0c1d63a} /* (4, 26, 27) {real, imag} */,
  {32'hc1a2dcb0, 32'h411ad7a4} /* (4, 26, 26) {real, imag} */,
  {32'h412255d4, 32'hc1340a5b} /* (4, 26, 25) {real, imag} */,
  {32'hc1aaf1fe, 32'h3f48a370} /* (4, 26, 24) {real, imag} */,
  {32'h40cf6151, 32'h3f319528} /* (4, 26, 23) {real, imag} */,
  {32'h3f3c4608, 32'h40493292} /* (4, 26, 22) {real, imag} */,
  {32'hc14d18c7, 32'hc0d4a510} /* (4, 26, 21) {real, imag} */,
  {32'h40ecc65e, 32'hc0658426} /* (4, 26, 20) {real, imag} */,
  {32'h4180fb91, 32'h407e01a6} /* (4, 26, 19) {real, imag} */,
  {32'hbfcd22e8, 32'h4145f147} /* (4, 26, 18) {real, imag} */,
  {32'hbed222a8, 32'hc007ce34} /* (4, 26, 17) {real, imag} */,
  {32'h400cfa67, 32'h4095ce90} /* (4, 26, 16) {real, imag} */,
  {32'h40f2f80c, 32'h4028b098} /* (4, 26, 15) {real, imag} */,
  {32'h407843ba, 32'hbf3136bc} /* (4, 26, 14) {real, imag} */,
  {32'hc0c69ca9, 32'h40912fe4} /* (4, 26, 13) {real, imag} */,
  {32'hc1a9831d, 32'hc0d13631} /* (4, 26, 12) {real, imag} */,
  {32'hc0f6a4e3, 32'h41a0ff26} /* (4, 26, 11) {real, imag} */,
  {32'hc0868bab, 32'hc1836a8e} /* (4, 26, 10) {real, imag} */,
  {32'hc16b0d7a, 32'h4098251d} /* (4, 26, 9) {real, imag} */,
  {32'hc1092ce3, 32'hc1474fc6} /* (4, 26, 8) {real, imag} */,
  {32'hbf4943f4, 32'h41125770} /* (4, 26, 7) {real, imag} */,
  {32'hbfde71a8, 32'h40ecfeaa} /* (4, 26, 6) {real, imag} */,
  {32'h3fb00010, 32'hc19e2a76} /* (4, 26, 5) {real, imag} */,
  {32'h400c20e0, 32'h3f883090} /* (4, 26, 4) {real, imag} */,
  {32'h41b2089d, 32'hbf3828b0} /* (4, 26, 3) {real, imag} */,
  {32'h415b9333, 32'hbec951e0} /* (4, 26, 2) {real, imag} */,
  {32'h418566bc, 32'hc1a71802} /* (4, 26, 1) {real, imag} */,
  {32'h4151757b, 32'h41926d0f} /* (4, 26, 0) {real, imag} */,
  {32'h3e229c00, 32'h41de5ed0} /* (4, 25, 31) {real, imag} */,
  {32'h4196639d, 32'hc1253c32} /* (4, 25, 30) {real, imag} */,
  {32'hbe76f0c0, 32'hc1067624} /* (4, 25, 29) {real, imag} */,
  {32'hc16db3c9, 32'h414112b2} /* (4, 25, 28) {real, imag} */,
  {32'h4209f01a, 32'hc1c63306} /* (4, 25, 27) {real, imag} */,
  {32'h411e4c54, 32'hc02cc3eb} /* (4, 25, 26) {real, imag} */,
  {32'hc1988057, 32'hc11e5b11} /* (4, 25, 25) {real, imag} */,
  {32'h40ae003e, 32'h3f775d50} /* (4, 25, 24) {real, imag} */,
  {32'h412b1276, 32'hc03bbd5c} /* (4, 25, 23) {real, imag} */,
  {32'h40a70dfa, 32'h40ca626a} /* (4, 25, 22) {real, imag} */,
  {32'hc0ae9a42, 32'hc1357e0f} /* (4, 25, 21) {real, imag} */,
  {32'hc1ade3e2, 32'hc0293420} /* (4, 25, 20) {real, imag} */,
  {32'hc19e20eb, 32'hc130b5a8} /* (4, 25, 19) {real, imag} */,
  {32'hc1714e8a, 32'h3f4ad230} /* (4, 25, 18) {real, imag} */,
  {32'hc1601659, 32'h418135a8} /* (4, 25, 17) {real, imag} */,
  {32'h4159987f, 32'h406a32b2} /* (4, 25, 16) {real, imag} */,
  {32'hbf603174, 32'hc1219cce} /* (4, 25, 15) {real, imag} */,
  {32'h417a3896, 32'h40d5b06f} /* (4, 25, 14) {real, imag} */,
  {32'hc0d06284, 32'hc1764ad2} /* (4, 25, 13) {real, imag} */,
  {32'h411cd558, 32'h40a34132} /* (4, 25, 12) {real, imag} */,
  {32'hc0a2fec1, 32'hc1807f1a} /* (4, 25, 11) {real, imag} */,
  {32'hbfe918f8, 32'h4125e41c} /* (4, 25, 10) {real, imag} */,
  {32'hbfbd584e, 32'hc1532650} /* (4, 25, 9) {real, imag} */,
  {32'hc1537006, 32'h4191a78a} /* (4, 25, 8) {real, imag} */,
  {32'h4078483a, 32'h40bd772a} /* (4, 25, 7) {real, imag} */,
  {32'h412e43f3, 32'h40e014c9} /* (4, 25, 6) {real, imag} */,
  {32'h41a061da, 32'hc0dc7b8c} /* (4, 25, 5) {real, imag} */,
  {32'hc18f8df0, 32'h41b938dc} /* (4, 25, 4) {real, imag} */,
  {32'hc1150396, 32'h41357b46} /* (4, 25, 3) {real, imag} */,
  {32'hc098814a, 32'hc1dac3cc} /* (4, 25, 2) {real, imag} */,
  {32'hc1dc7086, 32'h3f37d3cc} /* (4, 25, 1) {real, imag} */,
  {32'hc1c6088a, 32'h411a5c4a} /* (4, 25, 0) {real, imag} */,
  {32'hbff1f918, 32'hc165830c} /* (4, 24, 31) {real, imag} */,
  {32'hc1a86cd2, 32'h4190e353} /* (4, 24, 30) {real, imag} */,
  {32'hbfc31862, 32'hbfc46f18} /* (4, 24, 29) {real, imag} */,
  {32'hc0865ddb, 32'h3f86cc7c} /* (4, 24, 28) {real, imag} */,
  {32'hbe8eb100, 32'h418d97ea} /* (4, 24, 27) {real, imag} */,
  {32'hc0c8d5a6, 32'hc149d87e} /* (4, 24, 26) {real, imag} */,
  {32'hc0b40eec, 32'hc027aa38} /* (4, 24, 25) {real, imag} */,
  {32'hc10a4634, 32'hc0ebaaee} /* (4, 24, 24) {real, imag} */,
  {32'h414cecfc, 32'hc19ba022} /* (4, 24, 23) {real, imag} */,
  {32'h418e1ac9, 32'h3fe0d3f0} /* (4, 24, 22) {real, imag} */,
  {32'hc104945a, 32'h3c70ea00} /* (4, 24, 21) {real, imag} */,
  {32'hc05cd5b1, 32'hc08f38d0} /* (4, 24, 20) {real, imag} */,
  {32'h40b5ac29, 32'h415ccfc0} /* (4, 24, 19) {real, imag} */,
  {32'h41085a50, 32'hc189a7e1} /* (4, 24, 18) {real, imag} */,
  {32'hbfde8f66, 32'h3edd7da8} /* (4, 24, 17) {real, imag} */,
  {32'h3e19a478, 32'h410f44ca} /* (4, 24, 16) {real, imag} */,
  {32'h4119801e, 32'hc04fb8c2} /* (4, 24, 15) {real, imag} */,
  {32'h40406782, 32'hc018b7ca} /* (4, 24, 14) {real, imag} */,
  {32'hc124bbd2, 32'hc117fa5e} /* (4, 24, 13) {real, imag} */,
  {32'h413f15fd, 32'h4175e13e} /* (4, 24, 12) {real, imag} */,
  {32'h3f7a9ac8, 32'hc156ecc7} /* (4, 24, 11) {real, imag} */,
  {32'hc151cd81, 32'hc1206be6} /* (4, 24, 10) {real, imag} */,
  {32'hc1a4db44, 32'h41080e71} /* (4, 24, 9) {real, imag} */,
  {32'hc19d6e1d, 32'h40aba6a3} /* (4, 24, 8) {real, imag} */,
  {32'hc1377614, 32'hc0aac088} /* (4, 24, 7) {real, imag} */,
  {32'h40d6a198, 32'h411450e8} /* (4, 24, 6) {real, imag} */,
  {32'h40da4f68, 32'h414aa07c} /* (4, 24, 5) {real, imag} */,
  {32'h415cc0f6, 32'h403013d6} /* (4, 24, 4) {real, imag} */,
  {32'h409e0f20, 32'hc0d504e2} /* (4, 24, 3) {real, imag} */,
  {32'hc20c18a4, 32'h414378a6} /* (4, 24, 2) {real, imag} */,
  {32'h423e96a6, 32'hc10b7fcf} /* (4, 24, 1) {real, imag} */,
  {32'h41af95a3, 32'hc2092d0c} /* (4, 24, 0) {real, imag} */,
  {32'hc16a0e35, 32'h40cd133a} /* (4, 23, 31) {real, imag} */,
  {32'h3fac7528, 32'hc03cf69b} /* (4, 23, 30) {real, imag} */,
  {32'h4138de7e, 32'hc1bdc7bc} /* (4, 23, 29) {real, imag} */,
  {32'h401deec0, 32'h416bca74} /* (4, 23, 28) {real, imag} */,
  {32'hc07974ac, 32'h411b95cb} /* (4, 23, 27) {real, imag} */,
  {32'hbff954a6, 32'hc1034225} /* (4, 23, 26) {real, imag} */,
  {32'h40505204, 32'hc094f5f6} /* (4, 23, 25) {real, imag} */,
  {32'hc0169ac7, 32'h3e0840c0} /* (4, 23, 24) {real, imag} */,
  {32'hc0f45db9, 32'hc092ba80} /* (4, 23, 23) {real, imag} */,
  {32'h4160bf4a, 32'h417882b2} /* (4, 23, 22) {real, imag} */,
  {32'hc163b1f2, 32'h411cfedb} /* (4, 23, 21) {real, imag} */,
  {32'hc02f059b, 32'h416f5fd4} /* (4, 23, 20) {real, imag} */,
  {32'hc068e66c, 32'hbe652670} /* (4, 23, 19) {real, imag} */,
  {32'hc09cbca8, 32'h3febb618} /* (4, 23, 18) {real, imag} */,
  {32'hc001b6be, 32'h408684ca} /* (4, 23, 17) {real, imag} */,
  {32'hc13b66d0, 32'h41862175} /* (4, 23, 16) {real, imag} */,
  {32'h408d9339, 32'hc0e942b7} /* (4, 23, 15) {real, imag} */,
  {32'hc08b90d4, 32'hc0fc0f7f} /* (4, 23, 14) {real, imag} */,
  {32'hc19d4502, 32'hbfdd1250} /* (4, 23, 13) {real, imag} */,
  {32'h40eca350, 32'hc192c51f} /* (4, 23, 12) {real, imag} */,
  {32'hc08a4ea4, 32'h413c2587} /* (4, 23, 11) {real, imag} */,
  {32'hc0bc7260, 32'h417998b5} /* (4, 23, 10) {real, imag} */,
  {32'hc160d8c3, 32'h41b468e2} /* (4, 23, 9) {real, imag} */,
  {32'hc080a85d, 32'hc08702c8} /* (4, 23, 8) {real, imag} */,
  {32'hc0d5a559, 32'hc15f8cf1} /* (4, 23, 7) {real, imag} */,
  {32'h41a8c2ad, 32'hc001ea50} /* (4, 23, 6) {real, imag} */,
  {32'h41b1bbc6, 32'hc181be5f} /* (4, 23, 5) {real, imag} */,
  {32'h4082b1e6, 32'h40e508a4} /* (4, 23, 4) {real, imag} */,
  {32'hc07576c4, 32'h415560b5} /* (4, 23, 3) {real, imag} */,
  {32'h4048b4a4, 32'h3fda6310} /* (4, 23, 2) {real, imag} */,
  {32'h410b6442, 32'h3f7435d0} /* (4, 23, 1) {real, imag} */,
  {32'hc0ace468, 32'hc174ddbd} /* (4, 23, 0) {real, imag} */,
  {32'hc1597c3b, 32'h3fa88c3e} /* (4, 22, 31) {real, imag} */,
  {32'h419c9715, 32'hc11a3eb5} /* (4, 22, 30) {real, imag} */,
  {32'hc0d99177, 32'h40f0a243} /* (4, 22, 29) {real, imag} */,
  {32'hbf90d1b0, 32'h40e468db} /* (4, 22, 28) {real, imag} */,
  {32'h410ae95b, 32'h41964c3e} /* (4, 22, 27) {real, imag} */,
  {32'h418101bf, 32'hc13a6e1c} /* (4, 22, 26) {real, imag} */,
  {32'hc12cfcfa, 32'hc10abef6} /* (4, 22, 25) {real, imag} */,
  {32'hc10be33c, 32'hc1034964} /* (4, 22, 24) {real, imag} */,
  {32'hbea9cb40, 32'hc16fd94e} /* (4, 22, 23) {real, imag} */,
  {32'h411c961c, 32'h4111d848} /* (4, 22, 22) {real, imag} */,
  {32'h41a4c715, 32'hc0f5e8d0} /* (4, 22, 21) {real, imag} */,
  {32'h4198d087, 32'h40d41000} /* (4, 22, 20) {real, imag} */,
  {32'hbffd0e64, 32'hc0ca823c} /* (4, 22, 19) {real, imag} */,
  {32'hc0ab5cd8, 32'hc0eeacd3} /* (4, 22, 18) {real, imag} */,
  {32'h408e69dd, 32'h408bf8c9} /* (4, 22, 17) {real, imag} */,
  {32'h40150843, 32'hc14d3674} /* (4, 22, 16) {real, imag} */,
  {32'h3fb4f966, 32'hc0c29718} /* (4, 22, 15) {real, imag} */,
  {32'hc018bdc8, 32'hc0943618} /* (4, 22, 14) {real, imag} */,
  {32'hbfc2e5b0, 32'hc001ef3a} /* (4, 22, 13) {real, imag} */,
  {32'h4163d019, 32'hc0b8ee5a} /* (4, 22, 12) {real, imag} */,
  {32'hc0d0fc34, 32'h414e4c9a} /* (4, 22, 11) {real, imag} */,
  {32'hc110e90c, 32'hc1490885} /* (4, 22, 10) {real, imag} */,
  {32'h404da5a8, 32'h3fb5c26f} /* (4, 22, 9) {real, imag} */,
  {32'hc114c565, 32'hc1b6e4c9} /* (4, 22, 8) {real, imag} */,
  {32'hc0a6dc0e, 32'h40a58dfe} /* (4, 22, 7) {real, imag} */,
  {32'h411f318c, 32'h40cdbfd4} /* (4, 22, 6) {real, imag} */,
  {32'h41c2bee3, 32'hc15f7075} /* (4, 22, 5) {real, imag} */,
  {32'hc049591a, 32'hbfeb2b8c} /* (4, 22, 4) {real, imag} */,
  {32'hc1989a9f, 32'hc1a23602} /* (4, 22, 3) {real, imag} */,
  {32'h3fa1578a, 32'h4129f866} /* (4, 22, 2) {real, imag} */,
  {32'h4176bb58, 32'h4139fcc1} /* (4, 22, 1) {real, imag} */,
  {32'hc183c667, 32'h41a92d22} /* (4, 22, 0) {real, imag} */,
  {32'hc000a81a, 32'hc21cb290} /* (4, 21, 31) {real, imag} */,
  {32'hc0618118, 32'h415d7304} /* (4, 21, 30) {real, imag} */,
  {32'hc1b5d760, 32'h40b7a610} /* (4, 21, 29) {real, imag} */,
  {32'hbfceb084, 32'h4118016b} /* (4, 21, 28) {real, imag} */,
  {32'hc140be68, 32'hc07c301c} /* (4, 21, 27) {real, imag} */,
  {32'h41a50f17, 32'hc0e324a2} /* (4, 21, 26) {real, imag} */,
  {32'h416fe189, 32'hbe4dcc80} /* (4, 21, 25) {real, imag} */,
  {32'hc106a89a, 32'h405365a8} /* (4, 21, 24) {real, imag} */,
  {32'hc1361251, 32'hc0d591b2} /* (4, 21, 23) {real, imag} */,
  {32'hc128364b, 32'hc07d36ed} /* (4, 21, 22) {real, imag} */,
  {32'hc11466bd, 32'h413f53b6} /* (4, 21, 21) {real, imag} */,
  {32'hc15dd17f, 32'h4118d912} /* (4, 21, 20) {real, imag} */,
  {32'hc076f52d, 32'h412551cf} /* (4, 21, 19) {real, imag} */,
  {32'h41a1c805, 32'h40941a42} /* (4, 21, 18) {real, imag} */,
  {32'hbeaccc60, 32'hc0f1afcc} /* (4, 21, 17) {real, imag} */,
  {32'h40ecb998, 32'hc01648f4} /* (4, 21, 16) {real, imag} */,
  {32'hc0a86992, 32'h4167172c} /* (4, 21, 15) {real, imag} */,
  {32'hc1595252, 32'hc0fde3e4} /* (4, 21, 14) {real, imag} */,
  {32'hc0216326, 32'hc000c008} /* (4, 21, 13) {real, imag} */,
  {32'h4106405e, 32'h4064a1c0} /* (4, 21, 12) {real, imag} */,
  {32'hc128abac, 32'h3f783dd8} /* (4, 21, 11) {real, imag} */,
  {32'hc10a2ce6, 32'hc11dcb7a} /* (4, 21, 10) {real, imag} */,
  {32'h3f0a7eac, 32'h411a53f4} /* (4, 21, 9) {real, imag} */,
  {32'hc0a0a292, 32'hc0be1d1a} /* (4, 21, 8) {real, imag} */,
  {32'h4117809e, 32'hc0005c28} /* (4, 21, 7) {real, imag} */,
  {32'hc0c1eb7a, 32'hc07c5a1c} /* (4, 21, 6) {real, imag} */,
  {32'hc08294f9, 32'h4168d502} /* (4, 21, 5) {real, imag} */,
  {32'h40d3e39a, 32'hbffe3264} /* (4, 21, 4) {real, imag} */,
  {32'hc16f962b, 32'hc07cf4a6} /* (4, 21, 3) {real, imag} */,
  {32'hc1650f46, 32'h41104dd9} /* (4, 21, 2) {real, imag} */,
  {32'h40fbe16f, 32'hc1942e25} /* (4, 21, 1) {real, imag} */,
  {32'h420660cc, 32'hc0f62072} /* (4, 21, 0) {real, imag} */,
  {32'h4059867b, 32'h40d77070} /* (4, 20, 31) {real, imag} */,
  {32'h402535a3, 32'hc0b45999} /* (4, 20, 30) {real, imag} */,
  {32'hc126fb48, 32'h40d0cad7} /* (4, 20, 29) {real, imag} */,
  {32'hc10eb760, 32'hc159936b} /* (4, 20, 28) {real, imag} */,
  {32'h40fcbcdc, 32'h41b6f8ff} /* (4, 20, 27) {real, imag} */,
  {32'h40d2346c, 32'hc08a482a} /* (4, 20, 26) {real, imag} */,
  {32'h40a8c94b, 32'h3f831de0} /* (4, 20, 25) {real, imag} */,
  {32'h415b36f0, 32'hc176469d} /* (4, 20, 24) {real, imag} */,
  {32'h41234800, 32'hc0732792} /* (4, 20, 23) {real, imag} */,
  {32'hc1960b06, 32'h40af4732} /* (4, 20, 22) {real, imag} */,
  {32'h408b461e, 32'h4033efdf} /* (4, 20, 21) {real, imag} */,
  {32'h4168d0a4, 32'hc115f91b} /* (4, 20, 20) {real, imag} */,
  {32'hc0b31ccc, 32'hc112a0fc} /* (4, 20, 19) {real, imag} */,
  {32'h4139f0cf, 32'hc03b215c} /* (4, 20, 18) {real, imag} */,
  {32'hc18d3e21, 32'hc05fc7d6} /* (4, 20, 17) {real, imag} */,
  {32'hbdc6f680, 32'h3f6bf288} /* (4, 20, 16) {real, imag} */,
  {32'h41559e90, 32'hc098a8d2} /* (4, 20, 15) {real, imag} */,
  {32'h40ecb76b, 32'hc0abb938} /* (4, 20, 14) {real, imag} */,
  {32'h419c222a, 32'h403256e8} /* (4, 20, 13) {real, imag} */,
  {32'hc11566e1, 32'h3fbe69f4} /* (4, 20, 12) {real, imag} */,
  {32'h3b816000, 32'hc188e4d9} /* (4, 20, 11) {real, imag} */,
  {32'h41758f7e, 32'h41be8e2a} /* (4, 20, 10) {real, imag} */,
  {32'hc11ddc40, 32'h3f0bfca0} /* (4, 20, 9) {real, imag} */,
  {32'h40e8b00e, 32'h3fb359f4} /* (4, 20, 8) {real, imag} */,
  {32'hc0472cac, 32'h41a54263} /* (4, 20, 7) {real, imag} */,
  {32'hc1766a56, 32'h408d9a7e} /* (4, 20, 6) {real, imag} */,
  {32'h4114ae47, 32'h40affd42} /* (4, 20, 5) {real, imag} */,
  {32'h41069960, 32'hc00170a0} /* (4, 20, 4) {real, imag} */,
  {32'hc13f797f, 32'hc0b66946} /* (4, 20, 3) {real, imag} */,
  {32'hc10c0730, 32'hc16b5854} /* (4, 20, 2) {real, imag} */,
  {32'hc092be58, 32'hc061b2b9} /* (4, 20, 1) {real, imag} */,
  {32'hc100a0d0, 32'hbe83ff10} /* (4, 20, 0) {real, imag} */,
  {32'h4111592d, 32'h411b3ebe} /* (4, 19, 31) {real, imag} */,
  {32'h40c5f5c0, 32'hc11386b2} /* (4, 19, 30) {real, imag} */,
  {32'hc00b7f01, 32'h40d72df0} /* (4, 19, 29) {real, imag} */,
  {32'hc107b390, 32'h40ab80d3} /* (4, 19, 28) {real, imag} */,
  {32'hc1383d48, 32'hc0b5f46f} /* (4, 19, 27) {real, imag} */,
  {32'hc11a9d6b, 32'h416d9c43} /* (4, 19, 26) {real, imag} */,
  {32'hc18f7b47, 32'h4150524d} /* (4, 19, 25) {real, imag} */,
  {32'hc0805535, 32'hc1a8e5b8} /* (4, 19, 24) {real, imag} */,
  {32'h4114b8cc, 32'hbd465fc0} /* (4, 19, 23) {real, imag} */,
  {32'hc16302b2, 32'hc050da09} /* (4, 19, 22) {real, imag} */,
  {32'h40b1df36, 32'h40a0080a} /* (4, 19, 21) {real, imag} */,
  {32'h40bd52d2, 32'hc083ca20} /* (4, 19, 20) {real, imag} */,
  {32'hc0fdda77, 32'hc19649ec} /* (4, 19, 19) {real, imag} */,
  {32'hc0c43ee4, 32'hbffaeee6} /* (4, 19, 18) {real, imag} */,
  {32'h411e907c, 32'h419a865a} /* (4, 19, 17) {real, imag} */,
  {32'h4040963c, 32'h4048b7de} /* (4, 19, 16) {real, imag} */,
  {32'hc0cb41bc, 32'h4107c172} /* (4, 19, 15) {real, imag} */,
  {32'h3fa3191c, 32'h412d724b} /* (4, 19, 14) {real, imag} */,
  {32'hc12f2e17, 32'h4019b804} /* (4, 19, 13) {real, imag} */,
  {32'hc158cec0, 32'h4114864b} /* (4, 19, 12) {real, imag} */,
  {32'h41a0011e, 32'hc0a60d2a} /* (4, 19, 11) {real, imag} */,
  {32'h3f8d87ea, 32'h4111e0fb} /* (4, 19, 10) {real, imag} */,
  {32'hc152ef3e, 32'hc180729b} /* (4, 19, 9) {real, imag} */,
  {32'h41389654, 32'h3fabfe5a} /* (4, 19, 8) {real, imag} */,
  {32'h40a09502, 32'hc16f0977} /* (4, 19, 7) {real, imag} */,
  {32'hc10c9da8, 32'h40beee28} /* (4, 19, 6) {real, imag} */,
  {32'hc0af39b6, 32'h410a70b6} /* (4, 19, 5) {real, imag} */,
  {32'h3f056927, 32'h3f1bd0c4} /* (4, 19, 4) {real, imag} */,
  {32'h400be66a, 32'h41776306} /* (4, 19, 3) {real, imag} */,
  {32'h407cea61, 32'hbf368af6} /* (4, 19, 2) {real, imag} */,
  {32'hc160b363, 32'h40b7e0a3} /* (4, 19, 1) {real, imag} */,
  {32'hc0c33b5f, 32'hc09027fc} /* (4, 19, 0) {real, imag} */,
  {32'hc18a05a3, 32'h40e0aee1} /* (4, 18, 31) {real, imag} */,
  {32'hc02af6bd, 32'h3e8213c0} /* (4, 18, 30) {real, imag} */,
  {32'h4038bb9c, 32'h3fe8c250} /* (4, 18, 29) {real, imag} */,
  {32'h4104afd4, 32'hc125e6fa} /* (4, 18, 28) {real, imag} */,
  {32'h40471f62, 32'h409e4bd3} /* (4, 18, 27) {real, imag} */,
  {32'h3fd78dca, 32'hbf82e044} /* (4, 18, 26) {real, imag} */,
  {32'hc09d71e9, 32'h4146baf8} /* (4, 18, 25) {real, imag} */,
  {32'hc026c327, 32'h40ea7a70} /* (4, 18, 24) {real, imag} */,
  {32'h419e105c, 32'h410493b0} /* (4, 18, 23) {real, imag} */,
  {32'hc07bd376, 32'h40650202} /* (4, 18, 22) {real, imag} */,
  {32'h3fba54bc, 32'hc1590d88} /* (4, 18, 21) {real, imag} */,
  {32'hc0957404, 32'h409ec32d} /* (4, 18, 20) {real, imag} */,
  {32'hc0ce4b89, 32'hbfadfac0} /* (4, 18, 19) {real, imag} */,
  {32'hbfa54628, 32'hc0553c6d} /* (4, 18, 18) {real, imag} */,
  {32'hc12e5476, 32'h3f8adf76} /* (4, 18, 17) {real, imag} */,
  {32'hbfe0d194, 32'h403e6cdf} /* (4, 18, 16) {real, imag} */,
  {32'h4044b6a1, 32'h40108d10} /* (4, 18, 15) {real, imag} */,
  {32'h401ec598, 32'h418b9cac} /* (4, 18, 14) {real, imag} */,
  {32'hc134b0c8, 32'hc004bc37} /* (4, 18, 13) {real, imag} */,
  {32'h3ff33c53, 32'h3f8ab9f6} /* (4, 18, 12) {real, imag} */,
  {32'h40ea2bc0, 32'hc1608db6} /* (4, 18, 11) {real, imag} */,
  {32'h3fc48ec6, 32'hbf429cbc} /* (4, 18, 10) {real, imag} */,
  {32'h3ff35d00, 32'h4136083b} /* (4, 18, 9) {real, imag} */,
  {32'h4102b6af, 32'hc0b7f8ff} /* (4, 18, 8) {real, imag} */,
  {32'h408baa91, 32'hbe0d7200} /* (4, 18, 7) {real, imag} */,
  {32'hc0a8bfca, 32'hc1181029} /* (4, 18, 6) {real, imag} */,
  {32'h40a0ec51, 32'h414b2452} /* (4, 18, 5) {real, imag} */,
  {32'hc0ea904e, 32'hbfa0bdac} /* (4, 18, 4) {real, imag} */,
  {32'h40d20597, 32'h416fc10b} /* (4, 18, 3) {real, imag} */,
  {32'hc093a2fb, 32'h3f0aa980} /* (4, 18, 2) {real, imag} */,
  {32'h413de1f4, 32'hc1557bf3} /* (4, 18, 1) {real, imag} */,
  {32'h3f29b15e, 32'hc0dedb95} /* (4, 18, 0) {real, imag} */,
  {32'hc0ce915e, 32'h412ad585} /* (4, 17, 31) {real, imag} */,
  {32'hc09e7fbf, 32'hc1320965} /* (4, 17, 30) {real, imag} */,
  {32'h410b052b, 32'h410388e3} /* (4, 17, 29) {real, imag} */,
  {32'h40d5bcfd, 32'h3fbce4e8} /* (4, 17, 28) {real, imag} */,
  {32'hc190df56, 32'hbe2d5d40} /* (4, 17, 27) {real, imag} */,
  {32'h40c202ed, 32'h3feb4678} /* (4, 17, 26) {real, imag} */,
  {32'h3e83eda0, 32'hbf0a4d10} /* (4, 17, 25) {real, imag} */,
  {32'hc04ed95c, 32'hc02fb7ec} /* (4, 17, 24) {real, imag} */,
  {32'h4145e632, 32'h411853f9} /* (4, 17, 23) {real, imag} */,
  {32'hbf4c1b28, 32'hbf254784} /* (4, 17, 22) {real, imag} */,
  {32'hc04d0397, 32'h4112d95f} /* (4, 17, 21) {real, imag} */,
  {32'h40c216bc, 32'hbea571e8} /* (4, 17, 20) {real, imag} */,
  {32'h413a046b, 32'h4070409d} /* (4, 17, 19) {real, imag} */,
  {32'hc0f3638c, 32'h4126615b} /* (4, 17, 18) {real, imag} */,
  {32'h3fe5a899, 32'hc12ee702} /* (4, 17, 17) {real, imag} */,
  {32'h40d385fb, 32'h3ff6b002} /* (4, 17, 16) {real, imag} */,
  {32'hc0f0028f, 32'hc0078ec2} /* (4, 17, 15) {real, imag} */,
  {32'h41229559, 32'hc0acea4b} /* (4, 17, 14) {real, imag} */,
  {32'h4162ad1a, 32'hc12d88ec} /* (4, 17, 13) {real, imag} */,
  {32'h41381c9f, 32'hc0896874} /* (4, 17, 12) {real, imag} */,
  {32'hc0975db5, 32'hc107388f} /* (4, 17, 11) {real, imag} */,
  {32'hc1276710, 32'h40e4d1de} /* (4, 17, 10) {real, imag} */,
  {32'hc09b4556, 32'h41058ba0} /* (4, 17, 9) {real, imag} */,
  {32'hc0c76142, 32'h3ef0f058} /* (4, 17, 8) {real, imag} */,
  {32'h4000417a, 32'h411a65e8} /* (4, 17, 7) {real, imag} */,
  {32'h4134265a, 32'h40cde41e} /* (4, 17, 6) {real, imag} */,
  {32'h408f970e, 32'h406ffe47} /* (4, 17, 5) {real, imag} */,
  {32'hc08b4a0f, 32'hbf5f786a} /* (4, 17, 4) {real, imag} */,
  {32'hc0ada9ab, 32'hc0eb0174} /* (4, 17, 3) {real, imag} */,
  {32'hc06232dc, 32'hc02afca2} /* (4, 17, 2) {real, imag} */,
  {32'h406d84ea, 32'h41730ca4} /* (4, 17, 1) {real, imag} */,
  {32'hc0809e79, 32'h41a2b519} /* (4, 17, 0) {real, imag} */,
  {32'hc0db38cf, 32'hc0f61d66} /* (4, 16, 31) {real, imag} */,
  {32'hc0c23126, 32'hbfe881d1} /* (4, 16, 30) {real, imag} */,
  {32'hc0af5818, 32'hbf52d4c8} /* (4, 16, 29) {real, imag} */,
  {32'h40c96e2b, 32'hc1167279} /* (4, 16, 28) {real, imag} */,
  {32'h40e262ac, 32'hc10d45fb} /* (4, 16, 27) {real, imag} */,
  {32'h3fcfb3e2, 32'h3ec603a0} /* (4, 16, 26) {real, imag} */,
  {32'hc06635f8, 32'hc150ec38} /* (4, 16, 25) {real, imag} */,
  {32'h405b328b, 32'hc09227fa} /* (4, 16, 24) {real, imag} */,
  {32'hbf7e2158, 32'h4008556e} /* (4, 16, 23) {real, imag} */,
  {32'hc1295421, 32'hc13f21c7} /* (4, 16, 22) {real, imag} */,
  {32'hc101bf54, 32'hc0005d54} /* (4, 16, 21) {real, imag} */,
  {32'h4045a84b, 32'hc071e326} /* (4, 16, 20) {real, imag} */,
  {32'h40816963, 32'hc0ceb01b} /* (4, 16, 19) {real, imag} */,
  {32'hc0ecf7f7, 32'hbfb073a4} /* (4, 16, 18) {real, imag} */,
  {32'hbb68f000, 32'hbfe8c78a} /* (4, 16, 17) {real, imag} */,
  {32'hc040580e, 32'h00000000} /* (4, 16, 16) {real, imag} */,
  {32'hbb68f000, 32'h3fe8c78a} /* (4, 16, 15) {real, imag} */,
  {32'hc0ecf7f7, 32'h3fb073a4} /* (4, 16, 14) {real, imag} */,
  {32'h40816963, 32'h40ceb01b} /* (4, 16, 13) {real, imag} */,
  {32'h4045a84b, 32'h4071e326} /* (4, 16, 12) {real, imag} */,
  {32'hc101bf54, 32'h40005d54} /* (4, 16, 11) {real, imag} */,
  {32'hc1295421, 32'h413f21c7} /* (4, 16, 10) {real, imag} */,
  {32'hbf7e2158, 32'hc008556e} /* (4, 16, 9) {real, imag} */,
  {32'h405b328b, 32'h409227fa} /* (4, 16, 8) {real, imag} */,
  {32'hc06635f8, 32'h4150ec38} /* (4, 16, 7) {real, imag} */,
  {32'h3fcfb3e2, 32'hbec603a0} /* (4, 16, 6) {real, imag} */,
  {32'h40e262ac, 32'h410d45fb} /* (4, 16, 5) {real, imag} */,
  {32'h40c96e2b, 32'h41167279} /* (4, 16, 4) {real, imag} */,
  {32'hc0af5818, 32'h3f52d4c8} /* (4, 16, 3) {real, imag} */,
  {32'hc0c23126, 32'h3fe881d1} /* (4, 16, 2) {real, imag} */,
  {32'hc0db38cf, 32'h40f61d66} /* (4, 16, 1) {real, imag} */,
  {32'h401871fc, 32'h00000000} /* (4, 16, 0) {real, imag} */,
  {32'h406d84ea, 32'hc1730ca4} /* (4, 15, 31) {real, imag} */,
  {32'hc06232dc, 32'h402afca2} /* (4, 15, 30) {real, imag} */,
  {32'hc0ada9ab, 32'h40eb0174} /* (4, 15, 29) {real, imag} */,
  {32'hc08b4a0f, 32'h3f5f786a} /* (4, 15, 28) {real, imag} */,
  {32'h408f970e, 32'hc06ffe47} /* (4, 15, 27) {real, imag} */,
  {32'h4134265a, 32'hc0cde41e} /* (4, 15, 26) {real, imag} */,
  {32'h4000417a, 32'hc11a65e8} /* (4, 15, 25) {real, imag} */,
  {32'hc0c76142, 32'hbef0f058} /* (4, 15, 24) {real, imag} */,
  {32'hc09b4556, 32'hc1058ba0} /* (4, 15, 23) {real, imag} */,
  {32'hc1276710, 32'hc0e4d1de} /* (4, 15, 22) {real, imag} */,
  {32'hc0975db5, 32'h4107388f} /* (4, 15, 21) {real, imag} */,
  {32'h41381c9f, 32'h40896874} /* (4, 15, 20) {real, imag} */,
  {32'h4162ad1a, 32'h412d88ec} /* (4, 15, 19) {real, imag} */,
  {32'h41229559, 32'h40acea4b} /* (4, 15, 18) {real, imag} */,
  {32'hc0f0028f, 32'h40078ec2} /* (4, 15, 17) {real, imag} */,
  {32'h40d385fb, 32'hbff6b002} /* (4, 15, 16) {real, imag} */,
  {32'h3fe5a899, 32'h412ee702} /* (4, 15, 15) {real, imag} */,
  {32'hc0f3638c, 32'hc126615b} /* (4, 15, 14) {real, imag} */,
  {32'h413a046b, 32'hc070409d} /* (4, 15, 13) {real, imag} */,
  {32'h40c216bc, 32'h3ea571e8} /* (4, 15, 12) {real, imag} */,
  {32'hc04d0397, 32'hc112d95f} /* (4, 15, 11) {real, imag} */,
  {32'hbf4c1b28, 32'h3f254784} /* (4, 15, 10) {real, imag} */,
  {32'h4145e632, 32'hc11853f9} /* (4, 15, 9) {real, imag} */,
  {32'hc04ed95c, 32'h402fb7ec} /* (4, 15, 8) {real, imag} */,
  {32'h3e83eda0, 32'h3f0a4d10} /* (4, 15, 7) {real, imag} */,
  {32'h40c202ed, 32'hbfeb4678} /* (4, 15, 6) {real, imag} */,
  {32'hc190df56, 32'h3e2d5d40} /* (4, 15, 5) {real, imag} */,
  {32'h40d5bcfd, 32'hbfbce4e8} /* (4, 15, 4) {real, imag} */,
  {32'h410b052b, 32'hc10388e3} /* (4, 15, 3) {real, imag} */,
  {32'hc09e7fbf, 32'h41320965} /* (4, 15, 2) {real, imag} */,
  {32'hc0ce915e, 32'hc12ad585} /* (4, 15, 1) {real, imag} */,
  {32'hc0809e79, 32'hc1a2b519} /* (4, 15, 0) {real, imag} */,
  {32'h413de1f4, 32'h41557bf3} /* (4, 14, 31) {real, imag} */,
  {32'hc093a2fb, 32'hbf0aa980} /* (4, 14, 30) {real, imag} */,
  {32'h40d20597, 32'hc16fc10b} /* (4, 14, 29) {real, imag} */,
  {32'hc0ea904e, 32'h3fa0bdac} /* (4, 14, 28) {real, imag} */,
  {32'h40a0ec51, 32'hc14b2452} /* (4, 14, 27) {real, imag} */,
  {32'hc0a8bfca, 32'h41181029} /* (4, 14, 26) {real, imag} */,
  {32'h408baa91, 32'h3e0d7200} /* (4, 14, 25) {real, imag} */,
  {32'h4102b6af, 32'h40b7f8ff} /* (4, 14, 24) {real, imag} */,
  {32'h3ff35d00, 32'hc136083b} /* (4, 14, 23) {real, imag} */,
  {32'h3fc48ec6, 32'h3f429cbc} /* (4, 14, 22) {real, imag} */,
  {32'h40ea2bc0, 32'h41608db6} /* (4, 14, 21) {real, imag} */,
  {32'h3ff33c53, 32'hbf8ab9f6} /* (4, 14, 20) {real, imag} */,
  {32'hc134b0c8, 32'h4004bc37} /* (4, 14, 19) {real, imag} */,
  {32'h401ec598, 32'hc18b9cac} /* (4, 14, 18) {real, imag} */,
  {32'h4044b6a1, 32'hc0108d10} /* (4, 14, 17) {real, imag} */,
  {32'hbfe0d194, 32'hc03e6cdf} /* (4, 14, 16) {real, imag} */,
  {32'hc12e5476, 32'hbf8adf76} /* (4, 14, 15) {real, imag} */,
  {32'hbfa54628, 32'h40553c6d} /* (4, 14, 14) {real, imag} */,
  {32'hc0ce4b89, 32'h3fadfac0} /* (4, 14, 13) {real, imag} */,
  {32'hc0957404, 32'hc09ec32d} /* (4, 14, 12) {real, imag} */,
  {32'h3fba54bc, 32'h41590d88} /* (4, 14, 11) {real, imag} */,
  {32'hc07bd376, 32'hc0650202} /* (4, 14, 10) {real, imag} */,
  {32'h419e105c, 32'hc10493b0} /* (4, 14, 9) {real, imag} */,
  {32'hc026c327, 32'hc0ea7a70} /* (4, 14, 8) {real, imag} */,
  {32'hc09d71e9, 32'hc146baf8} /* (4, 14, 7) {real, imag} */,
  {32'h3fd78dca, 32'h3f82e044} /* (4, 14, 6) {real, imag} */,
  {32'h40471f62, 32'hc09e4bd3} /* (4, 14, 5) {real, imag} */,
  {32'h4104afd4, 32'h4125e6fa} /* (4, 14, 4) {real, imag} */,
  {32'h4038bb9c, 32'hbfe8c250} /* (4, 14, 3) {real, imag} */,
  {32'hc02af6bd, 32'hbe8213c0} /* (4, 14, 2) {real, imag} */,
  {32'hc18a05a3, 32'hc0e0aee1} /* (4, 14, 1) {real, imag} */,
  {32'h3f29b15e, 32'h40dedb95} /* (4, 14, 0) {real, imag} */,
  {32'hc160b363, 32'hc0b7e0a3} /* (4, 13, 31) {real, imag} */,
  {32'h407cea61, 32'h3f368af6} /* (4, 13, 30) {real, imag} */,
  {32'h400be66a, 32'hc1776306} /* (4, 13, 29) {real, imag} */,
  {32'h3f056927, 32'hbf1bd0c4} /* (4, 13, 28) {real, imag} */,
  {32'hc0af39b6, 32'hc10a70b6} /* (4, 13, 27) {real, imag} */,
  {32'hc10c9da8, 32'hc0beee28} /* (4, 13, 26) {real, imag} */,
  {32'h40a09502, 32'h416f0977} /* (4, 13, 25) {real, imag} */,
  {32'h41389654, 32'hbfabfe5a} /* (4, 13, 24) {real, imag} */,
  {32'hc152ef3e, 32'h4180729b} /* (4, 13, 23) {real, imag} */,
  {32'h3f8d87ea, 32'hc111e0fb} /* (4, 13, 22) {real, imag} */,
  {32'h41a0011e, 32'h40a60d2a} /* (4, 13, 21) {real, imag} */,
  {32'hc158cec0, 32'hc114864b} /* (4, 13, 20) {real, imag} */,
  {32'hc12f2e17, 32'hc019b804} /* (4, 13, 19) {real, imag} */,
  {32'h3fa3191c, 32'hc12d724b} /* (4, 13, 18) {real, imag} */,
  {32'hc0cb41bc, 32'hc107c172} /* (4, 13, 17) {real, imag} */,
  {32'h4040963c, 32'hc048b7de} /* (4, 13, 16) {real, imag} */,
  {32'h411e907c, 32'hc19a865a} /* (4, 13, 15) {real, imag} */,
  {32'hc0c43ee4, 32'h3ffaeee6} /* (4, 13, 14) {real, imag} */,
  {32'hc0fdda77, 32'h419649ec} /* (4, 13, 13) {real, imag} */,
  {32'h40bd52d2, 32'h4083ca20} /* (4, 13, 12) {real, imag} */,
  {32'h40b1df36, 32'hc0a0080a} /* (4, 13, 11) {real, imag} */,
  {32'hc16302b2, 32'h4050da09} /* (4, 13, 10) {real, imag} */,
  {32'h4114b8cc, 32'h3d465fc0} /* (4, 13, 9) {real, imag} */,
  {32'hc0805535, 32'h41a8e5b8} /* (4, 13, 8) {real, imag} */,
  {32'hc18f7b47, 32'hc150524d} /* (4, 13, 7) {real, imag} */,
  {32'hc11a9d6b, 32'hc16d9c43} /* (4, 13, 6) {real, imag} */,
  {32'hc1383d48, 32'h40b5f46f} /* (4, 13, 5) {real, imag} */,
  {32'hc107b390, 32'hc0ab80d3} /* (4, 13, 4) {real, imag} */,
  {32'hc00b7f01, 32'hc0d72df0} /* (4, 13, 3) {real, imag} */,
  {32'h40c5f5c0, 32'h411386b2} /* (4, 13, 2) {real, imag} */,
  {32'h4111592d, 32'hc11b3ebe} /* (4, 13, 1) {real, imag} */,
  {32'hc0c33b5f, 32'h409027fc} /* (4, 13, 0) {real, imag} */,
  {32'hc092be58, 32'h4061b2b9} /* (4, 12, 31) {real, imag} */,
  {32'hc10c0730, 32'h416b5854} /* (4, 12, 30) {real, imag} */,
  {32'hc13f797f, 32'h40b66946} /* (4, 12, 29) {real, imag} */,
  {32'h41069960, 32'h400170a0} /* (4, 12, 28) {real, imag} */,
  {32'h4114ae47, 32'hc0affd42} /* (4, 12, 27) {real, imag} */,
  {32'hc1766a56, 32'hc08d9a7e} /* (4, 12, 26) {real, imag} */,
  {32'hc0472cac, 32'hc1a54263} /* (4, 12, 25) {real, imag} */,
  {32'h40e8b00e, 32'hbfb359f4} /* (4, 12, 24) {real, imag} */,
  {32'hc11ddc40, 32'hbf0bfca0} /* (4, 12, 23) {real, imag} */,
  {32'h41758f7e, 32'hc1be8e2a} /* (4, 12, 22) {real, imag} */,
  {32'h3b816000, 32'h4188e4d9} /* (4, 12, 21) {real, imag} */,
  {32'hc11566e1, 32'hbfbe69f4} /* (4, 12, 20) {real, imag} */,
  {32'h419c222a, 32'hc03256e8} /* (4, 12, 19) {real, imag} */,
  {32'h40ecb76b, 32'h40abb938} /* (4, 12, 18) {real, imag} */,
  {32'h41559e90, 32'h4098a8d2} /* (4, 12, 17) {real, imag} */,
  {32'hbdc6f680, 32'hbf6bf288} /* (4, 12, 16) {real, imag} */,
  {32'hc18d3e21, 32'h405fc7d6} /* (4, 12, 15) {real, imag} */,
  {32'h4139f0cf, 32'h403b215c} /* (4, 12, 14) {real, imag} */,
  {32'hc0b31ccc, 32'h4112a0fc} /* (4, 12, 13) {real, imag} */,
  {32'h4168d0a4, 32'h4115f91b} /* (4, 12, 12) {real, imag} */,
  {32'h408b461e, 32'hc033efdf} /* (4, 12, 11) {real, imag} */,
  {32'hc1960b06, 32'hc0af4732} /* (4, 12, 10) {real, imag} */,
  {32'h41234800, 32'h40732792} /* (4, 12, 9) {real, imag} */,
  {32'h415b36f0, 32'h4176469d} /* (4, 12, 8) {real, imag} */,
  {32'h40a8c94b, 32'hbf831de0} /* (4, 12, 7) {real, imag} */,
  {32'h40d2346c, 32'h408a482a} /* (4, 12, 6) {real, imag} */,
  {32'h40fcbcdc, 32'hc1b6f8ff} /* (4, 12, 5) {real, imag} */,
  {32'hc10eb760, 32'h4159936b} /* (4, 12, 4) {real, imag} */,
  {32'hc126fb48, 32'hc0d0cad7} /* (4, 12, 3) {real, imag} */,
  {32'h402535a3, 32'h40b45999} /* (4, 12, 2) {real, imag} */,
  {32'h4059867b, 32'hc0d77070} /* (4, 12, 1) {real, imag} */,
  {32'hc100a0d0, 32'h3e83ff10} /* (4, 12, 0) {real, imag} */,
  {32'h40fbe16f, 32'h41942e25} /* (4, 11, 31) {real, imag} */,
  {32'hc1650f46, 32'hc1104dd9} /* (4, 11, 30) {real, imag} */,
  {32'hc16f962b, 32'h407cf4a6} /* (4, 11, 29) {real, imag} */,
  {32'h40d3e39a, 32'h3ffe3264} /* (4, 11, 28) {real, imag} */,
  {32'hc08294f9, 32'hc168d502} /* (4, 11, 27) {real, imag} */,
  {32'hc0c1eb7a, 32'h407c5a1c} /* (4, 11, 26) {real, imag} */,
  {32'h4117809e, 32'h40005c28} /* (4, 11, 25) {real, imag} */,
  {32'hc0a0a292, 32'h40be1d1a} /* (4, 11, 24) {real, imag} */,
  {32'h3f0a7eac, 32'hc11a53f4} /* (4, 11, 23) {real, imag} */,
  {32'hc10a2ce6, 32'h411dcb7a} /* (4, 11, 22) {real, imag} */,
  {32'hc128abac, 32'hbf783dd8} /* (4, 11, 21) {real, imag} */,
  {32'h4106405e, 32'hc064a1c0} /* (4, 11, 20) {real, imag} */,
  {32'hc0216326, 32'h4000c008} /* (4, 11, 19) {real, imag} */,
  {32'hc1595252, 32'h40fde3e4} /* (4, 11, 18) {real, imag} */,
  {32'hc0a86992, 32'hc167172c} /* (4, 11, 17) {real, imag} */,
  {32'h40ecb998, 32'h401648f4} /* (4, 11, 16) {real, imag} */,
  {32'hbeaccc60, 32'h40f1afcc} /* (4, 11, 15) {real, imag} */,
  {32'h41a1c805, 32'hc0941a42} /* (4, 11, 14) {real, imag} */,
  {32'hc076f52d, 32'hc12551cf} /* (4, 11, 13) {real, imag} */,
  {32'hc15dd17f, 32'hc118d912} /* (4, 11, 12) {real, imag} */,
  {32'hc11466bd, 32'hc13f53b6} /* (4, 11, 11) {real, imag} */,
  {32'hc128364b, 32'h407d36ed} /* (4, 11, 10) {real, imag} */,
  {32'hc1361251, 32'h40d591b2} /* (4, 11, 9) {real, imag} */,
  {32'hc106a89a, 32'hc05365a8} /* (4, 11, 8) {real, imag} */,
  {32'h416fe189, 32'h3e4dcc80} /* (4, 11, 7) {real, imag} */,
  {32'h41a50f17, 32'h40e324a2} /* (4, 11, 6) {real, imag} */,
  {32'hc140be68, 32'h407c301c} /* (4, 11, 5) {real, imag} */,
  {32'hbfceb084, 32'hc118016b} /* (4, 11, 4) {real, imag} */,
  {32'hc1b5d760, 32'hc0b7a610} /* (4, 11, 3) {real, imag} */,
  {32'hc0618118, 32'hc15d7304} /* (4, 11, 2) {real, imag} */,
  {32'hc000a81a, 32'h421cb290} /* (4, 11, 1) {real, imag} */,
  {32'h420660cc, 32'h40f62072} /* (4, 11, 0) {real, imag} */,
  {32'h4176bb58, 32'hc139fcc1} /* (4, 10, 31) {real, imag} */,
  {32'h3fa1578a, 32'hc129f866} /* (4, 10, 30) {real, imag} */,
  {32'hc1989a9f, 32'h41a23602} /* (4, 10, 29) {real, imag} */,
  {32'hc049591a, 32'h3feb2b8c} /* (4, 10, 28) {real, imag} */,
  {32'h41c2bee3, 32'h415f7075} /* (4, 10, 27) {real, imag} */,
  {32'h411f318c, 32'hc0cdbfd4} /* (4, 10, 26) {real, imag} */,
  {32'hc0a6dc0e, 32'hc0a58dfe} /* (4, 10, 25) {real, imag} */,
  {32'hc114c565, 32'h41b6e4c9} /* (4, 10, 24) {real, imag} */,
  {32'h404da5a8, 32'hbfb5c26f} /* (4, 10, 23) {real, imag} */,
  {32'hc110e90c, 32'h41490885} /* (4, 10, 22) {real, imag} */,
  {32'hc0d0fc34, 32'hc14e4c9a} /* (4, 10, 21) {real, imag} */,
  {32'h4163d019, 32'h40b8ee5a} /* (4, 10, 20) {real, imag} */,
  {32'hbfc2e5b0, 32'h4001ef3a} /* (4, 10, 19) {real, imag} */,
  {32'hc018bdc8, 32'h40943618} /* (4, 10, 18) {real, imag} */,
  {32'h3fb4f966, 32'h40c29718} /* (4, 10, 17) {real, imag} */,
  {32'h40150843, 32'h414d3674} /* (4, 10, 16) {real, imag} */,
  {32'h408e69dd, 32'hc08bf8c9} /* (4, 10, 15) {real, imag} */,
  {32'hc0ab5cd8, 32'h40eeacd3} /* (4, 10, 14) {real, imag} */,
  {32'hbffd0e64, 32'h40ca823c} /* (4, 10, 13) {real, imag} */,
  {32'h4198d087, 32'hc0d41000} /* (4, 10, 12) {real, imag} */,
  {32'h41a4c715, 32'h40f5e8d0} /* (4, 10, 11) {real, imag} */,
  {32'h411c961c, 32'hc111d848} /* (4, 10, 10) {real, imag} */,
  {32'hbea9cb40, 32'h416fd94e} /* (4, 10, 9) {real, imag} */,
  {32'hc10be33c, 32'h41034964} /* (4, 10, 8) {real, imag} */,
  {32'hc12cfcfa, 32'h410abef6} /* (4, 10, 7) {real, imag} */,
  {32'h418101bf, 32'h413a6e1c} /* (4, 10, 6) {real, imag} */,
  {32'h410ae95b, 32'hc1964c3e} /* (4, 10, 5) {real, imag} */,
  {32'hbf90d1b0, 32'hc0e468db} /* (4, 10, 4) {real, imag} */,
  {32'hc0d99177, 32'hc0f0a243} /* (4, 10, 3) {real, imag} */,
  {32'h419c9715, 32'h411a3eb5} /* (4, 10, 2) {real, imag} */,
  {32'hc1597c3b, 32'hbfa88c3e} /* (4, 10, 1) {real, imag} */,
  {32'hc183c667, 32'hc1a92d22} /* (4, 10, 0) {real, imag} */,
  {32'h410b6442, 32'hbf7435d0} /* (4, 9, 31) {real, imag} */,
  {32'h4048b4a4, 32'hbfda6310} /* (4, 9, 30) {real, imag} */,
  {32'hc07576c4, 32'hc15560b5} /* (4, 9, 29) {real, imag} */,
  {32'h4082b1e6, 32'hc0e508a4} /* (4, 9, 28) {real, imag} */,
  {32'h41b1bbc6, 32'h4181be5f} /* (4, 9, 27) {real, imag} */,
  {32'h41a8c2ad, 32'h4001ea50} /* (4, 9, 26) {real, imag} */,
  {32'hc0d5a559, 32'h415f8cf1} /* (4, 9, 25) {real, imag} */,
  {32'hc080a85d, 32'h408702c8} /* (4, 9, 24) {real, imag} */,
  {32'hc160d8c3, 32'hc1b468e2} /* (4, 9, 23) {real, imag} */,
  {32'hc0bc7260, 32'hc17998b5} /* (4, 9, 22) {real, imag} */,
  {32'hc08a4ea4, 32'hc13c2587} /* (4, 9, 21) {real, imag} */,
  {32'h40eca350, 32'h4192c51f} /* (4, 9, 20) {real, imag} */,
  {32'hc19d4502, 32'h3fdd1250} /* (4, 9, 19) {real, imag} */,
  {32'hc08b90d4, 32'h40fc0f7f} /* (4, 9, 18) {real, imag} */,
  {32'h408d9339, 32'h40e942b7} /* (4, 9, 17) {real, imag} */,
  {32'hc13b66d0, 32'hc1862175} /* (4, 9, 16) {real, imag} */,
  {32'hc001b6be, 32'hc08684ca} /* (4, 9, 15) {real, imag} */,
  {32'hc09cbca8, 32'hbfebb618} /* (4, 9, 14) {real, imag} */,
  {32'hc068e66c, 32'h3e652670} /* (4, 9, 13) {real, imag} */,
  {32'hc02f059b, 32'hc16f5fd4} /* (4, 9, 12) {real, imag} */,
  {32'hc163b1f2, 32'hc11cfedb} /* (4, 9, 11) {real, imag} */,
  {32'h4160bf4a, 32'hc17882b2} /* (4, 9, 10) {real, imag} */,
  {32'hc0f45db9, 32'h4092ba80} /* (4, 9, 9) {real, imag} */,
  {32'hc0169ac7, 32'hbe0840c0} /* (4, 9, 8) {real, imag} */,
  {32'h40505204, 32'h4094f5f6} /* (4, 9, 7) {real, imag} */,
  {32'hbff954a6, 32'h41034225} /* (4, 9, 6) {real, imag} */,
  {32'hc07974ac, 32'hc11b95cb} /* (4, 9, 5) {real, imag} */,
  {32'h401deec0, 32'hc16bca74} /* (4, 9, 4) {real, imag} */,
  {32'h4138de7e, 32'h41bdc7bc} /* (4, 9, 3) {real, imag} */,
  {32'h3fac7528, 32'h403cf69b} /* (4, 9, 2) {real, imag} */,
  {32'hc16a0e35, 32'hc0cd133a} /* (4, 9, 1) {real, imag} */,
  {32'hc0ace468, 32'h4174ddbd} /* (4, 9, 0) {real, imag} */,
  {32'h423e96a6, 32'h410b7fcf} /* (4, 8, 31) {real, imag} */,
  {32'hc20c18a4, 32'hc14378a6} /* (4, 8, 30) {real, imag} */,
  {32'h409e0f20, 32'h40d504e2} /* (4, 8, 29) {real, imag} */,
  {32'h415cc0f6, 32'hc03013d6} /* (4, 8, 28) {real, imag} */,
  {32'h40da4f68, 32'hc14aa07c} /* (4, 8, 27) {real, imag} */,
  {32'h40d6a198, 32'hc11450e8} /* (4, 8, 26) {real, imag} */,
  {32'hc1377614, 32'h40aac088} /* (4, 8, 25) {real, imag} */,
  {32'hc19d6e1d, 32'hc0aba6a3} /* (4, 8, 24) {real, imag} */,
  {32'hc1a4db44, 32'hc1080e71} /* (4, 8, 23) {real, imag} */,
  {32'hc151cd81, 32'h41206be6} /* (4, 8, 22) {real, imag} */,
  {32'h3f7a9ac8, 32'h4156ecc7} /* (4, 8, 21) {real, imag} */,
  {32'h413f15fd, 32'hc175e13e} /* (4, 8, 20) {real, imag} */,
  {32'hc124bbd2, 32'h4117fa5e} /* (4, 8, 19) {real, imag} */,
  {32'h40406782, 32'h4018b7ca} /* (4, 8, 18) {real, imag} */,
  {32'h4119801e, 32'h404fb8c2} /* (4, 8, 17) {real, imag} */,
  {32'h3e19a478, 32'hc10f44ca} /* (4, 8, 16) {real, imag} */,
  {32'hbfde8f66, 32'hbedd7da8} /* (4, 8, 15) {real, imag} */,
  {32'h41085a50, 32'h4189a7e1} /* (4, 8, 14) {real, imag} */,
  {32'h40b5ac29, 32'hc15ccfc0} /* (4, 8, 13) {real, imag} */,
  {32'hc05cd5b1, 32'h408f38d0} /* (4, 8, 12) {real, imag} */,
  {32'hc104945a, 32'hbc70ea00} /* (4, 8, 11) {real, imag} */,
  {32'h418e1ac9, 32'hbfe0d3f0} /* (4, 8, 10) {real, imag} */,
  {32'h414cecfc, 32'h419ba022} /* (4, 8, 9) {real, imag} */,
  {32'hc10a4634, 32'h40ebaaee} /* (4, 8, 8) {real, imag} */,
  {32'hc0b40eec, 32'h4027aa38} /* (4, 8, 7) {real, imag} */,
  {32'hc0c8d5a6, 32'h4149d87e} /* (4, 8, 6) {real, imag} */,
  {32'hbe8eb100, 32'hc18d97ea} /* (4, 8, 5) {real, imag} */,
  {32'hc0865ddb, 32'hbf86cc7c} /* (4, 8, 4) {real, imag} */,
  {32'hbfc31862, 32'h3fc46f18} /* (4, 8, 3) {real, imag} */,
  {32'hc1a86cd2, 32'hc190e353} /* (4, 8, 2) {real, imag} */,
  {32'hbff1f918, 32'h4165830c} /* (4, 8, 1) {real, imag} */,
  {32'h41af95a3, 32'h42092d0c} /* (4, 8, 0) {real, imag} */,
  {32'hc1dc7086, 32'hbf37d3cc} /* (4, 7, 31) {real, imag} */,
  {32'hc098814a, 32'h41dac3cc} /* (4, 7, 30) {real, imag} */,
  {32'hc1150396, 32'hc1357b46} /* (4, 7, 29) {real, imag} */,
  {32'hc18f8df0, 32'hc1b938dc} /* (4, 7, 28) {real, imag} */,
  {32'h41a061da, 32'h40dc7b8c} /* (4, 7, 27) {real, imag} */,
  {32'h412e43f3, 32'hc0e014c9} /* (4, 7, 26) {real, imag} */,
  {32'h4078483a, 32'hc0bd772a} /* (4, 7, 25) {real, imag} */,
  {32'hc1537006, 32'hc191a78a} /* (4, 7, 24) {real, imag} */,
  {32'hbfbd584e, 32'h41532650} /* (4, 7, 23) {real, imag} */,
  {32'hbfe918f8, 32'hc125e41c} /* (4, 7, 22) {real, imag} */,
  {32'hc0a2fec1, 32'h41807f1a} /* (4, 7, 21) {real, imag} */,
  {32'h411cd558, 32'hc0a34132} /* (4, 7, 20) {real, imag} */,
  {32'hc0d06284, 32'h41764ad2} /* (4, 7, 19) {real, imag} */,
  {32'h417a3896, 32'hc0d5b06f} /* (4, 7, 18) {real, imag} */,
  {32'hbf603174, 32'h41219cce} /* (4, 7, 17) {real, imag} */,
  {32'h4159987f, 32'hc06a32b2} /* (4, 7, 16) {real, imag} */,
  {32'hc1601659, 32'hc18135a8} /* (4, 7, 15) {real, imag} */,
  {32'hc1714e8a, 32'hbf4ad230} /* (4, 7, 14) {real, imag} */,
  {32'hc19e20eb, 32'h4130b5a8} /* (4, 7, 13) {real, imag} */,
  {32'hc1ade3e2, 32'h40293420} /* (4, 7, 12) {real, imag} */,
  {32'hc0ae9a42, 32'h41357e0f} /* (4, 7, 11) {real, imag} */,
  {32'h40a70dfa, 32'hc0ca626a} /* (4, 7, 10) {real, imag} */,
  {32'h412b1276, 32'h403bbd5c} /* (4, 7, 9) {real, imag} */,
  {32'h40ae003e, 32'hbf775d50} /* (4, 7, 8) {real, imag} */,
  {32'hc1988057, 32'h411e5b11} /* (4, 7, 7) {real, imag} */,
  {32'h411e4c54, 32'h402cc3eb} /* (4, 7, 6) {real, imag} */,
  {32'h4209f01a, 32'h41c63306} /* (4, 7, 5) {real, imag} */,
  {32'hc16db3c9, 32'hc14112b2} /* (4, 7, 4) {real, imag} */,
  {32'hbe76f0c0, 32'h41067624} /* (4, 7, 3) {real, imag} */,
  {32'h4196639d, 32'h41253c32} /* (4, 7, 2) {real, imag} */,
  {32'h3e229c00, 32'hc1de5ed0} /* (4, 7, 1) {real, imag} */,
  {32'hc1c6088a, 32'hc11a5c4a} /* (4, 7, 0) {real, imag} */,
  {32'h418566bc, 32'h41a71802} /* (4, 6, 31) {real, imag} */,
  {32'h415b9333, 32'h3ec951e0} /* (4, 6, 30) {real, imag} */,
  {32'h41b2089d, 32'h3f3828b0} /* (4, 6, 29) {real, imag} */,
  {32'h400c20e0, 32'hbf883090} /* (4, 6, 28) {real, imag} */,
  {32'h3fb00010, 32'h419e2a76} /* (4, 6, 27) {real, imag} */,
  {32'hbfde71a8, 32'hc0ecfeaa} /* (4, 6, 26) {real, imag} */,
  {32'hbf4943f4, 32'hc1125770} /* (4, 6, 25) {real, imag} */,
  {32'hc1092ce3, 32'h41474fc6} /* (4, 6, 24) {real, imag} */,
  {32'hc16b0d7a, 32'hc098251d} /* (4, 6, 23) {real, imag} */,
  {32'hc0868bab, 32'h41836a8e} /* (4, 6, 22) {real, imag} */,
  {32'hc0f6a4e3, 32'hc1a0ff26} /* (4, 6, 21) {real, imag} */,
  {32'hc1a9831d, 32'h40d13631} /* (4, 6, 20) {real, imag} */,
  {32'hc0c69ca9, 32'hc0912fe4} /* (4, 6, 19) {real, imag} */,
  {32'h407843ba, 32'h3f3136bc} /* (4, 6, 18) {real, imag} */,
  {32'h40f2f80c, 32'hc028b098} /* (4, 6, 17) {real, imag} */,
  {32'h400cfa67, 32'hc095ce90} /* (4, 6, 16) {real, imag} */,
  {32'hbed222a8, 32'h4007ce34} /* (4, 6, 15) {real, imag} */,
  {32'hbfcd22e8, 32'hc145f147} /* (4, 6, 14) {real, imag} */,
  {32'h4180fb91, 32'hc07e01a6} /* (4, 6, 13) {real, imag} */,
  {32'h40ecc65e, 32'h40658426} /* (4, 6, 12) {real, imag} */,
  {32'hc14d18c7, 32'h40d4a510} /* (4, 6, 11) {real, imag} */,
  {32'h3f3c4608, 32'hc0493292} /* (4, 6, 10) {real, imag} */,
  {32'h40cf6151, 32'hbf319528} /* (4, 6, 9) {real, imag} */,
  {32'hc1aaf1fe, 32'hbf48a370} /* (4, 6, 8) {real, imag} */,
  {32'h412255d4, 32'h41340a5b} /* (4, 6, 7) {real, imag} */,
  {32'hc1a2dcb0, 32'hc11ad7a4} /* (4, 6, 6) {real, imag} */,
  {32'hc09d9fa9, 32'h40c1d63a} /* (4, 6, 5) {real, imag} */,
  {32'hc0b9af60, 32'hc11a5db0} /* (4, 6, 4) {real, imag} */,
  {32'hc134a0be, 32'h40c159b7} /* (4, 6, 3) {real, imag} */,
  {32'hc1ae8ad9, 32'hc0891fca} /* (4, 6, 2) {real, imag} */,
  {32'h4188b211, 32'h4144fc49} /* (4, 6, 1) {real, imag} */,
  {32'h4151757b, 32'hc1926d0f} /* (4, 6, 0) {real, imag} */,
  {32'h425a6421, 32'h41b24c80} /* (4, 5, 31) {real, imag} */,
  {32'hc22feab3, 32'hc14d9c0a} /* (4, 5, 30) {real, imag} */,
  {32'hc03b7eaa, 32'hc13b7e25} /* (4, 5, 29) {real, imag} */,
  {32'h41ba9428, 32'hc1af9882} /* (4, 5, 28) {real, imag} */,
  {32'hc1a819a3, 32'hc0999575} /* (4, 5, 27) {real, imag} */,
  {32'hc11a5dea, 32'h41295625} /* (4, 5, 26) {real, imag} */,
  {32'h41c45c7e, 32'h4127cbc8} /* (4, 5, 25) {real, imag} */,
  {32'hc10a68f8, 32'hbfcbb67e} /* (4, 5, 24) {real, imag} */,
  {32'h40b5de95, 32'hc1610bf2} /* (4, 5, 23) {real, imag} */,
  {32'hc0076fa0, 32'h3f15ce48} /* (4, 5, 22) {real, imag} */,
  {32'hc10a65c0, 32'h41e962b4} /* (4, 5, 21) {real, imag} */,
  {32'hc0ede98c, 32'h408eaf0e} /* (4, 5, 20) {real, imag} */,
  {32'hc13a10a6, 32'h3fa54dc0} /* (4, 5, 19) {real, imag} */,
  {32'h412fd40e, 32'h40e0cafe} /* (4, 5, 18) {real, imag} */,
  {32'hc0e1e64c, 32'h40f4062e} /* (4, 5, 17) {real, imag} */,
  {32'hc007ff72, 32'h41024680} /* (4, 5, 16) {real, imag} */,
  {32'h40e91b94, 32'hc0a48f20} /* (4, 5, 15) {real, imag} */,
  {32'h412a229e, 32'hc0df34f4} /* (4, 5, 14) {real, imag} */,
  {32'hc050a042, 32'hc12a4d8f} /* (4, 5, 13) {real, imag} */,
  {32'hc0984681, 32'h404bee1c} /* (4, 5, 12) {real, imag} */,
  {32'hc055cc9e, 32'hc1d22e0e} /* (4, 5, 11) {real, imag} */,
  {32'h40dbab23, 32'h418dbbd8} /* (4, 5, 10) {real, imag} */,
  {32'hbed7a1f0, 32'h3fb3ff90} /* (4, 5, 9) {real, imag} */,
  {32'h404c4244, 32'hc048e5ae} /* (4, 5, 8) {real, imag} */,
  {32'hbf94a736, 32'h409b60f2} /* (4, 5, 7) {real, imag} */,
  {32'hc12a11f4, 32'hc15aaea5} /* (4, 5, 6) {real, imag} */,
  {32'hc1cd0fde, 32'hc1f5e207} /* (4, 5, 5) {real, imag} */,
  {32'h418ac180, 32'hc0f32361} /* (4, 5, 4) {real, imag} */,
  {32'h41a8b277, 32'h40641184} /* (4, 5, 3) {real, imag} */,
  {32'h40f9080c, 32'h41c62afb} /* (4, 5, 2) {real, imag} */,
  {32'h42a47c5e, 32'h42217a40} /* (4, 5, 1) {real, imag} */,
  {32'h42a3bf55, 32'hc0b2cd1c} /* (4, 5, 0) {real, imag} */,
  {32'hc2223b39, 32'hc2a4f48e} /* (4, 4, 31) {real, imag} */,
  {32'h42291cb5, 32'h42b9daec} /* (4, 4, 30) {real, imag} */,
  {32'hc0c83d1a, 32'h40f2d4fc} /* (4, 4, 29) {real, imag} */,
  {32'hc18fc2ba, 32'h40f3c6e3} /* (4, 4, 28) {real, imag} */,
  {32'h3faa71c2, 32'hc16c7ef0} /* (4, 4, 27) {real, imag} */,
  {32'hc223cb80, 32'hc1398b2c} /* (4, 4, 26) {real, imag} */,
  {32'h4113b0b0, 32'h3e09ec20} /* (4, 4, 25) {real, imag} */,
  {32'h4116f687, 32'hbeb75778} /* (4, 4, 24) {real, imag} */,
  {32'h3fa460c8, 32'h407ec0db} /* (4, 4, 23) {real, imag} */,
  {32'h412dcdbb, 32'hc057924f} /* (4, 4, 22) {real, imag} */,
  {32'h41f2c0ca, 32'hc0fdac7d} /* (4, 4, 21) {real, imag} */,
  {32'hc091bdc4, 32'h4089679a} /* (4, 4, 20) {real, imag} */,
  {32'h40d7c127, 32'hc0aafcbc} /* (4, 4, 19) {real, imag} */,
  {32'h3d8bd940, 32'h40d4eab6} /* (4, 4, 18) {real, imag} */,
  {32'hc03e688e, 32'h413b3a58} /* (4, 4, 17) {real, imag} */,
  {32'hc0cf493b, 32'hc0fd1e16} /* (4, 4, 16) {real, imag} */,
  {32'hc0fb58e8, 32'hbfa74958} /* (4, 4, 15) {real, imag} */,
  {32'hc0479f21, 32'h41515276} /* (4, 4, 14) {real, imag} */,
  {32'hc08385e5, 32'hc01add16} /* (4, 4, 13) {real, imag} */,
  {32'hbf28b274, 32'hbeeca9c0} /* (4, 4, 12) {real, imag} */,
  {32'hbedfd01c, 32'hc128f18f} /* (4, 4, 11) {real, imag} */,
  {32'h4144f75c, 32'hc159ae4a} /* (4, 4, 10) {real, imag} */,
  {32'hbefef2d0, 32'h4156adb8} /* (4, 4, 9) {real, imag} */,
  {32'h40348c1a, 32'h410dd106} /* (4, 4, 8) {real, imag} */,
  {32'hc1a56632, 32'h40d1664a} /* (4, 4, 7) {real, imag} */,
  {32'h405ecf00, 32'hc12c1a5e} /* (4, 4, 6) {real, imag} */,
  {32'h41a74907, 32'hc0bdd40c} /* (4, 4, 5) {real, imag} */,
  {32'h41b820bc, 32'hc1875424} /* (4, 4, 4) {real, imag} */,
  {32'hc19e1673, 32'h41e59480} /* (4, 4, 3) {real, imag} */,
  {32'h42b21df1, 32'h424393a6} /* (4, 4, 2) {real, imag} */,
  {32'hc318991c, 32'hc24626ac} /* (4, 4, 1) {real, imag} */,
  {32'hc237cfd6, 32'hc1204cc8} /* (4, 4, 0) {real, imag} */,
  {32'h42a89fe7, 32'hc2597180} /* (4, 3, 31) {real, imag} */,
  {32'hc23ae113, 32'h420d1e00} /* (4, 3, 30) {real, imag} */,
  {32'hbef56a00, 32'h410f23ed} /* (4, 3, 29) {real, imag} */,
  {32'hc1cb52c6, 32'hc138f8bd} /* (4, 3, 28) {real, imag} */,
  {32'h42017646, 32'hc1c49091} /* (4, 3, 27) {real, imag} */,
  {32'hc0fd5344, 32'hc16bf55c} /* (4, 3, 26) {real, imag} */,
  {32'hc0f9a733, 32'h4151590e} /* (4, 3, 25) {real, imag} */,
  {32'h4078f89e, 32'h41b2c1a8} /* (4, 3, 24) {real, imag} */,
  {32'hc0a0fa2c, 32'hc1979d86} /* (4, 3, 23) {real, imag} */,
  {32'h41301c06, 32'hc17bac9d} /* (4, 3, 22) {real, imag} */,
  {32'hc1273458, 32'hc0fa333c} /* (4, 3, 21) {real, imag} */,
  {32'h3fcae430, 32'hbe49e8f4} /* (4, 3, 20) {real, imag} */,
  {32'hc0f9d999, 32'hc0d17123} /* (4, 3, 19) {real, imag} */,
  {32'hc196f64a, 32'hc0631ac6} /* (4, 3, 18) {real, imag} */,
  {32'h411d0c24, 32'h4037d1b9} /* (4, 3, 17) {real, imag} */,
  {32'h411a36fe, 32'hc128093b} /* (4, 3, 16) {real, imag} */,
  {32'h4096a47c, 32'h3e8ec6a8} /* (4, 3, 15) {real, imag} */,
  {32'hbfb58f34, 32'h4152fef7} /* (4, 3, 14) {real, imag} */,
  {32'h411d5c2e, 32'h404cbda8} /* (4, 3, 13) {real, imag} */,
  {32'h411e4222, 32'hc11d30db} /* (4, 3, 12) {real, imag} */,
  {32'hc1704451, 32'hc084d772} /* (4, 3, 11) {real, imag} */,
  {32'h3f945574, 32'hc08afe0c} /* (4, 3, 10) {real, imag} */,
  {32'hc0aa23b5, 32'hc052ad2c} /* (4, 3, 9) {real, imag} */,
  {32'h3f552ca8, 32'h41670325} /* (4, 3, 8) {real, imag} */,
  {32'hc091466c, 32'hc1f8531c} /* (4, 3, 7) {real, imag} */,
  {32'h3e685580, 32'hc126a326} /* (4, 3, 6) {real, imag} */,
  {32'hc1daba0f, 32'hc11c7bec} /* (4, 3, 5) {real, imag} */,
  {32'h41d50140, 32'hc1be00e3} /* (4, 3, 4) {real, imag} */,
  {32'hc10f8a99, 32'hc18e8801} /* (4, 3, 3) {real, imag} */,
  {32'h415b17d7, 32'h42e13b1e} /* (4, 3, 2) {real, imag} */,
  {32'hc2978967, 32'h412990d8} /* (4, 3, 1) {real, imag} */,
  {32'h4153a6a1, 32'h41ccb1aa} /* (4, 3, 0) {real, imag} */,
  {32'h43eccb8f, 32'h41e09371} /* (4, 2, 31) {real, imag} */,
  {32'hc36d9e45, 32'h424bfea8} /* (4, 2, 30) {real, imag} */,
  {32'h3f76fe20, 32'h41f4cdb0} /* (4, 2, 29) {real, imag} */,
  {32'h411b3a96, 32'hc28ba956} /* (4, 2, 28) {real, imag} */,
  {32'hc2477ed0, 32'h41a7ce8e} /* (4, 2, 27) {real, imag} */,
  {32'hc1d336de, 32'h41ff7bee} /* (4, 2, 26) {real, imag} */,
  {32'h410819cc, 32'hc20ac40f} /* (4, 2, 25) {real, imag} */,
  {32'hc121c3ec, 32'h427ee26a} /* (4, 2, 24) {real, imag} */,
  {32'hc122c4dc, 32'h40a27409} /* (4, 2, 23) {real, imag} */,
  {32'h3f00fd80, 32'h4124ad02} /* (4, 2, 22) {real, imag} */,
  {32'hc1276fd4, 32'h41a028fa} /* (4, 2, 21) {real, imag} */,
  {32'h412518f8, 32'hc0616509} /* (4, 2, 20) {real, imag} */,
  {32'hc0667f96, 32'hc10bb15a} /* (4, 2, 19) {real, imag} */,
  {32'h409776e0, 32'h40690e34} /* (4, 2, 18) {real, imag} */,
  {32'hbfa36e56, 32'hc18d98d2} /* (4, 2, 17) {real, imag} */,
  {32'h40e6aef0, 32'hc0d2a889} /* (4, 2, 16) {real, imag} */,
  {32'h409adc31, 32'h413aa487} /* (4, 2, 15) {real, imag} */,
  {32'hc098bb90, 32'hc19c22a7} /* (4, 2, 14) {real, imag} */,
  {32'hc0bd1688, 32'hc08bf04b} /* (4, 2, 13) {real, imag} */,
  {32'h41347e97, 32'h411c15f8} /* (4, 2, 12) {real, imag} */,
  {32'hc11bf068, 32'hc12c79e1} /* (4, 2, 11) {real, imag} */,
  {32'h410ce546, 32'h41ad22cf} /* (4, 2, 10) {real, imag} */,
  {32'h40bc9e98, 32'h409f63ce} /* (4, 2, 9) {real, imag} */,
  {32'hc1f238c7, 32'hc146e651} /* (4, 2, 8) {real, imag} */,
  {32'h41b1302c, 32'hc0e13a6d} /* (4, 2, 7) {real, imag} */,
  {32'h4138a4d6, 32'h418b1eda} /* (4, 2, 6) {real, imag} */,
  {32'hc1a71aba, 32'hc2713038} /* (4, 2, 5) {real, imag} */,
  {32'h42b5abc9, 32'h40a026fe} /* (4, 2, 4) {real, imag} */,
  {32'hc17a7a2c, 32'h4114b956} /* (4, 2, 3) {real, imag} */,
  {32'hc3631e4d, 32'h42f92c8a} /* (4, 2, 2) {real, imag} */,
  {32'h4389ad3f, 32'h3fe65600} /* (4, 2, 1) {real, imag} */,
  {32'h432f23e6, 32'h410f84c4} /* (4, 2, 0) {real, imag} */,
  {32'hc3931668, 32'h419a93d0} /* (4, 1, 31) {real, imag} */,
  {32'h43268dc8, 32'h41fc72eb} /* (4, 1, 30) {real, imag} */,
  {32'h42482ec2, 32'hc220f71e} /* (4, 1, 29) {real, imag} */,
  {32'hc25eee70, 32'hc28f469a} /* (4, 1, 28) {real, imag} */,
  {32'h42cb796e, 32'h40a90a2e} /* (4, 1, 27) {real, imag} */,
  {32'h4176b5ca, 32'hc18101b6} /* (4, 1, 26) {real, imag} */,
  {32'hc1c1b6c6, 32'hc07e6a5a} /* (4, 1, 25) {real, imag} */,
  {32'h41bacac0, 32'hc14b082a} /* (4, 1, 24) {real, imag} */,
  {32'hc088855e, 32'h401f0d88} /* (4, 1, 23) {real, imag} */,
  {32'hc0ad9324, 32'hc18bf683} /* (4, 1, 22) {real, imag} */,
  {32'h41bf87c2, 32'hc10fe028} /* (4, 1, 21) {real, imag} */,
  {32'h40614bda, 32'h405941ec} /* (4, 1, 20) {real, imag} */,
  {32'h40b40592, 32'hc0c212ce} /* (4, 1, 19) {real, imag} */,
  {32'h4096341b, 32'hc18e4304} /* (4, 1, 18) {real, imag} */,
  {32'h411b17d8, 32'h4127b11e} /* (4, 1, 17) {real, imag} */,
  {32'hc1563d96, 32'hc107be28} /* (4, 1, 16) {real, imag} */,
  {32'h4139a562, 32'h401c5e2a} /* (4, 1, 15) {real, imag} */,
  {32'hc1c63230, 32'h4191c066} /* (4, 1, 14) {real, imag} */,
  {32'h40b73c2e, 32'hc05aeacf} /* (4, 1, 13) {real, imag} */,
  {32'hc06e09ec, 32'hc0ad394b} /* (4, 1, 12) {real, imag} */,
  {32'hc0bbadc9, 32'h418922e1} /* (4, 1, 11) {real, imag} */,
  {32'h4100b80e, 32'h4071e4ad} /* (4, 1, 10) {real, imag} */,
  {32'hc1aba055, 32'h4185b886} /* (4, 1, 9) {real, imag} */,
  {32'h3f874130, 32'h42164f38} /* (4, 1, 8) {real, imag} */,
  {32'hc16b9284, 32'hc0351bf0} /* (4, 1, 7) {real, imag} */,
  {32'hc1b11f6b, 32'hc1cbc0dd} /* (4, 1, 6) {real, imag} */,
  {32'h4278e9ef, 32'h41d3ca10} /* (4, 1, 5) {real, imag} */,
  {32'h409f04c4, 32'hc223ec2c} /* (4, 1, 4) {real, imag} */,
  {32'h414bffd6, 32'hc24b2118} /* (4, 1, 3) {real, imag} */,
  {32'h436356ee, 32'h433bd49a} /* (4, 1, 2) {real, imag} */,
  {32'hc3bb4b8d, 32'hc3ad18d3} /* (4, 1, 1) {real, imag} */,
  {32'hc1a2e928, 32'h425fb30c} /* (4, 1, 0) {real, imag} */,
  {32'hc3002b48, 32'h428b010e} /* (4, 0, 31) {real, imag} */,
  {32'h42b178a0, 32'hc20606a2} /* (4, 0, 30) {real, imag} */,
  {32'h42abe6c6, 32'hc241d192} /* (4, 0, 29) {real, imag} */,
  {32'hc15b2781, 32'hc292e12e} /* (4, 0, 28) {real, imag} */,
  {32'h4235b418, 32'hc0469068} /* (4, 0, 27) {real, imag} */,
  {32'h42127170, 32'h41191dd9} /* (4, 0, 26) {real, imag} */,
  {32'hc0477c15, 32'h41157b5c} /* (4, 0, 25) {real, imag} */,
  {32'hc1b2e364, 32'hc1ad7932} /* (4, 0, 24) {real, imag} */,
  {32'h4031fdf6, 32'hc110a344} /* (4, 0, 23) {real, imag} */,
  {32'hc141cffa, 32'hc12c7ff3} /* (4, 0, 22) {real, imag} */,
  {32'hc123e3a0, 32'hbdcf8200} /* (4, 0, 21) {real, imag} */,
  {32'hc149125f, 32'h40ad5d7f} /* (4, 0, 20) {real, imag} */,
  {32'h41631407, 32'hbfab79c4} /* (4, 0, 19) {real, imag} */,
  {32'h410c9958, 32'hc0ba2333} /* (4, 0, 18) {real, imag} */,
  {32'h3f0a8574, 32'h40e0d6f9} /* (4, 0, 17) {real, imag} */,
  {32'hc0b04bee, 32'h00000000} /* (4, 0, 16) {real, imag} */,
  {32'h3f0a8574, 32'hc0e0d6f9} /* (4, 0, 15) {real, imag} */,
  {32'h410c9958, 32'h40ba2333} /* (4, 0, 14) {real, imag} */,
  {32'h41631407, 32'h3fab79c4} /* (4, 0, 13) {real, imag} */,
  {32'hc149125f, 32'hc0ad5d7f} /* (4, 0, 12) {real, imag} */,
  {32'hc123e3a0, 32'h3dcf8200} /* (4, 0, 11) {real, imag} */,
  {32'hc141cffa, 32'h412c7ff3} /* (4, 0, 10) {real, imag} */,
  {32'h4031fdf6, 32'h4110a344} /* (4, 0, 9) {real, imag} */,
  {32'hc1b2e364, 32'h41ad7932} /* (4, 0, 8) {real, imag} */,
  {32'hc0477c15, 32'hc1157b5c} /* (4, 0, 7) {real, imag} */,
  {32'h42127170, 32'hc1191dd9} /* (4, 0, 6) {real, imag} */,
  {32'h4235b418, 32'h40469068} /* (4, 0, 5) {real, imag} */,
  {32'hc15b2781, 32'h4292e12e} /* (4, 0, 4) {real, imag} */,
  {32'h42abe6c6, 32'h4241d192} /* (4, 0, 3) {real, imag} */,
  {32'h42b178a0, 32'h420606a2} /* (4, 0, 2) {real, imag} */,
  {32'hc3002b48, 32'hc28b010e} /* (4, 0, 1) {real, imag} */,
  {32'h43fd0662, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hc4444884, 32'h440832a4} /* (3, 31, 31) {real, imag} */,
  {32'h439a0f1a, 32'hc38021d2} /* (3, 31, 30) {real, imag} */,
  {32'h421b1624, 32'h41bd9cc4} /* (3, 31, 29) {real, imag} */,
  {32'hc203f346, 32'h41f47e24} /* (3, 31, 28) {real, imag} */,
  {32'h427f9bfe, 32'hc276da63} /* (3, 31, 27) {real, imag} */,
  {32'hc06fcfec, 32'h40dba976} /* (3, 31, 26) {real, imag} */,
  {32'hc0dd5c60, 32'h418e732e} /* (3, 31, 25) {real, imag} */,
  {32'h415d3728, 32'hc22ee7e5} /* (3, 31, 24) {real, imag} */,
  {32'hc142dda8, 32'hc074d03e} /* (3, 31, 23) {real, imag} */,
  {32'h4108b990, 32'hc14f17c0} /* (3, 31, 22) {real, imag} */,
  {32'h41717016, 32'hc1a7e156} /* (3, 31, 21) {real, imag} */,
  {32'hc10f4d6d, 32'hc02a845d} /* (3, 31, 20) {real, imag} */,
  {32'hbfec08e1, 32'h41154215} /* (3, 31, 19) {real, imag} */,
  {32'hc09c4f4c, 32'hc09673d0} /* (3, 31, 18) {real, imag} */,
  {32'h4120b3ae, 32'hc0b2bac3} /* (3, 31, 17) {real, imag} */,
  {32'h411d0f66, 32'hbed563e0} /* (3, 31, 16) {real, imag} */,
  {32'h40f64116, 32'hbfeefffc} /* (3, 31, 15) {real, imag} */,
  {32'hc0f6c315, 32'h416605fe} /* (3, 31, 14) {real, imag} */,
  {32'h3ffc7ecc, 32'h3ffe7eaa} /* (3, 31, 13) {real, imag} */,
  {32'hc0184bf1, 32'hc08f84c3} /* (3, 31, 12) {real, imag} */,
  {32'h41f3d926, 32'h41a0416a} /* (3, 31, 11) {real, imag} */,
  {32'hc0f5bda2, 32'hc0706ba6} /* (3, 31, 10) {real, imag} */,
  {32'hc0f88bdc, 32'h3fe695f0} /* (3, 31, 9) {real, imag} */,
  {32'h41ab861f, 32'h41c4082b} /* (3, 31, 8) {real, imag} */,
  {32'hc1a3b710, 32'hc1069f60} /* (3, 31, 7) {real, imag} */,
  {32'h4215c0bb, 32'h41480d04} /* (3, 31, 6) {real, imag} */,
  {32'h42fbad4c, 32'h40c5e14c} /* (3, 31, 5) {real, imag} */,
  {32'hc2b54e47, 32'h424cad5a} /* (3, 31, 4) {real, imag} */,
  {32'h425ce602, 32'h42227adc} /* (3, 31, 3) {real, imag} */,
  {32'h437b0f50, 32'hc22efbf8} /* (3, 31, 2) {real, imag} */,
  {32'hc4110235, 32'hc2bfa448} /* (3, 31, 1) {real, imag} */,
  {32'hc3a818e4, 32'hc205d494} /* (3, 31, 0) {real, imag} */,
  {32'h43c3a854, 32'h41585dc0} /* (3, 30, 31) {real, imag} */,
  {32'hc38d518a, 32'hc30a34a9} /* (3, 30, 30) {real, imag} */,
  {32'hc2169306, 32'hc08134c8} /* (3, 30, 29) {real, imag} */,
  {32'h42c8385c, 32'h40db6714} /* (3, 30, 28) {real, imag} */,
  {32'hc23ca142, 32'h4216aa0b} /* (3, 30, 27) {real, imag} */,
  {32'h412c336c, 32'hbf389968} /* (3, 30, 26) {real, imag} */,
  {32'h420a966e, 32'h412a65c0} /* (3, 30, 25) {real, imag} */,
  {32'hc1ea1dc3, 32'hbf1eed90} /* (3, 30, 24) {real, imag} */,
  {32'h40db206a, 32'h41481ca8} /* (3, 30, 23) {real, imag} */,
  {32'h417132e3, 32'hbdc7f600} /* (3, 30, 22) {real, imag} */,
  {32'hc14d68e3, 32'hc1540cdc} /* (3, 30, 21) {real, imag} */,
  {32'h41ae555e, 32'h3fdd6fe0} /* (3, 30, 20) {real, imag} */,
  {32'hc06b1114, 32'h4045d86c} /* (3, 30, 19) {real, imag} */,
  {32'h4019eede, 32'h41501514} /* (3, 30, 18) {real, imag} */,
  {32'h419017f2, 32'h413d9e46} /* (3, 30, 17) {real, imag} */,
  {32'h401a680a, 32'h3f951ce0} /* (3, 30, 16) {real, imag} */,
  {32'h4018a610, 32'hc10d610e} /* (3, 30, 15) {real, imag} */,
  {32'hc0630920, 32'hc1870199} /* (3, 30, 14) {real, imag} */,
  {32'hbffa1530, 32'hc124b86a} /* (3, 30, 13) {real, imag} */,
  {32'h400c8370, 32'h4121a997} /* (3, 30, 12) {real, imag} */,
  {32'hc130dc3a, 32'hc1eaa619} /* (3, 30, 11) {real, imag} */,
  {32'h418021a0, 32'h419acde5} /* (3, 30, 10) {real, imag} */,
  {32'hc1e1a859, 32'h411e5474} /* (3, 30, 9) {real, imag} */,
  {32'hc20256fc, 32'hc19dd252} /* (3, 30, 8) {real, imag} */,
  {32'h41c076aa, 32'h41a78db5} /* (3, 30, 7) {real, imag} */,
  {32'hc189978d, 32'hbf95b70c} /* (3, 30, 6) {real, imag} */,
  {32'hc246582c, 32'hc23746a4} /* (3, 30, 5) {real, imag} */,
  {32'h41f495c3, 32'h4285928a} /* (3, 30, 4) {real, imag} */,
  {32'h41c1b4d3, 32'hc2349180} /* (3, 30, 3) {real, imag} */,
  {32'hc3a7120c, 32'hc2bdd0ef} /* (3, 30, 2) {real, imag} */,
  {32'h44276ee7, 32'hc246afd1} /* (3, 30, 1) {real, imag} */,
  {32'h438ead27, 32'hc2a03054} /* (3, 30, 0) {real, imag} */,
  {32'hc2d74aea, 32'h41cdef58} /* (3, 29, 31) {real, imag} */,
  {32'hc15396bb, 32'hc30631b4} /* (3, 29, 30) {real, imag} */,
  {32'hc2239ca2, 32'h42361e24} /* (3, 29, 29) {real, imag} */,
  {32'h422999f5, 32'hc08b924e} /* (3, 29, 28) {real, imag} */,
  {32'hc21c85a2, 32'hc1bb0683} /* (3, 29, 27) {real, imag} */,
  {32'h3f83ae38, 32'h41f179c1} /* (3, 29, 26) {real, imag} */,
  {32'h40fb7fe4, 32'h41fdbab3} /* (3, 29, 25) {real, imag} */,
  {32'hc08270ca, 32'hc1789a55} /* (3, 29, 24) {real, imag} */,
  {32'h41d28e27, 32'hc0a75646} /* (3, 29, 23) {real, imag} */,
  {32'hbedf8084, 32'h410457ae} /* (3, 29, 22) {real, imag} */,
  {32'hc1b133de, 32'h41953ff2} /* (3, 29, 21) {real, imag} */,
  {32'hc08284ce, 32'hc0fcf968} /* (3, 29, 20) {real, imag} */,
  {32'hc1a6515f, 32'h3f0dd438} /* (3, 29, 19) {real, imag} */,
  {32'h4047d21b, 32'hc1b52ec5} /* (3, 29, 18) {real, imag} */,
  {32'hc0fa3db0, 32'h3f4ef150} /* (3, 29, 17) {real, imag} */,
  {32'hc0df8e05, 32'h409e2474} /* (3, 29, 16) {real, imag} */,
  {32'hc0e490de, 32'hbff1d8f6} /* (3, 29, 15) {real, imag} */,
  {32'hc0815074, 32'h3fb52572} /* (3, 29, 14) {real, imag} */,
  {32'h4119d8fd, 32'hbf500d48} /* (3, 29, 13) {real, imag} */,
  {32'hbf3e50f8, 32'hc0ff4ea1} /* (3, 29, 12) {real, imag} */,
  {32'h403f9ba4, 32'h4193fba6} /* (3, 29, 11) {real, imag} */,
  {32'h40da1afa, 32'hc11d646e} /* (3, 29, 10) {real, imag} */,
  {32'hc16c682b, 32'h4192afbf} /* (3, 29, 9) {real, imag} */,
  {32'hc00a957c, 32'hc204ae04} /* (3, 29, 8) {real, imag} */,
  {32'hc09dcb9f, 32'hc0404326} /* (3, 29, 7) {real, imag} */,
  {32'hc03e99dc, 32'hc0d98268} /* (3, 29, 6) {real, imag} */,
  {32'h42140c60, 32'h400b7768} /* (3, 29, 5) {real, imag} */,
  {32'hc146ea7d, 32'h411f9c17} /* (3, 29, 4) {real, imag} */,
  {32'hc0dd3dea, 32'h41d41960} /* (3, 29, 3) {real, imag} */,
  {32'hc279392a, 32'hc23e9b4f} /* (3, 29, 2) {real, imag} */,
  {32'h430d693c, 32'h4243905a} /* (3, 29, 1) {real, imag} */,
  {32'h41af1a47, 32'h41a46520} /* (3, 29, 0) {real, imag} */,
  {32'hc3290769, 32'h42763bdb} /* (3, 28, 31) {real, imag} */,
  {32'h42bd88de, 32'hc29a7d25} /* (3, 28, 30) {real, imag} */,
  {32'h40ee9915, 32'hc2164ecb} /* (3, 28, 29) {real, imag} */,
  {32'hc1eb9e66, 32'h414da3b2} /* (3, 28, 28) {real, imag} */,
  {32'h405c91a7, 32'hc1af52e0} /* (3, 28, 27) {real, imag} */,
  {32'h4142633a, 32'hc1313475} /* (3, 28, 26) {real, imag} */,
  {32'hbfa4c26c, 32'hc1512b39} /* (3, 28, 25) {real, imag} */,
  {32'h40d99c9a, 32'hc15528f3} /* (3, 28, 24) {real, imag} */,
  {32'h41750e6d, 32'h3cc58e00} /* (3, 28, 23) {real, imag} */,
  {32'hbf533949, 32'h410df6e2} /* (3, 28, 22) {real, imag} */,
  {32'hc0675d09, 32'hc085063c} /* (3, 28, 21) {real, imag} */,
  {32'hbfc56ce4, 32'h40189268} /* (3, 28, 20) {real, imag} */,
  {32'h407d4172, 32'hc17852bc} /* (3, 28, 19) {real, imag} */,
  {32'h408a91ea, 32'hc0cb3f46} /* (3, 28, 18) {real, imag} */,
  {32'h3ec74160, 32'hc0309dfa} /* (3, 28, 17) {real, imag} */,
  {32'h409c84eb, 32'h3f5fb802} /* (3, 28, 16) {real, imag} */,
  {32'hc066faed, 32'h406bf3dc} /* (3, 28, 15) {real, imag} */,
  {32'h41896b6d, 32'h410d1e38} /* (3, 28, 14) {real, imag} */,
  {32'hc05b2d97, 32'h41428c36} /* (3, 28, 13) {real, imag} */,
  {32'hc1382a31, 32'hc17951d0} /* (3, 28, 12) {real, imag} */,
  {32'h41ef032a, 32'h401e9408} /* (3, 28, 11) {real, imag} */,
  {32'hc1b79946, 32'h405549cf} /* (3, 28, 10) {real, imag} */,
  {32'hc1a22e48, 32'hc0ab3b33} /* (3, 28, 9) {real, imag} */,
  {32'hc12f5aba, 32'h416e86c6} /* (3, 28, 8) {real, imag} */,
  {32'h4024a93c, 32'h4166029e} /* (3, 28, 7) {real, imag} */,
  {32'hc124f123, 32'h41241377} /* (3, 28, 6) {real, imag} */,
  {32'h41dcb5ec, 32'h405b6954} /* (3, 28, 5) {real, imag} */,
  {32'hc0c8bb24, 32'h418ce2e6} /* (3, 28, 4) {real, imag} */,
  {32'hc17f6766, 32'hc20d0e7c} /* (3, 28, 3) {real, imag} */,
  {32'h41cfcfdd, 32'hc2bc406b} /* (3, 28, 2) {real, imag} */,
  {32'hc23f4fee, 32'h42b59c6e} /* (3, 28, 1) {real, imag} */,
  {32'hc294b735, 32'h419912a0} /* (3, 28, 0) {real, imag} */,
  {32'h42ad387a, 32'hc2a13378} /* (3, 27, 31) {real, imag} */,
  {32'hc13bd2b8, 32'h414e01e2} /* (3, 27, 30) {real, imag} */,
  {32'hc18d44cc, 32'hc1415a4a} /* (3, 27, 29) {real, imag} */,
  {32'h41898b80, 32'hc06afea3} /* (3, 27, 28) {real, imag} */,
  {32'hc16268c2, 32'h41d169f8} /* (3, 27, 27) {real, imag} */,
  {32'hc1c6d7da, 32'h3f114be0} /* (3, 27, 26) {real, imag} */,
  {32'hc06fafa2, 32'h3f136170} /* (3, 27, 25) {real, imag} */,
  {32'hc0a6f0f7, 32'hc1040b32} /* (3, 27, 24) {real, imag} */,
  {32'h41a92b9c, 32'hc0de24e6} /* (3, 27, 23) {real, imag} */,
  {32'h41001ca2, 32'h40badf63} /* (3, 27, 22) {real, imag} */,
  {32'hc0bd1e5c, 32'h41481b5c} /* (3, 27, 21) {real, imag} */,
  {32'hc077577a, 32'hc0462f58} /* (3, 27, 20) {real, imag} */,
  {32'h4086db1a, 32'h41770352} /* (3, 27, 19) {real, imag} */,
  {32'h3f90a7da, 32'h403cb9af} /* (3, 27, 18) {real, imag} */,
  {32'hbff5f7d0, 32'h41a08712} /* (3, 27, 17) {real, imag} */,
  {32'hc13116d6, 32'hc0316ca3} /* (3, 27, 16) {real, imag} */,
  {32'hbf058400, 32'h4037161f} /* (3, 27, 15) {real, imag} */,
  {32'hc15c369e, 32'h40ca5b06} /* (3, 27, 14) {real, imag} */,
  {32'hbe47bff0, 32'hbea62428} /* (3, 27, 13) {real, imag} */,
  {32'h4013a400, 32'hc108234e} /* (3, 27, 12) {real, imag} */,
  {32'hc1bfe3c3, 32'hc0e6d764} /* (3, 27, 11) {real, imag} */,
  {32'hc16b317b, 32'hc10f51a2} /* (3, 27, 10) {real, imag} */,
  {32'hbfbc3498, 32'h400fd190} /* (3, 27, 9) {real, imag} */,
  {32'hc151bd33, 32'hc0387ddf} /* (3, 27, 8) {real, imag} */,
  {32'h4132d7c6, 32'hc12ab2f3} /* (3, 27, 7) {real, imag} */,
  {32'h405b8fba, 32'h40bf3041} /* (3, 27, 6) {real, imag} */,
  {32'hc1d2a943, 32'h3e106940} /* (3, 27, 5) {real, imag} */,
  {32'h414839a4, 32'h41d3533c} /* (3, 27, 4) {real, imag} */,
  {32'hc1901288, 32'h411af5fe} /* (3, 27, 3) {real, imag} */,
  {32'hc218ac70, 32'hc078793c} /* (3, 27, 2) {real, imag} */,
  {32'h42958132, 32'h411695ba} /* (3, 27, 1) {real, imag} */,
  {32'h42a529fb, 32'hc0b47bcc} /* (3, 27, 0) {real, imag} */,
  {32'h41b99064, 32'h416206e8} /* (3, 26, 31) {real, imag} */,
  {32'hc1b9221e, 32'hc14ae763} /* (3, 26, 30) {real, imag} */,
  {32'hc0785086, 32'hc10f9a78} /* (3, 26, 29) {real, imag} */,
  {32'h40c6cade, 32'h40ad7ddf} /* (3, 26, 28) {real, imag} */,
  {32'hc10cb9d0, 32'h4127a7ed} /* (3, 26, 27) {real, imag} */,
  {32'hc18b1ac1, 32'hc1a68040} /* (3, 26, 26) {real, imag} */,
  {32'h3f104cc0, 32'hc14b2459} /* (3, 26, 25) {real, imag} */,
  {32'hc08237e0, 32'h415dae3d} /* (3, 26, 24) {real, imag} */,
  {32'hc0bd4ef4, 32'hc1f60b21} /* (3, 26, 23) {real, imag} */,
  {32'h4106224c, 32'h4166339f} /* (3, 26, 22) {real, imag} */,
  {32'hc0ba49c6, 32'h41725f8d} /* (3, 26, 21) {real, imag} */,
  {32'hc12505c2, 32'h40285200} /* (3, 26, 20) {real, imag} */,
  {32'h40280080, 32'hc0afcbaf} /* (3, 26, 19) {real, imag} */,
  {32'h409d5838, 32'hc1bda12e} /* (3, 26, 18) {real, imag} */,
  {32'h40745eb3, 32'h4102141e} /* (3, 26, 17) {real, imag} */,
  {32'hc077445e, 32'h4152bf78} /* (3, 26, 16) {real, imag} */,
  {32'h409d6b26, 32'h40a50f48} /* (3, 26, 15) {real, imag} */,
  {32'h40cf3657, 32'hc0186a4f} /* (3, 26, 14) {real, imag} */,
  {32'hc0acd20b, 32'hc1c41508} /* (3, 26, 13) {real, imag} */,
  {32'h40e94d1f, 32'hc139d0e8} /* (3, 26, 12) {real, imag} */,
  {32'hc0d46c24, 32'h410d787e} /* (3, 26, 11) {real, imag} */,
  {32'h41455666, 32'hc0b2c313} /* (3, 26, 10) {real, imag} */,
  {32'h4122ae8b, 32'h412a042e} /* (3, 26, 9) {real, imag} */,
  {32'hc01bb2cb, 32'h405a1d24} /* (3, 26, 8) {real, imag} */,
  {32'h40103a40, 32'h418ba4ee} /* (3, 26, 7) {real, imag} */,
  {32'h40d357d8, 32'h3f40b7dc} /* (3, 26, 6) {real, imag} */,
  {32'hc127f426, 32'h407ca9d5} /* (3, 26, 5) {real, imag} */,
  {32'hc15e31f8, 32'h4189fed7} /* (3, 26, 4) {real, imag} */,
  {32'h403755d5, 32'h419f923e} /* (3, 26, 3) {real, imag} */,
  {32'hc0f59d0a, 32'hc080d8a4} /* (3, 26, 2) {real, imag} */,
  {32'h418875dc, 32'hc0d97d12} /* (3, 26, 1) {real, imag} */,
  {32'h40bfa0c0, 32'hc1921be8} /* (3, 26, 0) {real, imag} */,
  {32'hc1c52674, 32'h41a095c4} /* (3, 25, 31) {real, imag} */,
  {32'hc1b39dd0, 32'hc1aef548} /* (3, 25, 30) {real, imag} */,
  {32'h4055ab94, 32'hc0a91b0c} /* (3, 25, 29) {real, imag} */,
  {32'hc15666ca, 32'h415f1892} /* (3, 25, 28) {real, imag} */,
  {32'h410961e6, 32'hc0ee6ddc} /* (3, 25, 27) {real, imag} */,
  {32'h3fadb710, 32'h413eaf2e} /* (3, 25, 26) {real, imag} */,
  {32'h40b9ddc6, 32'hc0d70a64} /* (3, 25, 25) {real, imag} */,
  {32'h418ac668, 32'hc052764f} /* (3, 25, 24) {real, imag} */,
  {32'hc076bb98, 32'hc0f452f5} /* (3, 25, 23) {real, imag} */,
  {32'hc1209473, 32'hc02c2a0b} /* (3, 25, 22) {real, imag} */,
  {32'h40004150, 32'hbe0b8cc0} /* (3, 25, 21) {real, imag} */,
  {32'h409939c2, 32'hc0fbc9f3} /* (3, 25, 20) {real, imag} */,
  {32'hc0105cd0, 32'h3ded7910} /* (3, 25, 19) {real, imag} */,
  {32'h403db9ae, 32'h412ccbce} /* (3, 25, 18) {real, imag} */,
  {32'h40bacb01, 32'hc1799858} /* (3, 25, 17) {real, imag} */,
  {32'h409f9ba1, 32'hc11d8b2c} /* (3, 25, 16) {real, imag} */,
  {32'h408ca606, 32'hc1397b27} /* (3, 25, 15) {real, imag} */,
  {32'h3fec73e0, 32'h410a1bdf} /* (3, 25, 14) {real, imag} */,
  {32'hc1c0079e, 32'h3faadafa} /* (3, 25, 13) {real, imag} */,
  {32'hc03ae56e, 32'h41955723} /* (3, 25, 12) {real, imag} */,
  {32'hc18273e0, 32'h4024f8c4} /* (3, 25, 11) {real, imag} */,
  {32'h4188a7ee, 32'h40488598} /* (3, 25, 10) {real, imag} */,
  {32'hc10fae3d, 32'hc14ca355} /* (3, 25, 9) {real, imag} */,
  {32'hc061e0da, 32'hc13689b2} /* (3, 25, 8) {real, imag} */,
  {32'h4143d47f, 32'h41077fdc} /* (3, 25, 7) {real, imag} */,
  {32'h3e9838b8, 32'h416e68dd} /* (3, 25, 6) {real, imag} */,
  {32'h407f5c90, 32'hc21a7570} /* (3, 25, 5) {real, imag} */,
  {32'h40c45caa, 32'h4158006a} /* (3, 25, 4) {real, imag} */,
  {32'hc136d1c1, 32'hc133ad58} /* (3, 25, 3) {real, imag} */,
  {32'hc1a38152, 32'hc1111ebe} /* (3, 25, 2) {real, imag} */,
  {32'hc0ea2697, 32'hc0b9e3f5} /* (3, 25, 1) {real, imag} */,
  {32'h3f801530, 32'h41c2fbc8} /* (3, 25, 0) {real, imag} */,
  {32'h41d68b2c, 32'hc17f3716} /* (3, 24, 31) {real, imag} */,
  {32'hc0fc8e74, 32'h41669e65} /* (3, 24, 30) {real, imag} */,
  {32'hbeb9f5a0, 32'h40c613e7} /* (3, 24, 29) {real, imag} */,
  {32'hc03e2faa, 32'hc0fb362b} /* (3, 24, 28) {real, imag} */,
  {32'h4185b43c, 32'hc143507d} /* (3, 24, 27) {real, imag} */,
  {32'hc19b7d94, 32'h4164ab5c} /* (3, 24, 26) {real, imag} */,
  {32'hc1ab1071, 32'h4010b513} /* (3, 24, 25) {real, imag} */,
  {32'h407a66d0, 32'h408ae26a} /* (3, 24, 24) {real, imag} */,
  {32'hc1a17df1, 32'h413eaa35} /* (3, 24, 23) {real, imag} */,
  {32'h40c7d849, 32'h40e548f9} /* (3, 24, 22) {real, imag} */,
  {32'h40501dbe, 32'h41a045ca} /* (3, 24, 21) {real, imag} */,
  {32'h4072b496, 32'hc154dd65} /* (3, 24, 20) {real, imag} */,
  {32'h40eda44c, 32'hc144359d} /* (3, 24, 19) {real, imag} */,
  {32'hc1246025, 32'hc12b1fb1} /* (3, 24, 18) {real, imag} */,
  {32'hc0418874, 32'hc1477203} /* (3, 24, 17) {real, imag} */,
  {32'hc0124c6c, 32'h40980376} /* (3, 24, 16) {real, imag} */,
  {32'hc0b30534, 32'hc0aee2ed} /* (3, 24, 15) {real, imag} */,
  {32'h41757653, 32'hbfb84b90} /* (3, 24, 14) {real, imag} */,
  {32'h4138a4a5, 32'h4192a83c} /* (3, 24, 13) {real, imag} */,
  {32'hc19c18fc, 32'hc0b9d0db} /* (3, 24, 12) {real, imag} */,
  {32'hbe9addd0, 32'hc0da8a6c} /* (3, 24, 11) {real, imag} */,
  {32'hc185e9a2, 32'h416119ce} /* (3, 24, 10) {real, imag} */,
  {32'h405dffc0, 32'h3fa3e08a} /* (3, 24, 9) {real, imag} */,
  {32'hc18bd345, 32'hc053873a} /* (3, 24, 8) {real, imag} */,
  {32'hc02835a4, 32'hc1befe2a} /* (3, 24, 7) {real, imag} */,
  {32'h41280922, 32'hc01857fe} /* (3, 24, 6) {real, imag} */,
  {32'h3fe53d38, 32'h413dca90} /* (3, 24, 5) {real, imag} */,
  {32'h4146c75a, 32'hc0fc48c6} /* (3, 24, 4) {real, imag} */,
  {32'hc13d730f, 32'hbfc62678} /* (3, 24, 3) {real, imag} */,
  {32'hc1af06e6, 32'h40eb2454} /* (3, 24, 2) {real, imag} */,
  {32'h420a98e4, 32'hc19fbb66} /* (3, 24, 1) {real, imag} */,
  {32'h41ff2c6b, 32'h3fe0d17c} /* (3, 24, 0) {real, imag} */,
  {32'hc18a2e3a, 32'h413d4c96} /* (3, 23, 31) {real, imag} */,
  {32'hc18768a5, 32'h4185182e} /* (3, 23, 30) {real, imag} */,
  {32'hc0877ff0, 32'h405ec512} /* (3, 23, 29) {real, imag} */,
  {32'h40f902c4, 32'hc052e12c} /* (3, 23, 28) {real, imag} */,
  {32'hc0dd6d98, 32'h4124125c} /* (3, 23, 27) {real, imag} */,
  {32'hc0490815, 32'hc0a5dadb} /* (3, 23, 26) {real, imag} */,
  {32'hc140ffb4, 32'hc10b4001} /* (3, 23, 25) {real, imag} */,
  {32'h409b48cc, 32'h4125f5d1} /* (3, 23, 24) {real, imag} */,
  {32'hc16975fe, 32'hc11809f4} /* (3, 23, 23) {real, imag} */,
  {32'h415f4076, 32'h40b7cd06} /* (3, 23, 22) {real, imag} */,
  {32'hc09ccdee, 32'hc0c62345} /* (3, 23, 21) {real, imag} */,
  {32'h407374ea, 32'h40c2124e} /* (3, 23, 20) {real, imag} */,
  {32'hc155af34, 32'h4172dd10} /* (3, 23, 19) {real, imag} */,
  {32'hc13393e2, 32'hc1022eb7} /* (3, 23, 18) {real, imag} */,
  {32'h403444b7, 32'hc0fb7945} /* (3, 23, 17) {real, imag} */,
  {32'h418696a6, 32'h40504efe} /* (3, 23, 16) {real, imag} */,
  {32'h406bd1ce, 32'h41702bec} /* (3, 23, 15) {real, imag} */,
  {32'hc13bd9a7, 32'h3e1c6780} /* (3, 23, 14) {real, imag} */,
  {32'h412b68ae, 32'h4171a71d} /* (3, 23, 13) {real, imag} */,
  {32'h41399065, 32'h3f7ce810} /* (3, 23, 12) {real, imag} */,
  {32'h41837697, 32'h406f8a92} /* (3, 23, 11) {real, imag} */,
  {32'hc10ff34e, 32'h40f92fe1} /* (3, 23, 10) {real, imag} */,
  {32'hc18533b4, 32'h40e2feb2} /* (3, 23, 9) {real, imag} */,
  {32'h3e4b6a20, 32'hc07e1c7a} /* (3, 23, 8) {real, imag} */,
  {32'hc078b6cf, 32'h4158016a} /* (3, 23, 7) {real, imag} */,
  {32'h416daa92, 32'hbfa03998} /* (3, 23, 6) {real, imag} */,
  {32'hc007aff2, 32'hc1306dee} /* (3, 23, 5) {real, imag} */,
  {32'h414195fe, 32'h41137224} /* (3, 23, 4) {real, imag} */,
  {32'hc04f9f44, 32'h41740dad} /* (3, 23, 3) {real, imag} */,
  {32'h40fe2ed4, 32'hc1e9e4d9} /* (3, 23, 2) {real, imag} */,
  {32'hc0590cb8, 32'h3f1092f0} /* (3, 23, 1) {real, imag} */,
  {32'h3f4bb360, 32'h41276479} /* (3, 23, 0) {real, imag} */,
  {32'hc1a00e12, 32'h416e733d} /* (3, 22, 31) {real, imag} */,
  {32'h40be55c4, 32'hc119704c} /* (3, 22, 30) {real, imag} */,
  {32'h416bea81, 32'hc0b08406} /* (3, 22, 29) {real, imag} */,
  {32'h415a2cd6, 32'h4021855c} /* (3, 22, 28) {real, imag} */,
  {32'h40b1154a, 32'h3dcfb480} /* (3, 22, 27) {real, imag} */,
  {32'hc0b73321, 32'h40a950ee} /* (3, 22, 26) {real, imag} */,
  {32'h3e387920, 32'h40eb6fb7} /* (3, 22, 25) {real, imag} */,
  {32'h3e239060, 32'h403d7c9c} /* (3, 22, 24) {real, imag} */,
  {32'h3f17cc60, 32'hbffca512} /* (3, 22, 23) {real, imag} */,
  {32'hc0dea870, 32'hc10dac7f} /* (3, 22, 22) {real, imag} */,
  {32'hc03a28c2, 32'hc0df49b6} /* (3, 22, 21) {real, imag} */,
  {32'hc1381f01, 32'h3ebaef40} /* (3, 22, 20) {real, imag} */,
  {32'hc0f3d368, 32'h41c1df08} /* (3, 22, 19) {real, imag} */,
  {32'h418268fe, 32'hbfe726d4} /* (3, 22, 18) {real, imag} */,
  {32'h4049b26c, 32'hbf0ceb3c} /* (3, 22, 17) {real, imag} */,
  {32'h3eeb55b0, 32'h404d061e} /* (3, 22, 16) {real, imag} */,
  {32'hbfdfd0fe, 32'h4196e3be} /* (3, 22, 15) {real, imag} */,
  {32'hc15b6ddf, 32'h412f0b16} /* (3, 22, 14) {real, imag} */,
  {32'h411de6d0, 32'hc12f7530} /* (3, 22, 13) {real, imag} */,
  {32'hc1c731b5, 32'hc14d33c6} /* (3, 22, 12) {real, imag} */,
  {32'hc0014bd8, 32'h4114751e} /* (3, 22, 11) {real, imag} */,
  {32'h404f12ca, 32'hc10a3227} /* (3, 22, 10) {real, imag} */,
  {32'h3f2421a8, 32'hc055a9bd} /* (3, 22, 9) {real, imag} */,
  {32'h414889e6, 32'hc0c9cba8} /* (3, 22, 8) {real, imag} */,
  {32'hbf9fbf50, 32'hc09f18fb} /* (3, 22, 7) {real, imag} */,
  {32'h410ce39a, 32'h40a57569} /* (3, 22, 6) {real, imag} */,
  {32'h4090f64a, 32'h40228e2c} /* (3, 22, 5) {real, imag} */,
  {32'hc08f5abd, 32'hc19291a7} /* (3, 22, 4) {real, imag} */,
  {32'h3e774a40, 32'hbe17a280} /* (3, 22, 3) {real, imag} */,
  {32'hc00a837a, 32'hc120931d} /* (3, 22, 2) {real, imag} */,
  {32'h406968bc, 32'h40dc94ea} /* (3, 22, 1) {real, imag} */,
  {32'hbfae8794, 32'h416a89a4} /* (3, 22, 0) {real, imag} */,
  {32'hc0826c8d, 32'hc1917748} /* (3, 21, 31) {real, imag} */,
  {32'hc168f55e, 32'h4084d13a} /* (3, 21, 30) {real, imag} */,
  {32'h3da82cc0, 32'hc0f51122} /* (3, 21, 29) {real, imag} */,
  {32'hc153f8e0, 32'h416016bd} /* (3, 21, 28) {real, imag} */,
  {32'h411b4267, 32'h41924668} /* (3, 21, 27) {real, imag} */,
  {32'hc004b2d8, 32'h3e8ad390} /* (3, 21, 26) {real, imag} */,
  {32'hc07a530d, 32'hc1673cd8} /* (3, 21, 25) {real, imag} */,
  {32'h40f1db52, 32'h3f7b5f10} /* (3, 21, 24) {real, imag} */,
  {32'hc16a7a37, 32'h40b37583} /* (3, 21, 23) {real, imag} */,
  {32'hbf8b2d10, 32'hbef6a790} /* (3, 21, 22) {real, imag} */,
  {32'h410ddda0, 32'hc10c12f2} /* (3, 21, 21) {real, imag} */,
  {32'h40b18217, 32'h411a70ce} /* (3, 21, 20) {real, imag} */,
  {32'h3f93e7f0, 32'hc103ec52} /* (3, 21, 19) {real, imag} */,
  {32'hc04c2d51, 32'h40516b6c} /* (3, 21, 18) {real, imag} */,
  {32'h40ba1630, 32'h40164d2f} /* (3, 21, 17) {real, imag} */,
  {32'hc0b4f2b6, 32'h3f706112} /* (3, 21, 16) {real, imag} */,
  {32'h41abdfb8, 32'hc1205288} /* (3, 21, 15) {real, imag} */,
  {32'hc16c0ee8, 32'hc0740bba} /* (3, 21, 14) {real, imag} */,
  {32'hc0a38bd1, 32'h41a7837d} /* (3, 21, 13) {real, imag} */,
  {32'hbf7c7180, 32'h41acc6a0} /* (3, 21, 12) {real, imag} */,
  {32'h4061972c, 32'hc10a92a0} /* (3, 21, 11) {real, imag} */,
  {32'hc06347e0, 32'hbfbc25a0} /* (3, 21, 10) {real, imag} */,
  {32'hc07967b4, 32'hc08606eb} /* (3, 21, 9) {real, imag} */,
  {32'h4136aafc, 32'h41c2862e} /* (3, 21, 8) {real, imag} */,
  {32'h4124a3a4, 32'hc0c7cd29} /* (3, 21, 7) {real, imag} */,
  {32'h418d698a, 32'hc1777fef} /* (3, 21, 6) {real, imag} */,
  {32'h3fc7ecf0, 32'h40ad23c4} /* (3, 21, 5) {real, imag} */,
  {32'hc124719a, 32'h40c32178} /* (3, 21, 4) {real, imag} */,
  {32'hc1758f6c, 32'hbfd1f008} /* (3, 21, 3) {real, imag} */,
  {32'hc12c15c8, 32'h416d1399} /* (3, 21, 2) {real, imag} */,
  {32'h40dd762a, 32'hc0be8fb5} /* (3, 21, 1) {real, imag} */,
  {32'h41a6dd2d, 32'hc13aa684} /* (3, 21, 0) {real, imag} */,
  {32'h40e72c3d, 32'hc04c8274} /* (3, 20, 31) {real, imag} */,
  {32'h40eb3f40, 32'hc12b2879} /* (3, 20, 30) {real, imag} */,
  {32'hbfedf798, 32'hc083d550} /* (3, 20, 29) {real, imag} */,
  {32'hc0a133c4, 32'hbfe22198} /* (3, 20, 28) {real, imag} */,
  {32'h40c3ed76, 32'h41b2b0c6} /* (3, 20, 27) {real, imag} */,
  {32'h40676a85, 32'hc035bac1} /* (3, 20, 26) {real, imag} */,
  {32'h41c18ee1, 32'hbf343d30} /* (3, 20, 25) {real, imag} */,
  {32'hbc6b5400, 32'h4133360e} /* (3, 20, 24) {real, imag} */,
  {32'h411c4dce, 32'h416e7aa6} /* (3, 20, 23) {real, imag} */,
  {32'hc1100bc9, 32'hc12c7909} /* (3, 20, 22) {real, imag} */,
  {32'h40fe8c02, 32'h411a32da} /* (3, 20, 21) {real, imag} */,
  {32'hc09226d4, 32'hc0409794} /* (3, 20, 20) {real, imag} */,
  {32'h405ab282, 32'h415da2c4} /* (3, 20, 19) {real, imag} */,
  {32'h408eacf4, 32'hc104159c} /* (3, 20, 18) {real, imag} */,
  {32'h40531b00, 32'h4181cc01} /* (3, 20, 17) {real, imag} */,
  {32'h3ebe6c78, 32'hc0ba2447} /* (3, 20, 16) {real, imag} */,
  {32'hc0b12852, 32'h406d8388} /* (3, 20, 15) {real, imag} */,
  {32'h3efa6198, 32'hc0410f46} /* (3, 20, 14) {real, imag} */,
  {32'h3f4c4f93, 32'h41a96897} /* (3, 20, 13) {real, imag} */,
  {32'h40df4d6e, 32'h40f05337} /* (3, 20, 12) {real, imag} */,
  {32'hc0bf8e5c, 32'hbedc39f0} /* (3, 20, 11) {real, imag} */,
  {32'hc1477fd7, 32'h404e40b8} /* (3, 20, 10) {real, imag} */,
  {32'hc0bb21ac, 32'h3fe2d5aa} /* (3, 20, 9) {real, imag} */,
  {32'hc046a1d0, 32'h412cc927} /* (3, 20, 8) {real, imag} */,
  {32'hc0cb1d44, 32'h41a13274} /* (3, 20, 7) {real, imag} */,
  {32'hc1267c12, 32'hc0b69909} /* (3, 20, 6) {real, imag} */,
  {32'hc11420e1, 32'hc1672536} /* (3, 20, 5) {real, imag} */,
  {32'hc13d42d1, 32'hc0835657} /* (3, 20, 4) {real, imag} */,
  {32'h418d5465, 32'h40d909fd} /* (3, 20, 3) {real, imag} */,
  {32'hc124de64, 32'hc09953b4} /* (3, 20, 2) {real, imag} */,
  {32'h41989506, 32'hc0533bcc} /* (3, 20, 1) {real, imag} */,
  {32'hc165ed97, 32'hc0a58766} /* (3, 20, 0) {real, imag} */,
  {32'h40220d60, 32'h407b8b53} /* (3, 19, 31) {real, imag} */,
  {32'hbf50e952, 32'hc046ecd6} /* (3, 19, 30) {real, imag} */,
  {32'h40ca58db, 32'hbf55ed54} /* (3, 19, 29) {real, imag} */,
  {32'h409364ce, 32'h4102ab26} /* (3, 19, 28) {real, imag} */,
  {32'h414cc968, 32'hc11e8ad1} /* (3, 19, 27) {real, imag} */,
  {32'h414d4ec6, 32'h401f9374} /* (3, 19, 26) {real, imag} */,
  {32'h409b7cc4, 32'hc0ae12a2} /* (3, 19, 25) {real, imag} */,
  {32'h3f11b174, 32'h3f513f20} /* (3, 19, 24) {real, imag} */,
  {32'hc179c696, 32'h401f2d5e} /* (3, 19, 23) {real, imag} */,
  {32'h41175b80, 32'hc0a7ad02} /* (3, 19, 22) {real, imag} */,
  {32'hc1029d16, 32'hc11c4ecd} /* (3, 19, 21) {real, imag} */,
  {32'h41a72f9d, 32'hc060c1b2} /* (3, 19, 20) {real, imag} */,
  {32'hc0fff44b, 32'h4085812d} /* (3, 19, 19) {real, imag} */,
  {32'h400a2d0c, 32'h4037e304} /* (3, 19, 18) {real, imag} */,
  {32'hc0a2f203, 32'hc0859f36} /* (3, 19, 17) {real, imag} */,
  {32'hc16c9b28, 32'hc02f9e58} /* (3, 19, 16) {real, imag} */,
  {32'h4103c2ce, 32'h41436130} /* (3, 19, 15) {real, imag} */,
  {32'h3f2e3de8, 32'h41693b55} /* (3, 19, 14) {real, imag} */,
  {32'h41d5f08d, 32'hc15070a7} /* (3, 19, 13) {real, imag} */,
  {32'hc15ef586, 32'hc12b5ada} /* (3, 19, 12) {real, imag} */,
  {32'hc1713456, 32'hc0c16c70} /* (3, 19, 11) {real, imag} */,
  {32'hc02468d6, 32'h41399afa} /* (3, 19, 10) {real, imag} */,
  {32'hbf0b7f00, 32'hc0678680} /* (3, 19, 9) {real, imag} */,
  {32'hc10d8d51, 32'h3f98c112} /* (3, 19, 8) {real, imag} */,
  {32'h415de473, 32'hc06aba22} /* (3, 19, 7) {real, imag} */,
  {32'hc036bb0c, 32'hc19814e9} /* (3, 19, 6) {real, imag} */,
  {32'hc02aa1f5, 32'h400018ef} /* (3, 19, 5) {real, imag} */,
  {32'hc146581c, 32'hc00b62e6} /* (3, 19, 4) {real, imag} */,
  {32'hc0047644, 32'hc04dd59c} /* (3, 19, 3) {real, imag} */,
  {32'h3e935290, 32'hc0ae7bbe} /* (3, 19, 2) {real, imag} */,
  {32'hc155ed5b, 32'h4183d542} /* (3, 19, 1) {real, imag} */,
  {32'hc03d253c, 32'hc0d8081f} /* (3, 19, 0) {real, imag} */,
  {32'h40ace9e7, 32'hbfa9722c} /* (3, 18, 31) {real, imag} */,
  {32'h3f4785b0, 32'h4082e060} /* (3, 18, 30) {real, imag} */,
  {32'h41317464, 32'h408d9fce} /* (3, 18, 29) {real, imag} */,
  {32'h416d7627, 32'hc108927c} /* (3, 18, 28) {real, imag} */,
  {32'h40ecbd49, 32'h414a0f1b} /* (3, 18, 27) {real, imag} */,
  {32'hc0b51a2a, 32'h414a6ea9} /* (3, 18, 26) {real, imag} */,
  {32'hc0e6829c, 32'h4118d21e} /* (3, 18, 25) {real, imag} */,
  {32'h40d82e92, 32'h4128e378} /* (3, 18, 24) {real, imag} */,
  {32'hc1535f4e, 32'h3ee01300} /* (3, 18, 23) {real, imag} */,
  {32'hc1575152, 32'h4159f1fa} /* (3, 18, 22) {real, imag} */,
  {32'h3f510c34, 32'hc0fbad0c} /* (3, 18, 21) {real, imag} */,
  {32'h3f51e0e0, 32'hc008a746} /* (3, 18, 20) {real, imag} */,
  {32'hc024af24, 32'h40228e50} /* (3, 18, 19) {real, imag} */,
  {32'h40f157c9, 32'h3f8b86b6} /* (3, 18, 18) {real, imag} */,
  {32'h416c00a6, 32'hc14c3e6e} /* (3, 18, 17) {real, imag} */,
  {32'h40a47b0c, 32'h4093cb4f} /* (3, 18, 16) {real, imag} */,
  {32'hc107bef5, 32'h4094d477} /* (3, 18, 15) {real, imag} */,
  {32'h40a3a33c, 32'hc1562ba5} /* (3, 18, 14) {real, imag} */,
  {32'h3fc185ae, 32'h409884ea} /* (3, 18, 13) {real, imag} */,
  {32'h41a76336, 32'hc1c77922} /* (3, 18, 12) {real, imag} */,
  {32'h3f901b8f, 32'hc1181124} /* (3, 18, 11) {real, imag} */,
  {32'h3ff6e6ac, 32'h408bfcbe} /* (3, 18, 10) {real, imag} */,
  {32'hc00068a2, 32'hc0608108} /* (3, 18, 9) {real, imag} */,
  {32'h40c7ef51, 32'hc18742ab} /* (3, 18, 8) {real, imag} */,
  {32'hc022908c, 32'hc0344f16} /* (3, 18, 7) {real, imag} */,
  {32'hbff8c904, 32'h3f8ab0b0} /* (3, 18, 6) {real, imag} */,
  {32'hc0778222, 32'h404aad2a} /* (3, 18, 5) {real, imag} */,
  {32'h4174c9a7, 32'hc01d9d0c} /* (3, 18, 4) {real, imag} */,
  {32'h402b9bd0, 32'h40bb6606} /* (3, 18, 3) {real, imag} */,
  {32'hc145518f, 32'h413ca2c9} /* (3, 18, 2) {real, imag} */,
  {32'h415a6b83, 32'hc1237c83} /* (3, 18, 1) {real, imag} */,
  {32'h404b75d9, 32'hc10a9760} /* (3, 18, 0) {real, imag} */,
  {32'hc002bef5, 32'h40349e4c} /* (3, 17, 31) {real, imag} */,
  {32'h3fefadc3, 32'hc134bf0e} /* (3, 17, 30) {real, imag} */,
  {32'hc15137ce, 32'h40e51844} /* (3, 17, 29) {real, imag} */,
  {32'h40d3fe81, 32'h3fee4a48} /* (3, 17, 28) {real, imag} */,
  {32'hc06fb324, 32'hc02eea3c} /* (3, 17, 27) {real, imag} */,
  {32'h40dc1b06, 32'hbfc25ea8} /* (3, 17, 26) {real, imag} */,
  {32'h40e2e9ca, 32'hbe952eb0} /* (3, 17, 25) {real, imag} */,
  {32'h40192db4, 32'h3e9855c0} /* (3, 17, 24) {real, imag} */,
  {32'h412332ea, 32'h3e90d488} /* (3, 17, 23) {real, imag} */,
  {32'hc06f1fb4, 32'h40a1da3c} /* (3, 17, 22) {real, imag} */,
  {32'h40832e79, 32'h40de422c} /* (3, 17, 21) {real, imag} */,
  {32'hc06aae78, 32'hc0b4fc42} /* (3, 17, 20) {real, imag} */,
  {32'h3fd6a0ec, 32'h4163d199} /* (3, 17, 19) {real, imag} */,
  {32'h3fc57dee, 32'hc18fa455} /* (3, 17, 18) {real, imag} */,
  {32'hbeee2838, 32'h3fca274b} /* (3, 17, 17) {real, imag} */,
  {32'hc056c23e, 32'h40b581cf} /* (3, 17, 16) {real, imag} */,
  {32'hc15ece11, 32'hc15b097a} /* (3, 17, 15) {real, imag} */,
  {32'h40e51ebe, 32'h4094fab6} /* (3, 17, 14) {real, imag} */,
  {32'hc036e076, 32'h3e2512b0} /* (3, 17, 13) {real, imag} */,
  {32'hc144edd5, 32'h404d9698} /* (3, 17, 12) {real, imag} */,
  {32'hc01921ea, 32'hc0f531c2} /* (3, 17, 11) {real, imag} */,
  {32'h411ffe01, 32'hbd813ec0} /* (3, 17, 10) {real, imag} */,
  {32'hc13f4e4a, 32'hc0f11b7e} /* (3, 17, 9) {real, imag} */,
  {32'h403e3356, 32'hc15fb927} /* (3, 17, 8) {real, imag} */,
  {32'hc0de7f50, 32'h3ff5ffb2} /* (3, 17, 7) {real, imag} */,
  {32'h401b0ce0, 32'h41656b6a} /* (3, 17, 6) {real, imag} */,
  {32'hbfdc9790, 32'hc0af4da0} /* (3, 17, 5) {real, imag} */,
  {32'h41121fb2, 32'h40b45898} /* (3, 17, 4) {real, imag} */,
  {32'hbf50c874, 32'hc128899a} /* (3, 17, 3) {real, imag} */,
  {32'h4061ce5c, 32'hbfa8500f} /* (3, 17, 2) {real, imag} */,
  {32'h406e6316, 32'h40b30d33} /* (3, 17, 1) {real, imag} */,
  {32'h411d0d19, 32'h3f3b022c} /* (3, 17, 0) {real, imag} */,
  {32'h40e96a10, 32'hbf8e7800} /* (3, 16, 31) {real, imag} */,
  {32'hc05f4384, 32'h413fe7be} /* (3, 16, 30) {real, imag} */,
  {32'hbf3bdfc6, 32'h40ec09b6} /* (3, 16, 29) {real, imag} */,
  {32'h405361a9, 32'hc0601d82} /* (3, 16, 28) {real, imag} */,
  {32'hc0ce3961, 32'h4162aa68} /* (3, 16, 27) {real, imag} */,
  {32'h4090e393, 32'hc1353092} /* (3, 16, 26) {real, imag} */,
  {32'h3f3f0402, 32'h403a76aa} /* (3, 16, 25) {real, imag} */,
  {32'h40466056, 32'h3edad700} /* (3, 16, 24) {real, imag} */,
  {32'h40a5d198, 32'h402fe2c4} /* (3, 16, 23) {real, imag} */,
  {32'hbf2f0f28, 32'hc032d9fc} /* (3, 16, 22) {real, imag} */,
  {32'h410c88d6, 32'h40c6ed7c} /* (3, 16, 21) {real, imag} */,
  {32'h404b9e76, 32'h415a6a7e} /* (3, 16, 20) {real, imag} */,
  {32'hc169f72c, 32'h3fb227dd} /* (3, 16, 19) {real, imag} */,
  {32'hc0e4fda0, 32'h4020cc7e} /* (3, 16, 18) {real, imag} */,
  {32'hc0df95d6, 32'h409c711d} /* (3, 16, 17) {real, imag} */,
  {32'hc06cc3a2, 32'h00000000} /* (3, 16, 16) {real, imag} */,
  {32'hc0df95d6, 32'hc09c711d} /* (3, 16, 15) {real, imag} */,
  {32'hc0e4fda0, 32'hc020cc7e} /* (3, 16, 14) {real, imag} */,
  {32'hc169f72c, 32'hbfb227dd} /* (3, 16, 13) {real, imag} */,
  {32'h404b9e76, 32'hc15a6a7e} /* (3, 16, 12) {real, imag} */,
  {32'h410c88d6, 32'hc0c6ed7c} /* (3, 16, 11) {real, imag} */,
  {32'hbf2f0f28, 32'h4032d9fc} /* (3, 16, 10) {real, imag} */,
  {32'h40a5d198, 32'hc02fe2c4} /* (3, 16, 9) {real, imag} */,
  {32'h40466056, 32'hbedad700} /* (3, 16, 8) {real, imag} */,
  {32'h3f3f0402, 32'hc03a76aa} /* (3, 16, 7) {real, imag} */,
  {32'h4090e393, 32'h41353092} /* (3, 16, 6) {real, imag} */,
  {32'hc0ce3961, 32'hc162aa68} /* (3, 16, 5) {real, imag} */,
  {32'h405361a9, 32'h40601d82} /* (3, 16, 4) {real, imag} */,
  {32'hbf3bdfc6, 32'hc0ec09b6} /* (3, 16, 3) {real, imag} */,
  {32'hc05f4384, 32'hc13fe7be} /* (3, 16, 2) {real, imag} */,
  {32'h40e96a10, 32'h3f8e7800} /* (3, 16, 1) {real, imag} */,
  {32'hc0526ab0, 32'h00000000} /* (3, 16, 0) {real, imag} */,
  {32'h406e6316, 32'hc0b30d33} /* (3, 15, 31) {real, imag} */,
  {32'h4061ce5c, 32'h3fa8500f} /* (3, 15, 30) {real, imag} */,
  {32'hbf50c874, 32'h4128899a} /* (3, 15, 29) {real, imag} */,
  {32'h41121fb2, 32'hc0b45898} /* (3, 15, 28) {real, imag} */,
  {32'hbfdc9790, 32'h40af4da0} /* (3, 15, 27) {real, imag} */,
  {32'h401b0ce0, 32'hc1656b6a} /* (3, 15, 26) {real, imag} */,
  {32'hc0de7f50, 32'hbff5ffb2} /* (3, 15, 25) {real, imag} */,
  {32'h403e3356, 32'h415fb927} /* (3, 15, 24) {real, imag} */,
  {32'hc13f4e4a, 32'h40f11b7e} /* (3, 15, 23) {real, imag} */,
  {32'h411ffe01, 32'h3d813ec0} /* (3, 15, 22) {real, imag} */,
  {32'hc01921ea, 32'h40f531c2} /* (3, 15, 21) {real, imag} */,
  {32'hc144edd5, 32'hc04d9698} /* (3, 15, 20) {real, imag} */,
  {32'hc036e076, 32'hbe2512b0} /* (3, 15, 19) {real, imag} */,
  {32'h40e51ebe, 32'hc094fab6} /* (3, 15, 18) {real, imag} */,
  {32'hc15ece11, 32'h415b097a} /* (3, 15, 17) {real, imag} */,
  {32'hc056c23e, 32'hc0b581cf} /* (3, 15, 16) {real, imag} */,
  {32'hbeee2838, 32'hbfca274b} /* (3, 15, 15) {real, imag} */,
  {32'h3fc57dee, 32'h418fa455} /* (3, 15, 14) {real, imag} */,
  {32'h3fd6a0ec, 32'hc163d199} /* (3, 15, 13) {real, imag} */,
  {32'hc06aae78, 32'h40b4fc42} /* (3, 15, 12) {real, imag} */,
  {32'h40832e79, 32'hc0de422c} /* (3, 15, 11) {real, imag} */,
  {32'hc06f1fb4, 32'hc0a1da3c} /* (3, 15, 10) {real, imag} */,
  {32'h412332ea, 32'hbe90d488} /* (3, 15, 9) {real, imag} */,
  {32'h40192db4, 32'hbe9855c0} /* (3, 15, 8) {real, imag} */,
  {32'h40e2e9ca, 32'h3e952eb0} /* (3, 15, 7) {real, imag} */,
  {32'h40dc1b06, 32'h3fc25ea8} /* (3, 15, 6) {real, imag} */,
  {32'hc06fb324, 32'h402eea3c} /* (3, 15, 5) {real, imag} */,
  {32'h40d3fe81, 32'hbfee4a48} /* (3, 15, 4) {real, imag} */,
  {32'hc15137ce, 32'hc0e51844} /* (3, 15, 3) {real, imag} */,
  {32'h3fefadc3, 32'h4134bf0e} /* (3, 15, 2) {real, imag} */,
  {32'hc002bef5, 32'hc0349e4c} /* (3, 15, 1) {real, imag} */,
  {32'h411d0d19, 32'hbf3b022c} /* (3, 15, 0) {real, imag} */,
  {32'h415a6b83, 32'h41237c83} /* (3, 14, 31) {real, imag} */,
  {32'hc145518f, 32'hc13ca2c9} /* (3, 14, 30) {real, imag} */,
  {32'h402b9bd0, 32'hc0bb6606} /* (3, 14, 29) {real, imag} */,
  {32'h4174c9a7, 32'h401d9d0c} /* (3, 14, 28) {real, imag} */,
  {32'hc0778222, 32'hc04aad2a} /* (3, 14, 27) {real, imag} */,
  {32'hbff8c904, 32'hbf8ab0b0} /* (3, 14, 26) {real, imag} */,
  {32'hc022908c, 32'h40344f16} /* (3, 14, 25) {real, imag} */,
  {32'h40c7ef51, 32'h418742ab} /* (3, 14, 24) {real, imag} */,
  {32'hc00068a2, 32'h40608108} /* (3, 14, 23) {real, imag} */,
  {32'h3ff6e6ac, 32'hc08bfcbe} /* (3, 14, 22) {real, imag} */,
  {32'h3f901b8f, 32'h41181124} /* (3, 14, 21) {real, imag} */,
  {32'h41a76336, 32'h41c77922} /* (3, 14, 20) {real, imag} */,
  {32'h3fc185ae, 32'hc09884ea} /* (3, 14, 19) {real, imag} */,
  {32'h40a3a33c, 32'h41562ba5} /* (3, 14, 18) {real, imag} */,
  {32'hc107bef5, 32'hc094d477} /* (3, 14, 17) {real, imag} */,
  {32'h40a47b0c, 32'hc093cb4f} /* (3, 14, 16) {real, imag} */,
  {32'h416c00a6, 32'h414c3e6e} /* (3, 14, 15) {real, imag} */,
  {32'h40f157c9, 32'hbf8b86b6} /* (3, 14, 14) {real, imag} */,
  {32'hc024af24, 32'hc0228e50} /* (3, 14, 13) {real, imag} */,
  {32'h3f51e0e0, 32'h4008a746} /* (3, 14, 12) {real, imag} */,
  {32'h3f510c34, 32'h40fbad0c} /* (3, 14, 11) {real, imag} */,
  {32'hc1575152, 32'hc159f1fa} /* (3, 14, 10) {real, imag} */,
  {32'hc1535f4e, 32'hbee01300} /* (3, 14, 9) {real, imag} */,
  {32'h40d82e92, 32'hc128e378} /* (3, 14, 8) {real, imag} */,
  {32'hc0e6829c, 32'hc118d21e} /* (3, 14, 7) {real, imag} */,
  {32'hc0b51a2a, 32'hc14a6ea9} /* (3, 14, 6) {real, imag} */,
  {32'h40ecbd49, 32'hc14a0f1b} /* (3, 14, 5) {real, imag} */,
  {32'h416d7627, 32'h4108927c} /* (3, 14, 4) {real, imag} */,
  {32'h41317464, 32'hc08d9fce} /* (3, 14, 3) {real, imag} */,
  {32'h3f4785b0, 32'hc082e060} /* (3, 14, 2) {real, imag} */,
  {32'h40ace9e7, 32'h3fa9722c} /* (3, 14, 1) {real, imag} */,
  {32'h404b75d9, 32'h410a9760} /* (3, 14, 0) {real, imag} */,
  {32'hc155ed5b, 32'hc183d542} /* (3, 13, 31) {real, imag} */,
  {32'h3e935290, 32'h40ae7bbe} /* (3, 13, 30) {real, imag} */,
  {32'hc0047644, 32'h404dd59c} /* (3, 13, 29) {real, imag} */,
  {32'hc146581c, 32'h400b62e6} /* (3, 13, 28) {real, imag} */,
  {32'hc02aa1f5, 32'hc00018ef} /* (3, 13, 27) {real, imag} */,
  {32'hc036bb0c, 32'h419814e9} /* (3, 13, 26) {real, imag} */,
  {32'h415de473, 32'h406aba22} /* (3, 13, 25) {real, imag} */,
  {32'hc10d8d51, 32'hbf98c112} /* (3, 13, 24) {real, imag} */,
  {32'hbf0b7f00, 32'h40678680} /* (3, 13, 23) {real, imag} */,
  {32'hc02468d6, 32'hc1399afa} /* (3, 13, 22) {real, imag} */,
  {32'hc1713456, 32'h40c16c70} /* (3, 13, 21) {real, imag} */,
  {32'hc15ef586, 32'h412b5ada} /* (3, 13, 20) {real, imag} */,
  {32'h41d5f08d, 32'h415070a7} /* (3, 13, 19) {real, imag} */,
  {32'h3f2e3de8, 32'hc1693b55} /* (3, 13, 18) {real, imag} */,
  {32'h4103c2ce, 32'hc1436130} /* (3, 13, 17) {real, imag} */,
  {32'hc16c9b28, 32'h402f9e58} /* (3, 13, 16) {real, imag} */,
  {32'hc0a2f203, 32'h40859f36} /* (3, 13, 15) {real, imag} */,
  {32'h400a2d0c, 32'hc037e304} /* (3, 13, 14) {real, imag} */,
  {32'hc0fff44b, 32'hc085812d} /* (3, 13, 13) {real, imag} */,
  {32'h41a72f9d, 32'h4060c1b2} /* (3, 13, 12) {real, imag} */,
  {32'hc1029d16, 32'h411c4ecd} /* (3, 13, 11) {real, imag} */,
  {32'h41175b80, 32'h40a7ad02} /* (3, 13, 10) {real, imag} */,
  {32'hc179c696, 32'hc01f2d5e} /* (3, 13, 9) {real, imag} */,
  {32'h3f11b174, 32'hbf513f20} /* (3, 13, 8) {real, imag} */,
  {32'h409b7cc4, 32'h40ae12a2} /* (3, 13, 7) {real, imag} */,
  {32'h414d4ec6, 32'hc01f9374} /* (3, 13, 6) {real, imag} */,
  {32'h414cc968, 32'h411e8ad1} /* (3, 13, 5) {real, imag} */,
  {32'h409364ce, 32'hc102ab26} /* (3, 13, 4) {real, imag} */,
  {32'h40ca58db, 32'h3f55ed54} /* (3, 13, 3) {real, imag} */,
  {32'hbf50e952, 32'h4046ecd6} /* (3, 13, 2) {real, imag} */,
  {32'h40220d60, 32'hc07b8b53} /* (3, 13, 1) {real, imag} */,
  {32'hc03d253c, 32'h40d8081f} /* (3, 13, 0) {real, imag} */,
  {32'h41989506, 32'h40533bcc} /* (3, 12, 31) {real, imag} */,
  {32'hc124de64, 32'h409953b4} /* (3, 12, 30) {real, imag} */,
  {32'h418d5465, 32'hc0d909fd} /* (3, 12, 29) {real, imag} */,
  {32'hc13d42d1, 32'h40835657} /* (3, 12, 28) {real, imag} */,
  {32'hc11420e1, 32'h41672536} /* (3, 12, 27) {real, imag} */,
  {32'hc1267c12, 32'h40b69909} /* (3, 12, 26) {real, imag} */,
  {32'hc0cb1d44, 32'hc1a13274} /* (3, 12, 25) {real, imag} */,
  {32'hc046a1d0, 32'hc12cc927} /* (3, 12, 24) {real, imag} */,
  {32'hc0bb21ac, 32'hbfe2d5aa} /* (3, 12, 23) {real, imag} */,
  {32'hc1477fd7, 32'hc04e40b8} /* (3, 12, 22) {real, imag} */,
  {32'hc0bf8e5c, 32'h3edc39f0} /* (3, 12, 21) {real, imag} */,
  {32'h40df4d6e, 32'hc0f05337} /* (3, 12, 20) {real, imag} */,
  {32'h3f4c4f93, 32'hc1a96897} /* (3, 12, 19) {real, imag} */,
  {32'h3efa6198, 32'h40410f46} /* (3, 12, 18) {real, imag} */,
  {32'hc0b12852, 32'hc06d8388} /* (3, 12, 17) {real, imag} */,
  {32'h3ebe6c78, 32'h40ba2447} /* (3, 12, 16) {real, imag} */,
  {32'h40531b00, 32'hc181cc01} /* (3, 12, 15) {real, imag} */,
  {32'h408eacf4, 32'h4104159c} /* (3, 12, 14) {real, imag} */,
  {32'h405ab282, 32'hc15da2c4} /* (3, 12, 13) {real, imag} */,
  {32'hc09226d4, 32'h40409794} /* (3, 12, 12) {real, imag} */,
  {32'h40fe8c02, 32'hc11a32da} /* (3, 12, 11) {real, imag} */,
  {32'hc1100bc9, 32'h412c7909} /* (3, 12, 10) {real, imag} */,
  {32'h411c4dce, 32'hc16e7aa6} /* (3, 12, 9) {real, imag} */,
  {32'hbc6b5400, 32'hc133360e} /* (3, 12, 8) {real, imag} */,
  {32'h41c18ee1, 32'h3f343d30} /* (3, 12, 7) {real, imag} */,
  {32'h40676a85, 32'h4035bac1} /* (3, 12, 6) {real, imag} */,
  {32'h40c3ed76, 32'hc1b2b0c6} /* (3, 12, 5) {real, imag} */,
  {32'hc0a133c4, 32'h3fe22198} /* (3, 12, 4) {real, imag} */,
  {32'hbfedf798, 32'h4083d550} /* (3, 12, 3) {real, imag} */,
  {32'h40eb3f40, 32'h412b2879} /* (3, 12, 2) {real, imag} */,
  {32'h40e72c3d, 32'h404c8274} /* (3, 12, 1) {real, imag} */,
  {32'hc165ed97, 32'h40a58766} /* (3, 12, 0) {real, imag} */,
  {32'h40dd762a, 32'h40be8fb5} /* (3, 11, 31) {real, imag} */,
  {32'hc12c15c8, 32'hc16d1399} /* (3, 11, 30) {real, imag} */,
  {32'hc1758f6c, 32'h3fd1f008} /* (3, 11, 29) {real, imag} */,
  {32'hc124719a, 32'hc0c32178} /* (3, 11, 28) {real, imag} */,
  {32'h3fc7ecf0, 32'hc0ad23c4} /* (3, 11, 27) {real, imag} */,
  {32'h418d698a, 32'h41777fef} /* (3, 11, 26) {real, imag} */,
  {32'h4124a3a4, 32'h40c7cd29} /* (3, 11, 25) {real, imag} */,
  {32'h4136aafc, 32'hc1c2862e} /* (3, 11, 24) {real, imag} */,
  {32'hc07967b4, 32'h408606eb} /* (3, 11, 23) {real, imag} */,
  {32'hc06347e0, 32'h3fbc25a0} /* (3, 11, 22) {real, imag} */,
  {32'h4061972c, 32'h410a92a0} /* (3, 11, 21) {real, imag} */,
  {32'hbf7c7180, 32'hc1acc6a0} /* (3, 11, 20) {real, imag} */,
  {32'hc0a38bd1, 32'hc1a7837d} /* (3, 11, 19) {real, imag} */,
  {32'hc16c0ee8, 32'h40740bba} /* (3, 11, 18) {real, imag} */,
  {32'h41abdfb8, 32'h41205288} /* (3, 11, 17) {real, imag} */,
  {32'hc0b4f2b6, 32'hbf706112} /* (3, 11, 16) {real, imag} */,
  {32'h40ba1630, 32'hc0164d2f} /* (3, 11, 15) {real, imag} */,
  {32'hc04c2d51, 32'hc0516b6c} /* (3, 11, 14) {real, imag} */,
  {32'h3f93e7f0, 32'h4103ec52} /* (3, 11, 13) {real, imag} */,
  {32'h40b18217, 32'hc11a70ce} /* (3, 11, 12) {real, imag} */,
  {32'h410ddda0, 32'h410c12f2} /* (3, 11, 11) {real, imag} */,
  {32'hbf8b2d10, 32'h3ef6a790} /* (3, 11, 10) {real, imag} */,
  {32'hc16a7a37, 32'hc0b37583} /* (3, 11, 9) {real, imag} */,
  {32'h40f1db52, 32'hbf7b5f10} /* (3, 11, 8) {real, imag} */,
  {32'hc07a530d, 32'h41673cd8} /* (3, 11, 7) {real, imag} */,
  {32'hc004b2d8, 32'hbe8ad390} /* (3, 11, 6) {real, imag} */,
  {32'h411b4267, 32'hc1924668} /* (3, 11, 5) {real, imag} */,
  {32'hc153f8e0, 32'hc16016bd} /* (3, 11, 4) {real, imag} */,
  {32'h3da82cc0, 32'h40f51122} /* (3, 11, 3) {real, imag} */,
  {32'hc168f55e, 32'hc084d13a} /* (3, 11, 2) {real, imag} */,
  {32'hc0826c8d, 32'h41917748} /* (3, 11, 1) {real, imag} */,
  {32'h41a6dd2d, 32'h413aa684} /* (3, 11, 0) {real, imag} */,
  {32'h406968bc, 32'hc0dc94ea} /* (3, 10, 31) {real, imag} */,
  {32'hc00a837a, 32'h4120931d} /* (3, 10, 30) {real, imag} */,
  {32'h3e774a40, 32'h3e17a280} /* (3, 10, 29) {real, imag} */,
  {32'hc08f5abd, 32'h419291a7} /* (3, 10, 28) {real, imag} */,
  {32'h4090f64a, 32'hc0228e2c} /* (3, 10, 27) {real, imag} */,
  {32'h410ce39a, 32'hc0a57569} /* (3, 10, 26) {real, imag} */,
  {32'hbf9fbf50, 32'h409f18fb} /* (3, 10, 25) {real, imag} */,
  {32'h414889e6, 32'h40c9cba8} /* (3, 10, 24) {real, imag} */,
  {32'h3f2421a8, 32'h4055a9bd} /* (3, 10, 23) {real, imag} */,
  {32'h404f12ca, 32'h410a3227} /* (3, 10, 22) {real, imag} */,
  {32'hc0014bd8, 32'hc114751e} /* (3, 10, 21) {real, imag} */,
  {32'hc1c731b5, 32'h414d33c6} /* (3, 10, 20) {real, imag} */,
  {32'h411de6d0, 32'h412f7530} /* (3, 10, 19) {real, imag} */,
  {32'hc15b6ddf, 32'hc12f0b16} /* (3, 10, 18) {real, imag} */,
  {32'hbfdfd0fe, 32'hc196e3be} /* (3, 10, 17) {real, imag} */,
  {32'h3eeb55b0, 32'hc04d061e} /* (3, 10, 16) {real, imag} */,
  {32'h4049b26c, 32'h3f0ceb3c} /* (3, 10, 15) {real, imag} */,
  {32'h418268fe, 32'h3fe726d4} /* (3, 10, 14) {real, imag} */,
  {32'hc0f3d368, 32'hc1c1df08} /* (3, 10, 13) {real, imag} */,
  {32'hc1381f01, 32'hbebaef40} /* (3, 10, 12) {real, imag} */,
  {32'hc03a28c2, 32'h40df49b6} /* (3, 10, 11) {real, imag} */,
  {32'hc0dea870, 32'h410dac7f} /* (3, 10, 10) {real, imag} */,
  {32'h3f17cc60, 32'h3ffca512} /* (3, 10, 9) {real, imag} */,
  {32'h3e239060, 32'hc03d7c9c} /* (3, 10, 8) {real, imag} */,
  {32'h3e387920, 32'hc0eb6fb7} /* (3, 10, 7) {real, imag} */,
  {32'hc0b73321, 32'hc0a950ee} /* (3, 10, 6) {real, imag} */,
  {32'h40b1154a, 32'hbdcfb480} /* (3, 10, 5) {real, imag} */,
  {32'h415a2cd6, 32'hc021855c} /* (3, 10, 4) {real, imag} */,
  {32'h416bea81, 32'h40b08406} /* (3, 10, 3) {real, imag} */,
  {32'h40be55c4, 32'h4119704c} /* (3, 10, 2) {real, imag} */,
  {32'hc1a00e12, 32'hc16e733d} /* (3, 10, 1) {real, imag} */,
  {32'hbfae8794, 32'hc16a89a4} /* (3, 10, 0) {real, imag} */,
  {32'hc0590cb8, 32'hbf1092f0} /* (3, 9, 31) {real, imag} */,
  {32'h40fe2ed4, 32'h41e9e4d9} /* (3, 9, 30) {real, imag} */,
  {32'hc04f9f44, 32'hc1740dad} /* (3, 9, 29) {real, imag} */,
  {32'h414195fe, 32'hc1137224} /* (3, 9, 28) {real, imag} */,
  {32'hc007aff2, 32'h41306dee} /* (3, 9, 27) {real, imag} */,
  {32'h416daa92, 32'h3fa03998} /* (3, 9, 26) {real, imag} */,
  {32'hc078b6cf, 32'hc158016a} /* (3, 9, 25) {real, imag} */,
  {32'h3e4b6a20, 32'h407e1c7a} /* (3, 9, 24) {real, imag} */,
  {32'hc18533b4, 32'hc0e2feb2} /* (3, 9, 23) {real, imag} */,
  {32'hc10ff34e, 32'hc0f92fe1} /* (3, 9, 22) {real, imag} */,
  {32'h41837697, 32'hc06f8a92} /* (3, 9, 21) {real, imag} */,
  {32'h41399065, 32'hbf7ce810} /* (3, 9, 20) {real, imag} */,
  {32'h412b68ae, 32'hc171a71d} /* (3, 9, 19) {real, imag} */,
  {32'hc13bd9a7, 32'hbe1c6780} /* (3, 9, 18) {real, imag} */,
  {32'h406bd1ce, 32'hc1702bec} /* (3, 9, 17) {real, imag} */,
  {32'h418696a6, 32'hc0504efe} /* (3, 9, 16) {real, imag} */,
  {32'h403444b7, 32'h40fb7945} /* (3, 9, 15) {real, imag} */,
  {32'hc13393e2, 32'h41022eb7} /* (3, 9, 14) {real, imag} */,
  {32'hc155af34, 32'hc172dd10} /* (3, 9, 13) {real, imag} */,
  {32'h407374ea, 32'hc0c2124e} /* (3, 9, 12) {real, imag} */,
  {32'hc09ccdee, 32'h40c62345} /* (3, 9, 11) {real, imag} */,
  {32'h415f4076, 32'hc0b7cd06} /* (3, 9, 10) {real, imag} */,
  {32'hc16975fe, 32'h411809f4} /* (3, 9, 9) {real, imag} */,
  {32'h409b48cc, 32'hc125f5d1} /* (3, 9, 8) {real, imag} */,
  {32'hc140ffb4, 32'h410b4001} /* (3, 9, 7) {real, imag} */,
  {32'hc0490815, 32'h40a5dadb} /* (3, 9, 6) {real, imag} */,
  {32'hc0dd6d98, 32'hc124125c} /* (3, 9, 5) {real, imag} */,
  {32'h40f902c4, 32'h4052e12c} /* (3, 9, 4) {real, imag} */,
  {32'hc0877ff0, 32'hc05ec512} /* (3, 9, 3) {real, imag} */,
  {32'hc18768a5, 32'hc185182e} /* (3, 9, 2) {real, imag} */,
  {32'hc18a2e3a, 32'hc13d4c96} /* (3, 9, 1) {real, imag} */,
  {32'h3f4bb360, 32'hc1276479} /* (3, 9, 0) {real, imag} */,
  {32'h420a98e4, 32'h419fbb66} /* (3, 8, 31) {real, imag} */,
  {32'hc1af06e6, 32'hc0eb2454} /* (3, 8, 30) {real, imag} */,
  {32'hc13d730f, 32'h3fc62678} /* (3, 8, 29) {real, imag} */,
  {32'h4146c75a, 32'h40fc48c6} /* (3, 8, 28) {real, imag} */,
  {32'h3fe53d38, 32'hc13dca90} /* (3, 8, 27) {real, imag} */,
  {32'h41280922, 32'h401857fe} /* (3, 8, 26) {real, imag} */,
  {32'hc02835a4, 32'h41befe2a} /* (3, 8, 25) {real, imag} */,
  {32'hc18bd345, 32'h4053873a} /* (3, 8, 24) {real, imag} */,
  {32'h405dffc0, 32'hbfa3e08a} /* (3, 8, 23) {real, imag} */,
  {32'hc185e9a2, 32'hc16119ce} /* (3, 8, 22) {real, imag} */,
  {32'hbe9addd0, 32'h40da8a6c} /* (3, 8, 21) {real, imag} */,
  {32'hc19c18fc, 32'h40b9d0db} /* (3, 8, 20) {real, imag} */,
  {32'h4138a4a5, 32'hc192a83c} /* (3, 8, 19) {real, imag} */,
  {32'h41757653, 32'h3fb84b90} /* (3, 8, 18) {real, imag} */,
  {32'hc0b30534, 32'h40aee2ed} /* (3, 8, 17) {real, imag} */,
  {32'hc0124c6c, 32'hc0980376} /* (3, 8, 16) {real, imag} */,
  {32'hc0418874, 32'h41477203} /* (3, 8, 15) {real, imag} */,
  {32'hc1246025, 32'h412b1fb1} /* (3, 8, 14) {real, imag} */,
  {32'h40eda44c, 32'h4144359d} /* (3, 8, 13) {real, imag} */,
  {32'h4072b496, 32'h4154dd65} /* (3, 8, 12) {real, imag} */,
  {32'h40501dbe, 32'hc1a045ca} /* (3, 8, 11) {real, imag} */,
  {32'h40c7d849, 32'hc0e548f9} /* (3, 8, 10) {real, imag} */,
  {32'hc1a17df1, 32'hc13eaa35} /* (3, 8, 9) {real, imag} */,
  {32'h407a66d0, 32'hc08ae26a} /* (3, 8, 8) {real, imag} */,
  {32'hc1ab1071, 32'hc010b513} /* (3, 8, 7) {real, imag} */,
  {32'hc19b7d94, 32'hc164ab5c} /* (3, 8, 6) {real, imag} */,
  {32'h4185b43c, 32'h4143507d} /* (3, 8, 5) {real, imag} */,
  {32'hc03e2faa, 32'h40fb362b} /* (3, 8, 4) {real, imag} */,
  {32'hbeb9f5a0, 32'hc0c613e7} /* (3, 8, 3) {real, imag} */,
  {32'hc0fc8e74, 32'hc1669e65} /* (3, 8, 2) {real, imag} */,
  {32'h41d68b2c, 32'h417f3716} /* (3, 8, 1) {real, imag} */,
  {32'h41ff2c6b, 32'hbfe0d17c} /* (3, 8, 0) {real, imag} */,
  {32'hc0ea2697, 32'h40b9e3f5} /* (3, 7, 31) {real, imag} */,
  {32'hc1a38152, 32'h41111ebe} /* (3, 7, 30) {real, imag} */,
  {32'hc136d1c1, 32'h4133ad58} /* (3, 7, 29) {real, imag} */,
  {32'h40c45caa, 32'hc158006a} /* (3, 7, 28) {real, imag} */,
  {32'h407f5c90, 32'h421a7570} /* (3, 7, 27) {real, imag} */,
  {32'h3e9838b8, 32'hc16e68dd} /* (3, 7, 26) {real, imag} */,
  {32'h4143d47f, 32'hc1077fdc} /* (3, 7, 25) {real, imag} */,
  {32'hc061e0da, 32'h413689b2} /* (3, 7, 24) {real, imag} */,
  {32'hc10fae3d, 32'h414ca355} /* (3, 7, 23) {real, imag} */,
  {32'h4188a7ee, 32'hc0488598} /* (3, 7, 22) {real, imag} */,
  {32'hc18273e0, 32'hc024f8c4} /* (3, 7, 21) {real, imag} */,
  {32'hc03ae56e, 32'hc1955723} /* (3, 7, 20) {real, imag} */,
  {32'hc1c0079e, 32'hbfaadafa} /* (3, 7, 19) {real, imag} */,
  {32'h3fec73e0, 32'hc10a1bdf} /* (3, 7, 18) {real, imag} */,
  {32'h408ca606, 32'h41397b27} /* (3, 7, 17) {real, imag} */,
  {32'h409f9ba1, 32'h411d8b2c} /* (3, 7, 16) {real, imag} */,
  {32'h40bacb01, 32'h41799858} /* (3, 7, 15) {real, imag} */,
  {32'h403db9ae, 32'hc12ccbce} /* (3, 7, 14) {real, imag} */,
  {32'hc0105cd0, 32'hbded7910} /* (3, 7, 13) {real, imag} */,
  {32'h409939c2, 32'h40fbc9f3} /* (3, 7, 12) {real, imag} */,
  {32'h40004150, 32'h3e0b8cc0} /* (3, 7, 11) {real, imag} */,
  {32'hc1209473, 32'h402c2a0b} /* (3, 7, 10) {real, imag} */,
  {32'hc076bb98, 32'h40f452f5} /* (3, 7, 9) {real, imag} */,
  {32'h418ac668, 32'h4052764f} /* (3, 7, 8) {real, imag} */,
  {32'h40b9ddc6, 32'h40d70a64} /* (3, 7, 7) {real, imag} */,
  {32'h3fadb710, 32'hc13eaf2e} /* (3, 7, 6) {real, imag} */,
  {32'h410961e6, 32'h40ee6ddc} /* (3, 7, 5) {real, imag} */,
  {32'hc15666ca, 32'hc15f1892} /* (3, 7, 4) {real, imag} */,
  {32'h4055ab94, 32'h40a91b0c} /* (3, 7, 3) {real, imag} */,
  {32'hc1b39dd0, 32'h41aef548} /* (3, 7, 2) {real, imag} */,
  {32'hc1c52674, 32'hc1a095c4} /* (3, 7, 1) {real, imag} */,
  {32'h3f801530, 32'hc1c2fbc8} /* (3, 7, 0) {real, imag} */,
  {32'h418875dc, 32'h40d97d12} /* (3, 6, 31) {real, imag} */,
  {32'hc0f59d0a, 32'h4080d8a4} /* (3, 6, 30) {real, imag} */,
  {32'h403755d5, 32'hc19f923e} /* (3, 6, 29) {real, imag} */,
  {32'hc15e31f8, 32'hc189fed7} /* (3, 6, 28) {real, imag} */,
  {32'hc127f426, 32'hc07ca9d5} /* (3, 6, 27) {real, imag} */,
  {32'h40d357d8, 32'hbf40b7dc} /* (3, 6, 26) {real, imag} */,
  {32'h40103a40, 32'hc18ba4ee} /* (3, 6, 25) {real, imag} */,
  {32'hc01bb2cb, 32'hc05a1d24} /* (3, 6, 24) {real, imag} */,
  {32'h4122ae8b, 32'hc12a042e} /* (3, 6, 23) {real, imag} */,
  {32'h41455666, 32'h40b2c313} /* (3, 6, 22) {real, imag} */,
  {32'hc0d46c24, 32'hc10d787e} /* (3, 6, 21) {real, imag} */,
  {32'h40e94d1f, 32'h4139d0e8} /* (3, 6, 20) {real, imag} */,
  {32'hc0acd20b, 32'h41c41508} /* (3, 6, 19) {real, imag} */,
  {32'h40cf3657, 32'h40186a4f} /* (3, 6, 18) {real, imag} */,
  {32'h409d6b26, 32'hc0a50f48} /* (3, 6, 17) {real, imag} */,
  {32'hc077445e, 32'hc152bf78} /* (3, 6, 16) {real, imag} */,
  {32'h40745eb3, 32'hc102141e} /* (3, 6, 15) {real, imag} */,
  {32'h409d5838, 32'h41bda12e} /* (3, 6, 14) {real, imag} */,
  {32'h40280080, 32'h40afcbaf} /* (3, 6, 13) {real, imag} */,
  {32'hc12505c2, 32'hc0285200} /* (3, 6, 12) {real, imag} */,
  {32'hc0ba49c6, 32'hc1725f8d} /* (3, 6, 11) {real, imag} */,
  {32'h4106224c, 32'hc166339f} /* (3, 6, 10) {real, imag} */,
  {32'hc0bd4ef4, 32'h41f60b21} /* (3, 6, 9) {real, imag} */,
  {32'hc08237e0, 32'hc15dae3d} /* (3, 6, 8) {real, imag} */,
  {32'h3f104cc0, 32'h414b2459} /* (3, 6, 7) {real, imag} */,
  {32'hc18b1ac1, 32'h41a68040} /* (3, 6, 6) {real, imag} */,
  {32'hc10cb9d0, 32'hc127a7ed} /* (3, 6, 5) {real, imag} */,
  {32'h40c6cade, 32'hc0ad7ddf} /* (3, 6, 4) {real, imag} */,
  {32'hc0785086, 32'h410f9a78} /* (3, 6, 3) {real, imag} */,
  {32'hc1b9221e, 32'h414ae763} /* (3, 6, 2) {real, imag} */,
  {32'h41b99064, 32'hc16206e8} /* (3, 6, 1) {real, imag} */,
  {32'h40bfa0c0, 32'h41921be8} /* (3, 6, 0) {real, imag} */,
  {32'h42958132, 32'hc11695ba} /* (3, 5, 31) {real, imag} */,
  {32'hc218ac70, 32'h4078793c} /* (3, 5, 30) {real, imag} */,
  {32'hc1901288, 32'hc11af5fe} /* (3, 5, 29) {real, imag} */,
  {32'h414839a4, 32'hc1d3533c} /* (3, 5, 28) {real, imag} */,
  {32'hc1d2a943, 32'hbe106940} /* (3, 5, 27) {real, imag} */,
  {32'h405b8fba, 32'hc0bf3041} /* (3, 5, 26) {real, imag} */,
  {32'h4132d7c6, 32'h412ab2f3} /* (3, 5, 25) {real, imag} */,
  {32'hc151bd33, 32'h40387ddf} /* (3, 5, 24) {real, imag} */,
  {32'hbfbc3498, 32'hc00fd190} /* (3, 5, 23) {real, imag} */,
  {32'hc16b317b, 32'h410f51a2} /* (3, 5, 22) {real, imag} */,
  {32'hc1bfe3c3, 32'h40e6d764} /* (3, 5, 21) {real, imag} */,
  {32'h4013a400, 32'h4108234e} /* (3, 5, 20) {real, imag} */,
  {32'hbe47bff0, 32'h3ea62428} /* (3, 5, 19) {real, imag} */,
  {32'hc15c369e, 32'hc0ca5b06} /* (3, 5, 18) {real, imag} */,
  {32'hbf058400, 32'hc037161f} /* (3, 5, 17) {real, imag} */,
  {32'hc13116d6, 32'h40316ca3} /* (3, 5, 16) {real, imag} */,
  {32'hbff5f7d0, 32'hc1a08712} /* (3, 5, 15) {real, imag} */,
  {32'h3f90a7da, 32'hc03cb9af} /* (3, 5, 14) {real, imag} */,
  {32'h4086db1a, 32'hc1770352} /* (3, 5, 13) {real, imag} */,
  {32'hc077577a, 32'h40462f58} /* (3, 5, 12) {real, imag} */,
  {32'hc0bd1e5c, 32'hc1481b5c} /* (3, 5, 11) {real, imag} */,
  {32'h41001ca2, 32'hc0badf63} /* (3, 5, 10) {real, imag} */,
  {32'h41a92b9c, 32'h40de24e6} /* (3, 5, 9) {real, imag} */,
  {32'hc0a6f0f7, 32'h41040b32} /* (3, 5, 8) {real, imag} */,
  {32'hc06fafa2, 32'hbf136170} /* (3, 5, 7) {real, imag} */,
  {32'hc1c6d7da, 32'hbf114be0} /* (3, 5, 6) {real, imag} */,
  {32'hc16268c2, 32'hc1d169f8} /* (3, 5, 5) {real, imag} */,
  {32'h41898b80, 32'h406afea3} /* (3, 5, 4) {real, imag} */,
  {32'hc18d44cc, 32'h41415a4a} /* (3, 5, 3) {real, imag} */,
  {32'hc13bd2b8, 32'hc14e01e2} /* (3, 5, 2) {real, imag} */,
  {32'h42ad387a, 32'h42a13378} /* (3, 5, 1) {real, imag} */,
  {32'h42a529fb, 32'h40b47bcc} /* (3, 5, 0) {real, imag} */,
  {32'hc23f4fee, 32'hc2b59c6e} /* (3, 4, 31) {real, imag} */,
  {32'h41cfcfdd, 32'h42bc406b} /* (3, 4, 30) {real, imag} */,
  {32'hc17f6766, 32'h420d0e7c} /* (3, 4, 29) {real, imag} */,
  {32'hc0c8bb24, 32'hc18ce2e6} /* (3, 4, 28) {real, imag} */,
  {32'h41dcb5ec, 32'hc05b6954} /* (3, 4, 27) {real, imag} */,
  {32'hc124f123, 32'hc1241377} /* (3, 4, 26) {real, imag} */,
  {32'h4024a93c, 32'hc166029e} /* (3, 4, 25) {real, imag} */,
  {32'hc12f5aba, 32'hc16e86c6} /* (3, 4, 24) {real, imag} */,
  {32'hc1a22e48, 32'h40ab3b33} /* (3, 4, 23) {real, imag} */,
  {32'hc1b79946, 32'hc05549cf} /* (3, 4, 22) {real, imag} */,
  {32'h41ef032a, 32'hc01e9408} /* (3, 4, 21) {real, imag} */,
  {32'hc1382a31, 32'h417951d0} /* (3, 4, 20) {real, imag} */,
  {32'hc05b2d97, 32'hc1428c36} /* (3, 4, 19) {real, imag} */,
  {32'h41896b6d, 32'hc10d1e38} /* (3, 4, 18) {real, imag} */,
  {32'hc066faed, 32'hc06bf3dc} /* (3, 4, 17) {real, imag} */,
  {32'h409c84eb, 32'hbf5fb802} /* (3, 4, 16) {real, imag} */,
  {32'h3ec74160, 32'h40309dfa} /* (3, 4, 15) {real, imag} */,
  {32'h408a91ea, 32'h40cb3f46} /* (3, 4, 14) {real, imag} */,
  {32'h407d4172, 32'h417852bc} /* (3, 4, 13) {real, imag} */,
  {32'hbfc56ce4, 32'hc0189268} /* (3, 4, 12) {real, imag} */,
  {32'hc0675d09, 32'h4085063c} /* (3, 4, 11) {real, imag} */,
  {32'hbf533949, 32'hc10df6e2} /* (3, 4, 10) {real, imag} */,
  {32'h41750e6d, 32'hbcc58e00} /* (3, 4, 9) {real, imag} */,
  {32'h40d99c9a, 32'h415528f3} /* (3, 4, 8) {real, imag} */,
  {32'hbfa4c26c, 32'h41512b39} /* (3, 4, 7) {real, imag} */,
  {32'h4142633a, 32'h41313475} /* (3, 4, 6) {real, imag} */,
  {32'h405c91a7, 32'h41af52e0} /* (3, 4, 5) {real, imag} */,
  {32'hc1eb9e66, 32'hc14da3b2} /* (3, 4, 4) {real, imag} */,
  {32'h40ee9915, 32'h42164ecb} /* (3, 4, 3) {real, imag} */,
  {32'h42bd88de, 32'h429a7d25} /* (3, 4, 2) {real, imag} */,
  {32'hc3290769, 32'hc2763bdb} /* (3, 4, 1) {real, imag} */,
  {32'hc294b735, 32'hc19912a0} /* (3, 4, 0) {real, imag} */,
  {32'h430d693c, 32'hc243905a} /* (3, 3, 31) {real, imag} */,
  {32'hc279392a, 32'h423e9b4f} /* (3, 3, 30) {real, imag} */,
  {32'hc0dd3dea, 32'hc1d41960} /* (3, 3, 29) {real, imag} */,
  {32'hc146ea7d, 32'hc11f9c17} /* (3, 3, 28) {real, imag} */,
  {32'h42140c60, 32'hc00b7768} /* (3, 3, 27) {real, imag} */,
  {32'hc03e99dc, 32'h40d98268} /* (3, 3, 26) {real, imag} */,
  {32'hc09dcb9f, 32'h40404326} /* (3, 3, 25) {real, imag} */,
  {32'hc00a957c, 32'h4204ae04} /* (3, 3, 24) {real, imag} */,
  {32'hc16c682b, 32'hc192afbf} /* (3, 3, 23) {real, imag} */,
  {32'h40da1afa, 32'h411d646e} /* (3, 3, 22) {real, imag} */,
  {32'h403f9ba4, 32'hc193fba6} /* (3, 3, 21) {real, imag} */,
  {32'hbf3e50f8, 32'h40ff4ea1} /* (3, 3, 20) {real, imag} */,
  {32'h4119d8fd, 32'h3f500d48} /* (3, 3, 19) {real, imag} */,
  {32'hc0815074, 32'hbfb52572} /* (3, 3, 18) {real, imag} */,
  {32'hc0e490de, 32'h3ff1d8f6} /* (3, 3, 17) {real, imag} */,
  {32'hc0df8e05, 32'hc09e2474} /* (3, 3, 16) {real, imag} */,
  {32'hc0fa3db0, 32'hbf4ef150} /* (3, 3, 15) {real, imag} */,
  {32'h4047d21b, 32'h41b52ec5} /* (3, 3, 14) {real, imag} */,
  {32'hc1a6515f, 32'hbf0dd438} /* (3, 3, 13) {real, imag} */,
  {32'hc08284ce, 32'h40fcf968} /* (3, 3, 12) {real, imag} */,
  {32'hc1b133de, 32'hc1953ff2} /* (3, 3, 11) {real, imag} */,
  {32'hbedf8084, 32'hc10457ae} /* (3, 3, 10) {real, imag} */,
  {32'h41d28e27, 32'h40a75646} /* (3, 3, 9) {real, imag} */,
  {32'hc08270ca, 32'h41789a55} /* (3, 3, 8) {real, imag} */,
  {32'h40fb7fe4, 32'hc1fdbab3} /* (3, 3, 7) {real, imag} */,
  {32'h3f83ae38, 32'hc1f179c1} /* (3, 3, 6) {real, imag} */,
  {32'hc21c85a2, 32'h41bb0683} /* (3, 3, 5) {real, imag} */,
  {32'h422999f5, 32'h408b924e} /* (3, 3, 4) {real, imag} */,
  {32'hc2239ca2, 32'hc2361e24} /* (3, 3, 3) {real, imag} */,
  {32'hc15396bb, 32'h430631b4} /* (3, 3, 2) {real, imag} */,
  {32'hc2d74aea, 32'hc1cdef58} /* (3, 3, 1) {real, imag} */,
  {32'h41af1a47, 32'hc1a46520} /* (3, 3, 0) {real, imag} */,
  {32'h44276ee7, 32'h4246afd1} /* (3, 2, 31) {real, imag} */,
  {32'hc3a7120c, 32'h42bdd0ef} /* (3, 2, 30) {real, imag} */,
  {32'h41c1b4d3, 32'h42349180} /* (3, 2, 29) {real, imag} */,
  {32'h41f495c3, 32'hc285928a} /* (3, 2, 28) {real, imag} */,
  {32'hc246582c, 32'h423746a4} /* (3, 2, 27) {real, imag} */,
  {32'hc189978d, 32'h3f95b70c} /* (3, 2, 26) {real, imag} */,
  {32'h41c076aa, 32'hc1a78db5} /* (3, 2, 25) {real, imag} */,
  {32'hc20256fc, 32'h419dd252} /* (3, 2, 24) {real, imag} */,
  {32'hc1e1a859, 32'hc11e5474} /* (3, 2, 23) {real, imag} */,
  {32'h418021a0, 32'hc19acde5} /* (3, 2, 22) {real, imag} */,
  {32'hc130dc3a, 32'h41eaa619} /* (3, 2, 21) {real, imag} */,
  {32'h400c8370, 32'hc121a997} /* (3, 2, 20) {real, imag} */,
  {32'hbffa1530, 32'h4124b86a} /* (3, 2, 19) {real, imag} */,
  {32'hc0630920, 32'h41870199} /* (3, 2, 18) {real, imag} */,
  {32'h4018a610, 32'h410d610e} /* (3, 2, 17) {real, imag} */,
  {32'h401a680a, 32'hbf951ce0} /* (3, 2, 16) {real, imag} */,
  {32'h419017f2, 32'hc13d9e46} /* (3, 2, 15) {real, imag} */,
  {32'h4019eede, 32'hc1501514} /* (3, 2, 14) {real, imag} */,
  {32'hc06b1114, 32'hc045d86c} /* (3, 2, 13) {real, imag} */,
  {32'h41ae555e, 32'hbfdd6fe0} /* (3, 2, 12) {real, imag} */,
  {32'hc14d68e3, 32'h41540cdc} /* (3, 2, 11) {real, imag} */,
  {32'h417132e3, 32'h3dc7f600} /* (3, 2, 10) {real, imag} */,
  {32'h40db206a, 32'hc1481ca8} /* (3, 2, 9) {real, imag} */,
  {32'hc1ea1dc3, 32'h3f1eed90} /* (3, 2, 8) {real, imag} */,
  {32'h420a966e, 32'hc12a65c0} /* (3, 2, 7) {real, imag} */,
  {32'h412c336c, 32'h3f389968} /* (3, 2, 6) {real, imag} */,
  {32'hc23ca142, 32'hc216aa0b} /* (3, 2, 5) {real, imag} */,
  {32'h42c8385c, 32'hc0db6714} /* (3, 2, 4) {real, imag} */,
  {32'hc2169306, 32'h408134c8} /* (3, 2, 3) {real, imag} */,
  {32'hc38d518a, 32'h430a34a9} /* (3, 2, 2) {real, imag} */,
  {32'h43c3a854, 32'hc1585dc0} /* (3, 2, 1) {real, imag} */,
  {32'h438ead27, 32'h42a03054} /* (3, 2, 0) {real, imag} */,
  {32'hc4110235, 32'h42bfa448} /* (3, 1, 31) {real, imag} */,
  {32'h437b0f50, 32'h422efbf8} /* (3, 1, 30) {real, imag} */,
  {32'h425ce602, 32'hc2227adc} /* (3, 1, 29) {real, imag} */,
  {32'hc2b54e47, 32'hc24cad5a} /* (3, 1, 28) {real, imag} */,
  {32'h42fbad4c, 32'hc0c5e14c} /* (3, 1, 27) {real, imag} */,
  {32'h4215c0bb, 32'hc1480d04} /* (3, 1, 26) {real, imag} */,
  {32'hc1a3b710, 32'h41069f60} /* (3, 1, 25) {real, imag} */,
  {32'h41ab861f, 32'hc1c4082b} /* (3, 1, 24) {real, imag} */,
  {32'hc0f88bdc, 32'hbfe695f0} /* (3, 1, 23) {real, imag} */,
  {32'hc0f5bda2, 32'h40706ba6} /* (3, 1, 22) {real, imag} */,
  {32'h41f3d926, 32'hc1a0416a} /* (3, 1, 21) {real, imag} */,
  {32'hc0184bf1, 32'h408f84c3} /* (3, 1, 20) {real, imag} */,
  {32'h3ffc7ecc, 32'hbffe7eaa} /* (3, 1, 19) {real, imag} */,
  {32'hc0f6c315, 32'hc16605fe} /* (3, 1, 18) {real, imag} */,
  {32'h40f64116, 32'h3feefffc} /* (3, 1, 17) {real, imag} */,
  {32'h411d0f66, 32'h3ed563e0} /* (3, 1, 16) {real, imag} */,
  {32'h4120b3ae, 32'h40b2bac3} /* (3, 1, 15) {real, imag} */,
  {32'hc09c4f4c, 32'h409673d0} /* (3, 1, 14) {real, imag} */,
  {32'hbfec08e1, 32'hc1154215} /* (3, 1, 13) {real, imag} */,
  {32'hc10f4d6d, 32'h402a845d} /* (3, 1, 12) {real, imag} */,
  {32'h41717016, 32'h41a7e156} /* (3, 1, 11) {real, imag} */,
  {32'h4108b990, 32'h414f17c0} /* (3, 1, 10) {real, imag} */,
  {32'hc142dda8, 32'h4074d03e} /* (3, 1, 9) {real, imag} */,
  {32'h415d3728, 32'h422ee7e5} /* (3, 1, 8) {real, imag} */,
  {32'hc0dd5c60, 32'hc18e732e} /* (3, 1, 7) {real, imag} */,
  {32'hc06fcfec, 32'hc0dba976} /* (3, 1, 6) {real, imag} */,
  {32'h427f9bfe, 32'h4276da63} /* (3, 1, 5) {real, imag} */,
  {32'hc203f346, 32'hc1f47e24} /* (3, 1, 4) {real, imag} */,
  {32'h421b1624, 32'hc1bd9cc4} /* (3, 1, 3) {real, imag} */,
  {32'h439a0f1a, 32'h438021d2} /* (3, 1, 2) {real, imag} */,
  {32'hc4444884, 32'hc40832a4} /* (3, 1, 1) {real, imag} */,
  {32'hc3a818e4, 32'h4205d494} /* (3, 1, 0) {real, imag} */,
  {32'hc3a92762, 32'h43747352} /* (3, 0, 31) {real, imag} */,
  {32'h4299d169, 32'hc2a4c5ca} /* (3, 0, 30) {real, imag} */,
  {32'h42b0fd5c, 32'hc1ea1274} /* (3, 0, 29) {real, imag} */,
  {32'h40a47e74, 32'hc2aad320} /* (3, 0, 28) {real, imag} */,
  {32'h4288722f, 32'hc20cffe2} /* (3, 0, 27) {real, imag} */,
  {32'h414b2ff0, 32'h414b0d58} /* (3, 0, 26) {real, imag} */,
  {32'hc0bf1e92, 32'h415f3371} /* (3, 0, 25) {real, imag} */,
  {32'hbff9635e, 32'hc099c28b} /* (3, 0, 24) {real, imag} */,
  {32'h4205765f, 32'h40c00726} /* (3, 0, 23) {real, imag} */,
  {32'hc0310cea, 32'hc094ebd2} /* (3, 0, 22) {real, imag} */,
  {32'hc0d61730, 32'h404d512e} /* (3, 0, 21) {real, imag} */,
  {32'hc09e658d, 32'h408c61b5} /* (3, 0, 20) {real, imag} */,
  {32'hbfe20dfb, 32'hc1ba82a8} /* (3, 0, 19) {real, imag} */,
  {32'h40987b08, 32'h4195e7b8} /* (3, 0, 18) {real, imag} */,
  {32'h3ff2f5fb, 32'hc1385c4e} /* (3, 0, 17) {real, imag} */,
  {32'h3eba3178, 32'h00000000} /* (3, 0, 16) {real, imag} */,
  {32'h3ff2f5fb, 32'h41385c4e} /* (3, 0, 15) {real, imag} */,
  {32'h40987b08, 32'hc195e7b8} /* (3, 0, 14) {real, imag} */,
  {32'hbfe20dfb, 32'h41ba82a8} /* (3, 0, 13) {real, imag} */,
  {32'hc09e658d, 32'hc08c61b5} /* (3, 0, 12) {real, imag} */,
  {32'hc0d61730, 32'hc04d512e} /* (3, 0, 11) {real, imag} */,
  {32'hc0310cea, 32'h4094ebd2} /* (3, 0, 10) {real, imag} */,
  {32'h4205765f, 32'hc0c00726} /* (3, 0, 9) {real, imag} */,
  {32'hbff9635e, 32'h4099c28b} /* (3, 0, 8) {real, imag} */,
  {32'hc0bf1e92, 32'hc15f3371} /* (3, 0, 7) {real, imag} */,
  {32'h414b2ff0, 32'hc14b0d58} /* (3, 0, 6) {real, imag} */,
  {32'h4288722f, 32'h420cffe2} /* (3, 0, 5) {real, imag} */,
  {32'h40a47e74, 32'h42aad320} /* (3, 0, 4) {real, imag} */,
  {32'h42b0fd5c, 32'h41ea1274} /* (3, 0, 3) {real, imag} */,
  {32'h4299d169, 32'h42a4c5ca} /* (3, 0, 2) {real, imag} */,
  {32'hc3a92762, 32'hc3747352} /* (3, 0, 1) {real, imag} */,
  {32'h430d095b, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc46907cd, 32'h4413725e} /* (2, 31, 31) {real, imag} */,
  {32'h43a3d54f, 32'hc388fcd8} /* (2, 31, 30) {real, imag} */,
  {32'h425fb448, 32'h41a572b7} /* (2, 31, 29) {real, imag} */,
  {32'hc1422e86, 32'h41fc6dd4} /* (2, 31, 28) {real, imag} */,
  {32'h42529f59, 32'hc25bb22c} /* (2, 31, 27) {real, imag} */,
  {32'hc004efc0, 32'hbea8db40} /* (2, 31, 26) {real, imag} */,
  {32'hc0d8990b, 32'h41bc837d} /* (2, 31, 25) {real, imag} */,
  {32'h41b34014, 32'hc1e84d50} /* (2, 31, 24) {real, imag} */,
  {32'hc0421ad4, 32'h40526afe} /* (2, 31, 23) {real, imag} */,
  {32'h415a6014, 32'h408ffaf9} /* (2, 31, 22) {real, imag} */,
  {32'h4174ad1b, 32'hc14c2a32} /* (2, 31, 21) {real, imag} */,
  {32'h417b333c, 32'h3fedfbac} /* (2, 31, 20) {real, imag} */,
  {32'hc01c7f60, 32'h4178d327} /* (2, 31, 19) {real, imag} */,
  {32'hbfd2ac05, 32'hc107a08e} /* (2, 31, 18) {real, imag} */,
  {32'h4021b65a, 32'h4097137f} /* (2, 31, 17) {real, imag} */,
  {32'hc1123ff8, 32'hc076a105} /* (2, 31, 16) {real, imag} */,
  {32'hc04c8e17, 32'h414be896} /* (2, 31, 15) {real, imag} */,
  {32'hc0da80d5, 32'h409335a7} /* (2, 31, 14) {real, imag} */,
  {32'hc140ea95, 32'h41228405} /* (2, 31, 13) {real, imag} */,
  {32'hc0656644, 32'hc180bf32} /* (2, 31, 12) {real, imag} */,
  {32'h4218df18, 32'h4172fb38} /* (2, 31, 11) {real, imag} */,
  {32'hc14762d8, 32'hc11302f3} /* (2, 31, 10) {real, imag} */,
  {32'h40c952ea, 32'h409471c9} /* (2, 31, 9) {real, imag} */,
  {32'h41e5e12a, 32'h40c913ce} /* (2, 31, 8) {real, imag} */,
  {32'hc018bdc8, 32'hc0b9249a} /* (2, 31, 7) {real, imag} */,
  {32'h4217b59e, 32'h417a58a0} /* (2, 31, 6) {real, imag} */,
  {32'h4304ef9c, 32'h405fabef} /* (2, 31, 5) {real, imag} */,
  {32'hc2bafd8c, 32'h423203bd} /* (2, 31, 4) {real, imag} */,
  {32'h424721b1, 32'h4222b064} /* (2, 31, 3) {real, imag} */,
  {32'h4376d04c, 32'hc200fcee} /* (2, 31, 2) {real, imag} */,
  {32'hc41f114e, 32'hc2d8475e} /* (2, 31, 1) {real, imag} */,
  {32'hc3ff6ad2, 32'hc26409e0} /* (2, 31, 0) {real, imag} */,
  {32'h43b44612, 32'h40bd3590} /* (2, 30, 31) {real, imag} */,
  {32'hc37f12ef, 32'hc3188f98} /* (2, 30, 30) {real, imag} */,
  {32'hc20ddc1e, 32'h41f3b55d} /* (2, 30, 29) {real, imag} */,
  {32'h42cdc345, 32'hc1d35bdc} /* (2, 30, 28) {real, imag} */,
  {32'hc245dc90, 32'h423a7fcf} /* (2, 30, 27) {real, imag} */,
  {32'hc1a3c7fa, 32'h416df2fa} /* (2, 30, 26) {real, imag} */,
  {32'hbdca1c60, 32'hc0b19e9c} /* (2, 30, 25) {real, imag} */,
  {32'hc1eabcf3, 32'hc1475f89} /* (2, 30, 24) {real, imag} */,
  {32'h400c895c, 32'hc0ba4594} /* (2, 30, 23) {real, imag} */,
  {32'h41e2c600, 32'hc1d51546} /* (2, 30, 22) {real, imag} */,
  {32'hbf7416b0, 32'h411a876e} /* (2, 30, 21) {real, imag} */,
  {32'h40e155bc, 32'hc18125af} /* (2, 30, 20) {real, imag} */,
  {32'h40df7c14, 32'h3eb7d33c} /* (2, 30, 19) {real, imag} */,
  {32'hbf61e188, 32'h416e348c} /* (2, 30, 18) {real, imag} */,
  {32'hc05e694b, 32'h4129fd95} /* (2, 30, 17) {real, imag} */,
  {32'hc01b6993, 32'h413e64ba} /* (2, 30, 16) {real, imag} */,
  {32'h40766859, 32'h41199c0a} /* (2, 30, 15) {real, imag} */,
  {32'hc11f2aeb, 32'hbf887d60} /* (2, 30, 14) {real, imag} */,
  {32'hc0d6a184, 32'hc03b0f18} /* (2, 30, 13) {real, imag} */,
  {32'h40fe08b0, 32'hc06e65f0} /* (2, 30, 12) {real, imag} */,
  {32'hc0c6ffd5, 32'hc1c55133} /* (2, 30, 11) {real, imag} */,
  {32'hc109b59e, 32'h41a3d72c} /* (2, 30, 10) {real, imag} */,
  {32'hc122e60a, 32'h41001244} /* (2, 30, 9) {real, imag} */,
  {32'hc226c5cf, 32'hc1fa9ce7} /* (2, 30, 8) {real, imag} */,
  {32'h40ba5829, 32'h41217e15} /* (2, 30, 7) {real, imag} */,
  {32'h408bec05, 32'h413cc014} /* (2, 30, 6) {real, imag} */,
  {32'hc206e118, 32'hc25cccc6} /* (2, 30, 5) {real, imag} */,
  {32'h424eb7cb, 32'h423cfc89} /* (2, 30, 4) {real, imag} */,
  {32'h424ee380, 32'hc1d3104c} /* (2, 30, 3) {real, imag} */,
  {32'hc3b249c6, 32'hc29af864} /* (2, 30, 2) {real, imag} */,
  {32'h4434eca6, 32'hc28fcaa9} /* (2, 30, 1) {real, imag} */,
  {32'h43a2e7b4, 32'hc2da7243} /* (2, 30, 0) {real, imag} */,
  {32'hc2b82e10, 32'h4207d672} /* (2, 29, 31) {real, imag} */,
  {32'hc18db9a5, 32'hc3161d4e} /* (2, 29, 30) {real, imag} */,
  {32'hc24c7612, 32'h420b7d8f} /* (2, 29, 29) {real, imag} */,
  {32'h41e42d9d, 32'hc147f2b6} /* (2, 29, 28) {real, imag} */,
  {32'hc1dbc29f, 32'hc2152930} /* (2, 29, 27) {real, imag} */,
  {32'hc1b8addb, 32'hc0597af5} /* (2, 29, 26) {real, imag} */,
  {32'h41835836, 32'h41716260} /* (2, 29, 25) {real, imag} */,
  {32'hc023ce2b, 32'hc17aed6a} /* (2, 29, 24) {real, imag} */,
  {32'h4004f7df, 32'h3dd59fc0} /* (2, 29, 23) {real, imag} */,
  {32'h419c9116, 32'hc1480c61} /* (2, 29, 22) {real, imag} */,
  {32'hc034dfe4, 32'h415f0747} /* (2, 29, 21) {real, imag} */,
  {32'h4190bf80, 32'h40abe3f5} /* (2, 29, 20) {real, imag} */,
  {32'h3d119280, 32'hc0e4f9c9} /* (2, 29, 19) {real, imag} */,
  {32'h40fbec9c, 32'hc1a23d2e} /* (2, 29, 18) {real, imag} */,
  {32'h40a5ce7a, 32'h414bbb35} /* (2, 29, 17) {real, imag} */,
  {32'hc0aea740, 32'h40cd155c} /* (2, 29, 16) {real, imag} */,
  {32'h412d34a8, 32'h410ebe38} /* (2, 29, 15) {real, imag} */,
  {32'h4045b7aa, 32'h3f67d948} /* (2, 29, 14) {real, imag} */,
  {32'hbff28ede, 32'hc0e0d55c} /* (2, 29, 13) {real, imag} */,
  {32'hc0ea4bf8, 32'hc191a97e} /* (2, 29, 12) {real, imag} */,
  {32'hbf84c948, 32'h40dd0195} /* (2, 29, 11) {real, imag} */,
  {32'hbf1c84b2, 32'hc0bcbd52} /* (2, 29, 10) {real, imag} */,
  {32'hc1304b02, 32'h4207833b} /* (2, 29, 9) {real, imag} */,
  {32'hc0f16765, 32'hc1baff6c} /* (2, 29, 8) {real, imag} */,
  {32'hc1101cc3, 32'hc0ef7cab} /* (2, 29, 7) {real, imag} */,
  {32'h40c3fa4c, 32'hc15da79e} /* (2, 29, 6) {real, imag} */,
  {32'h403d9806, 32'hc0ec0c68} /* (2, 29, 5) {real, imag} */,
  {32'hc053c17c, 32'h412f335c} /* (2, 29, 4) {real, imag} */,
  {32'hc227278c, 32'h41db0308} /* (2, 29, 3) {real, imag} */,
  {32'hc2973cba, 32'hc28ef77f} /* (2, 29, 2) {real, imag} */,
  {32'h431f3a08, 32'h42b44ce4} /* (2, 29, 1) {real, imag} */,
  {32'h420173f0, 32'h41fa2460} /* (2, 29, 0) {real, imag} */,
  {32'hc3343598, 32'h424adba7} /* (2, 28, 31) {real, imag} */,
  {32'h42cfc2b9, 32'hc2e4f8c0} /* (2, 28, 30) {real, imag} */,
  {32'h3f3979d8, 32'hc18945fd} /* (2, 28, 29) {real, imag} */,
  {32'hbff76008, 32'h407663f8} /* (2, 28, 28) {real, imag} */,
  {32'hc0fd19a4, 32'hc034b3c8} /* (2, 28, 27) {real, imag} */,
  {32'h410d8a5e, 32'hc119e61c} /* (2, 28, 26) {real, imag} */,
  {32'hc19b42ef, 32'hc0ab6100} /* (2, 28, 25) {real, imag} */,
  {32'hc0e594d2, 32'hc19eab97} /* (2, 28, 24) {real, imag} */,
  {32'h410ee724, 32'h407dff68} /* (2, 28, 23) {real, imag} */,
  {32'hc0781cf6, 32'h3f535630} /* (2, 28, 22) {real, imag} */,
  {32'hc0a35982, 32'hc0de1908} /* (2, 28, 21) {real, imag} */,
  {32'h40e6bf48, 32'hc0877e5e} /* (2, 28, 20) {real, imag} */,
  {32'h416a7e04, 32'hc120ecc4} /* (2, 28, 19) {real, imag} */,
  {32'h41432590, 32'hbf63aff8} /* (2, 28, 18) {real, imag} */,
  {32'h409db033, 32'h405db040} /* (2, 28, 17) {real, imag} */,
  {32'h40b5f934, 32'hc08b0111} /* (2, 28, 16) {real, imag} */,
  {32'hc0370de8, 32'h40e665e8} /* (2, 28, 15) {real, imag} */,
  {32'hc1461abe, 32'h41218f56} /* (2, 28, 14) {real, imag} */,
  {32'hc187d80d, 32'h3e7ef6f0} /* (2, 28, 13) {real, imag} */,
  {32'h405d6d09, 32'h412a590e} /* (2, 28, 12) {real, imag} */,
  {32'h41ce5102, 32'h40eda2c0} /* (2, 28, 11) {real, imag} */,
  {32'hc0f42a00, 32'hc1398fe1} /* (2, 28, 10) {real, imag} */,
  {32'hc12cb2fe, 32'h41123672} /* (2, 28, 9) {real, imag} */,
  {32'h40639b4b, 32'h4183ca5a} /* (2, 28, 8) {real, imag} */,
  {32'hc10b6d49, 32'h419ae8d8} /* (2, 28, 7) {real, imag} */,
  {32'h41498ca3, 32'h41a3b74d} /* (2, 28, 6) {real, imag} */,
  {32'h41e21601, 32'hc16a027e} /* (2, 28, 5) {real, imag} */,
  {32'hc1fad8bc, 32'h41d225da} /* (2, 28, 4) {real, imag} */,
  {32'hc162ad07, 32'hc0c40cc0} /* (2, 28, 3) {real, imag} */,
  {32'h41895e18, 32'hc2adbd78} /* (2, 28, 2) {real, imag} */,
  {32'hc2841c49, 32'h428e6902} /* (2, 28, 1) {real, imag} */,
  {32'hc28863b4, 32'h41a68f73} /* (2, 28, 0) {real, imag} */,
  {32'h4291edd5, 32'hc2ca7164} /* (2, 27, 31) {real, imag} */,
  {32'h3fa36350, 32'h4176ef05} /* (2, 27, 30) {real, imag} */,
  {32'hc0330576, 32'h410a9a44} /* (2, 27, 29) {real, imag} */,
  {32'hc0ccd964, 32'h40d1a49e} /* (2, 27, 28) {real, imag} */,
  {32'hc19e7668, 32'h41b2d0ee} /* (2, 27, 27) {real, imag} */,
  {32'h402bcdac, 32'h40c0f16b} /* (2, 27, 26) {real, imag} */,
  {32'hc1e51ffa, 32'hc0fd9fb2} /* (2, 27, 25) {real, imag} */,
  {32'hbf962258, 32'h4116aa06} /* (2, 27, 24) {real, imag} */,
  {32'hc102b1ad, 32'hc11ed95f} /* (2, 27, 23) {real, imag} */,
  {32'h40caf08c, 32'h3fd80a00} /* (2, 27, 22) {real, imag} */,
  {32'hc0527d98, 32'hc098d8da} /* (2, 27, 21) {real, imag} */,
  {32'hc0472d94, 32'h404ae2e4} /* (2, 27, 20) {real, imag} */,
  {32'h410012bd, 32'hc1348675} /* (2, 27, 19) {real, imag} */,
  {32'hbf5f6284, 32'h41353fc7} /* (2, 27, 18) {real, imag} */,
  {32'hc1086afb, 32'hc0c7f49f} /* (2, 27, 17) {real, imag} */,
  {32'h4111e5e0, 32'h40d6248c} /* (2, 27, 16) {real, imag} */,
  {32'hc051213a, 32'hc0811b00} /* (2, 27, 15) {real, imag} */,
  {32'hc18e74c7, 32'hc0630a50} /* (2, 27, 14) {real, imag} */,
  {32'h402e8e9a, 32'hbecb9d50} /* (2, 27, 13) {real, imag} */,
  {32'hc0fc73f5, 32'h3ff3d980} /* (2, 27, 12) {real, imag} */,
  {32'hc0f4f15c, 32'hc0f24d09} /* (2, 27, 11) {real, imag} */,
  {32'hc0c7007e, 32'h40792480} /* (2, 27, 10) {real, imag} */,
  {32'hc0f8e73d, 32'hc145bba7} /* (2, 27, 9) {real, imag} */,
  {32'h3fc4bdd4, 32'hc1d24eee} /* (2, 27, 8) {real, imag} */,
  {32'hc0aa7ce8, 32'hc0150796} /* (2, 27, 7) {real, imag} */,
  {32'h412ddb16, 32'h41789de1} /* (2, 27, 6) {real, imag} */,
  {32'hc1f852a9, 32'hc0872b6d} /* (2, 27, 5) {real, imag} */,
  {32'h41135a02, 32'h4132de17} /* (2, 27, 4) {real, imag} */,
  {32'hc09d0e2e, 32'hc1435bb5} /* (2, 27, 3) {real, imag} */,
  {32'hc24d1080, 32'h41bcd08a} /* (2, 27, 2) {real, imag} */,
  {32'h42c374f4, 32'hc0e2deb0} /* (2, 27, 1) {real, imag} */,
  {32'h42b1a711, 32'hc1b409b8} /* (2, 27, 0) {real, imag} */,
  {32'h40de2112, 32'h413a4cd4} /* (2, 26, 31) {real, imag} */,
  {32'hc0f4f1c0, 32'h41bae389} /* (2, 26, 30) {real, imag} */,
  {32'hba404000, 32'h3fa8bd04} /* (2, 26, 29) {real, imag} */,
  {32'h40a6ed69, 32'h4088ef7d} /* (2, 26, 28) {real, imag} */,
  {32'h405ca074, 32'h3ed403c0} /* (2, 26, 27) {real, imag} */,
  {32'hc10756ac, 32'hc0993721} /* (2, 26, 26) {real, imag} */,
  {32'hc09e0792, 32'hc1842dd0} /* (2, 26, 25) {real, imag} */,
  {32'hc10830ee, 32'h40b92f8c} /* (2, 26, 24) {real, imag} */,
  {32'hbe04da00, 32'hc1aa2bf2} /* (2, 26, 23) {real, imag} */,
  {32'h419efe4b, 32'h402df6e0} /* (2, 26, 22) {real, imag} */,
  {32'h4149d4e2, 32'h409715d6} /* (2, 26, 21) {real, imag} */,
  {32'hc1867ea1, 32'h415555f3} /* (2, 26, 20) {real, imag} */,
  {32'hc1074c1c, 32'hc0fd7acb} /* (2, 26, 19) {real, imag} */,
  {32'hbff8361a, 32'h413d399a} /* (2, 26, 18) {real, imag} */,
  {32'h3fd5a3c0, 32'h4040acfd} /* (2, 26, 17) {real, imag} */,
  {32'h3ea766e0, 32'h411d811d} /* (2, 26, 16) {real, imag} */,
  {32'hc0edd045, 32'hc04a342e} /* (2, 26, 15) {real, imag} */,
  {32'hc07b883a, 32'h411c2f56} /* (2, 26, 14) {real, imag} */,
  {32'h40f5d092, 32'hbbd5fc00} /* (2, 26, 13) {real, imag} */,
  {32'h411db68c, 32'hc12b7e73} /* (2, 26, 12) {real, imag} */,
  {32'hbfba5e68, 32'hc0a0e058} /* (2, 26, 11) {real, imag} */,
  {32'h416c288f, 32'h4134ecea} /* (2, 26, 10) {real, imag} */,
  {32'hc14a77ae, 32'hc086a392} /* (2, 26, 9) {real, imag} */,
  {32'hc0b83389, 32'hc19d6487} /* (2, 26, 8) {real, imag} */,
  {32'hc11718a6, 32'h404fb7dc} /* (2, 26, 7) {real, imag} */,
  {32'h40a3e206, 32'h4118681d} /* (2, 26, 6) {real, imag} */,
  {32'h3fcf3b7e, 32'h41e48fdc} /* (2, 26, 5) {real, imag} */,
  {32'hc1c4d0d5, 32'h41c0d341} /* (2, 26, 4) {real, imag} */,
  {32'h412a4c3a, 32'hc112bf4c} /* (2, 26, 3) {real, imag} */,
  {32'hbf946e00, 32'h40fda365} /* (2, 26, 2) {real, imag} */,
  {32'hc1215b1a, 32'hc18164d5} /* (2, 26, 1) {real, imag} */,
  {32'h4187d9f9, 32'hc11d8f51} /* (2, 26, 0) {real, imag} */,
  {32'hc1825b20, 32'h41325113} /* (2, 25, 31) {real, imag} */,
  {32'hc1420da0, 32'hc16273dc} /* (2, 25, 30) {real, imag} */,
  {32'h41540ffa, 32'hc05f7ff5} /* (2, 25, 29) {real, imag} */,
  {32'hc0eaa11a, 32'h416703ce} /* (2, 25, 28) {real, imag} */,
  {32'hbeb8ad50, 32'hc16d54a2} /* (2, 25, 27) {real, imag} */,
  {32'hc0c600fe, 32'h40a677f6} /* (2, 25, 26) {real, imag} */,
  {32'h40acf734, 32'hc059a068} /* (2, 25, 25) {real, imag} */,
  {32'hc092352e, 32'h4123e63d} /* (2, 25, 24) {real, imag} */,
  {32'h4136064f, 32'hc16f7157} /* (2, 25, 23) {real, imag} */,
  {32'h4144f5cb, 32'hc1d67524} /* (2, 25, 22) {real, imag} */,
  {32'hc15772f4, 32'h4110dfd7} /* (2, 25, 21) {real, imag} */,
  {32'h3fdd95f0, 32'h402bb37a} /* (2, 25, 20) {real, imag} */,
  {32'h40653529, 32'hc105883c} /* (2, 25, 19) {real, imag} */,
  {32'hc166df53, 32'h41591c12} /* (2, 25, 18) {real, imag} */,
  {32'h41419d14, 32'h3fd35672} /* (2, 25, 17) {real, imag} */,
  {32'hc0b7e982, 32'hc08d246c} /* (2, 25, 16) {real, imag} */,
  {32'h40f06de8, 32'h40e9b89e} /* (2, 25, 15) {real, imag} */,
  {32'hc1351c5b, 32'hc02e3b68} /* (2, 25, 14) {real, imag} */,
  {32'h41515753, 32'h40b4edfa} /* (2, 25, 13) {real, imag} */,
  {32'h3f57bca0, 32'h4042dc70} /* (2, 25, 12) {real, imag} */,
  {32'h40df7bbe, 32'hc0b37c92} /* (2, 25, 11) {real, imag} */,
  {32'hc17d8217, 32'hc13aff4a} /* (2, 25, 10) {real, imag} */,
  {32'hc1bc1c48, 32'hc0e2cba6} /* (2, 25, 9) {real, imag} */,
  {32'h401ac684, 32'hbfc4d5a2} /* (2, 25, 8) {real, imag} */,
  {32'hc1643679, 32'hc1b07d50} /* (2, 25, 7) {real, imag} */,
  {32'hbfbaaf78, 32'hc10a8f43} /* (2, 25, 6) {real, imag} */,
  {32'h3f8119c0, 32'hc1595507} /* (2, 25, 5) {real, imag} */,
  {32'hc181c744, 32'hc0442776} /* (2, 25, 4) {real, imag} */,
  {32'hc1acc2b0, 32'h4145907c} /* (2, 25, 3) {real, imag} */,
  {32'hbfa69134, 32'h40ea0951} /* (2, 25, 2) {real, imag} */,
  {32'hc0c26dd5, 32'hc04963f4} /* (2, 25, 1) {real, imag} */,
  {32'h3f96af50, 32'h41553c41} /* (2, 25, 0) {real, imag} */,
  {32'h416902b0, 32'hc1f50973} /* (2, 24, 31) {real, imag} */,
  {32'h40a734a7, 32'h41c54375} /* (2, 24, 30) {real, imag} */,
  {32'hc04dde4a, 32'h3f52aa68} /* (2, 24, 29) {real, imag} */,
  {32'h400c1e7c, 32'hc00461c4} /* (2, 24, 28) {real, imag} */,
  {32'h400b8650, 32'h405ba5de} /* (2, 24, 27) {real, imag} */,
  {32'hc13af802, 32'h41f0b3d3} /* (2, 24, 26) {real, imag} */,
  {32'hc1a9fc84, 32'h41541de4} /* (2, 24, 25) {real, imag} */,
  {32'hc0698978, 32'h3e118130} /* (2, 24, 24) {real, imag} */,
  {32'hc16676e3, 32'hc1c07b0d} /* (2, 24, 23) {real, imag} */,
  {32'hbec7f550, 32'hc12a5696} /* (2, 24, 22) {real, imag} */,
  {32'hc1127c2a, 32'h41c461f6} /* (2, 24, 21) {real, imag} */,
  {32'h4192fbcb, 32'h403da9a6} /* (2, 24, 20) {real, imag} */,
  {32'hc0a4a334, 32'h41360167} /* (2, 24, 19) {real, imag} */,
  {32'hbfd336d8, 32'h411dd96e} /* (2, 24, 18) {real, imag} */,
  {32'h4091d26a, 32'hc15b532d} /* (2, 24, 17) {real, imag} */,
  {32'h40149860, 32'hc18a1288} /* (2, 24, 16) {real, imag} */,
  {32'h40c68b38, 32'h40c97ef6} /* (2, 24, 15) {real, imag} */,
  {32'h3de3d300, 32'h40a7d313} /* (2, 24, 14) {real, imag} */,
  {32'hc019d4fa, 32'hc19023ba} /* (2, 24, 13) {real, imag} */,
  {32'h4133342d, 32'h40e8bfe0} /* (2, 24, 12) {real, imag} */,
  {32'h4082e90b, 32'h41533d32} /* (2, 24, 11) {real, imag} */,
  {32'hc00cda56, 32'h41ea78f4} /* (2, 24, 10) {real, imag} */,
  {32'h41bf32c0, 32'hc0fbc8dc} /* (2, 24, 9) {real, imag} */,
  {32'h40901ce9, 32'hc1a225b7} /* (2, 24, 8) {real, imag} */,
  {32'h418faff6, 32'hc1cdd8e2} /* (2, 24, 7) {real, imag} */,
  {32'h413d1d6f, 32'hc16f7384} /* (2, 24, 6) {real, imag} */,
  {32'hbf86ab10, 32'h409bc73a} /* (2, 24, 5) {real, imag} */,
  {32'h3fbb2d59, 32'hc1c9c9f2} /* (2, 24, 4) {real, imag} */,
  {32'hc19fb35e, 32'h418e88a5} /* (2, 24, 3) {real, imag} */,
  {32'hc20cfa02, 32'hc1e694d0} /* (2, 24, 2) {real, imag} */,
  {32'h423fe59d, 32'hc19a4594} /* (2, 24, 1) {real, imag} */,
  {32'h40faa4c2, 32'hc00992f0} /* (2, 24, 0) {real, imag} */,
  {32'hc19094c7, 32'h41de04b6} /* (2, 23, 31) {real, imag} */,
  {32'h4092d7fa, 32'h4147a555} /* (2, 23, 30) {real, imag} */,
  {32'hc1bba9c5, 32'hc17c9595} /* (2, 23, 29) {real, imag} */,
  {32'hc12039f0, 32'h41557300} /* (2, 23, 28) {real, imag} */,
  {32'hc122f81e, 32'h41ae8e61} /* (2, 23, 27) {real, imag} */,
  {32'hc01f40ed, 32'hc1b7eaa1} /* (2, 23, 26) {real, imag} */,
  {32'hbfaaa3ec, 32'h40b2d79c} /* (2, 23, 25) {real, imag} */,
  {32'hc14d9aeb, 32'h3f83aaf6} /* (2, 23, 24) {real, imag} */,
  {32'h41326b84, 32'hc0a4bb01} /* (2, 23, 23) {real, imag} */,
  {32'hc1187cda, 32'h3f501440} /* (2, 23, 22) {real, imag} */,
  {32'hc0aa84de, 32'hc1860715} /* (2, 23, 21) {real, imag} */,
  {32'hc1abb034, 32'hc10a4675} /* (2, 23, 20) {real, imag} */,
  {32'h412baef6, 32'h40307e73} /* (2, 23, 19) {real, imag} */,
  {32'hc1547af4, 32'hc1299f77} /* (2, 23, 18) {real, imag} */,
  {32'hc155590c, 32'hc13e7896} /* (2, 23, 17) {real, imag} */,
  {32'h40a3887c, 32'hc114810c} /* (2, 23, 16) {real, imag} */,
  {32'hc10a31cd, 32'h40dac8f3} /* (2, 23, 15) {real, imag} */,
  {32'h41d158db, 32'h4002c7c2} /* (2, 23, 14) {real, imag} */,
  {32'hc1181f7c, 32'hc07661ab} /* (2, 23, 13) {real, imag} */,
  {32'hc18f57a3, 32'h40ae70ea} /* (2, 23, 12) {real, imag} */,
  {32'hc0de5bd8, 32'hc189042c} /* (2, 23, 11) {real, imag} */,
  {32'h3fbe1a2a, 32'hbf7b5d38} /* (2, 23, 10) {real, imag} */,
  {32'h400433e4, 32'h400d001e} /* (2, 23, 9) {real, imag} */,
  {32'hc143e457, 32'hc045fdf8} /* (2, 23, 8) {real, imag} */,
  {32'hc05afe68, 32'h3fc38a10} /* (2, 23, 7) {real, imag} */,
  {32'h4120bcd6, 32'h4005d455} /* (2, 23, 6) {real, imag} */,
  {32'h419f648f, 32'hc11d3858} /* (2, 23, 5) {real, imag} */,
  {32'h40aedf54, 32'hc03ee195} /* (2, 23, 4) {real, imag} */,
  {32'hbf087320, 32'h40fe949e} /* (2, 23, 3) {real, imag} */,
  {32'h415e5689, 32'hc1d5a3cb} /* (2, 23, 2) {real, imag} */,
  {32'h41618f6c, 32'hc0a36b1b} /* (2, 23, 1) {real, imag} */,
  {32'hc15ba0ba, 32'h418a62da} /* (2, 23, 0) {real, imag} */,
  {32'hc1a35a44, 32'h413e38d8} /* (2, 22, 31) {real, imag} */,
  {32'hc16a6a0a, 32'hc198ed13} /* (2, 22, 30) {real, imag} */,
  {32'h41d1fe31, 32'hc01f0d0e} /* (2, 22, 29) {real, imag} */,
  {32'h3ef972a8, 32'hc120fe8f} /* (2, 22, 28) {real, imag} */,
  {32'h3e1514e0, 32'hc151916e} /* (2, 22, 27) {real, imag} */,
  {32'h4174b908, 32'h40c3f601} /* (2, 22, 26) {real, imag} */,
  {32'h4124ffbc, 32'hc0153900} /* (2, 22, 25) {real, imag} */,
  {32'hc15a52f2, 32'hc0a761d4} /* (2, 22, 24) {real, imag} */,
  {32'h40fd4cbf, 32'hc18818b2} /* (2, 22, 23) {real, imag} */,
  {32'h418e1da1, 32'hc060f4ee} /* (2, 22, 22) {real, imag} */,
  {32'hc0e962f4, 32'h4196297a} /* (2, 22, 21) {real, imag} */,
  {32'hc1548b1e, 32'h402e6715} /* (2, 22, 20) {real, imag} */,
  {32'h4080f4e8, 32'h41894c5c} /* (2, 22, 19) {real, imag} */,
  {32'h405b1868, 32'h3fe40ea8} /* (2, 22, 18) {real, imag} */,
  {32'h3ebd2228, 32'h40dd7372} /* (2, 22, 17) {real, imag} */,
  {32'h4115e3f7, 32'hc0bb5cc8} /* (2, 22, 16) {real, imag} */,
  {32'hc143f2f8, 32'h3ececd68} /* (2, 22, 15) {real, imag} */,
  {32'h4072225e, 32'hc13d9596} /* (2, 22, 14) {real, imag} */,
  {32'h412e2f0a, 32'h41a7b408} /* (2, 22, 13) {real, imag} */,
  {32'hc054028c, 32'hc0747258} /* (2, 22, 12) {real, imag} */,
  {32'hc02d610c, 32'h41a5b692} /* (2, 22, 11) {real, imag} */,
  {32'hc16ca7f2, 32'h3efcc3e0} /* (2, 22, 10) {real, imag} */,
  {32'hc0b6b027, 32'h411d074b} /* (2, 22, 9) {real, imag} */,
  {32'hc16505a2, 32'h40b7af91} /* (2, 22, 8) {real, imag} */,
  {32'hc0aab2c3, 32'h408dad3a} /* (2, 22, 7) {real, imag} */,
  {32'h40eaf2d5, 32'h40bbca7f} /* (2, 22, 6) {real, imag} */,
  {32'h408272f6, 32'h3fac3246} /* (2, 22, 5) {real, imag} */,
  {32'hc1a1e576, 32'h402b89c0} /* (2, 22, 4) {real, imag} */,
  {32'hc1967067, 32'hc0ed43c3} /* (2, 22, 3) {real, imag} */,
  {32'h4134688d, 32'hc1c52bea} /* (2, 22, 2) {real, imag} */,
  {32'h3fe40ef4, 32'h40940576} /* (2, 22, 1) {real, imag} */,
  {32'h417ee158, 32'h41228b36} /* (2, 22, 0) {real, imag} */,
  {32'h41150630, 32'hc1a42e12} /* (2, 21, 31) {real, imag} */,
  {32'hbf4124f0, 32'h418fba86} /* (2, 21, 30) {real, imag} */,
  {32'h401c9bb6, 32'hc15340b8} /* (2, 21, 29) {real, imag} */,
  {32'h40fe8260, 32'h41151a90} /* (2, 21, 28) {real, imag} */,
  {32'h41238fa2, 32'hbfbccc18} /* (2, 21, 27) {real, imag} */,
  {32'hbeb6be80, 32'h3f0b53d0} /* (2, 21, 26) {real, imag} */,
  {32'hc0b9bb5b, 32'h3f5d1108} /* (2, 21, 25) {real, imag} */,
  {32'h417a817c, 32'h4180c014} /* (2, 21, 24) {real, imag} */,
  {32'h412a1890, 32'h40d6139b} /* (2, 21, 23) {real, imag} */,
  {32'h3ff0c590, 32'h40758f2a} /* (2, 21, 22) {real, imag} */,
  {32'h40c3509c, 32'h4122aa90} /* (2, 21, 21) {real, imag} */,
  {32'h401f56b1, 32'h3fb609f4} /* (2, 21, 20) {real, imag} */,
  {32'hc11a8fa0, 32'h4042fc27} /* (2, 21, 19) {real, imag} */,
  {32'h40d7970c, 32'hc0df68fe} /* (2, 21, 18) {real, imag} */,
  {32'hbfeab7b8, 32'hc076ca36} /* (2, 21, 17) {real, imag} */,
  {32'hbfdb6788, 32'hc1319e82} /* (2, 21, 16) {real, imag} */,
  {32'hc08f21e6, 32'h407487d9} /* (2, 21, 15) {real, imag} */,
  {32'h41193444, 32'h3fc771e8} /* (2, 21, 14) {real, imag} */,
  {32'h3cc29e00, 32'hc0da7cd4} /* (2, 21, 13) {real, imag} */,
  {32'h40bb2d34, 32'hbf5bb608} /* (2, 21, 12) {real, imag} */,
  {32'hc0ae3806, 32'hc15eedac} /* (2, 21, 11) {real, imag} */,
  {32'h416d52aa, 32'hbf16f6d4} /* (2, 21, 10) {real, imag} */,
  {32'hc01560a0, 32'hc125ad45} /* (2, 21, 9) {real, imag} */,
  {32'h41247580, 32'h40619368} /* (2, 21, 8) {real, imag} */,
  {32'hc0efdc5e, 32'h40879e98} /* (2, 21, 7) {real, imag} */,
  {32'h3ff498f4, 32'hc110fb77} /* (2, 21, 6) {real, imag} */,
  {32'h411dc6fe, 32'hc0b8c42c} /* (2, 21, 5) {real, imag} */,
  {32'hc0edcd6c, 32'hbf4849c8} /* (2, 21, 4) {real, imag} */,
  {32'hc02e3c38, 32'h41220466} /* (2, 21, 3) {real, imag} */,
  {32'hc1ab3811, 32'hc0819c74} /* (2, 21, 2) {real, imag} */,
  {32'h4196ef36, 32'hc2122388} /* (2, 21, 1) {real, imag} */,
  {32'h413469dc, 32'hc1293396} /* (2, 21, 0) {real, imag} */,
  {32'hc03c6b0b, 32'h4060ab28} /* (2, 20, 31) {real, imag} */,
  {32'hc11f8386, 32'hbf8f6bde} /* (2, 20, 30) {real, imag} */,
  {32'hc01da997, 32'h400f896a} /* (2, 20, 29) {real, imag} */,
  {32'h3fccda0e, 32'hbede1908} /* (2, 20, 28) {real, imag} */,
  {32'hbfdc7068, 32'hbf2d4e88} /* (2, 20, 27) {real, imag} */,
  {32'hc0479020, 32'h40f131ba} /* (2, 20, 26) {real, imag} */,
  {32'hc1a5acc6, 32'hc0e8b30e} /* (2, 20, 25) {real, imag} */,
  {32'h40949283, 32'h41453686} /* (2, 20, 24) {real, imag} */,
  {32'h40514877, 32'h410f5550} /* (2, 20, 23) {real, imag} */,
  {32'h41759b44, 32'h4157f1b0} /* (2, 20, 22) {real, imag} */,
  {32'hc1441ed2, 32'h416e752c} /* (2, 20, 21) {real, imag} */,
  {32'hc0755008, 32'hbfc0e9b6} /* (2, 20, 20) {real, imag} */,
  {32'hc13c8b41, 32'hc1b99c3b} /* (2, 20, 19) {real, imag} */,
  {32'hc110827b, 32'h3fed0518} /* (2, 20, 18) {real, imag} */,
  {32'hbfb08ad7, 32'hc1868468} /* (2, 20, 17) {real, imag} */,
  {32'h3ffec3eb, 32'hc162345c} /* (2, 20, 16) {real, imag} */,
  {32'hc1181faa, 32'hc17a7d9a} /* (2, 20, 15) {real, imag} */,
  {32'hc115a57c, 32'hc19794f4} /* (2, 20, 14) {real, imag} */,
  {32'hc15bbd3a, 32'hc129b239} /* (2, 20, 13) {real, imag} */,
  {32'h418eb4a7, 32'hc0bc2441} /* (2, 20, 12) {real, imag} */,
  {32'h41323823, 32'h409c4437} /* (2, 20, 11) {real, imag} */,
  {32'h4026977c, 32'h40f338b4} /* (2, 20, 10) {real, imag} */,
  {32'h40ee8af4, 32'h3f9d3ac2} /* (2, 20, 9) {real, imag} */,
  {32'hc06658fb, 32'hc0e7bbda} /* (2, 20, 8) {real, imag} */,
  {32'h4124e712, 32'h413265a9} /* (2, 20, 7) {real, imag} */,
  {32'h409bc772, 32'hc1381e78} /* (2, 20, 6) {real, imag} */,
  {32'h414b292f, 32'h411180f5} /* (2, 20, 5) {real, imag} */,
  {32'h40cbb529, 32'hc09215a5} /* (2, 20, 4) {real, imag} */,
  {32'h41640260, 32'h414de44a} /* (2, 20, 3) {real, imag} */,
  {32'h405c449c, 32'hbe4d1c00} /* (2, 20, 2) {real, imag} */,
  {32'h4170e490, 32'h415bdf4a} /* (2, 20, 1) {real, imag} */,
  {32'h40f16628, 32'h4114c54f} /* (2, 20, 0) {real, imag} */,
  {32'h40ef7810, 32'hc13bfd7e} /* (2, 19, 31) {real, imag} */,
  {32'h3f819a4c, 32'hc0c28f84} /* (2, 19, 30) {real, imag} */,
  {32'hbfd2f394, 32'hc138a80e} /* (2, 19, 29) {real, imag} */,
  {32'hc1aa6816, 32'hc1458ec1} /* (2, 19, 28) {real, imag} */,
  {32'h41684603, 32'h40caa200} /* (2, 19, 27) {real, imag} */,
  {32'hc0438270, 32'h412f16e2} /* (2, 19, 26) {real, imag} */,
  {32'hc11ff6e7, 32'hc084d333} /* (2, 19, 25) {real, imag} */,
  {32'hc16e1339, 32'hc13f2640} /* (2, 19, 24) {real, imag} */,
  {32'h40d6e36a, 32'h41914560} /* (2, 19, 23) {real, imag} */,
  {32'hc165cde0, 32'hc0ad3300} /* (2, 19, 22) {real, imag} */,
  {32'hc0dedf98, 32'h41851b42} /* (2, 19, 21) {real, imag} */,
  {32'hc0fb67b8, 32'h410393ec} /* (2, 19, 20) {real, imag} */,
  {32'hbfc21e2c, 32'h3fd3e811} /* (2, 19, 19) {real, imag} */,
  {32'hc1273eb3, 32'hc1a5edd2} /* (2, 19, 18) {real, imag} */,
  {32'h400bc480, 32'h3fff4fa8} /* (2, 19, 17) {real, imag} */,
  {32'hc11b85b5, 32'h4018817a} /* (2, 19, 16) {real, imag} */,
  {32'hbf8f46cc, 32'hc149d364} /* (2, 19, 15) {real, imag} */,
  {32'h4140b11e, 32'h4119b99c} /* (2, 19, 14) {real, imag} */,
  {32'hc19a3f60, 32'hc10a7fa4} /* (2, 19, 13) {real, imag} */,
  {32'hbfbbeefe, 32'h407f0648} /* (2, 19, 12) {real, imag} */,
  {32'hbf8fe33e, 32'hc05703f4} /* (2, 19, 11) {real, imag} */,
  {32'hbfff01e4, 32'h410ec673} /* (2, 19, 10) {real, imag} */,
  {32'hc1051097, 32'h407e5f90} /* (2, 19, 9) {real, imag} */,
  {32'h413198b7, 32'h3da47140} /* (2, 19, 8) {real, imag} */,
  {32'h40e872aa, 32'hc11c3797} /* (2, 19, 7) {real, imag} */,
  {32'hbfe72312, 32'h3ea97e40} /* (2, 19, 6) {real, imag} */,
  {32'hc0a50985, 32'h3f3dd89c} /* (2, 19, 5) {real, imag} */,
  {32'hc0aa4ce2, 32'h3ff06b86} /* (2, 19, 4) {real, imag} */,
  {32'hc02d0beb, 32'hc09f769b} /* (2, 19, 3) {real, imag} */,
  {32'h407ccfd0, 32'h410f5806} /* (2, 19, 2) {real, imag} */,
  {32'hc15f89ee, 32'h4151069c} /* (2, 19, 1) {real, imag} */,
  {32'hc1181e2c, 32'h416da6e7} /* (2, 19, 0) {real, imag} */,
  {32'h413b3896, 32'hc0a53f58} /* (2, 18, 31) {real, imag} */,
  {32'hc103baef, 32'hc00d0212} /* (2, 18, 30) {real, imag} */,
  {32'hc0de521f, 32'hbfb1053c} /* (2, 18, 29) {real, imag} */,
  {32'h405679a6, 32'hbfe802a4} /* (2, 18, 28) {real, imag} */,
  {32'hbff436f4, 32'h4145ea9a} /* (2, 18, 27) {real, imag} */,
  {32'h4022065c, 32'hc0dd0cd6} /* (2, 18, 26) {real, imag} */,
  {32'hc1181398, 32'hc1b688f7} /* (2, 18, 25) {real, imag} */,
  {32'hc1475721, 32'hc09cf1c8} /* (2, 18, 24) {real, imag} */,
  {32'h419832ab, 32'hc19ad2be} /* (2, 18, 23) {real, imag} */,
  {32'hc1482816, 32'hc07e589a} /* (2, 18, 22) {real, imag} */,
  {32'h41833589, 32'h4151827f} /* (2, 18, 21) {real, imag} */,
  {32'h407ba27e, 32'h416cef91} /* (2, 18, 20) {real, imag} */,
  {32'h4070356a, 32'h41ab96d4} /* (2, 18, 19) {real, imag} */,
  {32'hc054b400, 32'h4068e0a8} /* (2, 18, 18) {real, imag} */,
  {32'h412b93a1, 32'hc05e86b9} /* (2, 18, 17) {real, imag} */,
  {32'hc121e99a, 32'h40aa8c38} /* (2, 18, 16) {real, imag} */,
  {32'h40ad576a, 32'hc0d50b62} /* (2, 18, 15) {real, imag} */,
  {32'hc10f9e87, 32'hc0dac9da} /* (2, 18, 14) {real, imag} */,
  {32'hbf5a2604, 32'hbfc0c930} /* (2, 18, 13) {real, imag} */,
  {32'hc0f8bda5, 32'h41a1dab2} /* (2, 18, 12) {real, imag} */,
  {32'hc04cdf7a, 32'h41a12ffd} /* (2, 18, 11) {real, imag} */,
  {32'h40b485ba, 32'hc178ba26} /* (2, 18, 10) {real, imag} */,
  {32'hc1d4a70c, 32'h4018bfa4} /* (2, 18, 9) {real, imag} */,
  {32'hc0dfdadc, 32'hc06b5801} /* (2, 18, 8) {real, imag} */,
  {32'hbc086000, 32'hc11f29b1} /* (2, 18, 7) {real, imag} */,
  {32'h406af564, 32'h410d6366} /* (2, 18, 6) {real, imag} */,
  {32'hc0a7f9c1, 32'hbfcf33ac} /* (2, 18, 5) {real, imag} */,
  {32'h41810098, 32'hc137ddf6} /* (2, 18, 4) {real, imag} */,
  {32'h4107526f, 32'h4119e75c} /* (2, 18, 3) {real, imag} */,
  {32'hc0569866, 32'h411bee80} /* (2, 18, 2) {real, imag} */,
  {32'h3f96bee4, 32'hc1b6e4a8} /* (2, 18, 1) {real, imag} */,
  {32'hc02335c2, 32'h403c2b16} /* (2, 18, 0) {real, imag} */,
  {32'h40850424, 32'h4167f44e} /* (2, 17, 31) {real, imag} */,
  {32'hc0d9381c, 32'hc0b62eac} /* (2, 17, 30) {real, imag} */,
  {32'h407f4cd4, 32'hc09550e2} /* (2, 17, 29) {real, imag} */,
  {32'h41179a10, 32'hc0c2257c} /* (2, 17, 28) {real, imag} */,
  {32'hc0b7ea58, 32'h409850a3} /* (2, 17, 27) {real, imag} */,
  {32'h40c9ae36, 32'hc1095caf} /* (2, 17, 26) {real, imag} */,
  {32'h40aa3227, 32'h402d37dd} /* (2, 17, 25) {real, imag} */,
  {32'hc0f5700a, 32'hc05851be} /* (2, 17, 24) {real, imag} */,
  {32'hc15dcc0b, 32'hc0a62cb2} /* (2, 17, 23) {real, imag} */,
  {32'h41407082, 32'hc020d6bb} /* (2, 17, 22) {real, imag} */,
  {32'hc091caf8, 32'h417fb04e} /* (2, 17, 21) {real, imag} */,
  {32'h40adbdbd, 32'hc08bb1b2} /* (2, 17, 20) {real, imag} */,
  {32'hc10a0bab, 32'hc0a027f4} /* (2, 17, 19) {real, imag} */,
  {32'hc0f3958f, 32'h3fedeb6c} /* (2, 17, 18) {real, imag} */,
  {32'hc08fb784, 32'h400774a4} /* (2, 17, 17) {real, imag} */,
  {32'h40f23a0f, 32'h4104618b} /* (2, 17, 16) {real, imag} */,
  {32'hc0aeac21, 32'h3fc07d54} /* (2, 17, 15) {real, imag} */,
  {32'hc0bc6c8e, 32'hc093338e} /* (2, 17, 14) {real, imag} */,
  {32'h3eec7c80, 32'h41a5c8b3} /* (2, 17, 13) {real, imag} */,
  {32'h404109e3, 32'hc168077a} /* (2, 17, 12) {real, imag} */,
  {32'h41749654, 32'hbdadd580} /* (2, 17, 11) {real, imag} */,
  {32'h405cafee, 32'hc0caae3e} /* (2, 17, 10) {real, imag} */,
  {32'h4105bd25, 32'hc1339f98} /* (2, 17, 9) {real, imag} */,
  {32'h4186f1f6, 32'h412681b7} /* (2, 17, 8) {real, imag} */,
  {32'hc0b2404f, 32'hc17c9060} /* (2, 17, 7) {real, imag} */,
  {32'h408485f8, 32'hc00991a5} /* (2, 17, 6) {real, imag} */,
  {32'h41817b3a, 32'h414ab793} /* (2, 17, 5) {real, imag} */,
  {32'hc049e498, 32'h40ab07c4} /* (2, 17, 4) {real, imag} */,
  {32'hc0a62469, 32'h402b9b77} /* (2, 17, 3) {real, imag} */,
  {32'hc0d48bf0, 32'hbf9184a0} /* (2, 17, 2) {real, imag} */,
  {32'hc0ca0338, 32'h4102f1aa} /* (2, 17, 1) {real, imag} */,
  {32'hc0e8dfd4, 32'h3ee55a88} /* (2, 17, 0) {real, imag} */,
  {32'h402eef54, 32'h4073060d} /* (2, 16, 31) {real, imag} */,
  {32'h4098ae3f, 32'h40b38c2c} /* (2, 16, 30) {real, imag} */,
  {32'hc137959d, 32'h419dd25c} /* (2, 16, 29) {real, imag} */,
  {32'h409d9bd3, 32'h41071093} /* (2, 16, 28) {real, imag} */,
  {32'h409497b6, 32'hc07d1a38} /* (2, 16, 27) {real, imag} */,
  {32'h3fe885fa, 32'h40d5665a} /* (2, 16, 26) {real, imag} */,
  {32'hc03a188e, 32'hbfd1fd80} /* (2, 16, 25) {real, imag} */,
  {32'hc1035dc0, 32'h4147dd90} /* (2, 16, 24) {real, imag} */,
  {32'hc10b892e, 32'hc0fa6985} /* (2, 16, 23) {real, imag} */,
  {32'h3f912fa4, 32'hc10ec5ce} /* (2, 16, 22) {real, imag} */,
  {32'hc094e864, 32'h40ed4942} /* (2, 16, 21) {real, imag} */,
  {32'h410123b7, 32'hbf7f4288} /* (2, 16, 20) {real, imag} */,
  {32'h40bdf236, 32'hc13d7a9a} /* (2, 16, 19) {real, imag} */,
  {32'h40e0ddd1, 32'hbe329d00} /* (2, 16, 18) {real, imag} */,
  {32'hc0cb72b6, 32'hc0ecb332} /* (2, 16, 17) {real, imag} */,
  {32'hbf3147a8, 32'h00000000} /* (2, 16, 16) {real, imag} */,
  {32'hc0cb72b6, 32'h40ecb332} /* (2, 16, 15) {real, imag} */,
  {32'h40e0ddd1, 32'h3e329d00} /* (2, 16, 14) {real, imag} */,
  {32'h40bdf236, 32'h413d7a9a} /* (2, 16, 13) {real, imag} */,
  {32'h410123b7, 32'h3f7f4288} /* (2, 16, 12) {real, imag} */,
  {32'hc094e864, 32'hc0ed4942} /* (2, 16, 11) {real, imag} */,
  {32'h3f912fa4, 32'h410ec5ce} /* (2, 16, 10) {real, imag} */,
  {32'hc10b892e, 32'h40fa6985} /* (2, 16, 9) {real, imag} */,
  {32'hc1035dc0, 32'hc147dd90} /* (2, 16, 8) {real, imag} */,
  {32'hc03a188e, 32'h3fd1fd80} /* (2, 16, 7) {real, imag} */,
  {32'h3fe885fa, 32'hc0d5665a} /* (2, 16, 6) {real, imag} */,
  {32'h409497b6, 32'h407d1a38} /* (2, 16, 5) {real, imag} */,
  {32'h409d9bd3, 32'hc1071093} /* (2, 16, 4) {real, imag} */,
  {32'hc137959d, 32'hc19dd25c} /* (2, 16, 3) {real, imag} */,
  {32'h4098ae3f, 32'hc0b38c2c} /* (2, 16, 2) {real, imag} */,
  {32'h402eef54, 32'hc073060d} /* (2, 16, 1) {real, imag} */,
  {32'hc0a4dba6, 32'h00000000} /* (2, 16, 0) {real, imag} */,
  {32'hc0ca0338, 32'hc102f1aa} /* (2, 15, 31) {real, imag} */,
  {32'hc0d48bf0, 32'h3f9184a0} /* (2, 15, 30) {real, imag} */,
  {32'hc0a62469, 32'hc02b9b77} /* (2, 15, 29) {real, imag} */,
  {32'hc049e498, 32'hc0ab07c4} /* (2, 15, 28) {real, imag} */,
  {32'h41817b3a, 32'hc14ab793} /* (2, 15, 27) {real, imag} */,
  {32'h408485f8, 32'h400991a5} /* (2, 15, 26) {real, imag} */,
  {32'hc0b2404f, 32'h417c9060} /* (2, 15, 25) {real, imag} */,
  {32'h4186f1f6, 32'hc12681b7} /* (2, 15, 24) {real, imag} */,
  {32'h4105bd25, 32'h41339f98} /* (2, 15, 23) {real, imag} */,
  {32'h405cafee, 32'h40caae3e} /* (2, 15, 22) {real, imag} */,
  {32'h41749654, 32'h3dadd580} /* (2, 15, 21) {real, imag} */,
  {32'h404109e3, 32'h4168077a} /* (2, 15, 20) {real, imag} */,
  {32'h3eec7c80, 32'hc1a5c8b3} /* (2, 15, 19) {real, imag} */,
  {32'hc0bc6c8e, 32'h4093338e} /* (2, 15, 18) {real, imag} */,
  {32'hc0aeac21, 32'hbfc07d54} /* (2, 15, 17) {real, imag} */,
  {32'h40f23a0f, 32'hc104618b} /* (2, 15, 16) {real, imag} */,
  {32'hc08fb784, 32'hc00774a4} /* (2, 15, 15) {real, imag} */,
  {32'hc0f3958f, 32'hbfedeb6c} /* (2, 15, 14) {real, imag} */,
  {32'hc10a0bab, 32'h40a027f4} /* (2, 15, 13) {real, imag} */,
  {32'h40adbdbd, 32'h408bb1b2} /* (2, 15, 12) {real, imag} */,
  {32'hc091caf8, 32'hc17fb04e} /* (2, 15, 11) {real, imag} */,
  {32'h41407082, 32'h4020d6bb} /* (2, 15, 10) {real, imag} */,
  {32'hc15dcc0b, 32'h40a62cb2} /* (2, 15, 9) {real, imag} */,
  {32'hc0f5700a, 32'h405851be} /* (2, 15, 8) {real, imag} */,
  {32'h40aa3227, 32'hc02d37dd} /* (2, 15, 7) {real, imag} */,
  {32'h40c9ae36, 32'h41095caf} /* (2, 15, 6) {real, imag} */,
  {32'hc0b7ea58, 32'hc09850a3} /* (2, 15, 5) {real, imag} */,
  {32'h41179a10, 32'h40c2257c} /* (2, 15, 4) {real, imag} */,
  {32'h407f4cd4, 32'h409550e2} /* (2, 15, 3) {real, imag} */,
  {32'hc0d9381c, 32'h40b62eac} /* (2, 15, 2) {real, imag} */,
  {32'h40850424, 32'hc167f44e} /* (2, 15, 1) {real, imag} */,
  {32'hc0e8dfd4, 32'hbee55a88} /* (2, 15, 0) {real, imag} */,
  {32'h3f96bee4, 32'h41b6e4a8} /* (2, 14, 31) {real, imag} */,
  {32'hc0569866, 32'hc11bee80} /* (2, 14, 30) {real, imag} */,
  {32'h4107526f, 32'hc119e75c} /* (2, 14, 29) {real, imag} */,
  {32'h41810098, 32'h4137ddf6} /* (2, 14, 28) {real, imag} */,
  {32'hc0a7f9c1, 32'h3fcf33ac} /* (2, 14, 27) {real, imag} */,
  {32'h406af564, 32'hc10d6366} /* (2, 14, 26) {real, imag} */,
  {32'hbc086000, 32'h411f29b1} /* (2, 14, 25) {real, imag} */,
  {32'hc0dfdadc, 32'h406b5801} /* (2, 14, 24) {real, imag} */,
  {32'hc1d4a70c, 32'hc018bfa4} /* (2, 14, 23) {real, imag} */,
  {32'h40b485ba, 32'h4178ba26} /* (2, 14, 22) {real, imag} */,
  {32'hc04cdf7a, 32'hc1a12ffd} /* (2, 14, 21) {real, imag} */,
  {32'hc0f8bda5, 32'hc1a1dab2} /* (2, 14, 20) {real, imag} */,
  {32'hbf5a2604, 32'h3fc0c930} /* (2, 14, 19) {real, imag} */,
  {32'hc10f9e87, 32'h40dac9da} /* (2, 14, 18) {real, imag} */,
  {32'h40ad576a, 32'h40d50b62} /* (2, 14, 17) {real, imag} */,
  {32'hc121e99a, 32'hc0aa8c38} /* (2, 14, 16) {real, imag} */,
  {32'h412b93a1, 32'h405e86b9} /* (2, 14, 15) {real, imag} */,
  {32'hc054b400, 32'hc068e0a8} /* (2, 14, 14) {real, imag} */,
  {32'h4070356a, 32'hc1ab96d4} /* (2, 14, 13) {real, imag} */,
  {32'h407ba27e, 32'hc16cef91} /* (2, 14, 12) {real, imag} */,
  {32'h41833589, 32'hc151827f} /* (2, 14, 11) {real, imag} */,
  {32'hc1482816, 32'h407e589a} /* (2, 14, 10) {real, imag} */,
  {32'h419832ab, 32'h419ad2be} /* (2, 14, 9) {real, imag} */,
  {32'hc1475721, 32'h409cf1c8} /* (2, 14, 8) {real, imag} */,
  {32'hc1181398, 32'h41b688f7} /* (2, 14, 7) {real, imag} */,
  {32'h4022065c, 32'h40dd0cd6} /* (2, 14, 6) {real, imag} */,
  {32'hbff436f4, 32'hc145ea9a} /* (2, 14, 5) {real, imag} */,
  {32'h405679a6, 32'h3fe802a4} /* (2, 14, 4) {real, imag} */,
  {32'hc0de521f, 32'h3fb1053c} /* (2, 14, 3) {real, imag} */,
  {32'hc103baef, 32'h400d0212} /* (2, 14, 2) {real, imag} */,
  {32'h413b3896, 32'h40a53f58} /* (2, 14, 1) {real, imag} */,
  {32'hc02335c2, 32'hc03c2b16} /* (2, 14, 0) {real, imag} */,
  {32'hc15f89ee, 32'hc151069c} /* (2, 13, 31) {real, imag} */,
  {32'h407ccfd0, 32'hc10f5806} /* (2, 13, 30) {real, imag} */,
  {32'hc02d0beb, 32'h409f769b} /* (2, 13, 29) {real, imag} */,
  {32'hc0aa4ce2, 32'hbff06b86} /* (2, 13, 28) {real, imag} */,
  {32'hc0a50985, 32'hbf3dd89c} /* (2, 13, 27) {real, imag} */,
  {32'hbfe72312, 32'hbea97e40} /* (2, 13, 26) {real, imag} */,
  {32'h40e872aa, 32'h411c3797} /* (2, 13, 25) {real, imag} */,
  {32'h413198b7, 32'hbda47140} /* (2, 13, 24) {real, imag} */,
  {32'hc1051097, 32'hc07e5f90} /* (2, 13, 23) {real, imag} */,
  {32'hbfff01e4, 32'hc10ec673} /* (2, 13, 22) {real, imag} */,
  {32'hbf8fe33e, 32'h405703f4} /* (2, 13, 21) {real, imag} */,
  {32'hbfbbeefe, 32'hc07f0648} /* (2, 13, 20) {real, imag} */,
  {32'hc19a3f60, 32'h410a7fa4} /* (2, 13, 19) {real, imag} */,
  {32'h4140b11e, 32'hc119b99c} /* (2, 13, 18) {real, imag} */,
  {32'hbf8f46cc, 32'h4149d364} /* (2, 13, 17) {real, imag} */,
  {32'hc11b85b5, 32'hc018817a} /* (2, 13, 16) {real, imag} */,
  {32'h400bc480, 32'hbfff4fa8} /* (2, 13, 15) {real, imag} */,
  {32'hc1273eb3, 32'h41a5edd2} /* (2, 13, 14) {real, imag} */,
  {32'hbfc21e2c, 32'hbfd3e811} /* (2, 13, 13) {real, imag} */,
  {32'hc0fb67b8, 32'hc10393ec} /* (2, 13, 12) {real, imag} */,
  {32'hc0dedf98, 32'hc1851b42} /* (2, 13, 11) {real, imag} */,
  {32'hc165cde0, 32'h40ad3300} /* (2, 13, 10) {real, imag} */,
  {32'h40d6e36a, 32'hc1914560} /* (2, 13, 9) {real, imag} */,
  {32'hc16e1339, 32'h413f2640} /* (2, 13, 8) {real, imag} */,
  {32'hc11ff6e7, 32'h4084d333} /* (2, 13, 7) {real, imag} */,
  {32'hc0438270, 32'hc12f16e2} /* (2, 13, 6) {real, imag} */,
  {32'h41684603, 32'hc0caa200} /* (2, 13, 5) {real, imag} */,
  {32'hc1aa6816, 32'h41458ec1} /* (2, 13, 4) {real, imag} */,
  {32'hbfd2f394, 32'h4138a80e} /* (2, 13, 3) {real, imag} */,
  {32'h3f819a4c, 32'h40c28f84} /* (2, 13, 2) {real, imag} */,
  {32'h40ef7810, 32'h413bfd7e} /* (2, 13, 1) {real, imag} */,
  {32'hc1181e2c, 32'hc16da6e7} /* (2, 13, 0) {real, imag} */,
  {32'h4170e490, 32'hc15bdf4a} /* (2, 12, 31) {real, imag} */,
  {32'h405c449c, 32'h3e4d1c00} /* (2, 12, 30) {real, imag} */,
  {32'h41640260, 32'hc14de44a} /* (2, 12, 29) {real, imag} */,
  {32'h40cbb529, 32'h409215a5} /* (2, 12, 28) {real, imag} */,
  {32'h414b292f, 32'hc11180f5} /* (2, 12, 27) {real, imag} */,
  {32'h409bc772, 32'h41381e78} /* (2, 12, 26) {real, imag} */,
  {32'h4124e712, 32'hc13265a9} /* (2, 12, 25) {real, imag} */,
  {32'hc06658fb, 32'h40e7bbda} /* (2, 12, 24) {real, imag} */,
  {32'h40ee8af4, 32'hbf9d3ac2} /* (2, 12, 23) {real, imag} */,
  {32'h4026977c, 32'hc0f338b4} /* (2, 12, 22) {real, imag} */,
  {32'h41323823, 32'hc09c4437} /* (2, 12, 21) {real, imag} */,
  {32'h418eb4a7, 32'h40bc2441} /* (2, 12, 20) {real, imag} */,
  {32'hc15bbd3a, 32'h4129b239} /* (2, 12, 19) {real, imag} */,
  {32'hc115a57c, 32'h419794f4} /* (2, 12, 18) {real, imag} */,
  {32'hc1181faa, 32'h417a7d9a} /* (2, 12, 17) {real, imag} */,
  {32'h3ffec3eb, 32'h4162345c} /* (2, 12, 16) {real, imag} */,
  {32'hbfb08ad7, 32'h41868468} /* (2, 12, 15) {real, imag} */,
  {32'hc110827b, 32'hbfed0518} /* (2, 12, 14) {real, imag} */,
  {32'hc13c8b41, 32'h41b99c3b} /* (2, 12, 13) {real, imag} */,
  {32'hc0755008, 32'h3fc0e9b6} /* (2, 12, 12) {real, imag} */,
  {32'hc1441ed2, 32'hc16e752c} /* (2, 12, 11) {real, imag} */,
  {32'h41759b44, 32'hc157f1b0} /* (2, 12, 10) {real, imag} */,
  {32'h40514877, 32'hc10f5550} /* (2, 12, 9) {real, imag} */,
  {32'h40949283, 32'hc1453686} /* (2, 12, 8) {real, imag} */,
  {32'hc1a5acc6, 32'h40e8b30e} /* (2, 12, 7) {real, imag} */,
  {32'hc0479020, 32'hc0f131ba} /* (2, 12, 6) {real, imag} */,
  {32'hbfdc7068, 32'h3f2d4e88} /* (2, 12, 5) {real, imag} */,
  {32'h3fccda0e, 32'h3ede1908} /* (2, 12, 4) {real, imag} */,
  {32'hc01da997, 32'hc00f896a} /* (2, 12, 3) {real, imag} */,
  {32'hc11f8386, 32'h3f8f6bde} /* (2, 12, 2) {real, imag} */,
  {32'hc03c6b0b, 32'hc060ab28} /* (2, 12, 1) {real, imag} */,
  {32'h40f16628, 32'hc114c54f} /* (2, 12, 0) {real, imag} */,
  {32'h4196ef36, 32'h42122388} /* (2, 11, 31) {real, imag} */,
  {32'hc1ab3811, 32'h40819c74} /* (2, 11, 30) {real, imag} */,
  {32'hc02e3c38, 32'hc1220466} /* (2, 11, 29) {real, imag} */,
  {32'hc0edcd6c, 32'h3f4849c8} /* (2, 11, 28) {real, imag} */,
  {32'h411dc6fe, 32'h40b8c42c} /* (2, 11, 27) {real, imag} */,
  {32'h3ff498f4, 32'h4110fb77} /* (2, 11, 26) {real, imag} */,
  {32'hc0efdc5e, 32'hc0879e98} /* (2, 11, 25) {real, imag} */,
  {32'h41247580, 32'hc0619368} /* (2, 11, 24) {real, imag} */,
  {32'hc01560a0, 32'h4125ad45} /* (2, 11, 23) {real, imag} */,
  {32'h416d52aa, 32'h3f16f6d4} /* (2, 11, 22) {real, imag} */,
  {32'hc0ae3806, 32'h415eedac} /* (2, 11, 21) {real, imag} */,
  {32'h40bb2d34, 32'h3f5bb608} /* (2, 11, 20) {real, imag} */,
  {32'h3cc29e00, 32'h40da7cd4} /* (2, 11, 19) {real, imag} */,
  {32'h41193444, 32'hbfc771e8} /* (2, 11, 18) {real, imag} */,
  {32'hc08f21e6, 32'hc07487d9} /* (2, 11, 17) {real, imag} */,
  {32'hbfdb6788, 32'h41319e82} /* (2, 11, 16) {real, imag} */,
  {32'hbfeab7b8, 32'h4076ca36} /* (2, 11, 15) {real, imag} */,
  {32'h40d7970c, 32'h40df68fe} /* (2, 11, 14) {real, imag} */,
  {32'hc11a8fa0, 32'hc042fc27} /* (2, 11, 13) {real, imag} */,
  {32'h401f56b1, 32'hbfb609f4} /* (2, 11, 12) {real, imag} */,
  {32'h40c3509c, 32'hc122aa90} /* (2, 11, 11) {real, imag} */,
  {32'h3ff0c590, 32'hc0758f2a} /* (2, 11, 10) {real, imag} */,
  {32'h412a1890, 32'hc0d6139b} /* (2, 11, 9) {real, imag} */,
  {32'h417a817c, 32'hc180c014} /* (2, 11, 8) {real, imag} */,
  {32'hc0b9bb5b, 32'hbf5d1108} /* (2, 11, 7) {real, imag} */,
  {32'hbeb6be80, 32'hbf0b53d0} /* (2, 11, 6) {real, imag} */,
  {32'h41238fa2, 32'h3fbccc18} /* (2, 11, 5) {real, imag} */,
  {32'h40fe8260, 32'hc1151a90} /* (2, 11, 4) {real, imag} */,
  {32'h401c9bb6, 32'h415340b8} /* (2, 11, 3) {real, imag} */,
  {32'hbf4124f0, 32'hc18fba86} /* (2, 11, 2) {real, imag} */,
  {32'h41150630, 32'h41a42e12} /* (2, 11, 1) {real, imag} */,
  {32'h413469dc, 32'h41293396} /* (2, 11, 0) {real, imag} */,
  {32'h3fe40ef4, 32'hc0940576} /* (2, 10, 31) {real, imag} */,
  {32'h4134688d, 32'h41c52bea} /* (2, 10, 30) {real, imag} */,
  {32'hc1967067, 32'h40ed43c3} /* (2, 10, 29) {real, imag} */,
  {32'hc1a1e576, 32'hc02b89c0} /* (2, 10, 28) {real, imag} */,
  {32'h408272f6, 32'hbfac3246} /* (2, 10, 27) {real, imag} */,
  {32'h40eaf2d5, 32'hc0bbca7f} /* (2, 10, 26) {real, imag} */,
  {32'hc0aab2c3, 32'hc08dad3a} /* (2, 10, 25) {real, imag} */,
  {32'hc16505a2, 32'hc0b7af91} /* (2, 10, 24) {real, imag} */,
  {32'hc0b6b027, 32'hc11d074b} /* (2, 10, 23) {real, imag} */,
  {32'hc16ca7f2, 32'hbefcc3e0} /* (2, 10, 22) {real, imag} */,
  {32'hc02d610c, 32'hc1a5b692} /* (2, 10, 21) {real, imag} */,
  {32'hc054028c, 32'h40747258} /* (2, 10, 20) {real, imag} */,
  {32'h412e2f0a, 32'hc1a7b408} /* (2, 10, 19) {real, imag} */,
  {32'h4072225e, 32'h413d9596} /* (2, 10, 18) {real, imag} */,
  {32'hc143f2f8, 32'hbececd68} /* (2, 10, 17) {real, imag} */,
  {32'h4115e3f7, 32'h40bb5cc8} /* (2, 10, 16) {real, imag} */,
  {32'h3ebd2228, 32'hc0dd7372} /* (2, 10, 15) {real, imag} */,
  {32'h405b1868, 32'hbfe40ea8} /* (2, 10, 14) {real, imag} */,
  {32'h4080f4e8, 32'hc1894c5c} /* (2, 10, 13) {real, imag} */,
  {32'hc1548b1e, 32'hc02e6715} /* (2, 10, 12) {real, imag} */,
  {32'hc0e962f4, 32'hc196297a} /* (2, 10, 11) {real, imag} */,
  {32'h418e1da1, 32'h4060f4ee} /* (2, 10, 10) {real, imag} */,
  {32'h40fd4cbf, 32'h418818b2} /* (2, 10, 9) {real, imag} */,
  {32'hc15a52f2, 32'h40a761d4} /* (2, 10, 8) {real, imag} */,
  {32'h4124ffbc, 32'h40153900} /* (2, 10, 7) {real, imag} */,
  {32'h4174b908, 32'hc0c3f601} /* (2, 10, 6) {real, imag} */,
  {32'h3e1514e0, 32'h4151916e} /* (2, 10, 5) {real, imag} */,
  {32'h3ef972a8, 32'h4120fe8f} /* (2, 10, 4) {real, imag} */,
  {32'h41d1fe31, 32'h401f0d0e} /* (2, 10, 3) {real, imag} */,
  {32'hc16a6a0a, 32'h4198ed13} /* (2, 10, 2) {real, imag} */,
  {32'hc1a35a44, 32'hc13e38d8} /* (2, 10, 1) {real, imag} */,
  {32'h417ee158, 32'hc1228b36} /* (2, 10, 0) {real, imag} */,
  {32'h41618f6c, 32'h40a36b1b} /* (2, 9, 31) {real, imag} */,
  {32'h415e5689, 32'h41d5a3cb} /* (2, 9, 30) {real, imag} */,
  {32'hbf087320, 32'hc0fe949e} /* (2, 9, 29) {real, imag} */,
  {32'h40aedf54, 32'h403ee195} /* (2, 9, 28) {real, imag} */,
  {32'h419f648f, 32'h411d3858} /* (2, 9, 27) {real, imag} */,
  {32'h4120bcd6, 32'hc005d455} /* (2, 9, 26) {real, imag} */,
  {32'hc05afe68, 32'hbfc38a10} /* (2, 9, 25) {real, imag} */,
  {32'hc143e457, 32'h4045fdf8} /* (2, 9, 24) {real, imag} */,
  {32'h400433e4, 32'hc00d001e} /* (2, 9, 23) {real, imag} */,
  {32'h3fbe1a2a, 32'h3f7b5d38} /* (2, 9, 22) {real, imag} */,
  {32'hc0de5bd8, 32'h4189042c} /* (2, 9, 21) {real, imag} */,
  {32'hc18f57a3, 32'hc0ae70ea} /* (2, 9, 20) {real, imag} */,
  {32'hc1181f7c, 32'h407661ab} /* (2, 9, 19) {real, imag} */,
  {32'h41d158db, 32'hc002c7c2} /* (2, 9, 18) {real, imag} */,
  {32'hc10a31cd, 32'hc0dac8f3} /* (2, 9, 17) {real, imag} */,
  {32'h40a3887c, 32'h4114810c} /* (2, 9, 16) {real, imag} */,
  {32'hc155590c, 32'h413e7896} /* (2, 9, 15) {real, imag} */,
  {32'hc1547af4, 32'h41299f77} /* (2, 9, 14) {real, imag} */,
  {32'h412baef6, 32'hc0307e73} /* (2, 9, 13) {real, imag} */,
  {32'hc1abb034, 32'h410a4675} /* (2, 9, 12) {real, imag} */,
  {32'hc0aa84de, 32'h41860715} /* (2, 9, 11) {real, imag} */,
  {32'hc1187cda, 32'hbf501440} /* (2, 9, 10) {real, imag} */,
  {32'h41326b84, 32'h40a4bb01} /* (2, 9, 9) {real, imag} */,
  {32'hc14d9aeb, 32'hbf83aaf6} /* (2, 9, 8) {real, imag} */,
  {32'hbfaaa3ec, 32'hc0b2d79c} /* (2, 9, 7) {real, imag} */,
  {32'hc01f40ed, 32'h41b7eaa1} /* (2, 9, 6) {real, imag} */,
  {32'hc122f81e, 32'hc1ae8e61} /* (2, 9, 5) {real, imag} */,
  {32'hc12039f0, 32'hc1557300} /* (2, 9, 4) {real, imag} */,
  {32'hc1bba9c5, 32'h417c9595} /* (2, 9, 3) {real, imag} */,
  {32'h4092d7fa, 32'hc147a555} /* (2, 9, 2) {real, imag} */,
  {32'hc19094c7, 32'hc1de04b6} /* (2, 9, 1) {real, imag} */,
  {32'hc15ba0ba, 32'hc18a62da} /* (2, 9, 0) {real, imag} */,
  {32'h423fe59d, 32'h419a4594} /* (2, 8, 31) {real, imag} */,
  {32'hc20cfa02, 32'h41e694d0} /* (2, 8, 30) {real, imag} */,
  {32'hc19fb35e, 32'hc18e88a5} /* (2, 8, 29) {real, imag} */,
  {32'h3fbb2d59, 32'h41c9c9f2} /* (2, 8, 28) {real, imag} */,
  {32'hbf86ab10, 32'hc09bc73a} /* (2, 8, 27) {real, imag} */,
  {32'h413d1d6f, 32'h416f7384} /* (2, 8, 26) {real, imag} */,
  {32'h418faff6, 32'h41cdd8e2} /* (2, 8, 25) {real, imag} */,
  {32'h40901ce9, 32'h41a225b7} /* (2, 8, 24) {real, imag} */,
  {32'h41bf32c0, 32'h40fbc8dc} /* (2, 8, 23) {real, imag} */,
  {32'hc00cda56, 32'hc1ea78f4} /* (2, 8, 22) {real, imag} */,
  {32'h4082e90b, 32'hc1533d32} /* (2, 8, 21) {real, imag} */,
  {32'h4133342d, 32'hc0e8bfe0} /* (2, 8, 20) {real, imag} */,
  {32'hc019d4fa, 32'h419023ba} /* (2, 8, 19) {real, imag} */,
  {32'h3de3d300, 32'hc0a7d313} /* (2, 8, 18) {real, imag} */,
  {32'h40c68b38, 32'hc0c97ef6} /* (2, 8, 17) {real, imag} */,
  {32'h40149860, 32'h418a1288} /* (2, 8, 16) {real, imag} */,
  {32'h4091d26a, 32'h415b532d} /* (2, 8, 15) {real, imag} */,
  {32'hbfd336d8, 32'hc11dd96e} /* (2, 8, 14) {real, imag} */,
  {32'hc0a4a334, 32'hc1360167} /* (2, 8, 13) {real, imag} */,
  {32'h4192fbcb, 32'hc03da9a6} /* (2, 8, 12) {real, imag} */,
  {32'hc1127c2a, 32'hc1c461f6} /* (2, 8, 11) {real, imag} */,
  {32'hbec7f550, 32'h412a5696} /* (2, 8, 10) {real, imag} */,
  {32'hc16676e3, 32'h41c07b0d} /* (2, 8, 9) {real, imag} */,
  {32'hc0698978, 32'hbe118130} /* (2, 8, 8) {real, imag} */,
  {32'hc1a9fc84, 32'hc1541de4} /* (2, 8, 7) {real, imag} */,
  {32'hc13af802, 32'hc1f0b3d3} /* (2, 8, 6) {real, imag} */,
  {32'h400b8650, 32'hc05ba5de} /* (2, 8, 5) {real, imag} */,
  {32'h400c1e7c, 32'h400461c4} /* (2, 8, 4) {real, imag} */,
  {32'hc04dde4a, 32'hbf52aa68} /* (2, 8, 3) {real, imag} */,
  {32'h40a734a7, 32'hc1c54375} /* (2, 8, 2) {real, imag} */,
  {32'h416902b0, 32'h41f50973} /* (2, 8, 1) {real, imag} */,
  {32'h40faa4c2, 32'h400992f0} /* (2, 8, 0) {real, imag} */,
  {32'hc0c26dd5, 32'h404963f4} /* (2, 7, 31) {real, imag} */,
  {32'hbfa69134, 32'hc0ea0951} /* (2, 7, 30) {real, imag} */,
  {32'hc1acc2b0, 32'hc145907c} /* (2, 7, 29) {real, imag} */,
  {32'hc181c744, 32'h40442776} /* (2, 7, 28) {real, imag} */,
  {32'h3f8119c0, 32'h41595507} /* (2, 7, 27) {real, imag} */,
  {32'hbfbaaf78, 32'h410a8f43} /* (2, 7, 26) {real, imag} */,
  {32'hc1643679, 32'h41b07d50} /* (2, 7, 25) {real, imag} */,
  {32'h401ac684, 32'h3fc4d5a2} /* (2, 7, 24) {real, imag} */,
  {32'hc1bc1c48, 32'h40e2cba6} /* (2, 7, 23) {real, imag} */,
  {32'hc17d8217, 32'h413aff4a} /* (2, 7, 22) {real, imag} */,
  {32'h40df7bbe, 32'h40b37c92} /* (2, 7, 21) {real, imag} */,
  {32'h3f57bca0, 32'hc042dc70} /* (2, 7, 20) {real, imag} */,
  {32'h41515753, 32'hc0b4edfa} /* (2, 7, 19) {real, imag} */,
  {32'hc1351c5b, 32'h402e3b68} /* (2, 7, 18) {real, imag} */,
  {32'h40f06de8, 32'hc0e9b89e} /* (2, 7, 17) {real, imag} */,
  {32'hc0b7e982, 32'h408d246c} /* (2, 7, 16) {real, imag} */,
  {32'h41419d14, 32'hbfd35672} /* (2, 7, 15) {real, imag} */,
  {32'hc166df53, 32'hc1591c12} /* (2, 7, 14) {real, imag} */,
  {32'h40653529, 32'h4105883c} /* (2, 7, 13) {real, imag} */,
  {32'h3fdd95f0, 32'hc02bb37a} /* (2, 7, 12) {real, imag} */,
  {32'hc15772f4, 32'hc110dfd7} /* (2, 7, 11) {real, imag} */,
  {32'h4144f5cb, 32'h41d67524} /* (2, 7, 10) {real, imag} */,
  {32'h4136064f, 32'h416f7157} /* (2, 7, 9) {real, imag} */,
  {32'hc092352e, 32'hc123e63d} /* (2, 7, 8) {real, imag} */,
  {32'h40acf734, 32'h4059a068} /* (2, 7, 7) {real, imag} */,
  {32'hc0c600fe, 32'hc0a677f6} /* (2, 7, 6) {real, imag} */,
  {32'hbeb8ad50, 32'h416d54a2} /* (2, 7, 5) {real, imag} */,
  {32'hc0eaa11a, 32'hc16703ce} /* (2, 7, 4) {real, imag} */,
  {32'h41540ffa, 32'h405f7ff5} /* (2, 7, 3) {real, imag} */,
  {32'hc1420da0, 32'h416273dc} /* (2, 7, 2) {real, imag} */,
  {32'hc1825b20, 32'hc1325113} /* (2, 7, 1) {real, imag} */,
  {32'h3f96af50, 32'hc1553c41} /* (2, 7, 0) {real, imag} */,
  {32'hc1215b1a, 32'h418164d5} /* (2, 6, 31) {real, imag} */,
  {32'hbf946e00, 32'hc0fda365} /* (2, 6, 30) {real, imag} */,
  {32'h412a4c3a, 32'h4112bf4c} /* (2, 6, 29) {real, imag} */,
  {32'hc1c4d0d5, 32'hc1c0d341} /* (2, 6, 28) {real, imag} */,
  {32'h3fcf3b7e, 32'hc1e48fdc} /* (2, 6, 27) {real, imag} */,
  {32'h40a3e206, 32'hc118681d} /* (2, 6, 26) {real, imag} */,
  {32'hc11718a6, 32'hc04fb7dc} /* (2, 6, 25) {real, imag} */,
  {32'hc0b83389, 32'h419d6487} /* (2, 6, 24) {real, imag} */,
  {32'hc14a77ae, 32'h4086a392} /* (2, 6, 23) {real, imag} */,
  {32'h416c288f, 32'hc134ecea} /* (2, 6, 22) {real, imag} */,
  {32'hbfba5e68, 32'h40a0e058} /* (2, 6, 21) {real, imag} */,
  {32'h411db68c, 32'h412b7e73} /* (2, 6, 20) {real, imag} */,
  {32'h40f5d092, 32'h3bd5fc00} /* (2, 6, 19) {real, imag} */,
  {32'hc07b883a, 32'hc11c2f56} /* (2, 6, 18) {real, imag} */,
  {32'hc0edd045, 32'h404a342e} /* (2, 6, 17) {real, imag} */,
  {32'h3ea766e0, 32'hc11d811d} /* (2, 6, 16) {real, imag} */,
  {32'h3fd5a3c0, 32'hc040acfd} /* (2, 6, 15) {real, imag} */,
  {32'hbff8361a, 32'hc13d399a} /* (2, 6, 14) {real, imag} */,
  {32'hc1074c1c, 32'h40fd7acb} /* (2, 6, 13) {real, imag} */,
  {32'hc1867ea1, 32'hc15555f3} /* (2, 6, 12) {real, imag} */,
  {32'h4149d4e2, 32'hc09715d6} /* (2, 6, 11) {real, imag} */,
  {32'h419efe4b, 32'hc02df6e0} /* (2, 6, 10) {real, imag} */,
  {32'hbe04da00, 32'h41aa2bf2} /* (2, 6, 9) {real, imag} */,
  {32'hc10830ee, 32'hc0b92f8c} /* (2, 6, 8) {real, imag} */,
  {32'hc09e0792, 32'h41842dd0} /* (2, 6, 7) {real, imag} */,
  {32'hc10756ac, 32'h40993721} /* (2, 6, 6) {real, imag} */,
  {32'h405ca074, 32'hbed403c0} /* (2, 6, 5) {real, imag} */,
  {32'h40a6ed69, 32'hc088ef7d} /* (2, 6, 4) {real, imag} */,
  {32'hba404000, 32'hbfa8bd04} /* (2, 6, 3) {real, imag} */,
  {32'hc0f4f1c0, 32'hc1bae389} /* (2, 6, 2) {real, imag} */,
  {32'h40de2112, 32'hc13a4cd4} /* (2, 6, 1) {real, imag} */,
  {32'h4187d9f9, 32'h411d8f51} /* (2, 6, 0) {real, imag} */,
  {32'h42c374f4, 32'h40e2deb0} /* (2, 5, 31) {real, imag} */,
  {32'hc24d1080, 32'hc1bcd08a} /* (2, 5, 30) {real, imag} */,
  {32'hc09d0e2e, 32'h41435bb5} /* (2, 5, 29) {real, imag} */,
  {32'h41135a02, 32'hc132de17} /* (2, 5, 28) {real, imag} */,
  {32'hc1f852a9, 32'h40872b6d} /* (2, 5, 27) {real, imag} */,
  {32'h412ddb16, 32'hc1789de1} /* (2, 5, 26) {real, imag} */,
  {32'hc0aa7ce8, 32'h40150796} /* (2, 5, 25) {real, imag} */,
  {32'h3fc4bdd4, 32'h41d24eee} /* (2, 5, 24) {real, imag} */,
  {32'hc0f8e73d, 32'h4145bba7} /* (2, 5, 23) {real, imag} */,
  {32'hc0c7007e, 32'hc0792480} /* (2, 5, 22) {real, imag} */,
  {32'hc0f4f15c, 32'h40f24d09} /* (2, 5, 21) {real, imag} */,
  {32'hc0fc73f5, 32'hbff3d980} /* (2, 5, 20) {real, imag} */,
  {32'h402e8e9a, 32'h3ecb9d50} /* (2, 5, 19) {real, imag} */,
  {32'hc18e74c7, 32'h40630a50} /* (2, 5, 18) {real, imag} */,
  {32'hc051213a, 32'h40811b00} /* (2, 5, 17) {real, imag} */,
  {32'h4111e5e0, 32'hc0d6248c} /* (2, 5, 16) {real, imag} */,
  {32'hc1086afb, 32'h40c7f49f} /* (2, 5, 15) {real, imag} */,
  {32'hbf5f6284, 32'hc1353fc7} /* (2, 5, 14) {real, imag} */,
  {32'h410012bd, 32'h41348675} /* (2, 5, 13) {real, imag} */,
  {32'hc0472d94, 32'hc04ae2e4} /* (2, 5, 12) {real, imag} */,
  {32'hc0527d98, 32'h4098d8da} /* (2, 5, 11) {real, imag} */,
  {32'h40caf08c, 32'hbfd80a00} /* (2, 5, 10) {real, imag} */,
  {32'hc102b1ad, 32'h411ed95f} /* (2, 5, 9) {real, imag} */,
  {32'hbf962258, 32'hc116aa06} /* (2, 5, 8) {real, imag} */,
  {32'hc1e51ffa, 32'h40fd9fb2} /* (2, 5, 7) {real, imag} */,
  {32'h402bcdac, 32'hc0c0f16b} /* (2, 5, 6) {real, imag} */,
  {32'hc19e7668, 32'hc1b2d0ee} /* (2, 5, 5) {real, imag} */,
  {32'hc0ccd964, 32'hc0d1a49e} /* (2, 5, 4) {real, imag} */,
  {32'hc0330576, 32'hc10a9a44} /* (2, 5, 3) {real, imag} */,
  {32'h3fa36350, 32'hc176ef05} /* (2, 5, 2) {real, imag} */,
  {32'h4291edd5, 32'h42ca7164} /* (2, 5, 1) {real, imag} */,
  {32'h42b1a711, 32'h41b409b8} /* (2, 5, 0) {real, imag} */,
  {32'hc2841c49, 32'hc28e6902} /* (2, 4, 31) {real, imag} */,
  {32'h41895e18, 32'h42adbd78} /* (2, 4, 30) {real, imag} */,
  {32'hc162ad07, 32'h40c40cc0} /* (2, 4, 29) {real, imag} */,
  {32'hc1fad8bc, 32'hc1d225da} /* (2, 4, 28) {real, imag} */,
  {32'h41e21601, 32'h416a027e} /* (2, 4, 27) {real, imag} */,
  {32'h41498ca3, 32'hc1a3b74d} /* (2, 4, 26) {real, imag} */,
  {32'hc10b6d49, 32'hc19ae8d8} /* (2, 4, 25) {real, imag} */,
  {32'h40639b4b, 32'hc183ca5a} /* (2, 4, 24) {real, imag} */,
  {32'hc12cb2fe, 32'hc1123672} /* (2, 4, 23) {real, imag} */,
  {32'hc0f42a00, 32'h41398fe1} /* (2, 4, 22) {real, imag} */,
  {32'h41ce5102, 32'hc0eda2c0} /* (2, 4, 21) {real, imag} */,
  {32'h405d6d09, 32'hc12a590e} /* (2, 4, 20) {real, imag} */,
  {32'hc187d80d, 32'hbe7ef6f0} /* (2, 4, 19) {real, imag} */,
  {32'hc1461abe, 32'hc1218f56} /* (2, 4, 18) {real, imag} */,
  {32'hc0370de8, 32'hc0e665e8} /* (2, 4, 17) {real, imag} */,
  {32'h40b5f934, 32'h408b0111} /* (2, 4, 16) {real, imag} */,
  {32'h409db033, 32'hc05db040} /* (2, 4, 15) {real, imag} */,
  {32'h41432590, 32'h3f63aff8} /* (2, 4, 14) {real, imag} */,
  {32'h416a7e04, 32'h4120ecc4} /* (2, 4, 13) {real, imag} */,
  {32'h40e6bf48, 32'h40877e5e} /* (2, 4, 12) {real, imag} */,
  {32'hc0a35982, 32'h40de1908} /* (2, 4, 11) {real, imag} */,
  {32'hc0781cf6, 32'hbf535630} /* (2, 4, 10) {real, imag} */,
  {32'h410ee724, 32'hc07dff68} /* (2, 4, 9) {real, imag} */,
  {32'hc0e594d2, 32'h419eab97} /* (2, 4, 8) {real, imag} */,
  {32'hc19b42ef, 32'h40ab6100} /* (2, 4, 7) {real, imag} */,
  {32'h410d8a5e, 32'h4119e61c} /* (2, 4, 6) {real, imag} */,
  {32'hc0fd19a4, 32'h4034b3c8} /* (2, 4, 5) {real, imag} */,
  {32'hbff76008, 32'hc07663f8} /* (2, 4, 4) {real, imag} */,
  {32'h3f3979d8, 32'h418945fd} /* (2, 4, 3) {real, imag} */,
  {32'h42cfc2b9, 32'h42e4f8c0} /* (2, 4, 2) {real, imag} */,
  {32'hc3343598, 32'hc24adba7} /* (2, 4, 1) {real, imag} */,
  {32'hc28863b4, 32'hc1a68f73} /* (2, 4, 0) {real, imag} */,
  {32'h431f3a08, 32'hc2b44ce4} /* (2, 3, 31) {real, imag} */,
  {32'hc2973cba, 32'h428ef77f} /* (2, 3, 30) {real, imag} */,
  {32'hc227278c, 32'hc1db0308} /* (2, 3, 29) {real, imag} */,
  {32'hc053c17c, 32'hc12f335c} /* (2, 3, 28) {real, imag} */,
  {32'h403d9806, 32'h40ec0c68} /* (2, 3, 27) {real, imag} */,
  {32'h40c3fa4c, 32'h415da79e} /* (2, 3, 26) {real, imag} */,
  {32'hc1101cc3, 32'h40ef7cab} /* (2, 3, 25) {real, imag} */,
  {32'hc0f16765, 32'h41baff6c} /* (2, 3, 24) {real, imag} */,
  {32'hc1304b02, 32'hc207833b} /* (2, 3, 23) {real, imag} */,
  {32'hbf1c84b2, 32'h40bcbd52} /* (2, 3, 22) {real, imag} */,
  {32'hbf84c948, 32'hc0dd0195} /* (2, 3, 21) {real, imag} */,
  {32'hc0ea4bf8, 32'h4191a97e} /* (2, 3, 20) {real, imag} */,
  {32'hbff28ede, 32'h40e0d55c} /* (2, 3, 19) {real, imag} */,
  {32'h4045b7aa, 32'hbf67d948} /* (2, 3, 18) {real, imag} */,
  {32'h412d34a8, 32'hc10ebe38} /* (2, 3, 17) {real, imag} */,
  {32'hc0aea740, 32'hc0cd155c} /* (2, 3, 16) {real, imag} */,
  {32'h40a5ce7a, 32'hc14bbb35} /* (2, 3, 15) {real, imag} */,
  {32'h40fbec9c, 32'h41a23d2e} /* (2, 3, 14) {real, imag} */,
  {32'h3d119280, 32'h40e4f9c9} /* (2, 3, 13) {real, imag} */,
  {32'h4190bf80, 32'hc0abe3f5} /* (2, 3, 12) {real, imag} */,
  {32'hc034dfe4, 32'hc15f0747} /* (2, 3, 11) {real, imag} */,
  {32'h419c9116, 32'h41480c61} /* (2, 3, 10) {real, imag} */,
  {32'h4004f7df, 32'hbdd59fc0} /* (2, 3, 9) {real, imag} */,
  {32'hc023ce2b, 32'h417aed6a} /* (2, 3, 8) {real, imag} */,
  {32'h41835836, 32'hc1716260} /* (2, 3, 7) {real, imag} */,
  {32'hc1b8addb, 32'h40597af5} /* (2, 3, 6) {real, imag} */,
  {32'hc1dbc29f, 32'h42152930} /* (2, 3, 5) {real, imag} */,
  {32'h41e42d9d, 32'h4147f2b6} /* (2, 3, 4) {real, imag} */,
  {32'hc24c7612, 32'hc20b7d8f} /* (2, 3, 3) {real, imag} */,
  {32'hc18db9a5, 32'h43161d4e} /* (2, 3, 2) {real, imag} */,
  {32'hc2b82e10, 32'hc207d672} /* (2, 3, 1) {real, imag} */,
  {32'h420173f0, 32'hc1fa2460} /* (2, 3, 0) {real, imag} */,
  {32'h4434eca6, 32'h428fcaa9} /* (2, 2, 31) {real, imag} */,
  {32'hc3b249c6, 32'h429af864} /* (2, 2, 30) {real, imag} */,
  {32'h424ee380, 32'h41d3104c} /* (2, 2, 29) {real, imag} */,
  {32'h424eb7cb, 32'hc23cfc89} /* (2, 2, 28) {real, imag} */,
  {32'hc206e118, 32'h425cccc6} /* (2, 2, 27) {real, imag} */,
  {32'h408bec05, 32'hc13cc014} /* (2, 2, 26) {real, imag} */,
  {32'h40ba5829, 32'hc1217e15} /* (2, 2, 25) {real, imag} */,
  {32'hc226c5cf, 32'h41fa9ce7} /* (2, 2, 24) {real, imag} */,
  {32'hc122e60a, 32'hc1001244} /* (2, 2, 23) {real, imag} */,
  {32'hc109b59e, 32'hc1a3d72c} /* (2, 2, 22) {real, imag} */,
  {32'hc0c6ffd5, 32'h41c55133} /* (2, 2, 21) {real, imag} */,
  {32'h40fe08b0, 32'h406e65f0} /* (2, 2, 20) {real, imag} */,
  {32'hc0d6a184, 32'h403b0f18} /* (2, 2, 19) {real, imag} */,
  {32'hc11f2aeb, 32'h3f887d60} /* (2, 2, 18) {real, imag} */,
  {32'h40766859, 32'hc1199c0a} /* (2, 2, 17) {real, imag} */,
  {32'hc01b6993, 32'hc13e64ba} /* (2, 2, 16) {real, imag} */,
  {32'hc05e694b, 32'hc129fd95} /* (2, 2, 15) {real, imag} */,
  {32'hbf61e188, 32'hc16e348c} /* (2, 2, 14) {real, imag} */,
  {32'h40df7c14, 32'hbeb7d33c} /* (2, 2, 13) {real, imag} */,
  {32'h40e155bc, 32'h418125af} /* (2, 2, 12) {real, imag} */,
  {32'hbf7416b0, 32'hc11a876e} /* (2, 2, 11) {real, imag} */,
  {32'h41e2c600, 32'h41d51546} /* (2, 2, 10) {real, imag} */,
  {32'h400c895c, 32'h40ba4594} /* (2, 2, 9) {real, imag} */,
  {32'hc1eabcf3, 32'h41475f89} /* (2, 2, 8) {real, imag} */,
  {32'hbdca1c60, 32'h40b19e9c} /* (2, 2, 7) {real, imag} */,
  {32'hc1a3c7fa, 32'hc16df2fa} /* (2, 2, 6) {real, imag} */,
  {32'hc245dc90, 32'hc23a7fcf} /* (2, 2, 5) {real, imag} */,
  {32'h42cdc345, 32'h41d35bdc} /* (2, 2, 4) {real, imag} */,
  {32'hc20ddc1e, 32'hc1f3b55d} /* (2, 2, 3) {real, imag} */,
  {32'hc37f12ef, 32'h43188f98} /* (2, 2, 2) {real, imag} */,
  {32'h43b44612, 32'hc0bd3590} /* (2, 2, 1) {real, imag} */,
  {32'h43a2e7b4, 32'h42da7243} /* (2, 2, 0) {real, imag} */,
  {32'hc41f114e, 32'h42d8475e} /* (2, 1, 31) {real, imag} */,
  {32'h4376d04c, 32'h4200fcee} /* (2, 1, 30) {real, imag} */,
  {32'h424721b1, 32'hc222b064} /* (2, 1, 29) {real, imag} */,
  {32'hc2bafd8c, 32'hc23203bd} /* (2, 1, 28) {real, imag} */,
  {32'h4304ef9c, 32'hc05fabef} /* (2, 1, 27) {real, imag} */,
  {32'h4217b59e, 32'hc17a58a0} /* (2, 1, 26) {real, imag} */,
  {32'hc018bdc8, 32'h40b9249a} /* (2, 1, 25) {real, imag} */,
  {32'h41e5e12a, 32'hc0c913ce} /* (2, 1, 24) {real, imag} */,
  {32'h40c952ea, 32'hc09471c9} /* (2, 1, 23) {real, imag} */,
  {32'hc14762d8, 32'h411302f3} /* (2, 1, 22) {real, imag} */,
  {32'h4218df18, 32'hc172fb38} /* (2, 1, 21) {real, imag} */,
  {32'hc0656644, 32'h4180bf32} /* (2, 1, 20) {real, imag} */,
  {32'hc140ea95, 32'hc1228405} /* (2, 1, 19) {real, imag} */,
  {32'hc0da80d5, 32'hc09335a7} /* (2, 1, 18) {real, imag} */,
  {32'hc04c8e17, 32'hc14be896} /* (2, 1, 17) {real, imag} */,
  {32'hc1123ff8, 32'h4076a105} /* (2, 1, 16) {real, imag} */,
  {32'h4021b65a, 32'hc097137f} /* (2, 1, 15) {real, imag} */,
  {32'hbfd2ac05, 32'h4107a08e} /* (2, 1, 14) {real, imag} */,
  {32'hc01c7f60, 32'hc178d327} /* (2, 1, 13) {real, imag} */,
  {32'h417b333c, 32'hbfedfbac} /* (2, 1, 12) {real, imag} */,
  {32'h4174ad1b, 32'h414c2a32} /* (2, 1, 11) {real, imag} */,
  {32'h415a6014, 32'hc08ffaf9} /* (2, 1, 10) {real, imag} */,
  {32'hc0421ad4, 32'hc0526afe} /* (2, 1, 9) {real, imag} */,
  {32'h41b34014, 32'h41e84d50} /* (2, 1, 8) {real, imag} */,
  {32'hc0d8990b, 32'hc1bc837d} /* (2, 1, 7) {real, imag} */,
  {32'hc004efc0, 32'h3ea8db40} /* (2, 1, 6) {real, imag} */,
  {32'h42529f59, 32'h425bb22c} /* (2, 1, 5) {real, imag} */,
  {32'hc1422e86, 32'hc1fc6dd4} /* (2, 1, 4) {real, imag} */,
  {32'h425fb448, 32'hc1a572b7} /* (2, 1, 3) {real, imag} */,
  {32'h43a3d54f, 32'h4388fcd8} /* (2, 1, 2) {real, imag} */,
  {32'hc46907cd, 32'hc413725e} /* (2, 1, 1) {real, imag} */,
  {32'hc3ff6ad2, 32'h426409e0} /* (2, 1, 0) {real, imag} */,
  {32'hc3dcc43f, 32'h438dbc6d} /* (2, 0, 31) {real, imag} */,
  {32'h4244186a, 32'hc2d9a97f} /* (2, 0, 30) {real, imag} */,
  {32'h425e9dc8, 32'hc23f6985} /* (2, 0, 29) {real, imag} */,
  {32'hc1c31f38, 32'hc2a140fc} /* (2, 0, 28) {real, imag} */,
  {32'h42495d5a, 32'hc17539ec} /* (2, 0, 27) {real, imag} */,
  {32'hc0ad891a, 32'h41a2a445} /* (2, 0, 26) {real, imag} */,
  {32'hbf8dd2e0, 32'h42015abd} /* (2, 0, 25) {real, imag} */,
  {32'h41b504e8, 32'hc198807d} /* (2, 0, 24) {real, imag} */,
  {32'h40c7f683, 32'hc0944859} /* (2, 0, 23) {real, imag} */,
  {32'h4182a5e5, 32'hc16cd5ec} /* (2, 0, 22) {real, imag} */,
  {32'h4114ceee, 32'hc19d0e7c} /* (2, 0, 21) {real, imag} */,
  {32'hc0236602, 32'h3fce0100} /* (2, 0, 20) {real, imag} */,
  {32'h4086c8c0, 32'h41017cc7} /* (2, 0, 19) {real, imag} */,
  {32'hc0d9c974, 32'hc036fda0} /* (2, 0, 18) {real, imag} */,
  {32'h4104ae48, 32'hc0b609ac} /* (2, 0, 17) {real, imag} */,
  {32'hbf8dcba4, 32'h00000000} /* (2, 0, 16) {real, imag} */,
  {32'h4104ae48, 32'h40b609ac} /* (2, 0, 15) {real, imag} */,
  {32'hc0d9c974, 32'h4036fda0} /* (2, 0, 14) {real, imag} */,
  {32'h4086c8c0, 32'hc1017cc7} /* (2, 0, 13) {real, imag} */,
  {32'hc0236602, 32'hbfce0100} /* (2, 0, 12) {real, imag} */,
  {32'h4114ceee, 32'h419d0e7c} /* (2, 0, 11) {real, imag} */,
  {32'h4182a5e5, 32'h416cd5ec} /* (2, 0, 10) {real, imag} */,
  {32'h40c7f683, 32'h40944859} /* (2, 0, 9) {real, imag} */,
  {32'h41b504e8, 32'h4198807d} /* (2, 0, 8) {real, imag} */,
  {32'hbf8dd2e0, 32'hc2015abd} /* (2, 0, 7) {real, imag} */,
  {32'hc0ad891a, 32'hc1a2a445} /* (2, 0, 6) {real, imag} */,
  {32'h42495d5a, 32'h417539ec} /* (2, 0, 5) {real, imag} */,
  {32'hc1c31f38, 32'h42a140fc} /* (2, 0, 4) {real, imag} */,
  {32'h425e9dc8, 32'h423f6985} /* (2, 0, 3) {real, imag} */,
  {32'h4244186a, 32'h42d9a97f} /* (2, 0, 2) {real, imag} */,
  {32'hc3dcc43f, 32'hc38dbc6d} /* (2, 0, 1) {real, imag} */,
  {32'hc2e389c6, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc4406709, 32'h43fa5546} /* (1, 31, 31) {real, imag} */,
  {32'h438ca72a, 32'hc367a1a0} /* (1, 31, 30) {real, imag} */,
  {32'h4272a66d, 32'hc0b6f578} /* (1, 31, 29) {real, imag} */,
  {32'h413ed3af, 32'h42288e11} /* (1, 31, 28) {real, imag} */,
  {32'h4271ea94, 32'hc213293c} /* (1, 31, 27) {real, imag} */,
  {32'h4132f384, 32'hc14ff0a1} /* (1, 31, 26) {real, imag} */,
  {32'hc166e3e4, 32'h42016cbe} /* (1, 31, 25) {real, imag} */,
  {32'h41678477, 32'hc169f1c1} /* (1, 31, 24) {real, imag} */,
  {32'hc0ee5500, 32'hc1c2b294} /* (1, 31, 23) {real, imag} */,
  {32'hc0fa3e6b, 32'h414d8960} /* (1, 31, 22) {real, imag} */,
  {32'hc10a07af, 32'hc075b93a} /* (1, 31, 21) {real, imag} */,
  {32'h4119a388, 32'h40985f5d} /* (1, 31, 20) {real, imag} */,
  {32'hc13885de, 32'hbfda0810} /* (1, 31, 19) {real, imag} */,
  {32'hc0ccf26a, 32'hc148672d} /* (1, 31, 18) {real, imag} */,
  {32'h40fbf15b, 32'h407bf001} /* (1, 31, 17) {real, imag} */,
  {32'hbdc65be0, 32'hbf9acad8} /* (1, 31, 16) {real, imag} */,
  {32'hc02598f4, 32'hc08488f5} /* (1, 31, 15) {real, imag} */,
  {32'hbf404404, 32'h3f829cc4} /* (1, 31, 14) {real, imag} */,
  {32'h40306312, 32'hbe08d180} /* (1, 31, 13) {real, imag} */,
  {32'hc0215bc4, 32'h40955167} /* (1, 31, 12) {real, imag} */,
  {32'h418e4ef0, 32'h41876ade} /* (1, 31, 11) {real, imag} */,
  {32'hc13c61bc, 32'h3feceea2} /* (1, 31, 10) {real, imag} */,
  {32'hc089ee3c, 32'h41af7294} /* (1, 31, 9) {real, imag} */,
  {32'h420fce5a, 32'h41c885b3} /* (1, 31, 8) {real, imag} */,
  {32'hc1abf0db, 32'h403b6654} /* (1, 31, 7) {real, imag} */,
  {32'h411ffd6c, 32'h41025ed4} /* (1, 31, 6) {real, imag} */,
  {32'h42edde0b, 32'h407a27d4} /* (1, 31, 5) {real, imag} */,
  {32'hc2a9ed83, 32'h41957882} /* (1, 31, 4) {real, imag} */,
  {32'h41db8bbf, 32'h41948293} /* (1, 31, 3) {real, imag} */,
  {32'h4330976e, 32'h4177ed99} /* (1, 31, 2) {real, imag} */,
  {32'hc403a91f, 32'hc26c4749} /* (1, 31, 1) {real, imag} */,
  {32'hc3f707f3, 32'hc2852fc4} /* (1, 31, 0) {real, imag} */,
  {32'h43820a3a, 32'hc04c3680} /* (1, 30, 31) {real, imag} */,
  {32'hc35ea3d9, 32'hc2e01cae} /* (1, 30, 30) {real, imag} */,
  {32'hbfb14b08, 32'h4221752f} /* (1, 30, 29) {real, imag} */,
  {32'h42d9c255, 32'hc1814f84} /* (1, 30, 28) {real, imag} */,
  {32'hc2343e4e, 32'h4216daa0} /* (1, 30, 27) {real, imag} */,
  {32'hc044de90, 32'hc0d4c3b8} /* (1, 30, 26) {real, imag} */,
  {32'h40fc76e6, 32'hc1c89424} /* (1, 30, 25) {real, imag} */,
  {32'hc230dda9, 32'h41d0ae8d} /* (1, 30, 24) {real, imag} */,
  {32'h408f55cc, 32'h40bd88ce} /* (1, 30, 23) {real, imag} */,
  {32'hbfbafe7c, 32'h402bc9de} /* (1, 30, 22) {real, imag} */,
  {32'hc1058d7c, 32'h418e832c} /* (1, 30, 21) {real, imag} */,
  {32'hc0be1710, 32'hc0ed7e51} /* (1, 30, 20) {real, imag} */,
  {32'h3e83dd34, 32'h3f1152d4} /* (1, 30, 19) {real, imag} */,
  {32'h41129baf, 32'h40a5698b} /* (1, 30, 18) {real, imag} */,
  {32'hbf1697ac, 32'hc032f798} /* (1, 30, 17) {real, imag} */,
  {32'hc04f1f28, 32'hc0963c10} /* (1, 30, 16) {real, imag} */,
  {32'h3ecc8e70, 32'h40880d63} /* (1, 30, 15) {real, imag} */,
  {32'hc0f2bc28, 32'h409c15e1} /* (1, 30, 14) {real, imag} */,
  {32'hc08ebab4, 32'h418e5fca} /* (1, 30, 13) {real, imag} */,
  {32'h405ab3fc, 32'hbf8af4f2} /* (1, 30, 12) {real, imag} */,
  {32'hc0d58bcb, 32'hc11e36ee} /* (1, 30, 11) {real, imag} */,
  {32'hc01d6ec2, 32'h41a495f4} /* (1, 30, 10) {real, imag} */,
  {32'hc11d502c, 32'hbf3fbcd8} /* (1, 30, 9) {real, imag} */,
  {32'hc204197a, 32'hc20f10a5} /* (1, 30, 8) {real, imag} */,
  {32'hbd877180, 32'h411fc5a6} /* (1, 30, 7) {real, imag} */,
  {32'h40d584f0, 32'h3f85f77c} /* (1, 30, 6) {real, imag} */,
  {32'hc20dfeb2, 32'hc258bd12} /* (1, 30, 5) {real, imag} */,
  {32'h422ede74, 32'h4190ddc8} /* (1, 30, 4) {real, imag} */,
  {32'h41eac239, 32'h41b057f4} /* (1, 30, 3) {real, imag} */,
  {32'hc3941f88, 32'hc1a755ad} /* (1, 30, 2) {real, imag} */,
  {32'h440f74bf, 32'hc27a5ecc} /* (1, 30, 1) {real, imag} */,
  {32'h437e832c, 32'hc2909d07} /* (1, 30, 0) {real, imag} */,
  {32'hc26040ab, 32'h4230f71b} /* (1, 29, 31) {real, imag} */,
  {32'hc16d933c, 32'hc3010ee2} /* (1, 29, 30) {real, imag} */,
  {32'hbf0ea8a0, 32'h42576169} /* (1, 29, 29) {real, imag} */,
  {32'h41cf4536, 32'hc1f6624c} /* (1, 29, 28) {real, imag} */,
  {32'hc20aa5ba, 32'hc1cc3352} /* (1, 29, 27) {real, imag} */,
  {32'hc1ec64a1, 32'h40e43823} /* (1, 29, 26) {real, imag} */,
  {32'hc137f387, 32'h41096234} /* (1, 29, 25) {real, imag} */,
  {32'hc1c80f7f, 32'hc0eac2d3} /* (1, 29, 24) {real, imag} */,
  {32'h412f9e06, 32'h40e396cd} /* (1, 29, 23) {real, imag} */,
  {32'h4171946d, 32'h408d1c7c} /* (1, 29, 22) {real, imag} */,
  {32'h3f3590bc, 32'hc083afda} /* (1, 29, 21) {real, imag} */,
  {32'h4203e9a2, 32'hc106bbfa} /* (1, 29, 20) {real, imag} */,
  {32'hbfcc04a8, 32'h3f839dfa} /* (1, 29, 19) {real, imag} */,
  {32'h40d17a24, 32'hbea00a20} /* (1, 29, 18) {real, imag} */,
  {32'hc0762f1f, 32'h40a5abd8} /* (1, 29, 17) {real, imag} */,
  {32'hc0a8feef, 32'h40a3aef1} /* (1, 29, 16) {real, imag} */,
  {32'h40ab0b36, 32'h40df740f} /* (1, 29, 15) {real, imag} */,
  {32'hc10159bf, 32'h40bb8e81} /* (1, 29, 14) {real, imag} */,
  {32'hc11d04f2, 32'h3d347c80} /* (1, 29, 13) {real, imag} */,
  {32'hc058362d, 32'h40e7449f} /* (1, 29, 12) {real, imag} */,
  {32'h40938120, 32'hbfeea84c} /* (1, 29, 11) {real, imag} */,
  {32'h402c2f60, 32'hc0ccea51} /* (1, 29, 10) {real, imag} */,
  {32'hc004dfec, 32'h40441726} /* (1, 29, 9) {real, imag} */,
  {32'h40a56d94, 32'hc1d6d76b} /* (1, 29, 8) {real, imag} */,
  {32'hc0e10c0c, 32'h3fdf7c08} /* (1, 29, 7) {real, imag} */,
  {32'hc16d045e, 32'h40b81de8} /* (1, 29, 6) {real, imag} */,
  {32'h418a60e2, 32'hc0c8ee59} /* (1, 29, 5) {real, imag} */,
  {32'hc1bd8d26, 32'h40e1d365} /* (1, 29, 4) {real, imag} */,
  {32'h407eba0c, 32'hc0e25ee6} /* (1, 29, 3) {real, imag} */,
  {32'hc23d3fcd, 32'hc29f93e2} /* (1, 29, 2) {real, imag} */,
  {32'h42f1bf5d, 32'h4266f6e8} /* (1, 29, 1) {real, imag} */,
  {32'h4203a094, 32'h40819160} /* (1, 29, 0) {real, imag} */,
  {32'hc30950b2, 32'h4188f442} /* (1, 28, 31) {real, imag} */,
  {32'h42795d7a, 32'hc2cce668} /* (1, 28, 30) {real, imag} */,
  {32'hc09bed98, 32'hc1e0093c} /* (1, 28, 29) {real, imag} */,
  {32'hc0c37dfe, 32'h407eace4} /* (1, 28, 28) {real, imag} */,
  {32'h415e9a6a, 32'h40efd804} /* (1, 28, 27) {real, imag} */,
  {32'h4122613e, 32'h410287ca} /* (1, 28, 26) {real, imag} */,
  {32'hc047fb76, 32'h41c1493c} /* (1, 28, 25) {real, imag} */,
  {32'h411a62b5, 32'hc14ed2bc} /* (1, 28, 24) {real, imag} */,
  {32'h41957666, 32'h404939f8} /* (1, 28, 23) {real, imag} */,
  {32'h418bf991, 32'h413d8b50} /* (1, 28, 22) {real, imag} */,
  {32'h4142196a, 32'hc1c1e220} /* (1, 28, 21) {real, imag} */,
  {32'h3f13d7b0, 32'h417c6572} /* (1, 28, 20) {real, imag} */,
  {32'hc02c4d18, 32'hc03d7285} /* (1, 28, 19) {real, imag} */,
  {32'hc13f8ab7, 32'hc1048f24} /* (1, 28, 18) {real, imag} */,
  {32'h40c19fd7, 32'h40eb5ae4} /* (1, 28, 17) {real, imag} */,
  {32'hbf97e2d1, 32'hc00ae2d4} /* (1, 28, 16) {real, imag} */,
  {32'hbff24d82, 32'h410b8125} /* (1, 28, 15) {real, imag} */,
  {32'h40664002, 32'hc0ba67af} /* (1, 28, 14) {real, imag} */,
  {32'hc0860f2a, 32'hc138a946} /* (1, 28, 13) {real, imag} */,
  {32'h3e3b6dc0, 32'hc163625f} /* (1, 28, 12) {real, imag} */,
  {32'h40caad7f, 32'hbf18db48} /* (1, 28, 11) {real, imag} */,
  {32'hc0f1c418, 32'h40c049ac} /* (1, 28, 10) {real, imag} */,
  {32'hc128a5ea, 32'h3f9d3c5e} /* (1, 28, 9) {real, imag} */,
  {32'hc0b0c3f8, 32'hc0d19bf0} /* (1, 28, 8) {real, imag} */,
  {32'hc15a273c, 32'h40e93c79} /* (1, 28, 7) {real, imag} */,
  {32'h413ffdc7, 32'h4164533c} /* (1, 28, 6) {real, imag} */,
  {32'h4186b53a, 32'h410bf7db} /* (1, 28, 5) {real, imag} */,
  {32'hc1c79f2d, 32'h4110a672} /* (1, 28, 4) {real, imag} */,
  {32'hc1a0dca4, 32'h41e57670} /* (1, 28, 3) {real, imag} */,
  {32'h4236463c, 32'hc2aa9da4} /* (1, 28, 2) {real, imag} */,
  {32'hc2815b13, 32'h4203face} /* (1, 28, 1) {real, imag} */,
  {32'hc0f36c28, 32'h416c282c} /* (1, 28, 0) {real, imag} */,
  {32'h4214f23c, 32'hc2998b9e} /* (1, 27, 31) {real, imag} */,
  {32'h41507e1a, 32'h419984ec} /* (1, 27, 30) {real, imag} */,
  {32'hc1282c4a, 32'h4133fcdf} /* (1, 27, 29) {real, imag} */,
  {32'hc03a54a4, 32'hc0f3e479} /* (1, 27, 28) {real, imag} */,
  {32'hc1af9810, 32'h41dca75e} /* (1, 27, 27) {real, imag} */,
  {32'hc0450b38, 32'h3fbaa5f8} /* (1, 27, 26) {real, imag} */,
  {32'h4103a914, 32'hc1a28b1a} /* (1, 27, 25) {real, imag} */,
  {32'hc123b4e2, 32'hc08c542b} /* (1, 27, 24) {real, imag} */,
  {32'h40b97122, 32'hc106fcf1} /* (1, 27, 23) {real, imag} */,
  {32'hc06429e1, 32'h40c20fee} /* (1, 27, 22) {real, imag} */,
  {32'hc05cc620, 32'h4047cae0} /* (1, 27, 21) {real, imag} */,
  {32'hc0ace988, 32'hc09df586} /* (1, 27, 20) {real, imag} */,
  {32'h41d46830, 32'hc115de7e} /* (1, 27, 19) {real, imag} */,
  {32'hc013eb5b, 32'hc02ba0ec} /* (1, 27, 18) {real, imag} */,
  {32'hc0991f49, 32'h405d1643} /* (1, 27, 17) {real, imag} */,
  {32'hc0d7aec0, 32'hc0cd419e} /* (1, 27, 16) {real, imag} */,
  {32'hc0fe8df4, 32'h3f3b0b80} /* (1, 27, 15) {real, imag} */,
  {32'h40ac25ed, 32'hc1a9d7fd} /* (1, 27, 14) {real, imag} */,
  {32'h41258f90, 32'hc00d1d31} /* (1, 27, 13) {real, imag} */,
  {32'h4159a23e, 32'h41adbab0} /* (1, 27, 12) {real, imag} */,
  {32'hbff4e636, 32'h40af373e} /* (1, 27, 11) {real, imag} */,
  {32'hc16f3ca9, 32'h405b2a3c} /* (1, 27, 10) {real, imag} */,
  {32'h40667237, 32'h40c235e6} /* (1, 27, 9) {real, imag} */,
  {32'h4160eb45, 32'h40a859c1} /* (1, 27, 8) {real, imag} */,
  {32'hc14a9a49, 32'hc04ac330} /* (1, 27, 7) {real, imag} */,
  {32'hc109540c, 32'h408659a0} /* (1, 27, 6) {real, imag} */,
  {32'h4094e870, 32'hc0f08b84} /* (1, 27, 5) {real, imag} */,
  {32'h40d00b12, 32'hc077c8c4} /* (1, 27, 4) {real, imag} */,
  {32'hc19c3c64, 32'hc17e0336} /* (1, 27, 3) {real, imag} */,
  {32'hc25200b2, 32'h40da0a54} /* (1, 27, 2) {real, imag} */,
  {32'h42ba7a75, 32'hc0a63c01} /* (1, 27, 1) {real, imag} */,
  {32'h4269f865, 32'hc1e2d3fc} /* (1, 27, 0) {real, imag} */,
  {32'hc0eb1d73, 32'hc178f41f} /* (1, 26, 31) {real, imag} */,
  {32'hbf93083a, 32'h415ae54e} /* (1, 26, 30) {real, imag} */,
  {32'hc092ce66, 32'h408a7b99} /* (1, 26, 29) {real, imag} */,
  {32'h413b8db3, 32'h40bf7a34} /* (1, 26, 28) {real, imag} */,
  {32'hc0ecd2ec, 32'hc0850018} /* (1, 26, 27) {real, imag} */,
  {32'hc12f52bc, 32'h412eacde} /* (1, 26, 26) {real, imag} */,
  {32'h418ed710, 32'h4169b823} /* (1, 26, 25) {real, imag} */,
  {32'h40cfa023, 32'h409d5f82} /* (1, 26, 24) {real, imag} */,
  {32'h413633a2, 32'hc1b7881c} /* (1, 26, 23) {real, imag} */,
  {32'h40d56ef7, 32'h409f2bea} /* (1, 26, 22) {real, imag} */,
  {32'hc0f10ea5, 32'h41971586} /* (1, 26, 21) {real, imag} */,
  {32'h3ff04aa6, 32'hbe8ce738} /* (1, 26, 20) {real, imag} */,
  {32'hc1498a73, 32'h40de144f} /* (1, 26, 19) {real, imag} */,
  {32'hbfcc8d94, 32'hc068828c} /* (1, 26, 18) {real, imag} */,
  {32'hc1072f8b, 32'h405f33f3} /* (1, 26, 17) {real, imag} */,
  {32'h40072552, 32'h3fd4d534} /* (1, 26, 16) {real, imag} */,
  {32'h40a85ce6, 32'h40c94e18} /* (1, 26, 15) {real, imag} */,
  {32'h3bf60f00, 32'h3ed447c0} /* (1, 26, 14) {real, imag} */,
  {32'h3fc664c8, 32'h412d85a8} /* (1, 26, 13) {real, imag} */,
  {32'h400c5642, 32'h3fa782f4} /* (1, 26, 12) {real, imag} */,
  {32'hc1540b4a, 32'h3f8ce6bc} /* (1, 26, 11) {real, imag} */,
  {32'h4083d81e, 32'h408a2866} /* (1, 26, 10) {real, imag} */,
  {32'hc18ffe2d, 32'hc1814d38} /* (1, 26, 9) {real, imag} */,
  {32'h3fee86fe, 32'hc072c71c} /* (1, 26, 8) {real, imag} */,
  {32'h40c3a154, 32'h3fc21e1b} /* (1, 26, 7) {real, imag} */,
  {32'h414bbdc4, 32'hc149a774} /* (1, 26, 6) {real, imag} */,
  {32'h41b4d0f1, 32'h41f2a08a} /* (1, 26, 5) {real, imag} */,
  {32'hc16fda0e, 32'h40e1da77} /* (1, 26, 4) {real, imag} */,
  {32'h4130fbe8, 32'h411f8ea8} /* (1, 26, 3) {real, imag} */,
  {32'hc1c789eb, 32'hc12017b4} /* (1, 26, 2) {real, imag} */,
  {32'hc144f184, 32'hc21b40b0} /* (1, 26, 1) {real, imag} */,
  {32'h418e5d0a, 32'h41e36aa2} /* (1, 26, 0) {real, imag} */,
  {32'h41d1151a, 32'h41a77e1e} /* (1, 25, 31) {real, imag} */,
  {32'hc1898137, 32'h41501e73} /* (1, 25, 30) {real, imag} */,
  {32'hc00dc441, 32'hc005942c} /* (1, 25, 29) {real, imag} */,
  {32'hc0217e03, 32'h408ebd06} /* (1, 25, 28) {real, imag} */,
  {32'hbf0f3640, 32'hc11815ef} /* (1, 25, 27) {real, imag} */,
  {32'hc1939ba1, 32'hc194fb68} /* (1, 25, 26) {real, imag} */,
  {32'hc140ddf4, 32'hc119bf2a} /* (1, 25, 25) {real, imag} */,
  {32'h409f2ec5, 32'hc06935d6} /* (1, 25, 24) {real, imag} */,
  {32'h41a2f6a7, 32'hc08d7394} /* (1, 25, 23) {real, imag} */,
  {32'h3e901f30, 32'hc17c68e1} /* (1, 25, 22) {real, imag} */,
  {32'h3fa2fd10, 32'hc130e3ca} /* (1, 25, 21) {real, imag} */,
  {32'hc09b811c, 32'h4196de2e} /* (1, 25, 20) {real, imag} */,
  {32'h3f8da13a, 32'hc127c5aa} /* (1, 25, 19) {real, imag} */,
  {32'h411d5ff9, 32'hc04141d7} /* (1, 25, 18) {real, imag} */,
  {32'h4093ccde, 32'h40c9dbf3} /* (1, 25, 17) {real, imag} */,
  {32'h3fc3da76, 32'hc1107443} /* (1, 25, 16) {real, imag} */,
  {32'h3ff91e88, 32'hc12f13bb} /* (1, 25, 15) {real, imag} */,
  {32'hc0ba4bcd, 32'hbf86f212} /* (1, 25, 14) {real, imag} */,
  {32'h3ef99620, 32'h409bcc8e} /* (1, 25, 13) {real, imag} */,
  {32'h402a86cc, 32'hc151c43b} /* (1, 25, 12) {real, imag} */,
  {32'hc10bd851, 32'hc124799c} /* (1, 25, 11) {real, imag} */,
  {32'hc0ad12c5, 32'hc0214859} /* (1, 25, 10) {real, imag} */,
  {32'hc0ff30e0, 32'hc1858c34} /* (1, 25, 9) {real, imag} */,
  {32'h418c6722, 32'h41904206} /* (1, 25, 8) {real, imag} */,
  {32'h41527864, 32'hc0ae0394} /* (1, 25, 7) {real, imag} */,
  {32'h4173035a, 32'hc0a18678} /* (1, 25, 6) {real, imag} */,
  {32'h40acac73, 32'h414a0fa9} /* (1, 25, 5) {real, imag} */,
  {32'hc198e080, 32'hc1f1ff0b} /* (1, 25, 4) {real, imag} */,
  {32'hc004dc1e, 32'h41050fda} /* (1, 25, 3) {real, imag} */,
  {32'h41201c43, 32'h40806194} /* (1, 25, 2) {real, imag} */,
  {32'hc1403e15, 32'hc12c4c32} /* (1, 25, 1) {real, imag} */,
  {32'h40824878, 32'h41438335} /* (1, 25, 0) {real, imag} */,
  {32'h419cd2fe, 32'hc1c01539} /* (1, 24, 31) {real, imag} */,
  {32'h40e13ea0, 32'hbfe8a410} /* (1, 24, 30) {real, imag} */,
  {32'hbfd17810, 32'hc0f00332} /* (1, 24, 29) {real, imag} */,
  {32'hc15b42a8, 32'hc1791a5c} /* (1, 24, 28) {real, imag} */,
  {32'hbc803180, 32'h4219c8b8} /* (1, 24, 27) {real, imag} */,
  {32'hc106b9b5, 32'h40913d61} /* (1, 24, 26) {real, imag} */,
  {32'h3fbb497f, 32'hc12d7771} /* (1, 24, 25) {real, imag} */,
  {32'h4096c6ec, 32'h418f1c30} /* (1, 24, 24) {real, imag} */,
  {32'h418db74a, 32'hc13ae5c8} /* (1, 24, 23) {real, imag} */,
  {32'h3df16b40, 32'hc1cd9fa6} /* (1, 24, 22) {real, imag} */,
  {32'h419fb2e6, 32'h410c34c1} /* (1, 24, 21) {real, imag} */,
  {32'hc09d7f00, 32'h418003a6} /* (1, 24, 20) {real, imag} */,
  {32'hc1476b29, 32'h417f3d72} /* (1, 24, 19) {real, imag} */,
  {32'h40bcf9d0, 32'h40bdc29b} /* (1, 24, 18) {real, imag} */,
  {32'h41160138, 32'hbf93f65a} /* (1, 24, 17) {real, imag} */,
  {32'hc12c6ca6, 32'hbec16e00} /* (1, 24, 16) {real, imag} */,
  {32'h409d2dd6, 32'hbfc24678} /* (1, 24, 15) {real, imag} */,
  {32'h408cc3fa, 32'hc0a0d0de} /* (1, 24, 14) {real, imag} */,
  {32'hc0e085cb, 32'h4197b956} /* (1, 24, 13) {real, imag} */,
  {32'hc15e279d, 32'hc13590d4} /* (1, 24, 12) {real, imag} */,
  {32'hbff68dac, 32'hc071b8b4} /* (1, 24, 11) {real, imag} */,
  {32'hc186bce8, 32'h41406f47} /* (1, 24, 10) {real, imag} */,
  {32'h41cb5f18, 32'hc09d946a} /* (1, 24, 9) {real, imag} */,
  {32'hc0bb3142, 32'hc1aaee09} /* (1, 24, 8) {real, imag} */,
  {32'h420aba94, 32'hc07d6eb3} /* (1, 24, 7) {real, imag} */,
  {32'hc02d3904, 32'hc15929c0} /* (1, 24, 6) {real, imag} */,
  {32'hbfcdf8dc, 32'hc10ff2a9} /* (1, 24, 5) {real, imag} */,
  {32'hc0886cff, 32'hc0c5847c} /* (1, 24, 4) {real, imag} */,
  {32'hc044f1d9, 32'h409179f8} /* (1, 24, 3) {real, imag} */,
  {32'hc2529dcf, 32'hc0cb78a6} /* (1, 24, 2) {real, imag} */,
  {32'h41f11a69, 32'hc1674c57} /* (1, 24, 1) {real, imag} */,
  {32'h413d11e8, 32'hc1e03a32} /* (1, 24, 0) {real, imag} */,
  {32'hc10e552b, 32'h40352514} /* (1, 23, 31) {real, imag} */,
  {32'h414125ce, 32'hc153bd05} /* (1, 23, 30) {real, imag} */,
  {32'hc13b5cc7, 32'hc1564c92} /* (1, 23, 29) {real, imag} */,
  {32'h41568702, 32'h41487c8b} /* (1, 23, 28) {real, imag} */,
  {32'hbf727446, 32'hbf82ba00} /* (1, 23, 27) {real, imag} */,
  {32'hc0eab588, 32'h412f42f8} /* (1, 23, 26) {real, imag} */,
  {32'hc066a554, 32'hc033650c} /* (1, 23, 25) {real, imag} */,
  {32'hc06bf525, 32'hbfe850dc} /* (1, 23, 24) {real, imag} */,
  {32'h4123a31c, 32'h3f1b3600} /* (1, 23, 23) {real, imag} */,
  {32'hc0f25d7b, 32'h3eb173b0} /* (1, 23, 22) {real, imag} */,
  {32'hc188f3f8, 32'h40dabfc4} /* (1, 23, 21) {real, imag} */,
  {32'h40a77d6e, 32'h40b9f892} /* (1, 23, 20) {real, imag} */,
  {32'h410361fd, 32'hc137fa8a} /* (1, 23, 19) {real, imag} */,
  {32'hc1071240, 32'h41d4cd14} /* (1, 23, 18) {real, imag} */,
  {32'hc0babfc1, 32'h40443745} /* (1, 23, 17) {real, imag} */,
  {32'h4137ba78, 32'hc17e5414} /* (1, 23, 16) {real, imag} */,
  {32'h41202ca9, 32'h40caf2c9} /* (1, 23, 15) {real, imag} */,
  {32'h41be3707, 32'hc0f5d65e} /* (1, 23, 14) {real, imag} */,
  {32'hc0de9e70, 32'hc06ec3e7} /* (1, 23, 13) {real, imag} */,
  {32'h403bc618, 32'h41b530d8} /* (1, 23, 12) {real, imag} */,
  {32'h40859c0c, 32'h3e55aaf0} /* (1, 23, 11) {real, imag} */,
  {32'h3f7499f0, 32'hc1283ca4} /* (1, 23, 10) {real, imag} */,
  {32'h4096b32a, 32'h40f27178} /* (1, 23, 9) {real, imag} */,
  {32'hbfe9bc28, 32'h411b5c50} /* (1, 23, 8) {real, imag} */,
  {32'hc129d2a1, 32'hc033779c} /* (1, 23, 7) {real, imag} */,
  {32'h4135482e, 32'h41684416} /* (1, 23, 6) {real, imag} */,
  {32'hc108f268, 32'h3fe878b4} /* (1, 23, 5) {real, imag} */,
  {32'hc08fa4fa, 32'h415b21b0} /* (1, 23, 4) {real, imag} */,
  {32'hc19aaf46, 32'h4163bcd9} /* (1, 23, 3) {real, imag} */,
  {32'h41244570, 32'hc1b205d8} /* (1, 23, 2) {real, imag} */,
  {32'h4062b852, 32'h40113358} /* (1, 23, 1) {real, imag} */,
  {32'hc18a8538, 32'h4092a964} /* (1, 23, 0) {real, imag} */,
  {32'h4124812f, 32'h40a20dbf} /* (1, 22, 31) {real, imag} */,
  {32'h4185fbdb, 32'hc1c09c35} /* (1, 22, 30) {real, imag} */,
  {32'h41abeed9, 32'h4074c832} /* (1, 22, 29) {real, imag} */,
  {32'h41388261, 32'hc01e7290} /* (1, 22, 28) {real, imag} */,
  {32'hc1370d5d, 32'h40bb5a28} /* (1, 22, 27) {real, imag} */,
  {32'hbfcc6432, 32'h412cfd34} /* (1, 22, 26) {real, imag} */,
  {32'h411007c5, 32'hbfd77bb0} /* (1, 22, 25) {real, imag} */,
  {32'hc106cf96, 32'h40635627} /* (1, 22, 24) {real, imag} */,
  {32'h41d539bd, 32'hbfc19654} /* (1, 22, 23) {real, imag} */,
  {32'h40e6bda4, 32'h3f319d40} /* (1, 22, 22) {real, imag} */,
  {32'hc0174a9a, 32'hc112cf26} /* (1, 22, 21) {real, imag} */,
  {32'hc17039fe, 32'h3fe73fb8} /* (1, 22, 20) {real, imag} */,
  {32'h40c7dd2e, 32'hc0afccbd} /* (1, 22, 19) {real, imag} */,
  {32'hc10a1818, 32'h41361ec6} /* (1, 22, 18) {real, imag} */,
  {32'hbfefd5d6, 32'hc0d69edb} /* (1, 22, 17) {real, imag} */,
  {32'h3ef39c9c, 32'hbe657490} /* (1, 22, 16) {real, imag} */,
  {32'h40c1586e, 32'h3fab7cf1} /* (1, 22, 15) {real, imag} */,
  {32'h3e40de80, 32'h3e588c80} /* (1, 22, 14) {real, imag} */,
  {32'h4114d66d, 32'hc0dc6843} /* (1, 22, 13) {real, imag} */,
  {32'hc06d2d71, 32'h4112f8aa} /* (1, 22, 12) {real, imag} */,
  {32'hc1a299eb, 32'hbfeabe00} /* (1, 22, 11) {real, imag} */,
  {32'h4037e58a, 32'hc1070906} /* (1, 22, 10) {real, imag} */,
  {32'h40b19b6c, 32'h410c05bb} /* (1, 22, 9) {real, imag} */,
  {32'h41938efc, 32'hc17740eb} /* (1, 22, 8) {real, imag} */,
  {32'hc1656ea3, 32'hbe780170} /* (1, 22, 7) {real, imag} */,
  {32'hc06c8cce, 32'hc06cba56} /* (1, 22, 6) {real, imag} */,
  {32'hc0da165a, 32'hc0b01014} /* (1, 22, 5) {real, imag} */,
  {32'hc098bc94, 32'h41bffd7a} /* (1, 22, 4) {real, imag} */,
  {32'hc14099ad, 32'h3f8339dc} /* (1, 22, 3) {real, imag} */,
  {32'hc0c42deb, 32'hc18f3aab} /* (1, 22, 2) {real, imag} */,
  {32'hc0a16149, 32'h418bf583} /* (1, 22, 1) {real, imag} */,
  {32'hc096715b, 32'h40740b1b} /* (1, 22, 0) {real, imag} */,
  {32'h4116c5a9, 32'hc1c648ba} /* (1, 21, 31) {real, imag} */,
  {32'h3ea38630, 32'h4107bf42} /* (1, 21, 30) {real, imag} */,
  {32'hc0f573c7, 32'h40e54a0e} /* (1, 21, 29) {real, imag} */,
  {32'h40a159ee, 32'h412d5863} /* (1, 21, 28) {real, imag} */,
  {32'hc184e76e, 32'h4054e9f2} /* (1, 21, 27) {real, imag} */,
  {32'h41361936, 32'h40cd924a} /* (1, 21, 26) {real, imag} */,
  {32'hc0374810, 32'h41555ec7} /* (1, 21, 25) {real, imag} */,
  {32'hc0925c6d, 32'hc0d715ce} /* (1, 21, 24) {real, imag} */,
  {32'hc0bab9c7, 32'h41192834} /* (1, 21, 23) {real, imag} */,
  {32'hc1a1cfdc, 32'h40a5002c} /* (1, 21, 22) {real, imag} */,
  {32'hc1d5a5ba, 32'h41570f54} /* (1, 21, 21) {real, imag} */,
  {32'hc0889dd6, 32'hc02dd05c} /* (1, 21, 20) {real, imag} */,
  {32'h40b69232, 32'h407f284b} /* (1, 21, 19) {real, imag} */,
  {32'hc09e9db6, 32'hc0bef119} /* (1, 21, 18) {real, imag} */,
  {32'hc0882d6a, 32'hbfbe56e0} /* (1, 21, 17) {real, imag} */,
  {32'h4109c370, 32'hc0220bdc} /* (1, 21, 16) {real, imag} */,
  {32'h41269198, 32'hbfdc752e} /* (1, 21, 15) {real, imag} */,
  {32'hc071b51a, 32'hbfc39730} /* (1, 21, 14) {real, imag} */,
  {32'hc091bad0, 32'h416fd6a0} /* (1, 21, 13) {real, imag} */,
  {32'hc1bf550b, 32'hc19f608a} /* (1, 21, 12) {real, imag} */,
  {32'h40bf6a4e, 32'h401f6de8} /* (1, 21, 11) {real, imag} */,
  {32'h4074b7d0, 32'hc14b9166} /* (1, 21, 10) {real, imag} */,
  {32'h41a0f686, 32'h41e4d2bc} /* (1, 21, 9) {real, imag} */,
  {32'h401c4ec0, 32'h3fca48ec} /* (1, 21, 8) {real, imag} */,
  {32'hc0d94781, 32'hc0ad65be} /* (1, 21, 7) {real, imag} */,
  {32'h416688b1, 32'hc0bb41a2} /* (1, 21, 6) {real, imag} */,
  {32'h3fa0cf58, 32'h41262851} /* (1, 21, 5) {real, imag} */,
  {32'h406b047d, 32'hc04eeba6} /* (1, 21, 4) {real, imag} */,
  {32'hc129e59b, 32'hc03d3033} /* (1, 21, 3) {real, imag} */,
  {32'h40091694, 32'h4202ebab} /* (1, 21, 2) {real, imag} */,
  {32'h417d130a, 32'hc168a13c} /* (1, 21, 1) {real, imag} */,
  {32'h4106cab6, 32'hbe4904c0} /* (1, 21, 0) {real, imag} */,
  {32'h415afe84, 32'h3fa78650} /* (1, 20, 31) {real, imag} */,
  {32'h40284aac, 32'h40b40a9f} /* (1, 20, 30) {real, imag} */,
  {32'hc0d596ab, 32'h40606392} /* (1, 20, 29) {real, imag} */,
  {32'h4127c00e, 32'h411d6d54} /* (1, 20, 28) {real, imag} */,
  {32'h4154e110, 32'h3d3b1200} /* (1, 20, 27) {real, imag} */,
  {32'h411ea700, 32'hbfa59c4c} /* (1, 20, 26) {real, imag} */,
  {32'hc185950c, 32'hc135006d} /* (1, 20, 25) {real, imag} */,
  {32'h4166a2ab, 32'h40a997a6} /* (1, 20, 24) {real, imag} */,
  {32'hbfdd60de, 32'hc1807a08} /* (1, 20, 23) {real, imag} */,
  {32'hc10c87b4, 32'h418a885e} /* (1, 20, 22) {real, imag} */,
  {32'h40201b1c, 32'hc0d9f333} /* (1, 20, 21) {real, imag} */,
  {32'hc134c4c5, 32'hc0a8c624} /* (1, 20, 20) {real, imag} */,
  {32'hc0a6bb34, 32'hbff504d3} /* (1, 20, 19) {real, imag} */,
  {32'h403c29ca, 32'hc1317393} /* (1, 20, 18) {real, imag} */,
  {32'h404c12c5, 32'hc0738f18} /* (1, 20, 17) {real, imag} */,
  {32'hc0f647b9, 32'h4146b940} /* (1, 20, 16) {real, imag} */,
  {32'hc0dc62fa, 32'hc0f995c8} /* (1, 20, 15) {real, imag} */,
  {32'h3f8aa540, 32'hc09df7e2} /* (1, 20, 14) {real, imag} */,
  {32'h40a31b11, 32'hc0bd6a6e} /* (1, 20, 13) {real, imag} */,
  {32'h413542f0, 32'hc1835dbf} /* (1, 20, 12) {real, imag} */,
  {32'hc118bac0, 32'hc1a98280} /* (1, 20, 11) {real, imag} */,
  {32'h41428a1a, 32'hc1aa89dc} /* (1, 20, 10) {real, imag} */,
  {32'h41153e57, 32'hc1773b13} /* (1, 20, 9) {real, imag} */,
  {32'hbe0c2fb0, 32'hbff305ec} /* (1, 20, 8) {real, imag} */,
  {32'h3ff80acc, 32'hbf445540} /* (1, 20, 7) {real, imag} */,
  {32'hbfdd55ae, 32'h418abd73} /* (1, 20, 6) {real, imag} */,
  {32'h4106f25d, 32'hc18b4dc0} /* (1, 20, 5) {real, imag} */,
  {32'hc0e2cd9b, 32'hc0c0ab02} /* (1, 20, 4) {real, imag} */,
  {32'hc0779448, 32'h414215a5} /* (1, 20, 3) {real, imag} */,
  {32'h41345048, 32'h410616d7} /* (1, 20, 2) {real, imag} */,
  {32'h4012b59a, 32'h4114729c} /* (1, 20, 1) {real, imag} */,
  {32'hbf762a40, 32'h414ad71e} /* (1, 20, 0) {real, imag} */,
  {32'hc0256825, 32'h41457fcc} /* (1, 19, 31) {real, imag} */,
  {32'h40becfec, 32'h400ac2fe} /* (1, 19, 30) {real, imag} */,
  {32'h3fe35e22, 32'h40b0e12a} /* (1, 19, 29) {real, imag} */,
  {32'hc1852c0b, 32'hbfd91d9e} /* (1, 19, 28) {real, imag} */,
  {32'hc0eaf962, 32'hc13e858a} /* (1, 19, 27) {real, imag} */,
  {32'hc144c908, 32'hc110ede7} /* (1, 19, 26) {real, imag} */,
  {32'hc0618e2d, 32'hc09dbc97} /* (1, 19, 25) {real, imag} */,
  {32'h3eb2db10, 32'h418073a7} /* (1, 19, 24) {real, imag} */,
  {32'h402ae28d, 32'hc1620a86} /* (1, 19, 23) {real, imag} */,
  {32'hc0a8e52d, 32'h3e89a218} /* (1, 19, 22) {real, imag} */,
  {32'h4141f3f6, 32'hc163ccfa} /* (1, 19, 21) {real, imag} */,
  {32'h3e97a974, 32'hbfd52c1f} /* (1, 19, 20) {real, imag} */,
  {32'h40abd1b6, 32'h40db6b62} /* (1, 19, 19) {real, imag} */,
  {32'hc015c139, 32'h407400e2} /* (1, 19, 18) {real, imag} */,
  {32'hc11ac91c, 32'h4101b6fa} /* (1, 19, 17) {real, imag} */,
  {32'h413ecef7, 32'h40d4aed0} /* (1, 19, 16) {real, imag} */,
  {32'h406b8420, 32'h407ba3c8} /* (1, 19, 15) {real, imag} */,
  {32'hc10aedc6, 32'h409f5051} /* (1, 19, 14) {real, imag} */,
  {32'hc07c8c1a, 32'h41420d1a} /* (1, 19, 13) {real, imag} */,
  {32'hc136a9cb, 32'hbffb5eb0} /* (1, 19, 12) {real, imag} */,
  {32'hc1104d76, 32'hc1474363} /* (1, 19, 11) {real, imag} */,
  {32'hc05cff03, 32'hc13d1363} /* (1, 19, 10) {real, imag} */,
  {32'h401c4b86, 32'h411dd876} /* (1, 19, 9) {real, imag} */,
  {32'h40fb1dbe, 32'hc12bd69a} /* (1, 19, 8) {real, imag} */,
  {32'hc032b49e, 32'hc13fe009} /* (1, 19, 7) {real, imag} */,
  {32'hbfa948a0, 32'h418028ad} /* (1, 19, 6) {real, imag} */,
  {32'h3fdbf183, 32'h3e1e4700} /* (1, 19, 5) {real, imag} */,
  {32'h4176cac0, 32'hc03ae56e} /* (1, 19, 4) {real, imag} */,
  {32'h40a27013, 32'hc00257f2} /* (1, 19, 3) {real, imag} */,
  {32'hc0e7591d, 32'hc0815fc4} /* (1, 19, 2) {real, imag} */,
  {32'h4106d454, 32'h418d5f76} /* (1, 19, 1) {real, imag} */,
  {32'h41299211, 32'h40950007} /* (1, 19, 0) {real, imag} */,
  {32'hc18f97df, 32'h40e67e3d} /* (1, 18, 31) {real, imag} */,
  {32'hc16690a8, 32'h40ae223c} /* (1, 18, 30) {real, imag} */,
  {32'h3dc72880, 32'hbf4b7c58} /* (1, 18, 29) {real, imag} */,
  {32'hc09df35c, 32'h40a8c910} /* (1, 18, 28) {real, imag} */,
  {32'hc0786e2a, 32'hc15b119c} /* (1, 18, 27) {real, imag} */,
  {32'h40e5c6d6, 32'hc0d2d583} /* (1, 18, 26) {real, imag} */,
  {32'hc035ac44, 32'h411ee528} /* (1, 18, 25) {real, imag} */,
  {32'h3ff0232d, 32'h402566aa} /* (1, 18, 24) {real, imag} */,
  {32'hc0d8c643, 32'h4090ac9e} /* (1, 18, 23) {real, imag} */,
  {32'h3fa0aed8, 32'hc0ab6368} /* (1, 18, 22) {real, imag} */,
  {32'hbfa19912, 32'h4124a12c} /* (1, 18, 21) {real, imag} */,
  {32'h40b00b71, 32'hc1525cce} /* (1, 18, 20) {real, imag} */,
  {32'hc1144026, 32'hc1431138} /* (1, 18, 19) {real, imag} */,
  {32'hc0765832, 32'hc039e6c6} /* (1, 18, 18) {real, imag} */,
  {32'h4094daf7, 32'hc03bc36c} /* (1, 18, 17) {real, imag} */,
  {32'h403a4766, 32'hc120ffc0} /* (1, 18, 16) {real, imag} */,
  {32'hbe0951c0, 32'hc12df99c} /* (1, 18, 15) {real, imag} */,
  {32'h40aa6b18, 32'h4092061e} /* (1, 18, 14) {real, imag} */,
  {32'h419f58e6, 32'h3fcba22c} /* (1, 18, 13) {real, imag} */,
  {32'h41732082, 32'h40f2a4eb} /* (1, 18, 12) {real, imag} */,
  {32'h4096d8f8, 32'hc19a86a9} /* (1, 18, 11) {real, imag} */,
  {32'hbf754428, 32'h414bf014} /* (1, 18, 10) {real, imag} */,
  {32'h3f955c7a, 32'h4090c694} /* (1, 18, 9) {real, imag} */,
  {32'h409ac114, 32'h4153aa40} /* (1, 18, 8) {real, imag} */,
  {32'h3e4006b8, 32'hbe947c20} /* (1, 18, 7) {real, imag} */,
  {32'h40b2eef9, 32'h4135b28e} /* (1, 18, 6) {real, imag} */,
  {32'hc14b91d7, 32'hc025fd93} /* (1, 18, 5) {real, imag} */,
  {32'hbfcecebc, 32'hc1116f43} /* (1, 18, 4) {real, imag} */,
  {32'h41318c83, 32'h40598260} /* (1, 18, 3) {real, imag} */,
  {32'hc178c550, 32'h402b7dfa} /* (1, 18, 2) {real, imag} */,
  {32'hc08c637c, 32'hbf136354} /* (1, 18, 1) {real, imag} */,
  {32'hc11e9437, 32'hc0059c86} /* (1, 18, 0) {real, imag} */,
  {32'h404129f3, 32'h4089e56e} /* (1, 17, 31) {real, imag} */,
  {32'h407b83ca, 32'h40ad8ce6} /* (1, 17, 30) {real, imag} */,
  {32'hc0d283ff, 32'hc0a69da9} /* (1, 17, 29) {real, imag} */,
  {32'hc02634c0, 32'hc087a5ed} /* (1, 17, 28) {real, imag} */,
  {32'hc1227820, 32'hc08823f7} /* (1, 17, 27) {real, imag} */,
  {32'hc0ddb638, 32'hc10bf850} /* (1, 17, 26) {real, imag} */,
  {32'h40f0b512, 32'hc0aba8cb} /* (1, 17, 25) {real, imag} */,
  {32'hc149de7b, 32'h4181a7f1} /* (1, 17, 24) {real, imag} */,
  {32'h4007361d, 32'h411afada} /* (1, 17, 23) {real, imag} */,
  {32'hc14e02ef, 32'hbf816590} /* (1, 17, 22) {real, imag} */,
  {32'h40317e18, 32'hc0a044e7} /* (1, 17, 21) {real, imag} */,
  {32'hc0581d0c, 32'hc0f3f267} /* (1, 17, 20) {real, imag} */,
  {32'h40a4b0fe, 32'h405ede74} /* (1, 17, 19) {real, imag} */,
  {32'hc0ecbc98, 32'hc086c5cd} /* (1, 17, 18) {real, imag} */,
  {32'h4118434c, 32'hc122723f} /* (1, 17, 17) {real, imag} */,
  {32'hc0ddf71c, 32'hc11930ad} /* (1, 17, 16) {real, imag} */,
  {32'hbf9440e4, 32'h4080c11c} /* (1, 17, 15) {real, imag} */,
  {32'hc145c9b6, 32'h407a9cce} /* (1, 17, 14) {real, imag} */,
  {32'hc1306334, 32'h400f6439} /* (1, 17, 13) {real, imag} */,
  {32'h408308a0, 32'h400c5857} /* (1, 17, 12) {real, imag} */,
  {32'hbf530078, 32'hc08231cf} /* (1, 17, 11) {real, imag} */,
  {32'hc03ec784, 32'hc119aece} /* (1, 17, 10) {real, imag} */,
  {32'h400d98cc, 32'h3fce759c} /* (1, 17, 9) {real, imag} */,
  {32'h40885084, 32'h4118e121} /* (1, 17, 8) {real, imag} */,
  {32'h4107e19e, 32'hc100fbdb} /* (1, 17, 7) {real, imag} */,
  {32'hbf2b1038, 32'h3e42db98} /* (1, 17, 6) {real, imag} */,
  {32'hc0152254, 32'h41176b9a} /* (1, 17, 5) {real, imag} */,
  {32'hbf2e7550, 32'h40e85883} /* (1, 17, 4) {real, imag} */,
  {32'hc174daee, 32'h3e8dada0} /* (1, 17, 3) {real, imag} */,
  {32'hc1256c5c, 32'hc084fd1c} /* (1, 17, 2) {real, imag} */,
  {32'h40c666a1, 32'h4094f99a} /* (1, 17, 1) {real, imag} */,
  {32'hbfcf956a, 32'hc12610be} /* (1, 17, 0) {real, imag} */,
  {32'h4074f4c2, 32'hbfdca2f2} /* (1, 16, 31) {real, imag} */,
  {32'hc0c65f0b, 32'h40a49a73} /* (1, 16, 30) {real, imag} */,
  {32'h4005a698, 32'hc033b368} /* (1, 16, 29) {real, imag} */,
  {32'hbe25c220, 32'hc1108f80} /* (1, 16, 28) {real, imag} */,
  {32'hc157f5c4, 32'hc15d6793} /* (1, 16, 27) {real, imag} */,
  {32'hbfd4d36c, 32'h409957e2} /* (1, 16, 26) {real, imag} */,
  {32'hc113012e, 32'hc07b8668} /* (1, 16, 25) {real, imag} */,
  {32'h40eca209, 32'h4051bad0} /* (1, 16, 24) {real, imag} */,
  {32'hc152891f, 32'hbfdef902} /* (1, 16, 23) {real, imag} */,
  {32'h407bf7f8, 32'h4151d192} /* (1, 16, 22) {real, imag} */,
  {32'hc1219b42, 32'hc00f6abe} /* (1, 16, 21) {real, imag} */,
  {32'hc0bb12d1, 32'h40028016} /* (1, 16, 20) {real, imag} */,
  {32'hbfd8a67a, 32'hc00fd57f} /* (1, 16, 19) {real, imag} */,
  {32'h410d3d59, 32'h40669eae} /* (1, 16, 18) {real, imag} */,
  {32'hc04a72b2, 32'h40097635} /* (1, 16, 17) {real, imag} */,
  {32'h41982cc1, 32'h00000000} /* (1, 16, 16) {real, imag} */,
  {32'hc04a72b2, 32'hc0097635} /* (1, 16, 15) {real, imag} */,
  {32'h410d3d59, 32'hc0669eae} /* (1, 16, 14) {real, imag} */,
  {32'hbfd8a67a, 32'h400fd57f} /* (1, 16, 13) {real, imag} */,
  {32'hc0bb12d1, 32'hc0028016} /* (1, 16, 12) {real, imag} */,
  {32'hc1219b42, 32'h400f6abe} /* (1, 16, 11) {real, imag} */,
  {32'h407bf7f8, 32'hc151d192} /* (1, 16, 10) {real, imag} */,
  {32'hc152891f, 32'h3fdef902} /* (1, 16, 9) {real, imag} */,
  {32'h40eca209, 32'hc051bad0} /* (1, 16, 8) {real, imag} */,
  {32'hc113012e, 32'h407b8668} /* (1, 16, 7) {real, imag} */,
  {32'hbfd4d36c, 32'hc09957e2} /* (1, 16, 6) {real, imag} */,
  {32'hc157f5c4, 32'h415d6793} /* (1, 16, 5) {real, imag} */,
  {32'hbe25c220, 32'h41108f80} /* (1, 16, 4) {real, imag} */,
  {32'h4005a698, 32'h4033b368} /* (1, 16, 3) {real, imag} */,
  {32'hc0c65f0b, 32'hc0a49a73} /* (1, 16, 2) {real, imag} */,
  {32'h4074f4c2, 32'h3fdca2f2} /* (1, 16, 1) {real, imag} */,
  {32'h4020d4a0, 32'h00000000} /* (1, 16, 0) {real, imag} */,
  {32'h40c666a1, 32'hc094f99a} /* (1, 15, 31) {real, imag} */,
  {32'hc1256c5c, 32'h4084fd1c} /* (1, 15, 30) {real, imag} */,
  {32'hc174daee, 32'hbe8dada0} /* (1, 15, 29) {real, imag} */,
  {32'hbf2e7550, 32'hc0e85883} /* (1, 15, 28) {real, imag} */,
  {32'hc0152254, 32'hc1176b9a} /* (1, 15, 27) {real, imag} */,
  {32'hbf2b1038, 32'hbe42db98} /* (1, 15, 26) {real, imag} */,
  {32'h4107e19e, 32'h4100fbdb} /* (1, 15, 25) {real, imag} */,
  {32'h40885084, 32'hc118e121} /* (1, 15, 24) {real, imag} */,
  {32'h400d98cc, 32'hbfce759c} /* (1, 15, 23) {real, imag} */,
  {32'hc03ec784, 32'h4119aece} /* (1, 15, 22) {real, imag} */,
  {32'hbf530078, 32'h408231cf} /* (1, 15, 21) {real, imag} */,
  {32'h408308a0, 32'hc00c5857} /* (1, 15, 20) {real, imag} */,
  {32'hc1306334, 32'hc00f6439} /* (1, 15, 19) {real, imag} */,
  {32'hc145c9b6, 32'hc07a9cce} /* (1, 15, 18) {real, imag} */,
  {32'hbf9440e4, 32'hc080c11c} /* (1, 15, 17) {real, imag} */,
  {32'hc0ddf71c, 32'h411930ad} /* (1, 15, 16) {real, imag} */,
  {32'h4118434c, 32'h4122723f} /* (1, 15, 15) {real, imag} */,
  {32'hc0ecbc98, 32'h4086c5cd} /* (1, 15, 14) {real, imag} */,
  {32'h40a4b0fe, 32'hc05ede74} /* (1, 15, 13) {real, imag} */,
  {32'hc0581d0c, 32'h40f3f267} /* (1, 15, 12) {real, imag} */,
  {32'h40317e18, 32'h40a044e7} /* (1, 15, 11) {real, imag} */,
  {32'hc14e02ef, 32'h3f816590} /* (1, 15, 10) {real, imag} */,
  {32'h4007361d, 32'hc11afada} /* (1, 15, 9) {real, imag} */,
  {32'hc149de7b, 32'hc181a7f1} /* (1, 15, 8) {real, imag} */,
  {32'h40f0b512, 32'h40aba8cb} /* (1, 15, 7) {real, imag} */,
  {32'hc0ddb638, 32'h410bf850} /* (1, 15, 6) {real, imag} */,
  {32'hc1227820, 32'h408823f7} /* (1, 15, 5) {real, imag} */,
  {32'hc02634c0, 32'h4087a5ed} /* (1, 15, 4) {real, imag} */,
  {32'hc0d283ff, 32'h40a69da9} /* (1, 15, 3) {real, imag} */,
  {32'h407b83ca, 32'hc0ad8ce6} /* (1, 15, 2) {real, imag} */,
  {32'h404129f3, 32'hc089e56e} /* (1, 15, 1) {real, imag} */,
  {32'hbfcf956a, 32'h412610be} /* (1, 15, 0) {real, imag} */,
  {32'hc08c637c, 32'h3f136354} /* (1, 14, 31) {real, imag} */,
  {32'hc178c550, 32'hc02b7dfa} /* (1, 14, 30) {real, imag} */,
  {32'h41318c83, 32'hc0598260} /* (1, 14, 29) {real, imag} */,
  {32'hbfcecebc, 32'h41116f43} /* (1, 14, 28) {real, imag} */,
  {32'hc14b91d7, 32'h4025fd93} /* (1, 14, 27) {real, imag} */,
  {32'h40b2eef9, 32'hc135b28e} /* (1, 14, 26) {real, imag} */,
  {32'h3e4006b8, 32'h3e947c20} /* (1, 14, 25) {real, imag} */,
  {32'h409ac114, 32'hc153aa40} /* (1, 14, 24) {real, imag} */,
  {32'h3f955c7a, 32'hc090c694} /* (1, 14, 23) {real, imag} */,
  {32'hbf754428, 32'hc14bf014} /* (1, 14, 22) {real, imag} */,
  {32'h4096d8f8, 32'h419a86a9} /* (1, 14, 21) {real, imag} */,
  {32'h41732082, 32'hc0f2a4eb} /* (1, 14, 20) {real, imag} */,
  {32'h419f58e6, 32'hbfcba22c} /* (1, 14, 19) {real, imag} */,
  {32'h40aa6b18, 32'hc092061e} /* (1, 14, 18) {real, imag} */,
  {32'hbe0951c0, 32'h412df99c} /* (1, 14, 17) {real, imag} */,
  {32'h403a4766, 32'h4120ffc0} /* (1, 14, 16) {real, imag} */,
  {32'h4094daf7, 32'h403bc36c} /* (1, 14, 15) {real, imag} */,
  {32'hc0765832, 32'h4039e6c6} /* (1, 14, 14) {real, imag} */,
  {32'hc1144026, 32'h41431138} /* (1, 14, 13) {real, imag} */,
  {32'h40b00b71, 32'h41525cce} /* (1, 14, 12) {real, imag} */,
  {32'hbfa19912, 32'hc124a12c} /* (1, 14, 11) {real, imag} */,
  {32'h3fa0aed8, 32'h40ab6368} /* (1, 14, 10) {real, imag} */,
  {32'hc0d8c643, 32'hc090ac9e} /* (1, 14, 9) {real, imag} */,
  {32'h3ff0232d, 32'hc02566aa} /* (1, 14, 8) {real, imag} */,
  {32'hc035ac44, 32'hc11ee528} /* (1, 14, 7) {real, imag} */,
  {32'h40e5c6d6, 32'h40d2d583} /* (1, 14, 6) {real, imag} */,
  {32'hc0786e2a, 32'h415b119c} /* (1, 14, 5) {real, imag} */,
  {32'hc09df35c, 32'hc0a8c910} /* (1, 14, 4) {real, imag} */,
  {32'h3dc72880, 32'h3f4b7c58} /* (1, 14, 3) {real, imag} */,
  {32'hc16690a8, 32'hc0ae223c} /* (1, 14, 2) {real, imag} */,
  {32'hc18f97df, 32'hc0e67e3d} /* (1, 14, 1) {real, imag} */,
  {32'hc11e9437, 32'h40059c86} /* (1, 14, 0) {real, imag} */,
  {32'h4106d454, 32'hc18d5f76} /* (1, 13, 31) {real, imag} */,
  {32'hc0e7591d, 32'h40815fc4} /* (1, 13, 30) {real, imag} */,
  {32'h40a27013, 32'h400257f2} /* (1, 13, 29) {real, imag} */,
  {32'h4176cac0, 32'h403ae56e} /* (1, 13, 28) {real, imag} */,
  {32'h3fdbf183, 32'hbe1e4700} /* (1, 13, 27) {real, imag} */,
  {32'hbfa948a0, 32'hc18028ad} /* (1, 13, 26) {real, imag} */,
  {32'hc032b49e, 32'h413fe009} /* (1, 13, 25) {real, imag} */,
  {32'h40fb1dbe, 32'h412bd69a} /* (1, 13, 24) {real, imag} */,
  {32'h401c4b86, 32'hc11dd876} /* (1, 13, 23) {real, imag} */,
  {32'hc05cff03, 32'h413d1363} /* (1, 13, 22) {real, imag} */,
  {32'hc1104d76, 32'h41474363} /* (1, 13, 21) {real, imag} */,
  {32'hc136a9cb, 32'h3ffb5eb0} /* (1, 13, 20) {real, imag} */,
  {32'hc07c8c1a, 32'hc1420d1a} /* (1, 13, 19) {real, imag} */,
  {32'hc10aedc6, 32'hc09f5051} /* (1, 13, 18) {real, imag} */,
  {32'h406b8420, 32'hc07ba3c8} /* (1, 13, 17) {real, imag} */,
  {32'h413ecef7, 32'hc0d4aed0} /* (1, 13, 16) {real, imag} */,
  {32'hc11ac91c, 32'hc101b6fa} /* (1, 13, 15) {real, imag} */,
  {32'hc015c139, 32'hc07400e2} /* (1, 13, 14) {real, imag} */,
  {32'h40abd1b6, 32'hc0db6b62} /* (1, 13, 13) {real, imag} */,
  {32'h3e97a974, 32'h3fd52c1f} /* (1, 13, 12) {real, imag} */,
  {32'h4141f3f6, 32'h4163ccfa} /* (1, 13, 11) {real, imag} */,
  {32'hc0a8e52d, 32'hbe89a218} /* (1, 13, 10) {real, imag} */,
  {32'h402ae28d, 32'h41620a86} /* (1, 13, 9) {real, imag} */,
  {32'h3eb2db10, 32'hc18073a7} /* (1, 13, 8) {real, imag} */,
  {32'hc0618e2d, 32'h409dbc97} /* (1, 13, 7) {real, imag} */,
  {32'hc144c908, 32'h4110ede7} /* (1, 13, 6) {real, imag} */,
  {32'hc0eaf962, 32'h413e858a} /* (1, 13, 5) {real, imag} */,
  {32'hc1852c0b, 32'h3fd91d9e} /* (1, 13, 4) {real, imag} */,
  {32'h3fe35e22, 32'hc0b0e12a} /* (1, 13, 3) {real, imag} */,
  {32'h40becfec, 32'hc00ac2fe} /* (1, 13, 2) {real, imag} */,
  {32'hc0256825, 32'hc1457fcc} /* (1, 13, 1) {real, imag} */,
  {32'h41299211, 32'hc0950007} /* (1, 13, 0) {real, imag} */,
  {32'h4012b59a, 32'hc114729c} /* (1, 12, 31) {real, imag} */,
  {32'h41345048, 32'hc10616d7} /* (1, 12, 30) {real, imag} */,
  {32'hc0779448, 32'hc14215a5} /* (1, 12, 29) {real, imag} */,
  {32'hc0e2cd9b, 32'h40c0ab02} /* (1, 12, 28) {real, imag} */,
  {32'h4106f25d, 32'h418b4dc0} /* (1, 12, 27) {real, imag} */,
  {32'hbfdd55ae, 32'hc18abd73} /* (1, 12, 26) {real, imag} */,
  {32'h3ff80acc, 32'h3f445540} /* (1, 12, 25) {real, imag} */,
  {32'hbe0c2fb0, 32'h3ff305ec} /* (1, 12, 24) {real, imag} */,
  {32'h41153e57, 32'h41773b13} /* (1, 12, 23) {real, imag} */,
  {32'h41428a1a, 32'h41aa89dc} /* (1, 12, 22) {real, imag} */,
  {32'hc118bac0, 32'h41a98280} /* (1, 12, 21) {real, imag} */,
  {32'h413542f0, 32'h41835dbf} /* (1, 12, 20) {real, imag} */,
  {32'h40a31b11, 32'h40bd6a6e} /* (1, 12, 19) {real, imag} */,
  {32'h3f8aa540, 32'h409df7e2} /* (1, 12, 18) {real, imag} */,
  {32'hc0dc62fa, 32'h40f995c8} /* (1, 12, 17) {real, imag} */,
  {32'hc0f647b9, 32'hc146b940} /* (1, 12, 16) {real, imag} */,
  {32'h404c12c5, 32'h40738f18} /* (1, 12, 15) {real, imag} */,
  {32'h403c29ca, 32'h41317393} /* (1, 12, 14) {real, imag} */,
  {32'hc0a6bb34, 32'h3ff504d3} /* (1, 12, 13) {real, imag} */,
  {32'hc134c4c5, 32'h40a8c624} /* (1, 12, 12) {real, imag} */,
  {32'h40201b1c, 32'h40d9f333} /* (1, 12, 11) {real, imag} */,
  {32'hc10c87b4, 32'hc18a885e} /* (1, 12, 10) {real, imag} */,
  {32'hbfdd60de, 32'h41807a08} /* (1, 12, 9) {real, imag} */,
  {32'h4166a2ab, 32'hc0a997a6} /* (1, 12, 8) {real, imag} */,
  {32'hc185950c, 32'h4135006d} /* (1, 12, 7) {real, imag} */,
  {32'h411ea700, 32'h3fa59c4c} /* (1, 12, 6) {real, imag} */,
  {32'h4154e110, 32'hbd3b1200} /* (1, 12, 5) {real, imag} */,
  {32'h4127c00e, 32'hc11d6d54} /* (1, 12, 4) {real, imag} */,
  {32'hc0d596ab, 32'hc0606392} /* (1, 12, 3) {real, imag} */,
  {32'h40284aac, 32'hc0b40a9f} /* (1, 12, 2) {real, imag} */,
  {32'h415afe84, 32'hbfa78650} /* (1, 12, 1) {real, imag} */,
  {32'hbf762a40, 32'hc14ad71e} /* (1, 12, 0) {real, imag} */,
  {32'h417d130a, 32'h4168a13c} /* (1, 11, 31) {real, imag} */,
  {32'h40091694, 32'hc202ebab} /* (1, 11, 30) {real, imag} */,
  {32'hc129e59b, 32'h403d3033} /* (1, 11, 29) {real, imag} */,
  {32'h406b047d, 32'h404eeba6} /* (1, 11, 28) {real, imag} */,
  {32'h3fa0cf58, 32'hc1262851} /* (1, 11, 27) {real, imag} */,
  {32'h416688b1, 32'h40bb41a2} /* (1, 11, 26) {real, imag} */,
  {32'hc0d94781, 32'h40ad65be} /* (1, 11, 25) {real, imag} */,
  {32'h401c4ec0, 32'hbfca48ec} /* (1, 11, 24) {real, imag} */,
  {32'h41a0f686, 32'hc1e4d2bc} /* (1, 11, 23) {real, imag} */,
  {32'h4074b7d0, 32'h414b9166} /* (1, 11, 22) {real, imag} */,
  {32'h40bf6a4e, 32'hc01f6de8} /* (1, 11, 21) {real, imag} */,
  {32'hc1bf550b, 32'h419f608a} /* (1, 11, 20) {real, imag} */,
  {32'hc091bad0, 32'hc16fd6a0} /* (1, 11, 19) {real, imag} */,
  {32'hc071b51a, 32'h3fc39730} /* (1, 11, 18) {real, imag} */,
  {32'h41269198, 32'h3fdc752e} /* (1, 11, 17) {real, imag} */,
  {32'h4109c370, 32'h40220bdc} /* (1, 11, 16) {real, imag} */,
  {32'hc0882d6a, 32'h3fbe56e0} /* (1, 11, 15) {real, imag} */,
  {32'hc09e9db6, 32'h40bef119} /* (1, 11, 14) {real, imag} */,
  {32'h40b69232, 32'hc07f284b} /* (1, 11, 13) {real, imag} */,
  {32'hc0889dd6, 32'h402dd05c} /* (1, 11, 12) {real, imag} */,
  {32'hc1d5a5ba, 32'hc1570f54} /* (1, 11, 11) {real, imag} */,
  {32'hc1a1cfdc, 32'hc0a5002c} /* (1, 11, 10) {real, imag} */,
  {32'hc0bab9c7, 32'hc1192834} /* (1, 11, 9) {real, imag} */,
  {32'hc0925c6d, 32'h40d715ce} /* (1, 11, 8) {real, imag} */,
  {32'hc0374810, 32'hc1555ec7} /* (1, 11, 7) {real, imag} */,
  {32'h41361936, 32'hc0cd924a} /* (1, 11, 6) {real, imag} */,
  {32'hc184e76e, 32'hc054e9f2} /* (1, 11, 5) {real, imag} */,
  {32'h40a159ee, 32'hc12d5863} /* (1, 11, 4) {real, imag} */,
  {32'hc0f573c7, 32'hc0e54a0e} /* (1, 11, 3) {real, imag} */,
  {32'h3ea38630, 32'hc107bf42} /* (1, 11, 2) {real, imag} */,
  {32'h4116c5a9, 32'h41c648ba} /* (1, 11, 1) {real, imag} */,
  {32'h4106cab6, 32'h3e4904c0} /* (1, 11, 0) {real, imag} */,
  {32'hc0a16149, 32'hc18bf583} /* (1, 10, 31) {real, imag} */,
  {32'hc0c42deb, 32'h418f3aab} /* (1, 10, 30) {real, imag} */,
  {32'hc14099ad, 32'hbf8339dc} /* (1, 10, 29) {real, imag} */,
  {32'hc098bc94, 32'hc1bffd7a} /* (1, 10, 28) {real, imag} */,
  {32'hc0da165a, 32'h40b01014} /* (1, 10, 27) {real, imag} */,
  {32'hc06c8cce, 32'h406cba56} /* (1, 10, 26) {real, imag} */,
  {32'hc1656ea3, 32'h3e780170} /* (1, 10, 25) {real, imag} */,
  {32'h41938efc, 32'h417740eb} /* (1, 10, 24) {real, imag} */,
  {32'h40b19b6c, 32'hc10c05bb} /* (1, 10, 23) {real, imag} */,
  {32'h4037e58a, 32'h41070906} /* (1, 10, 22) {real, imag} */,
  {32'hc1a299eb, 32'h3feabe00} /* (1, 10, 21) {real, imag} */,
  {32'hc06d2d71, 32'hc112f8aa} /* (1, 10, 20) {real, imag} */,
  {32'h4114d66d, 32'h40dc6843} /* (1, 10, 19) {real, imag} */,
  {32'h3e40de80, 32'hbe588c80} /* (1, 10, 18) {real, imag} */,
  {32'h40c1586e, 32'hbfab7cf1} /* (1, 10, 17) {real, imag} */,
  {32'h3ef39c9c, 32'h3e657490} /* (1, 10, 16) {real, imag} */,
  {32'hbfefd5d6, 32'h40d69edb} /* (1, 10, 15) {real, imag} */,
  {32'hc10a1818, 32'hc1361ec6} /* (1, 10, 14) {real, imag} */,
  {32'h40c7dd2e, 32'h40afccbd} /* (1, 10, 13) {real, imag} */,
  {32'hc17039fe, 32'hbfe73fb8} /* (1, 10, 12) {real, imag} */,
  {32'hc0174a9a, 32'h4112cf26} /* (1, 10, 11) {real, imag} */,
  {32'h40e6bda4, 32'hbf319d40} /* (1, 10, 10) {real, imag} */,
  {32'h41d539bd, 32'h3fc19654} /* (1, 10, 9) {real, imag} */,
  {32'hc106cf96, 32'hc0635627} /* (1, 10, 8) {real, imag} */,
  {32'h411007c5, 32'h3fd77bb0} /* (1, 10, 7) {real, imag} */,
  {32'hbfcc6432, 32'hc12cfd34} /* (1, 10, 6) {real, imag} */,
  {32'hc1370d5d, 32'hc0bb5a28} /* (1, 10, 5) {real, imag} */,
  {32'h41388261, 32'h401e7290} /* (1, 10, 4) {real, imag} */,
  {32'h41abeed9, 32'hc074c832} /* (1, 10, 3) {real, imag} */,
  {32'h4185fbdb, 32'h41c09c35} /* (1, 10, 2) {real, imag} */,
  {32'h4124812f, 32'hc0a20dbf} /* (1, 10, 1) {real, imag} */,
  {32'hc096715b, 32'hc0740b1b} /* (1, 10, 0) {real, imag} */,
  {32'h4062b852, 32'hc0113358} /* (1, 9, 31) {real, imag} */,
  {32'h41244570, 32'h41b205d8} /* (1, 9, 30) {real, imag} */,
  {32'hc19aaf46, 32'hc163bcd9} /* (1, 9, 29) {real, imag} */,
  {32'hc08fa4fa, 32'hc15b21b0} /* (1, 9, 28) {real, imag} */,
  {32'hc108f268, 32'hbfe878b4} /* (1, 9, 27) {real, imag} */,
  {32'h4135482e, 32'hc1684416} /* (1, 9, 26) {real, imag} */,
  {32'hc129d2a1, 32'h4033779c} /* (1, 9, 25) {real, imag} */,
  {32'hbfe9bc28, 32'hc11b5c50} /* (1, 9, 24) {real, imag} */,
  {32'h4096b32a, 32'hc0f27178} /* (1, 9, 23) {real, imag} */,
  {32'h3f7499f0, 32'h41283ca4} /* (1, 9, 22) {real, imag} */,
  {32'h40859c0c, 32'hbe55aaf0} /* (1, 9, 21) {real, imag} */,
  {32'h403bc618, 32'hc1b530d8} /* (1, 9, 20) {real, imag} */,
  {32'hc0de9e70, 32'h406ec3e7} /* (1, 9, 19) {real, imag} */,
  {32'h41be3707, 32'h40f5d65e} /* (1, 9, 18) {real, imag} */,
  {32'h41202ca9, 32'hc0caf2c9} /* (1, 9, 17) {real, imag} */,
  {32'h4137ba78, 32'h417e5414} /* (1, 9, 16) {real, imag} */,
  {32'hc0babfc1, 32'hc0443745} /* (1, 9, 15) {real, imag} */,
  {32'hc1071240, 32'hc1d4cd14} /* (1, 9, 14) {real, imag} */,
  {32'h410361fd, 32'h4137fa8a} /* (1, 9, 13) {real, imag} */,
  {32'h40a77d6e, 32'hc0b9f892} /* (1, 9, 12) {real, imag} */,
  {32'hc188f3f8, 32'hc0dabfc4} /* (1, 9, 11) {real, imag} */,
  {32'hc0f25d7b, 32'hbeb173b0} /* (1, 9, 10) {real, imag} */,
  {32'h4123a31c, 32'hbf1b3600} /* (1, 9, 9) {real, imag} */,
  {32'hc06bf525, 32'h3fe850dc} /* (1, 9, 8) {real, imag} */,
  {32'hc066a554, 32'h4033650c} /* (1, 9, 7) {real, imag} */,
  {32'hc0eab588, 32'hc12f42f8} /* (1, 9, 6) {real, imag} */,
  {32'hbf727446, 32'h3f82ba00} /* (1, 9, 5) {real, imag} */,
  {32'h41568702, 32'hc1487c8b} /* (1, 9, 4) {real, imag} */,
  {32'hc13b5cc7, 32'h41564c92} /* (1, 9, 3) {real, imag} */,
  {32'h414125ce, 32'h4153bd05} /* (1, 9, 2) {real, imag} */,
  {32'hc10e552b, 32'hc0352514} /* (1, 9, 1) {real, imag} */,
  {32'hc18a8538, 32'hc092a964} /* (1, 9, 0) {real, imag} */,
  {32'h41f11a69, 32'h41674c57} /* (1, 8, 31) {real, imag} */,
  {32'hc2529dcf, 32'h40cb78a6} /* (1, 8, 30) {real, imag} */,
  {32'hc044f1d9, 32'hc09179f8} /* (1, 8, 29) {real, imag} */,
  {32'hc0886cff, 32'h40c5847c} /* (1, 8, 28) {real, imag} */,
  {32'hbfcdf8dc, 32'h410ff2a9} /* (1, 8, 27) {real, imag} */,
  {32'hc02d3904, 32'h415929c0} /* (1, 8, 26) {real, imag} */,
  {32'h420aba94, 32'h407d6eb3} /* (1, 8, 25) {real, imag} */,
  {32'hc0bb3142, 32'h41aaee09} /* (1, 8, 24) {real, imag} */,
  {32'h41cb5f18, 32'h409d946a} /* (1, 8, 23) {real, imag} */,
  {32'hc186bce8, 32'hc1406f47} /* (1, 8, 22) {real, imag} */,
  {32'hbff68dac, 32'h4071b8b4} /* (1, 8, 21) {real, imag} */,
  {32'hc15e279d, 32'h413590d4} /* (1, 8, 20) {real, imag} */,
  {32'hc0e085cb, 32'hc197b956} /* (1, 8, 19) {real, imag} */,
  {32'h408cc3fa, 32'h40a0d0de} /* (1, 8, 18) {real, imag} */,
  {32'h409d2dd6, 32'h3fc24678} /* (1, 8, 17) {real, imag} */,
  {32'hc12c6ca6, 32'h3ec16e00} /* (1, 8, 16) {real, imag} */,
  {32'h41160138, 32'h3f93f65a} /* (1, 8, 15) {real, imag} */,
  {32'h40bcf9d0, 32'hc0bdc29b} /* (1, 8, 14) {real, imag} */,
  {32'hc1476b29, 32'hc17f3d72} /* (1, 8, 13) {real, imag} */,
  {32'hc09d7f00, 32'hc18003a6} /* (1, 8, 12) {real, imag} */,
  {32'h419fb2e6, 32'hc10c34c1} /* (1, 8, 11) {real, imag} */,
  {32'h3df16b40, 32'h41cd9fa6} /* (1, 8, 10) {real, imag} */,
  {32'h418db74a, 32'h413ae5c8} /* (1, 8, 9) {real, imag} */,
  {32'h4096c6ec, 32'hc18f1c30} /* (1, 8, 8) {real, imag} */,
  {32'h3fbb497f, 32'h412d7771} /* (1, 8, 7) {real, imag} */,
  {32'hc106b9b5, 32'hc0913d61} /* (1, 8, 6) {real, imag} */,
  {32'hbc803180, 32'hc219c8b8} /* (1, 8, 5) {real, imag} */,
  {32'hc15b42a8, 32'h41791a5c} /* (1, 8, 4) {real, imag} */,
  {32'hbfd17810, 32'h40f00332} /* (1, 8, 3) {real, imag} */,
  {32'h40e13ea0, 32'h3fe8a410} /* (1, 8, 2) {real, imag} */,
  {32'h419cd2fe, 32'h41c01539} /* (1, 8, 1) {real, imag} */,
  {32'h413d11e8, 32'h41e03a32} /* (1, 8, 0) {real, imag} */,
  {32'hc1403e15, 32'h412c4c32} /* (1, 7, 31) {real, imag} */,
  {32'h41201c43, 32'hc0806194} /* (1, 7, 30) {real, imag} */,
  {32'hc004dc1e, 32'hc1050fda} /* (1, 7, 29) {real, imag} */,
  {32'hc198e080, 32'h41f1ff0b} /* (1, 7, 28) {real, imag} */,
  {32'h40acac73, 32'hc14a0fa9} /* (1, 7, 27) {real, imag} */,
  {32'h4173035a, 32'h40a18678} /* (1, 7, 26) {real, imag} */,
  {32'h41527864, 32'h40ae0394} /* (1, 7, 25) {real, imag} */,
  {32'h418c6722, 32'hc1904206} /* (1, 7, 24) {real, imag} */,
  {32'hc0ff30e0, 32'h41858c34} /* (1, 7, 23) {real, imag} */,
  {32'hc0ad12c5, 32'h40214859} /* (1, 7, 22) {real, imag} */,
  {32'hc10bd851, 32'h4124799c} /* (1, 7, 21) {real, imag} */,
  {32'h402a86cc, 32'h4151c43b} /* (1, 7, 20) {real, imag} */,
  {32'h3ef99620, 32'hc09bcc8e} /* (1, 7, 19) {real, imag} */,
  {32'hc0ba4bcd, 32'h3f86f212} /* (1, 7, 18) {real, imag} */,
  {32'h3ff91e88, 32'h412f13bb} /* (1, 7, 17) {real, imag} */,
  {32'h3fc3da76, 32'h41107443} /* (1, 7, 16) {real, imag} */,
  {32'h4093ccde, 32'hc0c9dbf3} /* (1, 7, 15) {real, imag} */,
  {32'h411d5ff9, 32'h404141d7} /* (1, 7, 14) {real, imag} */,
  {32'h3f8da13a, 32'h4127c5aa} /* (1, 7, 13) {real, imag} */,
  {32'hc09b811c, 32'hc196de2e} /* (1, 7, 12) {real, imag} */,
  {32'h3fa2fd10, 32'h4130e3ca} /* (1, 7, 11) {real, imag} */,
  {32'h3e901f30, 32'h417c68e1} /* (1, 7, 10) {real, imag} */,
  {32'h41a2f6a7, 32'h408d7394} /* (1, 7, 9) {real, imag} */,
  {32'h409f2ec5, 32'h406935d6} /* (1, 7, 8) {real, imag} */,
  {32'hc140ddf4, 32'h4119bf2a} /* (1, 7, 7) {real, imag} */,
  {32'hc1939ba1, 32'h4194fb68} /* (1, 7, 6) {real, imag} */,
  {32'hbf0f3640, 32'h411815ef} /* (1, 7, 5) {real, imag} */,
  {32'hc0217e03, 32'hc08ebd06} /* (1, 7, 4) {real, imag} */,
  {32'hc00dc441, 32'h4005942c} /* (1, 7, 3) {real, imag} */,
  {32'hc1898137, 32'hc1501e73} /* (1, 7, 2) {real, imag} */,
  {32'h41d1151a, 32'hc1a77e1e} /* (1, 7, 1) {real, imag} */,
  {32'h40824878, 32'hc1438335} /* (1, 7, 0) {real, imag} */,
  {32'hc144f184, 32'h421b40b0} /* (1, 6, 31) {real, imag} */,
  {32'hc1c789eb, 32'h412017b4} /* (1, 6, 30) {real, imag} */,
  {32'h4130fbe8, 32'hc11f8ea8} /* (1, 6, 29) {real, imag} */,
  {32'hc16fda0e, 32'hc0e1da77} /* (1, 6, 28) {real, imag} */,
  {32'h41b4d0f1, 32'hc1f2a08a} /* (1, 6, 27) {real, imag} */,
  {32'h414bbdc4, 32'h4149a774} /* (1, 6, 26) {real, imag} */,
  {32'h40c3a154, 32'hbfc21e1b} /* (1, 6, 25) {real, imag} */,
  {32'h3fee86fe, 32'h4072c71c} /* (1, 6, 24) {real, imag} */,
  {32'hc18ffe2d, 32'h41814d38} /* (1, 6, 23) {real, imag} */,
  {32'h4083d81e, 32'hc08a2866} /* (1, 6, 22) {real, imag} */,
  {32'hc1540b4a, 32'hbf8ce6bc} /* (1, 6, 21) {real, imag} */,
  {32'h400c5642, 32'hbfa782f4} /* (1, 6, 20) {real, imag} */,
  {32'h3fc664c8, 32'hc12d85a8} /* (1, 6, 19) {real, imag} */,
  {32'h3bf60f00, 32'hbed447c0} /* (1, 6, 18) {real, imag} */,
  {32'h40a85ce6, 32'hc0c94e18} /* (1, 6, 17) {real, imag} */,
  {32'h40072552, 32'hbfd4d534} /* (1, 6, 16) {real, imag} */,
  {32'hc1072f8b, 32'hc05f33f3} /* (1, 6, 15) {real, imag} */,
  {32'hbfcc8d94, 32'h4068828c} /* (1, 6, 14) {real, imag} */,
  {32'hc1498a73, 32'hc0de144f} /* (1, 6, 13) {real, imag} */,
  {32'h3ff04aa6, 32'h3e8ce738} /* (1, 6, 12) {real, imag} */,
  {32'hc0f10ea5, 32'hc1971586} /* (1, 6, 11) {real, imag} */,
  {32'h40d56ef7, 32'hc09f2bea} /* (1, 6, 10) {real, imag} */,
  {32'h413633a2, 32'h41b7881c} /* (1, 6, 9) {real, imag} */,
  {32'h40cfa023, 32'hc09d5f82} /* (1, 6, 8) {real, imag} */,
  {32'h418ed710, 32'hc169b823} /* (1, 6, 7) {real, imag} */,
  {32'hc12f52bc, 32'hc12eacde} /* (1, 6, 6) {real, imag} */,
  {32'hc0ecd2ec, 32'h40850018} /* (1, 6, 5) {real, imag} */,
  {32'h413b8db3, 32'hc0bf7a34} /* (1, 6, 4) {real, imag} */,
  {32'hc092ce66, 32'hc08a7b99} /* (1, 6, 3) {real, imag} */,
  {32'hbf93083a, 32'hc15ae54e} /* (1, 6, 2) {real, imag} */,
  {32'hc0eb1d73, 32'h4178f41f} /* (1, 6, 1) {real, imag} */,
  {32'h418e5d0a, 32'hc1e36aa2} /* (1, 6, 0) {real, imag} */,
  {32'h42ba7a75, 32'h40a63c01} /* (1, 5, 31) {real, imag} */,
  {32'hc25200b2, 32'hc0da0a54} /* (1, 5, 30) {real, imag} */,
  {32'hc19c3c64, 32'h417e0336} /* (1, 5, 29) {real, imag} */,
  {32'h40d00b12, 32'h4077c8c4} /* (1, 5, 28) {real, imag} */,
  {32'h4094e870, 32'h40f08b84} /* (1, 5, 27) {real, imag} */,
  {32'hc109540c, 32'hc08659a0} /* (1, 5, 26) {real, imag} */,
  {32'hc14a9a49, 32'h404ac330} /* (1, 5, 25) {real, imag} */,
  {32'h4160eb45, 32'hc0a859c1} /* (1, 5, 24) {real, imag} */,
  {32'h40667237, 32'hc0c235e6} /* (1, 5, 23) {real, imag} */,
  {32'hc16f3ca9, 32'hc05b2a3c} /* (1, 5, 22) {real, imag} */,
  {32'hbff4e636, 32'hc0af373e} /* (1, 5, 21) {real, imag} */,
  {32'h4159a23e, 32'hc1adbab0} /* (1, 5, 20) {real, imag} */,
  {32'h41258f90, 32'h400d1d31} /* (1, 5, 19) {real, imag} */,
  {32'h40ac25ed, 32'h41a9d7fd} /* (1, 5, 18) {real, imag} */,
  {32'hc0fe8df4, 32'hbf3b0b80} /* (1, 5, 17) {real, imag} */,
  {32'hc0d7aec0, 32'h40cd419e} /* (1, 5, 16) {real, imag} */,
  {32'hc0991f49, 32'hc05d1643} /* (1, 5, 15) {real, imag} */,
  {32'hc013eb5b, 32'h402ba0ec} /* (1, 5, 14) {real, imag} */,
  {32'h41d46830, 32'h4115de7e} /* (1, 5, 13) {real, imag} */,
  {32'hc0ace988, 32'h409df586} /* (1, 5, 12) {real, imag} */,
  {32'hc05cc620, 32'hc047cae0} /* (1, 5, 11) {real, imag} */,
  {32'hc06429e1, 32'hc0c20fee} /* (1, 5, 10) {real, imag} */,
  {32'h40b97122, 32'h4106fcf1} /* (1, 5, 9) {real, imag} */,
  {32'hc123b4e2, 32'h408c542b} /* (1, 5, 8) {real, imag} */,
  {32'h4103a914, 32'h41a28b1a} /* (1, 5, 7) {real, imag} */,
  {32'hc0450b38, 32'hbfbaa5f8} /* (1, 5, 6) {real, imag} */,
  {32'hc1af9810, 32'hc1dca75e} /* (1, 5, 5) {real, imag} */,
  {32'hc03a54a4, 32'h40f3e479} /* (1, 5, 4) {real, imag} */,
  {32'hc1282c4a, 32'hc133fcdf} /* (1, 5, 3) {real, imag} */,
  {32'h41507e1a, 32'hc19984ec} /* (1, 5, 2) {real, imag} */,
  {32'h4214f23c, 32'h42998b9e} /* (1, 5, 1) {real, imag} */,
  {32'h4269f865, 32'h41e2d3fc} /* (1, 5, 0) {real, imag} */,
  {32'hc2815b13, 32'hc203face} /* (1, 4, 31) {real, imag} */,
  {32'h4236463c, 32'h42aa9da4} /* (1, 4, 30) {real, imag} */,
  {32'hc1a0dca4, 32'hc1e57670} /* (1, 4, 29) {real, imag} */,
  {32'hc1c79f2d, 32'hc110a672} /* (1, 4, 28) {real, imag} */,
  {32'h4186b53a, 32'hc10bf7db} /* (1, 4, 27) {real, imag} */,
  {32'h413ffdc7, 32'hc164533c} /* (1, 4, 26) {real, imag} */,
  {32'hc15a273c, 32'hc0e93c79} /* (1, 4, 25) {real, imag} */,
  {32'hc0b0c3f8, 32'h40d19bf0} /* (1, 4, 24) {real, imag} */,
  {32'hc128a5ea, 32'hbf9d3c5e} /* (1, 4, 23) {real, imag} */,
  {32'hc0f1c418, 32'hc0c049ac} /* (1, 4, 22) {real, imag} */,
  {32'h40caad7f, 32'h3f18db48} /* (1, 4, 21) {real, imag} */,
  {32'h3e3b6dc0, 32'h4163625f} /* (1, 4, 20) {real, imag} */,
  {32'hc0860f2a, 32'h4138a946} /* (1, 4, 19) {real, imag} */,
  {32'h40664002, 32'h40ba67af} /* (1, 4, 18) {real, imag} */,
  {32'hbff24d82, 32'hc10b8125} /* (1, 4, 17) {real, imag} */,
  {32'hbf97e2d1, 32'h400ae2d4} /* (1, 4, 16) {real, imag} */,
  {32'h40c19fd7, 32'hc0eb5ae4} /* (1, 4, 15) {real, imag} */,
  {32'hc13f8ab7, 32'h41048f24} /* (1, 4, 14) {real, imag} */,
  {32'hc02c4d18, 32'h403d7285} /* (1, 4, 13) {real, imag} */,
  {32'h3f13d7b0, 32'hc17c6572} /* (1, 4, 12) {real, imag} */,
  {32'h4142196a, 32'h41c1e220} /* (1, 4, 11) {real, imag} */,
  {32'h418bf991, 32'hc13d8b50} /* (1, 4, 10) {real, imag} */,
  {32'h41957666, 32'hc04939f8} /* (1, 4, 9) {real, imag} */,
  {32'h411a62b5, 32'h414ed2bc} /* (1, 4, 8) {real, imag} */,
  {32'hc047fb76, 32'hc1c1493c} /* (1, 4, 7) {real, imag} */,
  {32'h4122613e, 32'hc10287ca} /* (1, 4, 6) {real, imag} */,
  {32'h415e9a6a, 32'hc0efd804} /* (1, 4, 5) {real, imag} */,
  {32'hc0c37dfe, 32'hc07eace4} /* (1, 4, 4) {real, imag} */,
  {32'hc09bed98, 32'h41e0093c} /* (1, 4, 3) {real, imag} */,
  {32'h42795d7a, 32'h42cce668} /* (1, 4, 2) {real, imag} */,
  {32'hc30950b2, 32'hc188f442} /* (1, 4, 1) {real, imag} */,
  {32'hc0f36c28, 32'hc16c282c} /* (1, 4, 0) {real, imag} */,
  {32'h42f1bf5d, 32'hc266f6e8} /* (1, 3, 31) {real, imag} */,
  {32'hc23d3fcd, 32'h429f93e2} /* (1, 3, 30) {real, imag} */,
  {32'h407eba0c, 32'h40e25ee6} /* (1, 3, 29) {real, imag} */,
  {32'hc1bd8d26, 32'hc0e1d365} /* (1, 3, 28) {real, imag} */,
  {32'h418a60e2, 32'h40c8ee59} /* (1, 3, 27) {real, imag} */,
  {32'hc16d045e, 32'hc0b81de8} /* (1, 3, 26) {real, imag} */,
  {32'hc0e10c0c, 32'hbfdf7c08} /* (1, 3, 25) {real, imag} */,
  {32'h40a56d94, 32'h41d6d76b} /* (1, 3, 24) {real, imag} */,
  {32'hc004dfec, 32'hc0441726} /* (1, 3, 23) {real, imag} */,
  {32'h402c2f60, 32'h40ccea51} /* (1, 3, 22) {real, imag} */,
  {32'h40938120, 32'h3feea84c} /* (1, 3, 21) {real, imag} */,
  {32'hc058362d, 32'hc0e7449f} /* (1, 3, 20) {real, imag} */,
  {32'hc11d04f2, 32'hbd347c80} /* (1, 3, 19) {real, imag} */,
  {32'hc10159bf, 32'hc0bb8e81} /* (1, 3, 18) {real, imag} */,
  {32'h40ab0b36, 32'hc0df740f} /* (1, 3, 17) {real, imag} */,
  {32'hc0a8feef, 32'hc0a3aef1} /* (1, 3, 16) {real, imag} */,
  {32'hc0762f1f, 32'hc0a5abd8} /* (1, 3, 15) {real, imag} */,
  {32'h40d17a24, 32'h3ea00a20} /* (1, 3, 14) {real, imag} */,
  {32'hbfcc04a8, 32'hbf839dfa} /* (1, 3, 13) {real, imag} */,
  {32'h4203e9a2, 32'h4106bbfa} /* (1, 3, 12) {real, imag} */,
  {32'h3f3590bc, 32'h4083afda} /* (1, 3, 11) {real, imag} */,
  {32'h4171946d, 32'hc08d1c7c} /* (1, 3, 10) {real, imag} */,
  {32'h412f9e06, 32'hc0e396cd} /* (1, 3, 9) {real, imag} */,
  {32'hc1c80f7f, 32'h40eac2d3} /* (1, 3, 8) {real, imag} */,
  {32'hc137f387, 32'hc1096234} /* (1, 3, 7) {real, imag} */,
  {32'hc1ec64a1, 32'hc0e43823} /* (1, 3, 6) {real, imag} */,
  {32'hc20aa5ba, 32'h41cc3352} /* (1, 3, 5) {real, imag} */,
  {32'h41cf4536, 32'h41f6624c} /* (1, 3, 4) {real, imag} */,
  {32'hbf0ea8a0, 32'hc2576169} /* (1, 3, 3) {real, imag} */,
  {32'hc16d933c, 32'h43010ee2} /* (1, 3, 2) {real, imag} */,
  {32'hc26040ab, 32'hc230f71b} /* (1, 3, 1) {real, imag} */,
  {32'h4203a094, 32'hc0819160} /* (1, 3, 0) {real, imag} */,
  {32'h440f74bf, 32'h427a5ecc} /* (1, 2, 31) {real, imag} */,
  {32'hc3941f88, 32'h41a755ad} /* (1, 2, 30) {real, imag} */,
  {32'h41eac239, 32'hc1b057f4} /* (1, 2, 29) {real, imag} */,
  {32'h422ede74, 32'hc190ddc8} /* (1, 2, 28) {real, imag} */,
  {32'hc20dfeb2, 32'h4258bd12} /* (1, 2, 27) {real, imag} */,
  {32'h40d584f0, 32'hbf85f77c} /* (1, 2, 26) {real, imag} */,
  {32'hbd877180, 32'hc11fc5a6} /* (1, 2, 25) {real, imag} */,
  {32'hc204197a, 32'h420f10a5} /* (1, 2, 24) {real, imag} */,
  {32'hc11d502c, 32'h3f3fbcd8} /* (1, 2, 23) {real, imag} */,
  {32'hc01d6ec2, 32'hc1a495f4} /* (1, 2, 22) {real, imag} */,
  {32'hc0d58bcb, 32'h411e36ee} /* (1, 2, 21) {real, imag} */,
  {32'h405ab3fc, 32'h3f8af4f2} /* (1, 2, 20) {real, imag} */,
  {32'hc08ebab4, 32'hc18e5fca} /* (1, 2, 19) {real, imag} */,
  {32'hc0f2bc28, 32'hc09c15e1} /* (1, 2, 18) {real, imag} */,
  {32'h3ecc8e70, 32'hc0880d63} /* (1, 2, 17) {real, imag} */,
  {32'hc04f1f28, 32'h40963c10} /* (1, 2, 16) {real, imag} */,
  {32'hbf1697ac, 32'h4032f798} /* (1, 2, 15) {real, imag} */,
  {32'h41129baf, 32'hc0a5698b} /* (1, 2, 14) {real, imag} */,
  {32'h3e83dd34, 32'hbf1152d4} /* (1, 2, 13) {real, imag} */,
  {32'hc0be1710, 32'h40ed7e51} /* (1, 2, 12) {real, imag} */,
  {32'hc1058d7c, 32'hc18e832c} /* (1, 2, 11) {real, imag} */,
  {32'hbfbafe7c, 32'hc02bc9de} /* (1, 2, 10) {real, imag} */,
  {32'h408f55cc, 32'hc0bd88ce} /* (1, 2, 9) {real, imag} */,
  {32'hc230dda9, 32'hc1d0ae8d} /* (1, 2, 8) {real, imag} */,
  {32'h40fc76e6, 32'h41c89424} /* (1, 2, 7) {real, imag} */,
  {32'hc044de90, 32'h40d4c3b8} /* (1, 2, 6) {real, imag} */,
  {32'hc2343e4e, 32'hc216daa0} /* (1, 2, 5) {real, imag} */,
  {32'h42d9c255, 32'h41814f84} /* (1, 2, 4) {real, imag} */,
  {32'hbfb14b08, 32'hc221752f} /* (1, 2, 3) {real, imag} */,
  {32'hc35ea3d9, 32'h42e01cae} /* (1, 2, 2) {real, imag} */,
  {32'h43820a3a, 32'h404c3680} /* (1, 2, 1) {real, imag} */,
  {32'h437e832c, 32'h42909d07} /* (1, 2, 0) {real, imag} */,
  {32'hc403a91f, 32'h426c4749} /* (1, 1, 31) {real, imag} */,
  {32'h4330976e, 32'hc177ed99} /* (1, 1, 30) {real, imag} */,
  {32'h41db8bbf, 32'hc1948293} /* (1, 1, 29) {real, imag} */,
  {32'hc2a9ed83, 32'hc1957882} /* (1, 1, 28) {real, imag} */,
  {32'h42edde0b, 32'hc07a27d4} /* (1, 1, 27) {real, imag} */,
  {32'h411ffd6c, 32'hc1025ed4} /* (1, 1, 26) {real, imag} */,
  {32'hc1abf0db, 32'hc03b6654} /* (1, 1, 25) {real, imag} */,
  {32'h420fce5a, 32'hc1c885b3} /* (1, 1, 24) {real, imag} */,
  {32'hc089ee3c, 32'hc1af7294} /* (1, 1, 23) {real, imag} */,
  {32'hc13c61bc, 32'hbfeceea2} /* (1, 1, 22) {real, imag} */,
  {32'h418e4ef0, 32'hc1876ade} /* (1, 1, 21) {real, imag} */,
  {32'hc0215bc4, 32'hc0955167} /* (1, 1, 20) {real, imag} */,
  {32'h40306312, 32'h3e08d180} /* (1, 1, 19) {real, imag} */,
  {32'hbf404404, 32'hbf829cc4} /* (1, 1, 18) {real, imag} */,
  {32'hc02598f4, 32'h408488f5} /* (1, 1, 17) {real, imag} */,
  {32'hbdc65be0, 32'h3f9acad8} /* (1, 1, 16) {real, imag} */,
  {32'h40fbf15b, 32'hc07bf001} /* (1, 1, 15) {real, imag} */,
  {32'hc0ccf26a, 32'h4148672d} /* (1, 1, 14) {real, imag} */,
  {32'hc13885de, 32'h3fda0810} /* (1, 1, 13) {real, imag} */,
  {32'h4119a388, 32'hc0985f5d} /* (1, 1, 12) {real, imag} */,
  {32'hc10a07af, 32'h4075b93a} /* (1, 1, 11) {real, imag} */,
  {32'hc0fa3e6b, 32'hc14d8960} /* (1, 1, 10) {real, imag} */,
  {32'hc0ee5500, 32'h41c2b294} /* (1, 1, 9) {real, imag} */,
  {32'h41678477, 32'h4169f1c1} /* (1, 1, 8) {real, imag} */,
  {32'hc166e3e4, 32'hc2016cbe} /* (1, 1, 7) {real, imag} */,
  {32'h4132f384, 32'h414ff0a1} /* (1, 1, 6) {real, imag} */,
  {32'h4271ea94, 32'h4213293c} /* (1, 1, 5) {real, imag} */,
  {32'h413ed3af, 32'hc2288e11} /* (1, 1, 4) {real, imag} */,
  {32'h4272a66d, 32'h40b6f578} /* (1, 1, 3) {real, imag} */,
  {32'h438ca72a, 32'h4367a1a0} /* (1, 1, 2) {real, imag} */,
  {32'hc4406709, 32'hc3fa5546} /* (1, 1, 1) {real, imag} */,
  {32'hc3f707f3, 32'h42852fc4} /* (1, 1, 0) {real, imag} */,
  {32'hc3b20afc, 32'h435b72e7} /* (1, 0, 31) {real, imag} */,
  {32'h412f7d10, 32'hc28f4804} /* (1, 0, 30) {real, imag} */,
  {32'h4236ff0d, 32'hc1bf489c} /* (1, 0, 29) {real, imag} */,
  {32'hc1dbd2bf, 32'hc28369d2} /* (1, 0, 28) {real, imag} */,
  {32'h428f374c, 32'h418e43d0} /* (1, 0, 27) {real, imag} */,
  {32'h4112bbc5, 32'hc09a78e3} /* (1, 0, 26) {real, imag} */,
  {32'hc1900e2b, 32'h420e648c} /* (1, 0, 25) {real, imag} */,
  {32'hbfb69cb0, 32'hc1f51311} /* (1, 0, 24) {real, imag} */,
  {32'hc05b412c, 32'hc1724727} /* (1, 0, 23) {real, imag} */,
  {32'h4135bd18, 32'h41180ece} /* (1, 0, 22) {real, imag} */,
  {32'h41868c37, 32'hc07b6c40} /* (1, 0, 21) {real, imag} */,
  {32'h41295788, 32'h414a5be8} /* (1, 0, 20) {real, imag} */,
  {32'h41219658, 32'h41372024} /* (1, 0, 19) {real, imag} */,
  {32'hc055fe0a, 32'hc1ada58a} /* (1, 0, 18) {real, imag} */,
  {32'hc134423a, 32'h403bb1e4} /* (1, 0, 17) {real, imag} */,
  {32'h408ba361, 32'h00000000} /* (1, 0, 16) {real, imag} */,
  {32'hc134423a, 32'hc03bb1e4} /* (1, 0, 15) {real, imag} */,
  {32'hc055fe0a, 32'h41ada58a} /* (1, 0, 14) {real, imag} */,
  {32'h41219658, 32'hc1372024} /* (1, 0, 13) {real, imag} */,
  {32'h41295788, 32'hc14a5be8} /* (1, 0, 12) {real, imag} */,
  {32'h41868c37, 32'h407b6c40} /* (1, 0, 11) {real, imag} */,
  {32'h4135bd18, 32'hc1180ece} /* (1, 0, 10) {real, imag} */,
  {32'hc05b412c, 32'h41724727} /* (1, 0, 9) {real, imag} */,
  {32'hbfb69cb0, 32'h41f51311} /* (1, 0, 8) {real, imag} */,
  {32'hc1900e2b, 32'hc20e648c} /* (1, 0, 7) {real, imag} */,
  {32'h4112bbc5, 32'h409a78e3} /* (1, 0, 6) {real, imag} */,
  {32'h428f374c, 32'hc18e43d0} /* (1, 0, 5) {real, imag} */,
  {32'hc1dbd2bf, 32'h428369d2} /* (1, 0, 4) {real, imag} */,
  {32'h4236ff0d, 32'h41bf489c} /* (1, 0, 3) {real, imag} */,
  {32'h412f7d10, 32'h428f4804} /* (1, 0, 2) {real, imag} */,
  {32'hc3b20afc, 32'hc35b72e7} /* (1, 0, 1) {real, imag} */,
  {32'hc3489817, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hc3a10d46, 32'h4383b8de} /* (0, 31, 31) {real, imag} */,
  {32'h42b2ad2b, 32'hc258411c} /* (0, 31, 30) {real, imag} */,
  {32'h424ebd20, 32'h4029676e} /* (0, 31, 29) {real, imag} */,
  {32'h417fe53b, 32'h4182d502} /* (0, 31, 28) {real, imag} */,
  {32'h419b3910, 32'hc152d494} /* (0, 31, 27) {real, imag} */,
  {32'h417e81df, 32'hc0e8c852} /* (0, 31, 26) {real, imag} */,
  {32'hc0c92e41, 32'h40e13823} /* (0, 31, 25) {real, imag} */,
  {32'hc0495710, 32'hc18ae0d9} /* (0, 31, 24) {real, imag} */,
  {32'hc035966f, 32'h409c186a} /* (0, 31, 23) {real, imag} */,
  {32'hc0baef38, 32'h40e8e6e2} /* (0, 31, 22) {real, imag} */,
  {32'h417d81e2, 32'h3fca66d0} /* (0, 31, 21) {real, imag} */,
  {32'hc011da41, 32'h408e09c6} /* (0, 31, 20) {real, imag} */,
  {32'h40eb60be, 32'h40d65758} /* (0, 31, 19) {real, imag} */,
  {32'hc09b913e, 32'h40010da8} /* (0, 31, 18) {real, imag} */,
  {32'h40d1671a, 32'hbf635cb4} /* (0, 31, 17) {real, imag} */,
  {32'h40164b88, 32'h4045bb2c} /* (0, 31, 16) {real, imag} */,
  {32'h3fd3c3fc, 32'h40e56e7c} /* (0, 31, 15) {real, imag} */,
  {32'h40bec258, 32'h3fd84e8a} /* (0, 31, 14) {real, imag} */,
  {32'h3f0f7db8, 32'h40945df1} /* (0, 31, 13) {real, imag} */,
  {32'hbfb1340a, 32'hc15a5d96} /* (0, 31, 12) {real, imag} */,
  {32'h411387d7, 32'h4181534a} /* (0, 31, 11) {real, imag} */,
  {32'hc1026137, 32'hc12dc5ba} /* (0, 31, 10) {real, imag} */,
  {32'h41652414, 32'h4182562b} /* (0, 31, 9) {real, imag} */,
  {32'h408c6d49, 32'h41455d3b} /* (0, 31, 8) {real, imag} */,
  {32'hc0934e91, 32'h40eace5c} /* (0, 31, 7) {real, imag} */,
  {32'hbf181580, 32'hc0aac079} /* (0, 31, 6) {real, imag} */,
  {32'h427c6b5a, 32'hc152b368} /* (0, 31, 5) {real, imag} */,
  {32'hc20ab738, 32'h3fef9e20} /* (0, 31, 4) {real, imag} */,
  {32'h41ee39b6, 32'hbee5b580} /* (0, 31, 3) {real, imag} */,
  {32'h427d3b82, 32'h4152b7fe} /* (0, 31, 2) {real, imag} */,
  {32'hc340868e, 32'h40d4e948} /* (0, 31, 1) {real, imag} */,
  {32'hc35a7e04, 32'hc2a3a2bb} /* (0, 31, 0) {real, imag} */,
  {32'h42a05470, 32'hc1a1e13a} /* (0, 30, 31) {real, imag} */,
  {32'hc2ba574a, 32'hc25c7406} /* (0, 30, 30) {real, imag} */,
  {32'hc101ae78, 32'h41b2e1fd} /* (0, 30, 29) {real, imag} */,
  {32'h426b503f, 32'hc12b9a7c} /* (0, 30, 28) {real, imag} */,
  {32'hc1c14726, 32'h41fd7cca} /* (0, 30, 27) {real, imag} */,
  {32'h41865b1a, 32'hc13c831f} /* (0, 30, 26) {real, imag} */,
  {32'h41353c14, 32'hc00fd624} /* (0, 30, 25) {real, imag} */,
  {32'hc1d78e4e, 32'h41276c4c} /* (0, 30, 24) {real, imag} */,
  {32'hc0d7c989, 32'h4097beb0} /* (0, 30, 23) {real, imag} */,
  {32'hc09f318b, 32'h40f33898} /* (0, 30, 22) {real, imag} */,
  {32'hc029148e, 32'h419a7ce4} /* (0, 30, 21) {real, imag} */,
  {32'h40940a1a, 32'h4154c76c} /* (0, 30, 20) {real, imag} */,
  {32'hc12c2314, 32'h3dd147c0} /* (0, 30, 19) {real, imag} */,
  {32'hbfe4927c, 32'h40c22bf2} /* (0, 30, 18) {real, imag} */,
  {32'h41394f7b, 32'h4008a388} /* (0, 30, 17) {real, imag} */,
  {32'h40066a5d, 32'hbec2bb98} /* (0, 30, 16) {real, imag} */,
  {32'h3fa166da, 32'hc065dc8d} /* (0, 30, 15) {real, imag} */,
  {32'h3f98607a, 32'h3e950cc8} /* (0, 30, 14) {real, imag} */,
  {32'hc00fdfd8, 32'hbeab661c} /* (0, 30, 13) {real, imag} */,
  {32'hc10dc2ff, 32'hc015b914} /* (0, 30, 12) {real, imag} */,
  {32'hc0a5812b, 32'h40ab840c} /* (0, 30, 11) {real, imag} */,
  {32'h3fffac9e, 32'hbfd18d80} /* (0, 30, 10) {real, imag} */,
  {32'h3eaa9ca0, 32'hbffd2270} /* (0, 30, 9) {real, imag} */,
  {32'hc12c923b, 32'hc168ff5c} /* (0, 30, 8) {real, imag} */,
  {32'hbfa59288, 32'hc10f07cc} /* (0, 30, 7) {real, imag} */,
  {32'hc0ab37a6, 32'hc1475e7f} /* (0, 30, 6) {real, imag} */,
  {32'hc19ec512, 32'hc20ea3fe} /* (0, 30, 5) {real, imag} */,
  {32'h41561c24, 32'h40ce82a8} /* (0, 30, 4) {real, imag} */,
  {32'h4165c05c, 32'h41ddefee} /* (0, 30, 3) {real, imag} */,
  {32'hc2fbb0a2, 32'hc08d3768} /* (0, 30, 2) {real, imag} */,
  {32'h43744033, 32'hc1062dad} /* (0, 30, 1) {real, imag} */,
  {32'h42ad914c, 32'hc1b351a6} /* (0, 30, 0) {real, imag} */,
  {32'hc182c6cb, 32'h421ab240} /* (0, 29, 31) {real, imag} */,
  {32'hc1b70cdb, 32'hc25bd312} /* (0, 29, 30) {real, imag} */,
  {32'h412f456d, 32'h41db544e} /* (0, 29, 29) {real, imag} */,
  {32'h4196c8c0, 32'hc1ff74dc} /* (0, 29, 28) {real, imag} */,
  {32'hc10dcb31, 32'hc12c67e3} /* (0, 29, 27) {real, imag} */,
  {32'hc1337fe9, 32'h4174799d} /* (0, 29, 26) {real, imag} */,
  {32'hc1c57eec, 32'h4025fdee} /* (0, 29, 25) {real, imag} */,
  {32'h410c4836, 32'hbf43eca8} /* (0, 29, 24) {real, imag} */,
  {32'h3f97a1b0, 32'h411885db} /* (0, 29, 23) {real, imag} */,
  {32'h407fded0, 32'hbf8f6e84} /* (0, 29, 22) {real, imag} */,
  {32'h40c86d54, 32'hc09ab7b3} /* (0, 29, 21) {real, imag} */,
  {32'h41452218, 32'hbfdb2794} /* (0, 29, 20) {real, imag} */,
  {32'hc05d2074, 32'h40c56582} /* (0, 29, 19) {real, imag} */,
  {32'hc1203e7d, 32'h3e51d0b0} /* (0, 29, 18) {real, imag} */,
  {32'h405a3198, 32'h3f562a30} /* (0, 29, 17) {real, imag} */,
  {32'h3dd85e60, 32'hc0f64c0b} /* (0, 29, 16) {real, imag} */,
  {32'h4077e26c, 32'h4046c0ce} /* (0, 29, 15) {real, imag} */,
  {32'hc129fc0a, 32'hc04f693f} /* (0, 29, 14) {real, imag} */,
  {32'h3e27c4c0, 32'hc0f46267} /* (0, 29, 13) {real, imag} */,
  {32'hc108847e, 32'hc08f7f18} /* (0, 29, 12) {real, imag} */,
  {32'hc0b0606e, 32'hc0874786} /* (0, 29, 11) {real, imag} */,
  {32'hc0e5b4d7, 32'h408f8d13} /* (0, 29, 10) {real, imag} */,
  {32'hc0a74892, 32'hbcfd0b40} /* (0, 29, 9) {real, imag} */,
  {32'h40e592e6, 32'hc1432a4e} /* (0, 29, 8) {real, imag} */,
  {32'hbfbe1d08, 32'h413338ee} /* (0, 29, 7) {real, imag} */,
  {32'h3f68ed32, 32'hc08d7896} /* (0, 29, 6) {real, imag} */,
  {32'h41766c44, 32'h4180d3a8} /* (0, 29, 5) {real, imag} */,
  {32'hc144cc1f, 32'h40908fb3} /* (0, 29, 4) {real, imag} */,
  {32'h41a33db4, 32'hc14f82f2} /* (0, 29, 3) {real, imag} */,
  {32'hc19e0af6, 32'hc186614a} /* (0, 29, 2) {real, imag} */,
  {32'h4233a764, 32'h40e3c504} /* (0, 29, 1) {real, imag} */,
  {32'h41de95d2, 32'hc15052ca} /* (0, 29, 0) {real, imag} */,
  {32'hc23201f0, 32'hc142a4a8} /* (0, 28, 31) {real, imag} */,
  {32'h41a8f9f0, 32'hc1f9347e} /* (0, 28, 30) {real, imag} */,
  {32'h40f011c4, 32'hc2005571} /* (0, 28, 29) {real, imag} */,
  {32'h3e6f90c0, 32'hbf6e57e0} /* (0, 28, 28) {real, imag} */,
  {32'h411ecd13, 32'h3f108ab8} /* (0, 28, 27) {real, imag} */,
  {32'hc0601044, 32'hc042bed8} /* (0, 28, 26) {real, imag} */,
  {32'hc1248d1c, 32'h41874adc} /* (0, 28, 25) {real, imag} */,
  {32'h4128080e, 32'hbf0e2758} /* (0, 28, 24) {real, imag} */,
  {32'h40ba30ce, 32'hc0e4d338} /* (0, 28, 23) {real, imag} */,
  {32'h41662196, 32'hc0b933a0} /* (0, 28, 22) {real, imag} */,
  {32'hc08d3248, 32'hc137699d} /* (0, 28, 21) {real, imag} */,
  {32'h4044ab8b, 32'h40163b42} /* (0, 28, 20) {real, imag} */,
  {32'h3fecef18, 32'hbf28af5c} /* (0, 28, 19) {real, imag} */,
  {32'hc05a7a3a, 32'hc0eefe3a} /* (0, 28, 18) {real, imag} */,
  {32'hbf6f2788, 32'h3f88e8af} /* (0, 28, 17) {real, imag} */,
  {32'h40a7c95a, 32'h409e68fa} /* (0, 28, 16) {real, imag} */,
  {32'hc02ba366, 32'h404064af} /* (0, 28, 15) {real, imag} */,
  {32'h3fe51bad, 32'hc1303466} /* (0, 28, 14) {real, imag} */,
  {32'hc12a9756, 32'hc0ca0ea1} /* (0, 28, 13) {real, imag} */,
  {32'hc0ec5250, 32'hc0e6bfde} /* (0, 28, 12) {real, imag} */,
  {32'h40464a1a, 32'h4007eb44} /* (0, 28, 11) {real, imag} */,
  {32'hc0850e62, 32'hbf8eb1b6} /* (0, 28, 10) {real, imag} */,
  {32'hc191d060, 32'h416f9dcf} /* (0, 28, 9) {real, imag} */,
  {32'hc02f0890, 32'h418a6271} /* (0, 28, 8) {real, imag} */,
  {32'h41ccb336, 32'hc18bce38} /* (0, 28, 7) {real, imag} */,
  {32'h3fd66aa0, 32'h411ad78c} /* (0, 28, 6) {real, imag} */,
  {32'hbfc81890, 32'h40e1c18b} /* (0, 28, 5) {real, imag} */,
  {32'hc0a49ea4, 32'hc104c117} /* (0, 28, 4) {real, imag} */,
  {32'hc1363d48, 32'h4103d145} /* (0, 28, 3) {real, imag} */,
  {32'hc08e65d8, 32'hc228d210} /* (0, 28, 2) {real, imag} */,
  {32'hc1dafaea, 32'h41881c40} /* (0, 28, 1) {real, imag} */,
  {32'h41b44f1b, 32'h413f2c90} /* (0, 28, 0) {real, imag} */,
  {32'hc1198fdb, 32'hc1d7dc4d} /* (0, 27, 31) {real, imag} */,
  {32'h413ddea6, 32'h415cdc75} /* (0, 27, 30) {real, imag} */,
  {32'hc12ff2a9, 32'h411e4730} /* (0, 27, 29) {real, imag} */,
  {32'hc0bca84a, 32'hc16db3a4} /* (0, 27, 28) {real, imag} */,
  {32'h40b3d0be, 32'hc0bf2f64} /* (0, 27, 27) {real, imag} */,
  {32'hc1597cb2, 32'hc0b82e02} /* (0, 27, 26) {real, imag} */,
  {32'h41399b89, 32'hc02f1e4e} /* (0, 27, 25) {real, imag} */,
  {32'h3e9bd958, 32'hbdcc4700} /* (0, 27, 24) {real, imag} */,
  {32'h409e367b, 32'h4037d278} /* (0, 27, 23) {real, imag} */,
  {32'hc0c517f8, 32'hc0a691d6} /* (0, 27, 22) {real, imag} */,
  {32'hbe1c2280, 32'h412e8819} /* (0, 27, 21) {real, imag} */,
  {32'hc0c87ffa, 32'hbfcc1718} /* (0, 27, 20) {real, imag} */,
  {32'h409ef95f, 32'hc0df9f68} /* (0, 27, 19) {real, imag} */,
  {32'h40dc2cb4, 32'h406d3b7d} /* (0, 27, 18) {real, imag} */,
  {32'h40bb2a26, 32'h40a15a44} /* (0, 27, 17) {real, imag} */,
  {32'hbfd72b74, 32'hc0bf6484} /* (0, 27, 16) {real, imag} */,
  {32'hbfb2b73a, 32'h40860916} /* (0, 27, 15) {real, imag} */,
  {32'hc0e73106, 32'hc11b38c9} /* (0, 27, 14) {real, imag} */,
  {32'h40a9dc56, 32'hbf9396f8} /* (0, 27, 13) {real, imag} */,
  {32'hc0d93810, 32'h40b84952} /* (0, 27, 12) {real, imag} */,
  {32'hc1721631, 32'h409a8403} /* (0, 27, 11) {real, imag} */,
  {32'hc14a591c, 32'hc1084caf} /* (0, 27, 10) {real, imag} */,
  {32'h408373c4, 32'hbfe82520} /* (0, 27, 9) {real, imag} */,
  {32'hc03e4454, 32'h41563453} /* (0, 27, 8) {real, imag} */,
  {32'hc0b6de07, 32'hbe0e9f00} /* (0, 27, 7) {real, imag} */,
  {32'h412bec51, 32'hc08adcee} /* (0, 27, 6) {real, imag} */,
  {32'h4098191d, 32'hc108a1b4} /* (0, 27, 5) {real, imag} */,
  {32'h41423f02, 32'hbf9bbcb8} /* (0, 27, 4) {real, imag} */,
  {32'hc18b99ef, 32'hc14b6c8e} /* (0, 27, 3) {real, imag} */,
  {32'hc1ad3a30, 32'hc0e17768} /* (0, 27, 2) {real, imag} */,
  {32'h420ebaf4, 32'h413e497d} /* (0, 27, 1) {real, imag} */,
  {32'h41ef0010, 32'h403baf20} /* (0, 27, 0) {real, imag} */,
  {32'hc0eb36e7, 32'h40b0d796} /* (0, 26, 31) {real, imag} */,
  {32'hc05c1a98, 32'h40eeb2bc} /* (0, 26, 30) {real, imag} */,
  {32'h41550ada, 32'hc0345c6d} /* (0, 26, 29) {real, imag} */,
  {32'h418716b4, 32'h410eb088} /* (0, 26, 28) {real, imag} */,
  {32'hc0cce642, 32'h40264dfd} /* (0, 26, 27) {real, imag} */,
  {32'hc145b992, 32'hc0891e86} /* (0, 26, 26) {real, imag} */,
  {32'h40553024, 32'hc09c772a} /* (0, 26, 25) {real, imag} */,
  {32'h3f81fe79, 32'h410c96dc} /* (0, 26, 24) {real, imag} */,
  {32'h410145e6, 32'h408af1ed} /* (0, 26, 23) {real, imag} */,
  {32'hc0f15624, 32'hc1603869} /* (0, 26, 22) {real, imag} */,
  {32'hc00182cc, 32'hc103ac96} /* (0, 26, 21) {real, imag} */,
  {32'hbec7f460, 32'hc10c3284} /* (0, 26, 20) {real, imag} */,
  {32'h3f5b65c0, 32'h40c133c4} /* (0, 26, 19) {real, imag} */,
  {32'hc1399698, 32'hc145a30d} /* (0, 26, 18) {real, imag} */,
  {32'hc04f2eee, 32'h405bb8f9} /* (0, 26, 17) {real, imag} */,
  {32'h3fbf7191, 32'hc0bc1f6a} /* (0, 26, 16) {real, imag} */,
  {32'h40c17bbd, 32'hbe0a4338} /* (0, 26, 15) {real, imag} */,
  {32'h3fd86e88, 32'hbf456300} /* (0, 26, 14) {real, imag} */,
  {32'h40c2233c, 32'h40837bce} /* (0, 26, 13) {real, imag} */,
  {32'h40bae08d, 32'hbee32920} /* (0, 26, 12) {real, imag} */,
  {32'h41027bd2, 32'h3eea96f8} /* (0, 26, 11) {real, imag} */,
  {32'hc0418b20, 32'h40919bd7} /* (0, 26, 10) {real, imag} */,
  {32'h40fd5bbc, 32'h40283170} /* (0, 26, 9) {real, imag} */,
  {32'hbf7a254c, 32'h40a9e5ad} /* (0, 26, 8) {real, imag} */,
  {32'h412a21b2, 32'hc06a7ee0} /* (0, 26, 7) {real, imag} */,
  {32'h3ff95568, 32'hc0a5c11a} /* (0, 26, 6) {real, imag} */,
  {32'h41838458, 32'h40e5e4a5} /* (0, 26, 5) {real, imag} */,
  {32'hc0a96ee3, 32'hc15cf7c7} /* (0, 26, 4) {real, imag} */,
  {32'h410488b7, 32'h41e38a55} /* (0, 26, 3) {real, imag} */,
  {32'hc1ce89bd, 32'hc19e2916} /* (0, 26, 2) {real, imag} */,
  {32'hc0022fbc, 32'hc1819710} /* (0, 26, 1) {real, imag} */,
  {32'hc026a99e, 32'h41fc7d9c} /* (0, 26, 0) {real, imag} */,
  {32'h41d96da6, 32'h41c87663} /* (0, 25, 31) {real, imag} */,
  {32'hc174a89c, 32'h412e7ef2} /* (0, 25, 30) {real, imag} */,
  {32'h40c5e34e, 32'h4091ed56} /* (0, 25, 29) {real, imag} */,
  {32'h40bbdf66, 32'hbf769778} /* (0, 25, 28) {real, imag} */,
  {32'h4112a3c2, 32'hc129f5e2} /* (0, 25, 27) {real, imag} */,
  {32'hc1617a78, 32'hc110177a} /* (0, 25, 26) {real, imag} */,
  {32'hc11da280, 32'h4004d830} /* (0, 25, 25) {real, imag} */,
  {32'hc01e525e, 32'h40d60bf1} /* (0, 25, 24) {real, imag} */,
  {32'h40d18d0e, 32'hc0b54ca8} /* (0, 25, 23) {real, imag} */,
  {32'hc0bb40a9, 32'h40d4bbe8} /* (0, 25, 22) {real, imag} */,
  {32'h40d143f1, 32'hc0341e54} /* (0, 25, 21) {real, imag} */,
  {32'hc0b2a501, 32'hc112f19e} /* (0, 25, 20) {real, imag} */,
  {32'hbd895340, 32'hc1161296} /* (0, 25, 19) {real, imag} */,
  {32'h40d3a96e, 32'h4081df98} /* (0, 25, 18) {real, imag} */,
  {32'hbdf53800, 32'hc0780a80} /* (0, 25, 17) {real, imag} */,
  {32'hc0439498, 32'h410d5fe4} /* (0, 25, 16) {real, imag} */,
  {32'hc0aec7b8, 32'hc034d5c0} /* (0, 25, 15) {real, imag} */,
  {32'hc10ec66e, 32'h3fd05e94} /* (0, 25, 14) {real, imag} */,
  {32'hbea127e0, 32'hc0d5de2a} /* (0, 25, 13) {real, imag} */,
  {32'h3c23a800, 32'h3fd0d9da} /* (0, 25, 12) {real, imag} */,
  {32'h40c0076c, 32'h3f2f30f0} /* (0, 25, 11) {real, imag} */,
  {32'h405c391c, 32'h40b8618f} /* (0, 25, 10) {real, imag} */,
  {32'hbfe621b4, 32'h3f0ceee0} /* (0, 25, 9) {real, imag} */,
  {32'h4088ba00, 32'h4095ea24} /* (0, 25, 8) {real, imag} */,
  {32'h4049718e, 32'h3f058ea8} /* (0, 25, 7) {real, imag} */,
  {32'hc0ad4f6c, 32'hbf5dc930} /* (0, 25, 6) {real, imag} */,
  {32'hc0a52ca6, 32'h40439573} /* (0, 25, 5) {real, imag} */,
  {32'h4115bab6, 32'hc159c31b} /* (0, 25, 4) {real, imag} */,
  {32'hc0f7c858, 32'hc188692d} /* (0, 25, 3) {real, imag} */,
  {32'h4135eefe, 32'hbc7e4400} /* (0, 25, 2) {real, imag} */,
  {32'hc0a28002, 32'hc11cad96} /* (0, 25, 1) {real, imag} */,
  {32'hc057ffec, 32'h4120a24c} /* (0, 25, 0) {real, imag} */,
  {32'h3f9c3980, 32'hc1a15289} /* (0, 24, 31) {real, imag} */,
  {32'hc1895349, 32'hc0899336} /* (0, 24, 30) {real, imag} */,
  {32'hc181de38, 32'hc0847694} /* (0, 24, 29) {real, imag} */,
  {32'h401dca6a, 32'hc013c4b8} /* (0, 24, 28) {real, imag} */,
  {32'h40fd9973, 32'h40dd3c6a} /* (0, 24, 27) {real, imag} */,
  {32'hc1276a7e, 32'h41049026} /* (0, 24, 26) {real, imag} */,
  {32'h40e8aebc, 32'hc13c7027} /* (0, 24, 25) {real, imag} */,
  {32'h4062c7ba, 32'h3f503f30} /* (0, 24, 24) {real, imag} */,
  {32'hc00960bc, 32'h3f819d68} /* (0, 24, 23) {real, imag} */,
  {32'hc1363392, 32'hc0329500} /* (0, 24, 22) {real, imag} */,
  {32'h4110954c, 32'h40c322b9} /* (0, 24, 21) {real, imag} */,
  {32'hc0b5ab09, 32'h40ab1723} /* (0, 24, 20) {real, imag} */,
  {32'hc04350fc, 32'hc10e22ae} /* (0, 24, 19) {real, imag} */,
  {32'h40dc36e6, 32'hc152eba7} /* (0, 24, 18) {real, imag} */,
  {32'h405755f0, 32'hbf4c52b0} /* (0, 24, 17) {real, imag} */,
  {32'hbf31fc00, 32'h4135419e} /* (0, 24, 16) {real, imag} */,
  {32'hc0498d65, 32'h40147032} /* (0, 24, 15) {real, imag} */,
  {32'h412d80d0, 32'h408ca485} /* (0, 24, 14) {real, imag} */,
  {32'h40e87837, 32'hc0a1c36d} /* (0, 24, 13) {real, imag} */,
  {32'hc0bf7d6b, 32'h3fbea540} /* (0, 24, 12) {real, imag} */,
  {32'hc0a9e3f4, 32'hc13a7491} /* (0, 24, 11) {real, imag} */,
  {32'hc0fce8e5, 32'h41669015} /* (0, 24, 10) {real, imag} */,
  {32'h413c6d8b, 32'h408b0487} /* (0, 24, 9) {real, imag} */,
  {32'hc17cc5e2, 32'hc0b510ec} /* (0, 24, 8) {real, imag} */,
  {32'h410b3d56, 32'h4139ac7d} /* (0, 24, 7) {real, imag} */,
  {32'h40aeaff6, 32'hc01deacc} /* (0, 24, 6) {real, imag} */,
  {32'hc080034a, 32'h40ae6ea0} /* (0, 24, 5) {real, imag} */,
  {32'h417610dc, 32'h4096e9e6} /* (0, 24, 4) {real, imag} */,
  {32'hbf3cf3d8, 32'h409037e1} /* (0, 24, 3) {real, imag} */,
  {32'hc2064771, 32'h41069517} /* (0, 24, 2) {real, imag} */,
  {32'h40cc7b92, 32'hc18850e1} /* (0, 24, 1) {real, imag} */,
  {32'h41b1299e, 32'hc195be20} /* (0, 24, 0) {real, imag} */,
  {32'hc19d2422, 32'hc087ce90} /* (0, 23, 31) {real, imag} */,
  {32'h3fbe5a24, 32'hbf4c68c0} /* (0, 23, 30) {real, imag} */,
  {32'hbfe2ccbc, 32'h41384dc6} /* (0, 23, 29) {real, imag} */,
  {32'hc0191e32, 32'hc102cb4f} /* (0, 23, 28) {real, imag} */,
  {32'hbf58159a, 32'hc00fc468} /* (0, 23, 27) {real, imag} */,
  {32'h41215090, 32'hbfaaa520} /* (0, 23, 26) {real, imag} */,
  {32'h4056d538, 32'hbfc1c0f2} /* (0, 23, 25) {real, imag} */,
  {32'hbfdff710, 32'hc1485cc8} /* (0, 23, 24) {real, imag} */,
  {32'hc0dbfd9e, 32'h40063f86} /* (0, 23, 23) {real, imag} */,
  {32'h40fb4aa0, 32'hc114dc92} /* (0, 23, 22) {real, imag} */,
  {32'hc16ce180, 32'hbe624fc0} /* (0, 23, 21) {real, imag} */,
  {32'h411a2ed5, 32'hc1087a14} /* (0, 23, 20) {real, imag} */,
  {32'hbff37254, 32'hbed4f2a8} /* (0, 23, 19) {real, imag} */,
  {32'hc107b8ca, 32'hbdab0560} /* (0, 23, 18) {real, imag} */,
  {32'h3fcd0d20, 32'h401ec486} /* (0, 23, 17) {real, imag} */,
  {32'h4098bb41, 32'h3e808c40} /* (0, 23, 16) {real, imag} */,
  {32'hc065454f, 32'h40ca01d3} /* (0, 23, 15) {real, imag} */,
  {32'hc0c26d7d, 32'hc051c736} /* (0, 23, 14) {real, imag} */,
  {32'h40c5325c, 32'hbea42578} /* (0, 23, 13) {real, imag} */,
  {32'h3f67ee98, 32'h40c45ea4} /* (0, 23, 12) {real, imag} */,
  {32'hbf161320, 32'hbf71d198} /* (0, 23, 11) {real, imag} */,
  {32'hbda84880, 32'hc12560ce} /* (0, 23, 10) {real, imag} */,
  {32'h3fc91348, 32'hc056c3f6} /* (0, 23, 9) {real, imag} */,
  {32'h40af73ce, 32'h4128cbb5} /* (0, 23, 8) {real, imag} */,
  {32'h411bcfd6, 32'h3f14dd58} /* (0, 23, 7) {real, imag} */,
  {32'hbf7691a0, 32'h40dec45f} /* (0, 23, 6) {real, imag} */,
  {32'h40ecf843, 32'h3f273028} /* (0, 23, 5) {real, imag} */,
  {32'hc14ee360, 32'h418cf41b} /* (0, 23, 4) {real, imag} */,
  {32'hc1adc512, 32'hc141766c} /* (0, 23, 3) {real, imag} */,
  {32'h419e3a69, 32'hc182174f} /* (0, 23, 2) {real, imag} */,
  {32'h3edc3c28, 32'h408d45cf} /* (0, 23, 1) {real, imag} */,
  {32'hc14f06c5, 32'h4088554c} /* (0, 23, 0) {real, imag} */,
  {32'hc19a8a3c, 32'h3ea7da90} /* (0, 22, 31) {real, imag} */,
  {32'h4197403c, 32'hc1bef3a2} /* (0, 22, 30) {real, imag} */,
  {32'hbfc8e058, 32'hc026387b} /* (0, 22, 29) {real, imag} */,
  {32'h40885a68, 32'h410568ba} /* (0, 22, 28) {real, imag} */,
  {32'hc056b508, 32'h3eb34c28} /* (0, 22, 27) {real, imag} */,
  {32'hbff46e2c, 32'h3f663958} /* (0, 22, 26) {real, imag} */,
  {32'h408d32b6, 32'h40387fa8} /* (0, 22, 25) {real, imag} */,
  {32'h4098f172, 32'h404ffbb4} /* (0, 22, 24) {real, imag} */,
  {32'h3fd080fa, 32'h416af5ae} /* (0, 22, 23) {real, imag} */,
  {32'h41065f62, 32'h407ea096} /* (0, 22, 22) {real, imag} */,
  {32'h40a645f5, 32'h402f4698} /* (0, 22, 21) {real, imag} */,
  {32'hc15c6ba2, 32'h4168ca45} /* (0, 22, 20) {real, imag} */,
  {32'h41329ef4, 32'h400b6914} /* (0, 22, 19) {real, imag} */,
  {32'h40b0295c, 32'h408f237e} /* (0, 22, 18) {real, imag} */,
  {32'hc07cda8c, 32'hc0625f92} /* (0, 22, 17) {real, imag} */,
  {32'h4000c70a, 32'h40ad92bc} /* (0, 22, 16) {real, imag} */,
  {32'h3f4d43ec, 32'hbd8fbd00} /* (0, 22, 15) {real, imag} */,
  {32'hc0b12066, 32'h3feeb666} /* (0, 22, 14) {real, imag} */,
  {32'h409af9f8, 32'hbf274830} /* (0, 22, 13) {real, imag} */,
  {32'h404d83c4, 32'hc0f4f3b2} /* (0, 22, 12) {real, imag} */,
  {32'h404fbbfc, 32'h40e03e80} /* (0, 22, 11) {real, imag} */,
  {32'hc090570f, 32'h40c502aa} /* (0, 22, 10) {real, imag} */,
  {32'h40d88486, 32'h413b5b48} /* (0, 22, 9) {real, imag} */,
  {32'h416739a8, 32'h410964e2} /* (0, 22, 8) {real, imag} */,
  {32'h3f17c970, 32'h406a99db} /* (0, 22, 7) {real, imag} */,
  {32'hbf9dd44c, 32'hc12e7ede} /* (0, 22, 6) {real, imag} */,
  {32'h417420ec, 32'hc0a16d08} /* (0, 22, 5) {real, imag} */,
  {32'hc1197e51, 32'h4114e99f} /* (0, 22, 4) {real, imag} */,
  {32'hc089faa3, 32'h405393fd} /* (0, 22, 3) {real, imag} */,
  {32'hbf5e3410, 32'hc1082b57} /* (0, 22, 2) {real, imag} */,
  {32'hbf883304, 32'h40216f7e} /* (0, 22, 1) {real, imag} */,
  {32'h406d1ed8, 32'h4012ae52} /* (0, 22, 0) {real, imag} */,
  {32'h4086507f, 32'h40827d23} /* (0, 21, 31) {real, imag} */,
  {32'h4055c0b4, 32'h4140fcdd} /* (0, 21, 30) {real, imag} */,
  {32'h40d39569, 32'h40246088} /* (0, 21, 29) {real, imag} */,
  {32'hc0618ee6, 32'h412b2984} /* (0, 21, 28) {real, imag} */,
  {32'hc13c1c0e, 32'hc0dca805} /* (0, 21, 27) {real, imag} */,
  {32'h4052335c, 32'h403f15e8} /* (0, 21, 26) {real, imag} */,
  {32'h4084aa46, 32'h3f8404ad} /* (0, 21, 25) {real, imag} */,
  {32'hc014bec8, 32'hc0ec6655} /* (0, 21, 24) {real, imag} */,
  {32'h406c915e, 32'hc02091b0} /* (0, 21, 23) {real, imag} */,
  {32'hc1dbcabc, 32'h40a7c818} /* (0, 21, 22) {real, imag} */,
  {32'h4113d3dd, 32'h40788aaf} /* (0, 21, 21) {real, imag} */,
  {32'hc0bf1264, 32'hc19e6e4c} /* (0, 21, 20) {real, imag} */,
  {32'hbf9ed97c, 32'h4032b870} /* (0, 21, 19) {real, imag} */,
  {32'h415922de, 32'h406fb1ae} /* (0, 21, 18) {real, imag} */,
  {32'hc05e2b16, 32'hc0166295} /* (0, 21, 17) {real, imag} */,
  {32'hc04536e2, 32'hc08cdd56} /* (0, 21, 16) {real, imag} */,
  {32'hbf96fbdc, 32'h40e0963b} /* (0, 21, 15) {real, imag} */,
  {32'hc081069c, 32'hc11ac822} /* (0, 21, 14) {real, imag} */,
  {32'hc05d6290, 32'hc0e97720} /* (0, 21, 13) {real, imag} */,
  {32'h40d997b7, 32'hc08c1200} /* (0, 21, 12) {real, imag} */,
  {32'hc090e220, 32'h41cbfbb0} /* (0, 21, 11) {real, imag} */,
  {32'h3fd891e0, 32'hbf84e3e0} /* (0, 21, 10) {real, imag} */,
  {32'hc00379f0, 32'h403a598a} /* (0, 21, 9) {real, imag} */,
  {32'h40cd3e85, 32'hc12b0f0e} /* (0, 21, 8) {real, imag} */,
  {32'hc033ea35, 32'hc02dfd22} /* (0, 21, 7) {real, imag} */,
  {32'h412d1b80, 32'hc1103f66} /* (0, 21, 6) {real, imag} */,
  {32'hc02ca0d0, 32'h3eadc5e0} /* (0, 21, 5) {real, imag} */,
  {32'hc0fd3084, 32'h40be8708} /* (0, 21, 4) {real, imag} */,
  {32'hc10cd5c8, 32'hc12b2fb0} /* (0, 21, 3) {real, imag} */,
  {32'h4119aab3, 32'h408ab698} /* (0, 21, 2) {real, imag} */,
  {32'h413178fe, 32'hbf435440} /* (0, 21, 1) {real, imag} */,
  {32'hc03a6690, 32'hbf81b194} /* (0, 21, 0) {real, imag} */,
  {32'h410eb132, 32'h40d41659} /* (0, 20, 31) {real, imag} */,
  {32'h41295892, 32'hc0bea2dc} /* (0, 20, 30) {real, imag} */,
  {32'h3e604d40, 32'h3edaa400} /* (0, 20, 29) {real, imag} */,
  {32'hc0890d53, 32'hc112c8ac} /* (0, 20, 28) {real, imag} */,
  {32'hc09a7e45, 32'h412d2906} /* (0, 20, 27) {real, imag} */,
  {32'hc0caf0b4, 32'h4094d2d4} /* (0, 20, 26) {real, imag} */,
  {32'h40c3e9cb, 32'hc1311fae} /* (0, 20, 25) {real, imag} */,
  {32'h3e96a380, 32'h41239878} /* (0, 20, 24) {real, imag} */,
  {32'h4022b5da, 32'h3fa74ca4} /* (0, 20, 23) {real, imag} */,
  {32'h40b2803a, 32'h40a946ec} /* (0, 20, 22) {real, imag} */,
  {32'hc16376d2, 32'hbfb6d37d} /* (0, 20, 21) {real, imag} */,
  {32'h4081db02, 32'hc0f64178} /* (0, 20, 20) {real, imag} */,
  {32'h409d30c5, 32'h40ec944c} /* (0, 20, 19) {real, imag} */,
  {32'hc0b7dc10, 32'h411b09ea} /* (0, 20, 18) {real, imag} */,
  {32'h3fb87988, 32'h40fe05e2} /* (0, 20, 17) {real, imag} */,
  {32'hc036decc, 32'hc067f565} /* (0, 20, 16) {real, imag} */,
  {32'hc064950b, 32'hc0e66601} /* (0, 20, 15) {real, imag} */,
  {32'h40d90713, 32'h4009e298} /* (0, 20, 14) {real, imag} */,
  {32'h416955fa, 32'hc09a2e1f} /* (0, 20, 13) {real, imag} */,
  {32'h3ec0d330, 32'hbfe38e80} /* (0, 20, 12) {real, imag} */,
  {32'h40aee37a, 32'h40503379} /* (0, 20, 11) {real, imag} */,
  {32'h3fd792e7, 32'h3f07b970} /* (0, 20, 10) {real, imag} */,
  {32'hbfc2d440, 32'hc17317e6} /* (0, 20, 9) {real, imag} */,
  {32'hc0b29a89, 32'hc0ee6bc2} /* (0, 20, 8) {real, imag} */,
  {32'h4097d8c8, 32'h40845798} /* (0, 20, 7) {real, imag} */,
  {32'hc04d6beb, 32'h40eafc59} /* (0, 20, 6) {real, imag} */,
  {32'hc10cc4ce, 32'hbf7f5c10} /* (0, 20, 5) {real, imag} */,
  {32'hc0ff7558, 32'h3f981770} /* (0, 20, 4) {real, imag} */,
  {32'hc03f5527, 32'h412ea198} /* (0, 20, 3) {real, imag} */,
  {32'hc0776348, 32'h41091bc9} /* (0, 20, 2) {real, imag} */,
  {32'h4097eaae, 32'hc16fd661} /* (0, 20, 1) {real, imag} */,
  {32'h3f56b808, 32'h4115a892} /* (0, 20, 0) {real, imag} */,
  {32'h40f8e841, 32'hc00f6b7a} /* (0, 19, 31) {real, imag} */,
  {32'h3f27aac8, 32'h40bd4474} /* (0, 19, 30) {real, imag} */,
  {32'h4021bf94, 32'hc088b5f2} /* (0, 19, 29) {real, imag} */,
  {32'h3f54a6f0, 32'h41094a27} /* (0, 19, 28) {real, imag} */,
  {32'h3f8ac577, 32'hbfa01be2} /* (0, 19, 27) {real, imag} */,
  {32'h40135c45, 32'h40a30dc8} /* (0, 19, 26) {real, imag} */,
  {32'hc1315e52, 32'hc07f6773} /* (0, 19, 25) {real, imag} */,
  {32'h415633b8, 32'h412af2ad} /* (0, 19, 24) {real, imag} */,
  {32'hc0832715, 32'hc159868e} /* (0, 19, 23) {real, imag} */,
  {32'h416eaa25, 32'hbf870090} /* (0, 19, 22) {real, imag} */,
  {32'hc0e74fca, 32'hc024fbe2} /* (0, 19, 21) {real, imag} */,
  {32'hbf3a666c, 32'hbf8ab2bc} /* (0, 19, 20) {real, imag} */,
  {32'h40aae4e4, 32'h405d25f4} /* (0, 19, 19) {real, imag} */,
  {32'hc0f15950, 32'h40d1732c} /* (0, 19, 18) {real, imag} */,
  {32'h410931e8, 32'hbf853820} /* (0, 19, 17) {real, imag} */,
  {32'h40a9d8cc, 32'h3ff3633e} /* (0, 19, 16) {real, imag} */,
  {32'hc0782996, 32'hc106075f} /* (0, 19, 15) {real, imag} */,
  {32'hc12299ff, 32'hc14431a4} /* (0, 19, 14) {real, imag} */,
  {32'hc0e4ee0b, 32'hbffa5cfc} /* (0, 19, 13) {real, imag} */,
  {32'hc00d2450, 32'h3fd198c6} /* (0, 19, 12) {real, imag} */,
  {32'hc0d8370b, 32'h40ce7ddc} /* (0, 19, 11) {real, imag} */,
  {32'h40ed362e, 32'h40bc0318} /* (0, 19, 10) {real, imag} */,
  {32'h3fa3fc20, 32'hbfa04528} /* (0, 19, 9) {real, imag} */,
  {32'hbf7c21a8, 32'hc0d5211e} /* (0, 19, 8) {real, imag} */,
  {32'h40d44ec2, 32'hc0d1b25e} /* (0, 19, 7) {real, imag} */,
  {32'h40d547a3, 32'h40a184ae} /* (0, 19, 6) {real, imag} */,
  {32'hbc852a00, 32'h40a495a1} /* (0, 19, 5) {real, imag} */,
  {32'hc01f4ee0, 32'h4129aa18} /* (0, 19, 4) {real, imag} */,
  {32'hc13b4432, 32'hc0eb22b4} /* (0, 19, 3) {real, imag} */,
  {32'h41932189, 32'hc0ea3c26} /* (0, 19, 2) {real, imag} */,
  {32'hc06c0cf6, 32'h4124aa5b} /* (0, 19, 1) {real, imag} */,
  {32'hc150aa9e, 32'hc1120454} /* (0, 19, 0) {real, imag} */,
  {32'hc12dba82, 32'hc13069c2} /* (0, 18, 31) {real, imag} */,
  {32'hc0af8be0, 32'h40ebd1c5} /* (0, 18, 30) {real, imag} */,
  {32'h40dfe07b, 32'h40b1b8f0} /* (0, 18, 29) {real, imag} */,
  {32'h3fc91ffe, 32'hc0c211f3} /* (0, 18, 28) {real, imag} */,
  {32'hc06aed0e, 32'h412b82a8} /* (0, 18, 27) {real, imag} */,
  {32'h40896dd9, 32'hbfa15c56} /* (0, 18, 26) {real, imag} */,
  {32'h4109e1c8, 32'h40b9f2ac} /* (0, 18, 25) {real, imag} */,
  {32'h4011924d, 32'h4116d925} /* (0, 18, 24) {real, imag} */,
  {32'hc11cd7b3, 32'h40d6e5a6} /* (0, 18, 23) {real, imag} */,
  {32'hc0d480df, 32'hc0ca639c} /* (0, 18, 22) {real, imag} */,
  {32'h413951a8, 32'hc04a1988} /* (0, 18, 21) {real, imag} */,
  {32'h41277c65, 32'hc04319b0} /* (0, 18, 20) {real, imag} */,
  {32'h40b9f2cb, 32'h40903641} /* (0, 18, 19) {real, imag} */,
  {32'h4041fdda, 32'hbe49b6a0} /* (0, 18, 18) {real, imag} */,
  {32'hc007ce5a, 32'h40be04d2} /* (0, 18, 17) {real, imag} */,
  {32'h3f6acbd0, 32'h410dfeda} /* (0, 18, 16) {real, imag} */,
  {32'hc060cec8, 32'h40814057} /* (0, 18, 15) {real, imag} */,
  {32'h40b7c2e0, 32'hc10ec21c} /* (0, 18, 14) {real, imag} */,
  {32'hbf910ed8, 32'h3fc5e6d1} /* (0, 18, 13) {real, imag} */,
  {32'h40e677ec, 32'hbfca7e48} /* (0, 18, 12) {real, imag} */,
  {32'h406850ce, 32'hc055941a} /* (0, 18, 11) {real, imag} */,
  {32'hc04903ba, 32'h41a3fa4c} /* (0, 18, 10) {real, imag} */,
  {32'h4117543b, 32'hc0c72560} /* (0, 18, 9) {real, imag} */,
  {32'h3fabb6bc, 32'h409baf7f} /* (0, 18, 8) {real, imag} */,
  {32'hc02873ea, 32'h410dfeb8} /* (0, 18, 7) {real, imag} */,
  {32'hc08fd1b0, 32'hc067df2a} /* (0, 18, 6) {real, imag} */,
  {32'h400d82e9, 32'h4110bf2f} /* (0, 18, 5) {real, imag} */,
  {32'h40e568f4, 32'hc0e64bd6} /* (0, 18, 4) {real, imag} */,
  {32'hc07e843b, 32'hc0099d90} /* (0, 18, 3) {real, imag} */,
  {32'hc14f2ede, 32'h3cfa4140} /* (0, 18, 2) {real, imag} */,
  {32'hbfddee9d, 32'hbd6ce880} /* (0, 18, 1) {real, imag} */,
  {32'hbf973234, 32'hc0a82256} /* (0, 18, 0) {real, imag} */,
  {32'hc081b70a, 32'h408854c5} /* (0, 17, 31) {real, imag} */,
  {32'h4122d3ac, 32'hc11a5886} /* (0, 17, 30) {real, imag} */,
  {32'hc01f4d2c, 32'h3ff0c0e0} /* (0, 17, 29) {real, imag} */,
  {32'h3fa00d95, 32'h3ed35ac8} /* (0, 17, 28) {real, imag} */,
  {32'h3f464c90, 32'h3eee2a94} /* (0, 17, 27) {real, imag} */,
  {32'hc0cc0428, 32'hc02d6152} /* (0, 17, 26) {real, imag} */,
  {32'h40ba15dd, 32'h407be8f0} /* (0, 17, 25) {real, imag} */,
  {32'hc0102eea, 32'h40e03b9c} /* (0, 17, 24) {real, imag} */,
  {32'hc0af5d75, 32'h401eb344} /* (0, 17, 23) {real, imag} */,
  {32'h4118ebc2, 32'h40152545} /* (0, 17, 22) {real, imag} */,
  {32'hc08598f7, 32'hbfb17698} /* (0, 17, 21) {real, imag} */,
  {32'hc09926db, 32'h4129051f} /* (0, 17, 20) {real, imag} */,
  {32'h40f67076, 32'hc0c127a4} /* (0, 17, 19) {real, imag} */,
  {32'hbf518498, 32'h4040b6e1} /* (0, 17, 18) {real, imag} */,
  {32'hc07f0f10, 32'h3ed2ef60} /* (0, 17, 17) {real, imag} */,
  {32'hc0b881d8, 32'h3f98aabf} /* (0, 17, 16) {real, imag} */,
  {32'h40e17661, 32'h3ecb38f0} /* (0, 17, 15) {real, imag} */,
  {32'h40be0e12, 32'h40c1f5f7} /* (0, 17, 14) {real, imag} */,
  {32'hc0dbcc14, 32'hc0efb84e} /* (0, 17, 13) {real, imag} */,
  {32'hc06e8ea6, 32'h410d7cc4} /* (0, 17, 12) {real, imag} */,
  {32'hc08b652e, 32'hc106a54a} /* (0, 17, 11) {real, imag} */,
  {32'hc002f204, 32'h3f6e853c} /* (0, 17, 10) {real, imag} */,
  {32'h40d813b7, 32'h40e4c010} /* (0, 17, 9) {real, imag} */,
  {32'hc029cbb0, 32'hbfde1f86} /* (0, 17, 8) {real, imag} */,
  {32'h3ece0710, 32'hbe2d8780} /* (0, 17, 7) {real, imag} */,
  {32'h3fc9092c, 32'hc092264a} /* (0, 17, 6) {real, imag} */,
  {32'h403dcdc2, 32'hc0378610} /* (0, 17, 5) {real, imag} */,
  {32'hc08848c6, 32'hc00b5424} /* (0, 17, 4) {real, imag} */,
  {32'h401f3e45, 32'h3e8ec9d0} /* (0, 17, 3) {real, imag} */,
  {32'hbfa24610, 32'hc156b678} /* (0, 17, 2) {real, imag} */,
  {32'h4047ee00, 32'h41295790} /* (0, 17, 1) {real, imag} */,
  {32'hbe5cd958, 32'hc02991a8} /* (0, 17, 0) {real, imag} */,
  {32'hbfcc849f, 32'h3f3c5e48} /* (0, 16, 31) {real, imag} */,
  {32'h402d4e08, 32'h402f5ef0} /* (0, 16, 30) {real, imag} */,
  {32'hc05dcefa, 32'hbf1ff684} /* (0, 16, 29) {real, imag} */,
  {32'h3e143478, 32'h3fd68590} /* (0, 16, 28) {real, imag} */,
  {32'hbf8c2900, 32'hbc8d8e00} /* (0, 16, 27) {real, imag} */,
  {32'hc01444f2, 32'h3f69e3c8} /* (0, 16, 26) {real, imag} */,
  {32'hbeac0010, 32'h412ec518} /* (0, 16, 25) {real, imag} */,
  {32'h4072689c, 32'hbfca4df4} /* (0, 16, 24) {real, imag} */,
  {32'h41258d3c, 32'hbf871eba} /* (0, 16, 23) {real, imag} */,
  {32'hc02b123b, 32'h4062eccd} /* (0, 16, 22) {real, imag} */,
  {32'h3f3a52fa, 32'h40405df8} /* (0, 16, 21) {real, imag} */,
  {32'hc111ef80, 32'h407b6fd8} /* (0, 16, 20) {real, imag} */,
  {32'hbf01d956, 32'h41600c18} /* (0, 16, 19) {real, imag} */,
  {32'hc0257574, 32'h40125b1d} /* (0, 16, 18) {real, imag} */,
  {32'hbf61921a, 32'h408ac1e1} /* (0, 16, 17) {real, imag} */,
  {32'hbe2186f8, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hbf61921a, 32'hc08ac1e1} /* (0, 16, 15) {real, imag} */,
  {32'hc0257574, 32'hc0125b1d} /* (0, 16, 14) {real, imag} */,
  {32'hbf01d956, 32'hc1600c18} /* (0, 16, 13) {real, imag} */,
  {32'hc111ef80, 32'hc07b6fd8} /* (0, 16, 12) {real, imag} */,
  {32'h3f3a52fa, 32'hc0405df8} /* (0, 16, 11) {real, imag} */,
  {32'hc02b123b, 32'hc062eccd} /* (0, 16, 10) {real, imag} */,
  {32'h41258d3c, 32'h3f871eba} /* (0, 16, 9) {real, imag} */,
  {32'h4072689c, 32'h3fca4df4} /* (0, 16, 8) {real, imag} */,
  {32'hbeac0010, 32'hc12ec518} /* (0, 16, 7) {real, imag} */,
  {32'hc01444f2, 32'hbf69e3c8} /* (0, 16, 6) {real, imag} */,
  {32'hbf8c2900, 32'h3c8d8e00} /* (0, 16, 5) {real, imag} */,
  {32'h3e143478, 32'hbfd68590} /* (0, 16, 4) {real, imag} */,
  {32'hc05dcefa, 32'h3f1ff684} /* (0, 16, 3) {real, imag} */,
  {32'h402d4e08, 32'hc02f5ef0} /* (0, 16, 2) {real, imag} */,
  {32'hbfcc849f, 32'hbf3c5e48} /* (0, 16, 1) {real, imag} */,
  {32'h417765c6, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h4047ee00, 32'hc1295790} /* (0, 15, 31) {real, imag} */,
  {32'hbfa24610, 32'h4156b678} /* (0, 15, 30) {real, imag} */,
  {32'h401f3e45, 32'hbe8ec9d0} /* (0, 15, 29) {real, imag} */,
  {32'hc08848c6, 32'h400b5424} /* (0, 15, 28) {real, imag} */,
  {32'h403dcdc2, 32'h40378610} /* (0, 15, 27) {real, imag} */,
  {32'h3fc9092c, 32'h4092264a} /* (0, 15, 26) {real, imag} */,
  {32'h3ece0710, 32'h3e2d8780} /* (0, 15, 25) {real, imag} */,
  {32'hc029cbb0, 32'h3fde1f86} /* (0, 15, 24) {real, imag} */,
  {32'h40d813b7, 32'hc0e4c010} /* (0, 15, 23) {real, imag} */,
  {32'hc002f204, 32'hbf6e853c} /* (0, 15, 22) {real, imag} */,
  {32'hc08b652e, 32'h4106a54a} /* (0, 15, 21) {real, imag} */,
  {32'hc06e8ea6, 32'hc10d7cc4} /* (0, 15, 20) {real, imag} */,
  {32'hc0dbcc14, 32'h40efb84e} /* (0, 15, 19) {real, imag} */,
  {32'h40be0e12, 32'hc0c1f5f7} /* (0, 15, 18) {real, imag} */,
  {32'h40e17661, 32'hbecb38f0} /* (0, 15, 17) {real, imag} */,
  {32'hc0b881d8, 32'hbf98aabf} /* (0, 15, 16) {real, imag} */,
  {32'hc07f0f10, 32'hbed2ef60} /* (0, 15, 15) {real, imag} */,
  {32'hbf518498, 32'hc040b6e1} /* (0, 15, 14) {real, imag} */,
  {32'h40f67076, 32'h40c127a4} /* (0, 15, 13) {real, imag} */,
  {32'hc09926db, 32'hc129051f} /* (0, 15, 12) {real, imag} */,
  {32'hc08598f7, 32'h3fb17698} /* (0, 15, 11) {real, imag} */,
  {32'h4118ebc2, 32'hc0152545} /* (0, 15, 10) {real, imag} */,
  {32'hc0af5d75, 32'hc01eb344} /* (0, 15, 9) {real, imag} */,
  {32'hc0102eea, 32'hc0e03b9c} /* (0, 15, 8) {real, imag} */,
  {32'h40ba15dd, 32'hc07be8f0} /* (0, 15, 7) {real, imag} */,
  {32'hc0cc0428, 32'h402d6152} /* (0, 15, 6) {real, imag} */,
  {32'h3f464c90, 32'hbeee2a94} /* (0, 15, 5) {real, imag} */,
  {32'h3fa00d95, 32'hbed35ac8} /* (0, 15, 4) {real, imag} */,
  {32'hc01f4d2c, 32'hbff0c0e0} /* (0, 15, 3) {real, imag} */,
  {32'h4122d3ac, 32'h411a5886} /* (0, 15, 2) {real, imag} */,
  {32'hc081b70a, 32'hc08854c5} /* (0, 15, 1) {real, imag} */,
  {32'hbe5cd958, 32'h402991a8} /* (0, 15, 0) {real, imag} */,
  {32'hbfddee9d, 32'h3d6ce880} /* (0, 14, 31) {real, imag} */,
  {32'hc14f2ede, 32'hbcfa4140} /* (0, 14, 30) {real, imag} */,
  {32'hc07e843b, 32'h40099d90} /* (0, 14, 29) {real, imag} */,
  {32'h40e568f4, 32'h40e64bd6} /* (0, 14, 28) {real, imag} */,
  {32'h400d82e9, 32'hc110bf2f} /* (0, 14, 27) {real, imag} */,
  {32'hc08fd1b0, 32'h4067df2a} /* (0, 14, 26) {real, imag} */,
  {32'hc02873ea, 32'hc10dfeb8} /* (0, 14, 25) {real, imag} */,
  {32'h3fabb6bc, 32'hc09baf7f} /* (0, 14, 24) {real, imag} */,
  {32'h4117543b, 32'h40c72560} /* (0, 14, 23) {real, imag} */,
  {32'hc04903ba, 32'hc1a3fa4c} /* (0, 14, 22) {real, imag} */,
  {32'h406850ce, 32'h4055941a} /* (0, 14, 21) {real, imag} */,
  {32'h40e677ec, 32'h3fca7e48} /* (0, 14, 20) {real, imag} */,
  {32'hbf910ed8, 32'hbfc5e6d1} /* (0, 14, 19) {real, imag} */,
  {32'h40b7c2e0, 32'h410ec21c} /* (0, 14, 18) {real, imag} */,
  {32'hc060cec8, 32'hc0814057} /* (0, 14, 17) {real, imag} */,
  {32'h3f6acbd0, 32'hc10dfeda} /* (0, 14, 16) {real, imag} */,
  {32'hc007ce5a, 32'hc0be04d2} /* (0, 14, 15) {real, imag} */,
  {32'h4041fdda, 32'h3e49b6a0} /* (0, 14, 14) {real, imag} */,
  {32'h40b9f2cb, 32'hc0903641} /* (0, 14, 13) {real, imag} */,
  {32'h41277c65, 32'h404319b0} /* (0, 14, 12) {real, imag} */,
  {32'h413951a8, 32'h404a1988} /* (0, 14, 11) {real, imag} */,
  {32'hc0d480df, 32'h40ca639c} /* (0, 14, 10) {real, imag} */,
  {32'hc11cd7b3, 32'hc0d6e5a6} /* (0, 14, 9) {real, imag} */,
  {32'h4011924d, 32'hc116d925} /* (0, 14, 8) {real, imag} */,
  {32'h4109e1c8, 32'hc0b9f2ac} /* (0, 14, 7) {real, imag} */,
  {32'h40896dd9, 32'h3fa15c56} /* (0, 14, 6) {real, imag} */,
  {32'hc06aed0e, 32'hc12b82a8} /* (0, 14, 5) {real, imag} */,
  {32'h3fc91ffe, 32'h40c211f3} /* (0, 14, 4) {real, imag} */,
  {32'h40dfe07b, 32'hc0b1b8f0} /* (0, 14, 3) {real, imag} */,
  {32'hc0af8be0, 32'hc0ebd1c5} /* (0, 14, 2) {real, imag} */,
  {32'hc12dba82, 32'h413069c2} /* (0, 14, 1) {real, imag} */,
  {32'hbf973234, 32'h40a82256} /* (0, 14, 0) {real, imag} */,
  {32'hc06c0cf6, 32'hc124aa5b} /* (0, 13, 31) {real, imag} */,
  {32'h41932189, 32'h40ea3c26} /* (0, 13, 30) {real, imag} */,
  {32'hc13b4432, 32'h40eb22b4} /* (0, 13, 29) {real, imag} */,
  {32'hc01f4ee0, 32'hc129aa18} /* (0, 13, 28) {real, imag} */,
  {32'hbc852a00, 32'hc0a495a1} /* (0, 13, 27) {real, imag} */,
  {32'h40d547a3, 32'hc0a184ae} /* (0, 13, 26) {real, imag} */,
  {32'h40d44ec2, 32'h40d1b25e} /* (0, 13, 25) {real, imag} */,
  {32'hbf7c21a8, 32'h40d5211e} /* (0, 13, 24) {real, imag} */,
  {32'h3fa3fc20, 32'h3fa04528} /* (0, 13, 23) {real, imag} */,
  {32'h40ed362e, 32'hc0bc0318} /* (0, 13, 22) {real, imag} */,
  {32'hc0d8370b, 32'hc0ce7ddc} /* (0, 13, 21) {real, imag} */,
  {32'hc00d2450, 32'hbfd198c6} /* (0, 13, 20) {real, imag} */,
  {32'hc0e4ee0b, 32'h3ffa5cfc} /* (0, 13, 19) {real, imag} */,
  {32'hc12299ff, 32'h414431a4} /* (0, 13, 18) {real, imag} */,
  {32'hc0782996, 32'h4106075f} /* (0, 13, 17) {real, imag} */,
  {32'h40a9d8cc, 32'hbff3633e} /* (0, 13, 16) {real, imag} */,
  {32'h410931e8, 32'h3f853820} /* (0, 13, 15) {real, imag} */,
  {32'hc0f15950, 32'hc0d1732c} /* (0, 13, 14) {real, imag} */,
  {32'h40aae4e4, 32'hc05d25f4} /* (0, 13, 13) {real, imag} */,
  {32'hbf3a666c, 32'h3f8ab2bc} /* (0, 13, 12) {real, imag} */,
  {32'hc0e74fca, 32'h4024fbe2} /* (0, 13, 11) {real, imag} */,
  {32'h416eaa25, 32'h3f870090} /* (0, 13, 10) {real, imag} */,
  {32'hc0832715, 32'h4159868e} /* (0, 13, 9) {real, imag} */,
  {32'h415633b8, 32'hc12af2ad} /* (0, 13, 8) {real, imag} */,
  {32'hc1315e52, 32'h407f6773} /* (0, 13, 7) {real, imag} */,
  {32'h40135c45, 32'hc0a30dc8} /* (0, 13, 6) {real, imag} */,
  {32'h3f8ac577, 32'h3fa01be2} /* (0, 13, 5) {real, imag} */,
  {32'h3f54a6f0, 32'hc1094a27} /* (0, 13, 4) {real, imag} */,
  {32'h4021bf94, 32'h4088b5f2} /* (0, 13, 3) {real, imag} */,
  {32'h3f27aac8, 32'hc0bd4474} /* (0, 13, 2) {real, imag} */,
  {32'h40f8e841, 32'h400f6b7a} /* (0, 13, 1) {real, imag} */,
  {32'hc150aa9e, 32'h41120454} /* (0, 13, 0) {real, imag} */,
  {32'h4097eaae, 32'h416fd661} /* (0, 12, 31) {real, imag} */,
  {32'hc0776348, 32'hc1091bc9} /* (0, 12, 30) {real, imag} */,
  {32'hc03f5527, 32'hc12ea198} /* (0, 12, 29) {real, imag} */,
  {32'hc0ff7558, 32'hbf981770} /* (0, 12, 28) {real, imag} */,
  {32'hc10cc4ce, 32'h3f7f5c10} /* (0, 12, 27) {real, imag} */,
  {32'hc04d6beb, 32'hc0eafc59} /* (0, 12, 26) {real, imag} */,
  {32'h4097d8c8, 32'hc0845798} /* (0, 12, 25) {real, imag} */,
  {32'hc0b29a89, 32'h40ee6bc2} /* (0, 12, 24) {real, imag} */,
  {32'hbfc2d440, 32'h417317e6} /* (0, 12, 23) {real, imag} */,
  {32'h3fd792e7, 32'hbf07b970} /* (0, 12, 22) {real, imag} */,
  {32'h40aee37a, 32'hc0503379} /* (0, 12, 21) {real, imag} */,
  {32'h3ec0d330, 32'h3fe38e80} /* (0, 12, 20) {real, imag} */,
  {32'h416955fa, 32'h409a2e1f} /* (0, 12, 19) {real, imag} */,
  {32'h40d90713, 32'hc009e298} /* (0, 12, 18) {real, imag} */,
  {32'hc064950b, 32'h40e66601} /* (0, 12, 17) {real, imag} */,
  {32'hc036decc, 32'h4067f565} /* (0, 12, 16) {real, imag} */,
  {32'h3fb87988, 32'hc0fe05e2} /* (0, 12, 15) {real, imag} */,
  {32'hc0b7dc10, 32'hc11b09ea} /* (0, 12, 14) {real, imag} */,
  {32'h409d30c5, 32'hc0ec944c} /* (0, 12, 13) {real, imag} */,
  {32'h4081db02, 32'h40f64178} /* (0, 12, 12) {real, imag} */,
  {32'hc16376d2, 32'h3fb6d37d} /* (0, 12, 11) {real, imag} */,
  {32'h40b2803a, 32'hc0a946ec} /* (0, 12, 10) {real, imag} */,
  {32'h4022b5da, 32'hbfa74ca4} /* (0, 12, 9) {real, imag} */,
  {32'h3e96a380, 32'hc1239878} /* (0, 12, 8) {real, imag} */,
  {32'h40c3e9cb, 32'h41311fae} /* (0, 12, 7) {real, imag} */,
  {32'hc0caf0b4, 32'hc094d2d4} /* (0, 12, 6) {real, imag} */,
  {32'hc09a7e45, 32'hc12d2906} /* (0, 12, 5) {real, imag} */,
  {32'hc0890d53, 32'h4112c8ac} /* (0, 12, 4) {real, imag} */,
  {32'h3e604d40, 32'hbedaa400} /* (0, 12, 3) {real, imag} */,
  {32'h41295892, 32'h40bea2dc} /* (0, 12, 2) {real, imag} */,
  {32'h410eb132, 32'hc0d41659} /* (0, 12, 1) {real, imag} */,
  {32'h3f56b808, 32'hc115a892} /* (0, 12, 0) {real, imag} */,
  {32'h413178fe, 32'h3f435440} /* (0, 11, 31) {real, imag} */,
  {32'h4119aab3, 32'hc08ab698} /* (0, 11, 30) {real, imag} */,
  {32'hc10cd5c8, 32'h412b2fb0} /* (0, 11, 29) {real, imag} */,
  {32'hc0fd3084, 32'hc0be8708} /* (0, 11, 28) {real, imag} */,
  {32'hc02ca0d0, 32'hbeadc5e0} /* (0, 11, 27) {real, imag} */,
  {32'h412d1b80, 32'h41103f66} /* (0, 11, 26) {real, imag} */,
  {32'hc033ea35, 32'h402dfd22} /* (0, 11, 25) {real, imag} */,
  {32'h40cd3e85, 32'h412b0f0e} /* (0, 11, 24) {real, imag} */,
  {32'hc00379f0, 32'hc03a598a} /* (0, 11, 23) {real, imag} */,
  {32'h3fd891e0, 32'h3f84e3e0} /* (0, 11, 22) {real, imag} */,
  {32'hc090e220, 32'hc1cbfbb0} /* (0, 11, 21) {real, imag} */,
  {32'h40d997b7, 32'h408c1200} /* (0, 11, 20) {real, imag} */,
  {32'hc05d6290, 32'h40e97720} /* (0, 11, 19) {real, imag} */,
  {32'hc081069c, 32'h411ac822} /* (0, 11, 18) {real, imag} */,
  {32'hbf96fbdc, 32'hc0e0963b} /* (0, 11, 17) {real, imag} */,
  {32'hc04536e2, 32'h408cdd56} /* (0, 11, 16) {real, imag} */,
  {32'hc05e2b16, 32'h40166295} /* (0, 11, 15) {real, imag} */,
  {32'h415922de, 32'hc06fb1ae} /* (0, 11, 14) {real, imag} */,
  {32'hbf9ed97c, 32'hc032b870} /* (0, 11, 13) {real, imag} */,
  {32'hc0bf1264, 32'h419e6e4c} /* (0, 11, 12) {real, imag} */,
  {32'h4113d3dd, 32'hc0788aaf} /* (0, 11, 11) {real, imag} */,
  {32'hc1dbcabc, 32'hc0a7c818} /* (0, 11, 10) {real, imag} */,
  {32'h406c915e, 32'h402091b0} /* (0, 11, 9) {real, imag} */,
  {32'hc014bec8, 32'h40ec6655} /* (0, 11, 8) {real, imag} */,
  {32'h4084aa46, 32'hbf8404ad} /* (0, 11, 7) {real, imag} */,
  {32'h4052335c, 32'hc03f15e8} /* (0, 11, 6) {real, imag} */,
  {32'hc13c1c0e, 32'h40dca805} /* (0, 11, 5) {real, imag} */,
  {32'hc0618ee6, 32'hc12b2984} /* (0, 11, 4) {real, imag} */,
  {32'h40d39569, 32'hc0246088} /* (0, 11, 3) {real, imag} */,
  {32'h4055c0b4, 32'hc140fcdd} /* (0, 11, 2) {real, imag} */,
  {32'h4086507f, 32'hc0827d23} /* (0, 11, 1) {real, imag} */,
  {32'hc03a6690, 32'h3f81b194} /* (0, 11, 0) {real, imag} */,
  {32'hbf883304, 32'hc0216f7e} /* (0, 10, 31) {real, imag} */,
  {32'hbf5e3410, 32'h41082b57} /* (0, 10, 30) {real, imag} */,
  {32'hc089faa3, 32'hc05393fd} /* (0, 10, 29) {real, imag} */,
  {32'hc1197e51, 32'hc114e99f} /* (0, 10, 28) {real, imag} */,
  {32'h417420ec, 32'h40a16d08} /* (0, 10, 27) {real, imag} */,
  {32'hbf9dd44c, 32'h412e7ede} /* (0, 10, 26) {real, imag} */,
  {32'h3f17c970, 32'hc06a99db} /* (0, 10, 25) {real, imag} */,
  {32'h416739a8, 32'hc10964e2} /* (0, 10, 24) {real, imag} */,
  {32'h40d88486, 32'hc13b5b48} /* (0, 10, 23) {real, imag} */,
  {32'hc090570f, 32'hc0c502aa} /* (0, 10, 22) {real, imag} */,
  {32'h404fbbfc, 32'hc0e03e80} /* (0, 10, 21) {real, imag} */,
  {32'h404d83c4, 32'h40f4f3b2} /* (0, 10, 20) {real, imag} */,
  {32'h409af9f8, 32'h3f274830} /* (0, 10, 19) {real, imag} */,
  {32'hc0b12066, 32'hbfeeb666} /* (0, 10, 18) {real, imag} */,
  {32'h3f4d43ec, 32'h3d8fbd00} /* (0, 10, 17) {real, imag} */,
  {32'h4000c70a, 32'hc0ad92bc} /* (0, 10, 16) {real, imag} */,
  {32'hc07cda8c, 32'h40625f92} /* (0, 10, 15) {real, imag} */,
  {32'h40b0295c, 32'hc08f237e} /* (0, 10, 14) {real, imag} */,
  {32'h41329ef4, 32'hc00b6914} /* (0, 10, 13) {real, imag} */,
  {32'hc15c6ba2, 32'hc168ca45} /* (0, 10, 12) {real, imag} */,
  {32'h40a645f5, 32'hc02f4698} /* (0, 10, 11) {real, imag} */,
  {32'h41065f62, 32'hc07ea096} /* (0, 10, 10) {real, imag} */,
  {32'h3fd080fa, 32'hc16af5ae} /* (0, 10, 9) {real, imag} */,
  {32'h4098f172, 32'hc04ffbb4} /* (0, 10, 8) {real, imag} */,
  {32'h408d32b6, 32'hc0387fa8} /* (0, 10, 7) {real, imag} */,
  {32'hbff46e2c, 32'hbf663958} /* (0, 10, 6) {real, imag} */,
  {32'hc056b508, 32'hbeb34c28} /* (0, 10, 5) {real, imag} */,
  {32'h40885a68, 32'hc10568ba} /* (0, 10, 4) {real, imag} */,
  {32'hbfc8e058, 32'h4026387b} /* (0, 10, 3) {real, imag} */,
  {32'h4197403c, 32'h41bef3a2} /* (0, 10, 2) {real, imag} */,
  {32'hc19a8a3c, 32'hbea7da90} /* (0, 10, 1) {real, imag} */,
  {32'h406d1ed8, 32'hc012ae52} /* (0, 10, 0) {real, imag} */,
  {32'h3edc3c28, 32'hc08d45cf} /* (0, 9, 31) {real, imag} */,
  {32'h419e3a69, 32'h4182174f} /* (0, 9, 30) {real, imag} */,
  {32'hc1adc512, 32'h4141766c} /* (0, 9, 29) {real, imag} */,
  {32'hc14ee360, 32'hc18cf41b} /* (0, 9, 28) {real, imag} */,
  {32'h40ecf843, 32'hbf273028} /* (0, 9, 27) {real, imag} */,
  {32'hbf7691a0, 32'hc0dec45f} /* (0, 9, 26) {real, imag} */,
  {32'h411bcfd6, 32'hbf14dd58} /* (0, 9, 25) {real, imag} */,
  {32'h40af73ce, 32'hc128cbb5} /* (0, 9, 24) {real, imag} */,
  {32'h3fc91348, 32'h4056c3f6} /* (0, 9, 23) {real, imag} */,
  {32'hbda84880, 32'h412560ce} /* (0, 9, 22) {real, imag} */,
  {32'hbf161320, 32'h3f71d198} /* (0, 9, 21) {real, imag} */,
  {32'h3f67ee98, 32'hc0c45ea4} /* (0, 9, 20) {real, imag} */,
  {32'h40c5325c, 32'h3ea42578} /* (0, 9, 19) {real, imag} */,
  {32'hc0c26d7d, 32'h4051c736} /* (0, 9, 18) {real, imag} */,
  {32'hc065454f, 32'hc0ca01d3} /* (0, 9, 17) {real, imag} */,
  {32'h4098bb41, 32'hbe808c40} /* (0, 9, 16) {real, imag} */,
  {32'h3fcd0d20, 32'hc01ec486} /* (0, 9, 15) {real, imag} */,
  {32'hc107b8ca, 32'h3dab0560} /* (0, 9, 14) {real, imag} */,
  {32'hbff37254, 32'h3ed4f2a8} /* (0, 9, 13) {real, imag} */,
  {32'h411a2ed5, 32'h41087a14} /* (0, 9, 12) {real, imag} */,
  {32'hc16ce180, 32'h3e624fc0} /* (0, 9, 11) {real, imag} */,
  {32'h40fb4aa0, 32'h4114dc92} /* (0, 9, 10) {real, imag} */,
  {32'hc0dbfd9e, 32'hc0063f86} /* (0, 9, 9) {real, imag} */,
  {32'hbfdff710, 32'h41485cc8} /* (0, 9, 8) {real, imag} */,
  {32'h4056d538, 32'h3fc1c0f2} /* (0, 9, 7) {real, imag} */,
  {32'h41215090, 32'h3faaa520} /* (0, 9, 6) {real, imag} */,
  {32'hbf58159a, 32'h400fc468} /* (0, 9, 5) {real, imag} */,
  {32'hc0191e32, 32'h4102cb4f} /* (0, 9, 4) {real, imag} */,
  {32'hbfe2ccbc, 32'hc1384dc6} /* (0, 9, 3) {real, imag} */,
  {32'h3fbe5a24, 32'h3f4c68c0} /* (0, 9, 2) {real, imag} */,
  {32'hc19d2422, 32'h4087ce90} /* (0, 9, 1) {real, imag} */,
  {32'hc14f06c5, 32'hc088554c} /* (0, 9, 0) {real, imag} */,
  {32'h40cc7b92, 32'h418850e1} /* (0, 8, 31) {real, imag} */,
  {32'hc2064771, 32'hc1069517} /* (0, 8, 30) {real, imag} */,
  {32'hbf3cf3d8, 32'hc09037e1} /* (0, 8, 29) {real, imag} */,
  {32'h417610dc, 32'hc096e9e6} /* (0, 8, 28) {real, imag} */,
  {32'hc080034a, 32'hc0ae6ea0} /* (0, 8, 27) {real, imag} */,
  {32'h40aeaff6, 32'h401deacc} /* (0, 8, 26) {real, imag} */,
  {32'h410b3d56, 32'hc139ac7d} /* (0, 8, 25) {real, imag} */,
  {32'hc17cc5e2, 32'h40b510ec} /* (0, 8, 24) {real, imag} */,
  {32'h413c6d8b, 32'hc08b0487} /* (0, 8, 23) {real, imag} */,
  {32'hc0fce8e5, 32'hc1669015} /* (0, 8, 22) {real, imag} */,
  {32'hc0a9e3f4, 32'h413a7491} /* (0, 8, 21) {real, imag} */,
  {32'hc0bf7d6b, 32'hbfbea540} /* (0, 8, 20) {real, imag} */,
  {32'h40e87837, 32'h40a1c36d} /* (0, 8, 19) {real, imag} */,
  {32'h412d80d0, 32'hc08ca485} /* (0, 8, 18) {real, imag} */,
  {32'hc0498d65, 32'hc0147032} /* (0, 8, 17) {real, imag} */,
  {32'hbf31fc00, 32'hc135419e} /* (0, 8, 16) {real, imag} */,
  {32'h405755f0, 32'h3f4c52b0} /* (0, 8, 15) {real, imag} */,
  {32'h40dc36e6, 32'h4152eba7} /* (0, 8, 14) {real, imag} */,
  {32'hc04350fc, 32'h410e22ae} /* (0, 8, 13) {real, imag} */,
  {32'hc0b5ab09, 32'hc0ab1723} /* (0, 8, 12) {real, imag} */,
  {32'h4110954c, 32'hc0c322b9} /* (0, 8, 11) {real, imag} */,
  {32'hc1363392, 32'h40329500} /* (0, 8, 10) {real, imag} */,
  {32'hc00960bc, 32'hbf819d68} /* (0, 8, 9) {real, imag} */,
  {32'h4062c7ba, 32'hbf503f30} /* (0, 8, 8) {real, imag} */,
  {32'h40e8aebc, 32'h413c7027} /* (0, 8, 7) {real, imag} */,
  {32'hc1276a7e, 32'hc1049026} /* (0, 8, 6) {real, imag} */,
  {32'h40fd9973, 32'hc0dd3c6a} /* (0, 8, 5) {real, imag} */,
  {32'h401dca6a, 32'h4013c4b8} /* (0, 8, 4) {real, imag} */,
  {32'hc181de38, 32'h40847694} /* (0, 8, 3) {real, imag} */,
  {32'hc1895349, 32'h40899336} /* (0, 8, 2) {real, imag} */,
  {32'h3f9c3980, 32'h41a15289} /* (0, 8, 1) {real, imag} */,
  {32'h41b1299e, 32'h4195be20} /* (0, 8, 0) {real, imag} */,
  {32'hc0a28002, 32'h411cad96} /* (0, 7, 31) {real, imag} */,
  {32'h4135eefe, 32'h3c7e4400} /* (0, 7, 30) {real, imag} */,
  {32'hc0f7c858, 32'h4188692d} /* (0, 7, 29) {real, imag} */,
  {32'h4115bab6, 32'h4159c31b} /* (0, 7, 28) {real, imag} */,
  {32'hc0a52ca6, 32'hc0439573} /* (0, 7, 27) {real, imag} */,
  {32'hc0ad4f6c, 32'h3f5dc930} /* (0, 7, 26) {real, imag} */,
  {32'h4049718e, 32'hbf058ea8} /* (0, 7, 25) {real, imag} */,
  {32'h4088ba00, 32'hc095ea24} /* (0, 7, 24) {real, imag} */,
  {32'hbfe621b4, 32'hbf0ceee0} /* (0, 7, 23) {real, imag} */,
  {32'h405c391c, 32'hc0b8618f} /* (0, 7, 22) {real, imag} */,
  {32'h40c0076c, 32'hbf2f30f0} /* (0, 7, 21) {real, imag} */,
  {32'h3c23a800, 32'hbfd0d9da} /* (0, 7, 20) {real, imag} */,
  {32'hbea127e0, 32'h40d5de2a} /* (0, 7, 19) {real, imag} */,
  {32'hc10ec66e, 32'hbfd05e94} /* (0, 7, 18) {real, imag} */,
  {32'hc0aec7b8, 32'h4034d5c0} /* (0, 7, 17) {real, imag} */,
  {32'hc0439498, 32'hc10d5fe4} /* (0, 7, 16) {real, imag} */,
  {32'hbdf53800, 32'h40780a80} /* (0, 7, 15) {real, imag} */,
  {32'h40d3a96e, 32'hc081df98} /* (0, 7, 14) {real, imag} */,
  {32'hbd895340, 32'h41161296} /* (0, 7, 13) {real, imag} */,
  {32'hc0b2a501, 32'h4112f19e} /* (0, 7, 12) {real, imag} */,
  {32'h40d143f1, 32'h40341e54} /* (0, 7, 11) {real, imag} */,
  {32'hc0bb40a9, 32'hc0d4bbe8} /* (0, 7, 10) {real, imag} */,
  {32'h40d18d0e, 32'h40b54ca8} /* (0, 7, 9) {real, imag} */,
  {32'hc01e525e, 32'hc0d60bf1} /* (0, 7, 8) {real, imag} */,
  {32'hc11da280, 32'hc004d830} /* (0, 7, 7) {real, imag} */,
  {32'hc1617a78, 32'h4110177a} /* (0, 7, 6) {real, imag} */,
  {32'h4112a3c2, 32'h4129f5e2} /* (0, 7, 5) {real, imag} */,
  {32'h40bbdf66, 32'h3f769778} /* (0, 7, 4) {real, imag} */,
  {32'h40c5e34e, 32'hc091ed56} /* (0, 7, 3) {real, imag} */,
  {32'hc174a89c, 32'hc12e7ef2} /* (0, 7, 2) {real, imag} */,
  {32'h41d96da6, 32'hc1c87663} /* (0, 7, 1) {real, imag} */,
  {32'hc057ffec, 32'hc120a24c} /* (0, 7, 0) {real, imag} */,
  {32'hc0022fbc, 32'h41819710} /* (0, 6, 31) {real, imag} */,
  {32'hc1ce89bd, 32'h419e2916} /* (0, 6, 30) {real, imag} */,
  {32'h410488b7, 32'hc1e38a55} /* (0, 6, 29) {real, imag} */,
  {32'hc0a96ee3, 32'h415cf7c7} /* (0, 6, 28) {real, imag} */,
  {32'h41838458, 32'hc0e5e4a5} /* (0, 6, 27) {real, imag} */,
  {32'h3ff95568, 32'h40a5c11a} /* (0, 6, 26) {real, imag} */,
  {32'h412a21b2, 32'h406a7ee0} /* (0, 6, 25) {real, imag} */,
  {32'hbf7a254c, 32'hc0a9e5ad} /* (0, 6, 24) {real, imag} */,
  {32'h40fd5bbc, 32'hc0283170} /* (0, 6, 23) {real, imag} */,
  {32'hc0418b20, 32'hc0919bd7} /* (0, 6, 22) {real, imag} */,
  {32'h41027bd2, 32'hbeea96f8} /* (0, 6, 21) {real, imag} */,
  {32'h40bae08d, 32'h3ee32920} /* (0, 6, 20) {real, imag} */,
  {32'h40c2233c, 32'hc0837bce} /* (0, 6, 19) {real, imag} */,
  {32'h3fd86e88, 32'h3f456300} /* (0, 6, 18) {real, imag} */,
  {32'h40c17bbd, 32'h3e0a4338} /* (0, 6, 17) {real, imag} */,
  {32'h3fbf7191, 32'h40bc1f6a} /* (0, 6, 16) {real, imag} */,
  {32'hc04f2eee, 32'hc05bb8f9} /* (0, 6, 15) {real, imag} */,
  {32'hc1399698, 32'h4145a30d} /* (0, 6, 14) {real, imag} */,
  {32'h3f5b65c0, 32'hc0c133c4} /* (0, 6, 13) {real, imag} */,
  {32'hbec7f460, 32'h410c3284} /* (0, 6, 12) {real, imag} */,
  {32'hc00182cc, 32'h4103ac96} /* (0, 6, 11) {real, imag} */,
  {32'hc0f15624, 32'h41603869} /* (0, 6, 10) {real, imag} */,
  {32'h410145e6, 32'hc08af1ed} /* (0, 6, 9) {real, imag} */,
  {32'h3f81fe79, 32'hc10c96dc} /* (0, 6, 8) {real, imag} */,
  {32'h40553024, 32'h409c772a} /* (0, 6, 7) {real, imag} */,
  {32'hc145b992, 32'h40891e86} /* (0, 6, 6) {real, imag} */,
  {32'hc0cce642, 32'hc0264dfd} /* (0, 6, 5) {real, imag} */,
  {32'h418716b4, 32'hc10eb088} /* (0, 6, 4) {real, imag} */,
  {32'h41550ada, 32'h40345c6d} /* (0, 6, 3) {real, imag} */,
  {32'hc05c1a98, 32'hc0eeb2bc} /* (0, 6, 2) {real, imag} */,
  {32'hc0eb36e7, 32'hc0b0d796} /* (0, 6, 1) {real, imag} */,
  {32'hc026a99e, 32'hc1fc7d9c} /* (0, 6, 0) {real, imag} */,
  {32'h420ebaf4, 32'hc13e497d} /* (0, 5, 31) {real, imag} */,
  {32'hc1ad3a30, 32'h40e17768} /* (0, 5, 30) {real, imag} */,
  {32'hc18b99ef, 32'h414b6c8e} /* (0, 5, 29) {real, imag} */,
  {32'h41423f02, 32'h3f9bbcb8} /* (0, 5, 28) {real, imag} */,
  {32'h4098191d, 32'h4108a1b4} /* (0, 5, 27) {real, imag} */,
  {32'h412bec51, 32'h408adcee} /* (0, 5, 26) {real, imag} */,
  {32'hc0b6de07, 32'h3e0e9f00} /* (0, 5, 25) {real, imag} */,
  {32'hc03e4454, 32'hc1563453} /* (0, 5, 24) {real, imag} */,
  {32'h408373c4, 32'h3fe82520} /* (0, 5, 23) {real, imag} */,
  {32'hc14a591c, 32'h41084caf} /* (0, 5, 22) {real, imag} */,
  {32'hc1721631, 32'hc09a8403} /* (0, 5, 21) {real, imag} */,
  {32'hc0d93810, 32'hc0b84952} /* (0, 5, 20) {real, imag} */,
  {32'h40a9dc56, 32'h3f9396f8} /* (0, 5, 19) {real, imag} */,
  {32'hc0e73106, 32'h411b38c9} /* (0, 5, 18) {real, imag} */,
  {32'hbfb2b73a, 32'hc0860916} /* (0, 5, 17) {real, imag} */,
  {32'hbfd72b74, 32'h40bf6484} /* (0, 5, 16) {real, imag} */,
  {32'h40bb2a26, 32'hc0a15a44} /* (0, 5, 15) {real, imag} */,
  {32'h40dc2cb4, 32'hc06d3b7d} /* (0, 5, 14) {real, imag} */,
  {32'h409ef95f, 32'h40df9f68} /* (0, 5, 13) {real, imag} */,
  {32'hc0c87ffa, 32'h3fcc1718} /* (0, 5, 12) {real, imag} */,
  {32'hbe1c2280, 32'hc12e8819} /* (0, 5, 11) {real, imag} */,
  {32'hc0c517f8, 32'h40a691d6} /* (0, 5, 10) {real, imag} */,
  {32'h409e367b, 32'hc037d278} /* (0, 5, 9) {real, imag} */,
  {32'h3e9bd958, 32'h3dcc4700} /* (0, 5, 8) {real, imag} */,
  {32'h41399b89, 32'h402f1e4e} /* (0, 5, 7) {real, imag} */,
  {32'hc1597cb2, 32'h40b82e02} /* (0, 5, 6) {real, imag} */,
  {32'h40b3d0be, 32'h40bf2f64} /* (0, 5, 5) {real, imag} */,
  {32'hc0bca84a, 32'h416db3a4} /* (0, 5, 4) {real, imag} */,
  {32'hc12ff2a9, 32'hc11e4730} /* (0, 5, 3) {real, imag} */,
  {32'h413ddea6, 32'hc15cdc75} /* (0, 5, 2) {real, imag} */,
  {32'hc1198fdb, 32'h41d7dc4d} /* (0, 5, 1) {real, imag} */,
  {32'h41ef0010, 32'hc03baf20} /* (0, 5, 0) {real, imag} */,
  {32'hc1dafaea, 32'hc1881c40} /* (0, 4, 31) {real, imag} */,
  {32'hc08e65d8, 32'h4228d210} /* (0, 4, 30) {real, imag} */,
  {32'hc1363d48, 32'hc103d145} /* (0, 4, 29) {real, imag} */,
  {32'hc0a49ea4, 32'h4104c117} /* (0, 4, 28) {real, imag} */,
  {32'hbfc81890, 32'hc0e1c18b} /* (0, 4, 27) {real, imag} */,
  {32'h3fd66aa0, 32'hc11ad78c} /* (0, 4, 26) {real, imag} */,
  {32'h41ccb336, 32'h418bce38} /* (0, 4, 25) {real, imag} */,
  {32'hc02f0890, 32'hc18a6271} /* (0, 4, 24) {real, imag} */,
  {32'hc191d060, 32'hc16f9dcf} /* (0, 4, 23) {real, imag} */,
  {32'hc0850e62, 32'h3f8eb1b6} /* (0, 4, 22) {real, imag} */,
  {32'h40464a1a, 32'hc007eb44} /* (0, 4, 21) {real, imag} */,
  {32'hc0ec5250, 32'h40e6bfde} /* (0, 4, 20) {real, imag} */,
  {32'hc12a9756, 32'h40ca0ea1} /* (0, 4, 19) {real, imag} */,
  {32'h3fe51bad, 32'h41303466} /* (0, 4, 18) {real, imag} */,
  {32'hc02ba366, 32'hc04064af} /* (0, 4, 17) {real, imag} */,
  {32'h40a7c95a, 32'hc09e68fa} /* (0, 4, 16) {real, imag} */,
  {32'hbf6f2788, 32'hbf88e8af} /* (0, 4, 15) {real, imag} */,
  {32'hc05a7a3a, 32'h40eefe3a} /* (0, 4, 14) {real, imag} */,
  {32'h3fecef18, 32'h3f28af5c} /* (0, 4, 13) {real, imag} */,
  {32'h4044ab8b, 32'hc0163b42} /* (0, 4, 12) {real, imag} */,
  {32'hc08d3248, 32'h4137699d} /* (0, 4, 11) {real, imag} */,
  {32'h41662196, 32'h40b933a0} /* (0, 4, 10) {real, imag} */,
  {32'h40ba30ce, 32'h40e4d338} /* (0, 4, 9) {real, imag} */,
  {32'h4128080e, 32'h3f0e2758} /* (0, 4, 8) {real, imag} */,
  {32'hc1248d1c, 32'hc1874adc} /* (0, 4, 7) {real, imag} */,
  {32'hc0601044, 32'h4042bed8} /* (0, 4, 6) {real, imag} */,
  {32'h411ecd13, 32'hbf108ab8} /* (0, 4, 5) {real, imag} */,
  {32'h3e6f90c0, 32'h3f6e57e0} /* (0, 4, 4) {real, imag} */,
  {32'h40f011c4, 32'h42005571} /* (0, 4, 3) {real, imag} */,
  {32'h41a8f9f0, 32'h41f9347e} /* (0, 4, 2) {real, imag} */,
  {32'hc23201f0, 32'h4142a4a8} /* (0, 4, 1) {real, imag} */,
  {32'h41b44f1b, 32'hc13f2c90} /* (0, 4, 0) {real, imag} */,
  {32'h4233a764, 32'hc0e3c504} /* (0, 3, 31) {real, imag} */,
  {32'hc19e0af6, 32'h4186614a} /* (0, 3, 30) {real, imag} */,
  {32'h41a33db4, 32'h414f82f2} /* (0, 3, 29) {real, imag} */,
  {32'hc144cc1f, 32'hc0908fb3} /* (0, 3, 28) {real, imag} */,
  {32'h41766c44, 32'hc180d3a8} /* (0, 3, 27) {real, imag} */,
  {32'h3f68ed32, 32'h408d7896} /* (0, 3, 26) {real, imag} */,
  {32'hbfbe1d08, 32'hc13338ee} /* (0, 3, 25) {real, imag} */,
  {32'h40e592e6, 32'h41432a4e} /* (0, 3, 24) {real, imag} */,
  {32'hc0a74892, 32'h3cfd0b40} /* (0, 3, 23) {real, imag} */,
  {32'hc0e5b4d7, 32'hc08f8d13} /* (0, 3, 22) {real, imag} */,
  {32'hc0b0606e, 32'h40874786} /* (0, 3, 21) {real, imag} */,
  {32'hc108847e, 32'h408f7f18} /* (0, 3, 20) {real, imag} */,
  {32'h3e27c4c0, 32'h40f46267} /* (0, 3, 19) {real, imag} */,
  {32'hc129fc0a, 32'h404f693f} /* (0, 3, 18) {real, imag} */,
  {32'h4077e26c, 32'hc046c0ce} /* (0, 3, 17) {real, imag} */,
  {32'h3dd85e60, 32'h40f64c0b} /* (0, 3, 16) {real, imag} */,
  {32'h405a3198, 32'hbf562a30} /* (0, 3, 15) {real, imag} */,
  {32'hc1203e7d, 32'hbe51d0b0} /* (0, 3, 14) {real, imag} */,
  {32'hc05d2074, 32'hc0c56582} /* (0, 3, 13) {real, imag} */,
  {32'h41452218, 32'h3fdb2794} /* (0, 3, 12) {real, imag} */,
  {32'h40c86d54, 32'h409ab7b3} /* (0, 3, 11) {real, imag} */,
  {32'h407fded0, 32'h3f8f6e84} /* (0, 3, 10) {real, imag} */,
  {32'h3f97a1b0, 32'hc11885db} /* (0, 3, 9) {real, imag} */,
  {32'h410c4836, 32'h3f43eca8} /* (0, 3, 8) {real, imag} */,
  {32'hc1c57eec, 32'hc025fdee} /* (0, 3, 7) {real, imag} */,
  {32'hc1337fe9, 32'hc174799d} /* (0, 3, 6) {real, imag} */,
  {32'hc10dcb31, 32'h412c67e3} /* (0, 3, 5) {real, imag} */,
  {32'h4196c8c0, 32'h41ff74dc} /* (0, 3, 4) {real, imag} */,
  {32'h412f456d, 32'hc1db544e} /* (0, 3, 3) {real, imag} */,
  {32'hc1b70cdb, 32'h425bd312} /* (0, 3, 2) {real, imag} */,
  {32'hc182c6cb, 32'hc21ab240} /* (0, 3, 1) {real, imag} */,
  {32'h41de95d2, 32'h415052ca} /* (0, 3, 0) {real, imag} */,
  {32'h43744033, 32'h41062dad} /* (0, 2, 31) {real, imag} */,
  {32'hc2fbb0a2, 32'h408d3768} /* (0, 2, 30) {real, imag} */,
  {32'h4165c05c, 32'hc1ddefee} /* (0, 2, 29) {real, imag} */,
  {32'h41561c24, 32'hc0ce82a8} /* (0, 2, 28) {real, imag} */,
  {32'hc19ec512, 32'h420ea3fe} /* (0, 2, 27) {real, imag} */,
  {32'hc0ab37a6, 32'h41475e7f} /* (0, 2, 26) {real, imag} */,
  {32'hbfa59288, 32'h410f07cc} /* (0, 2, 25) {real, imag} */,
  {32'hc12c923b, 32'h4168ff5c} /* (0, 2, 24) {real, imag} */,
  {32'h3eaa9ca0, 32'h3ffd2270} /* (0, 2, 23) {real, imag} */,
  {32'h3fffac9e, 32'h3fd18d80} /* (0, 2, 22) {real, imag} */,
  {32'hc0a5812b, 32'hc0ab840c} /* (0, 2, 21) {real, imag} */,
  {32'hc10dc2ff, 32'h4015b914} /* (0, 2, 20) {real, imag} */,
  {32'hc00fdfd8, 32'h3eab661c} /* (0, 2, 19) {real, imag} */,
  {32'h3f98607a, 32'hbe950cc8} /* (0, 2, 18) {real, imag} */,
  {32'h3fa166da, 32'h4065dc8d} /* (0, 2, 17) {real, imag} */,
  {32'h40066a5d, 32'h3ec2bb98} /* (0, 2, 16) {real, imag} */,
  {32'h41394f7b, 32'hc008a388} /* (0, 2, 15) {real, imag} */,
  {32'hbfe4927c, 32'hc0c22bf2} /* (0, 2, 14) {real, imag} */,
  {32'hc12c2314, 32'hbdd147c0} /* (0, 2, 13) {real, imag} */,
  {32'h40940a1a, 32'hc154c76c} /* (0, 2, 12) {real, imag} */,
  {32'hc029148e, 32'hc19a7ce4} /* (0, 2, 11) {real, imag} */,
  {32'hc09f318b, 32'hc0f33898} /* (0, 2, 10) {real, imag} */,
  {32'hc0d7c989, 32'hc097beb0} /* (0, 2, 9) {real, imag} */,
  {32'hc1d78e4e, 32'hc1276c4c} /* (0, 2, 8) {real, imag} */,
  {32'h41353c14, 32'h400fd624} /* (0, 2, 7) {real, imag} */,
  {32'h41865b1a, 32'h413c831f} /* (0, 2, 6) {real, imag} */,
  {32'hc1c14726, 32'hc1fd7cca} /* (0, 2, 5) {real, imag} */,
  {32'h426b503f, 32'h412b9a7c} /* (0, 2, 4) {real, imag} */,
  {32'hc101ae78, 32'hc1b2e1fd} /* (0, 2, 3) {real, imag} */,
  {32'hc2ba574a, 32'h425c7406} /* (0, 2, 2) {real, imag} */,
  {32'h42a05470, 32'h41a1e13a} /* (0, 2, 1) {real, imag} */,
  {32'h42ad914c, 32'h41b351a6} /* (0, 2, 0) {real, imag} */,
  {32'hc340868e, 32'hc0d4e948} /* (0, 1, 31) {real, imag} */,
  {32'h427d3b82, 32'hc152b7fe} /* (0, 1, 30) {real, imag} */,
  {32'h41ee39b6, 32'h3ee5b580} /* (0, 1, 29) {real, imag} */,
  {32'hc20ab738, 32'hbfef9e20} /* (0, 1, 28) {real, imag} */,
  {32'h427c6b5a, 32'h4152b368} /* (0, 1, 27) {real, imag} */,
  {32'hbf181580, 32'h40aac079} /* (0, 1, 26) {real, imag} */,
  {32'hc0934e91, 32'hc0eace5c} /* (0, 1, 25) {real, imag} */,
  {32'h408c6d49, 32'hc1455d3b} /* (0, 1, 24) {real, imag} */,
  {32'h41652414, 32'hc182562b} /* (0, 1, 23) {real, imag} */,
  {32'hc1026137, 32'h412dc5ba} /* (0, 1, 22) {real, imag} */,
  {32'h411387d7, 32'hc181534a} /* (0, 1, 21) {real, imag} */,
  {32'hbfb1340a, 32'h415a5d96} /* (0, 1, 20) {real, imag} */,
  {32'h3f0f7db8, 32'hc0945df1} /* (0, 1, 19) {real, imag} */,
  {32'h40bec258, 32'hbfd84e8a} /* (0, 1, 18) {real, imag} */,
  {32'h3fd3c3fc, 32'hc0e56e7c} /* (0, 1, 17) {real, imag} */,
  {32'h40164b88, 32'hc045bb2c} /* (0, 1, 16) {real, imag} */,
  {32'h40d1671a, 32'h3f635cb4} /* (0, 1, 15) {real, imag} */,
  {32'hc09b913e, 32'hc0010da8} /* (0, 1, 14) {real, imag} */,
  {32'h40eb60be, 32'hc0d65758} /* (0, 1, 13) {real, imag} */,
  {32'hc011da41, 32'hc08e09c6} /* (0, 1, 12) {real, imag} */,
  {32'h417d81e2, 32'hbfca66d0} /* (0, 1, 11) {real, imag} */,
  {32'hc0baef38, 32'hc0e8e6e2} /* (0, 1, 10) {real, imag} */,
  {32'hc035966f, 32'hc09c186a} /* (0, 1, 9) {real, imag} */,
  {32'hc0495710, 32'h418ae0d9} /* (0, 1, 8) {real, imag} */,
  {32'hc0c92e41, 32'hc0e13823} /* (0, 1, 7) {real, imag} */,
  {32'h417e81df, 32'h40e8c852} /* (0, 1, 6) {real, imag} */,
  {32'h419b3910, 32'h4152d494} /* (0, 1, 5) {real, imag} */,
  {32'h417fe53b, 32'hc182d502} /* (0, 1, 4) {real, imag} */,
  {32'h424ebd20, 32'hc029676e} /* (0, 1, 3) {real, imag} */,
  {32'h42b2ad2b, 32'h4258411c} /* (0, 1, 2) {real, imag} */,
  {32'hc3a10d46, 32'hc383b8de} /* (0, 1, 1) {real, imag} */,
  {32'hc35a7e04, 32'h42a3a2bb} /* (0, 1, 0) {real, imag} */,
  {32'hc31d55bc, 32'h42bb5f38} /* (0, 0, 31) {real, imag} */,
  {32'hc1b20c7b, 32'h41c2d454} /* (0, 0, 30) {real, imag} */,
  {32'h4181198f, 32'h40bd7522} /* (0, 0, 29) {real, imag} */,
  {32'hc1962c74, 32'hc1e4475a} /* (0, 0, 28) {real, imag} */,
  {32'h425de962, 32'h409430e4} /* (0, 0, 27) {real, imag} */,
  {32'hc0ac66be, 32'hc177e7cb} /* (0, 0, 26) {real, imag} */,
  {32'hc19c3a57, 32'h4177d1f7} /* (0, 0, 25) {real, imag} */,
  {32'hbe0e3780, 32'hc14e46c3} /* (0, 0, 24) {real, imag} */,
  {32'h4121b702, 32'h4045463f} /* (0, 0, 23) {real, imag} */,
  {32'hc09c0618, 32'h41224160} /* (0, 0, 22) {real, imag} */,
  {32'h4050d97c, 32'h40648f5e} /* (0, 0, 21) {real, imag} */,
  {32'h40f4146c, 32'h41435b98} /* (0, 0, 20) {real, imag} */,
  {32'hc0f409a4, 32'hbfc8477d} /* (0, 0, 19) {real, imag} */,
  {32'h41029ec4, 32'hc1256217} /* (0, 0, 18) {real, imag} */,
  {32'hc0df606a, 32'hc04ad3e3} /* (0, 0, 17) {real, imag} */,
  {32'hbfd9867a, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'hc0df606a, 32'h404ad3e3} /* (0, 0, 15) {real, imag} */,
  {32'h41029ec4, 32'h41256217} /* (0, 0, 14) {real, imag} */,
  {32'hc0f409a4, 32'h3fc8477d} /* (0, 0, 13) {real, imag} */,
  {32'h40f4146c, 32'hc1435b98} /* (0, 0, 12) {real, imag} */,
  {32'h4050d97c, 32'hc0648f5e} /* (0, 0, 11) {real, imag} */,
  {32'hc09c0618, 32'hc1224160} /* (0, 0, 10) {real, imag} */,
  {32'h4121b702, 32'hc045463f} /* (0, 0, 9) {real, imag} */,
  {32'hbe0e3780, 32'h414e46c3} /* (0, 0, 8) {real, imag} */,
  {32'hc19c3a57, 32'hc177d1f7} /* (0, 0, 7) {real, imag} */,
  {32'hc0ac66be, 32'h4177e7cb} /* (0, 0, 6) {real, imag} */,
  {32'h425de962, 32'hc09430e4} /* (0, 0, 5) {real, imag} */,
  {32'hc1962c74, 32'h41e4475a} /* (0, 0, 4) {real, imag} */,
  {32'h4181198f, 32'hc0bd7522} /* (0, 0, 3) {real, imag} */,
  {32'hc1b20c7b, 32'hc1c2d454} /* (0, 0, 2) {real, imag} */,
  {32'hc31d55bc, 32'hc2bb5f38} /* (0, 0, 1) {real, imag} */,
  {32'hc3085967, 32'h00000000} /* (0, 0, 0) {real, imag} */};
