-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
J6mUXaCF2Yz6sBoNMHD80aMGWWxNBLXjuU6+pnRJpW6p6IaOqReJTLfS5/k9fkD+
3IEziAo6Ge+6Xq8LHZfOOX4KI+06BXBYacOWA2PSMiuNvxu55AqDFp4yi+HLAMQi
rIwVbD85oeeTf/T0VOsBn32isVr6k8qrxNGVz+8WGv1xtz+sWE3/cw==
--pragma protect end_key_block
--pragma protect digest_block
PlSv+B3kvSFvA15k6VhLM0shH28=
--pragma protect end_digest_block
--pragma protect data_block
tgVdyY9a2KrOTmXinviSUdh2DNWp4bPCc9+ilGXSwpMm8eFb01Q8feRlLksEDpbW
/6Xe/f3hXelPzf2R7V1r9UWXwBTyQ8ww3xIU4gf4Bb3gidQ6XPeWmRRbecIvsI6n
L+HXzKclcNiudj2xqPEsrk/CQ2MJSxXOUwoAaoCocYYMevZjmGuW2QluziS2qwUF
U11bCjVXTLrD8m4r627suMtfmSP5G/dbm2LXJO+2ozs/uAwi3Gonf8boEgOsKXZR
44u9B+p3bl1sKGpLJZxWbTnd4cR/WmW7bE0vUn5atByUpKpqmceoQ5E5Gqe2m9H+
3n7OuMEBizGIiKgFGBA2oCm7zLnk+6CM8dzugI5xBwrXaX0Q/uC//TXsjC+8+mb3
58mRfg2f2zFUE8Rexg/pzKidVmaWjoWptZzj0nqtyJfz1cH6rVHAx/SLCKs3m/bY
F1N0QtGp4NtmfzpOQvB8zbkZNCsbEpn3SvZGDO0zqI9L6FVj15j89REHpOfd8pdF
QNi53fKtW0svTNN0Sc/qA7nN/r2SwXtXrrK6h1MZjwSTJY4MrAI62y3S5unvUbiH
wvLBnduBPuavN4x1H+oRvEhs4RlDteGXBSFA0jXOH+nDnd5tcuRbspWWC+DXkRjT
V8NYOUE/V3GmzJDVpKCi0AjAKEP8qFX0zceP8C4iGlFlZWbUQEa3NzU0ghAEZ+2h
RvCH5l+K/+Is3oPEVH4AWwfWDBWAdUJh2V2jHvg/ssl5bVNYemp+kY8MMFCYIiMr
AqhhFzmRD9+BdcwqAxNXFhPrk7GESt2WAjjGzGDJht90s+hvV/C+C8t7dyTU/VmU
cJ4qm6Dhd0Viae7pCtH9kCX0ua0pBASCxWYVF5qBdpdadmWolpZKOeJ96fu4TZ4W
5+k0oZhSfhG+CPGcNllQLhA4HnhpxLXYncHItU4z8iJcUL+fGFb1eqd8aZSLDz06
ZRtPbP2HpKcjifJl3dZqr43umJltznOoMpZoY2Lga96WLIQYGEQfVD8gSfiHk5pK
mPW6+m47oGezMA3QQUecetgqZ9L7jCDGQk8ZA1DnstPYGyPLFumDFAgjsnGXISaQ
LjBXmMAUTBQep2GbsjHi2vUFrda8ZrqAqXs6lvbddNINT98emesQUWCHNCjSSy3U
VhzzfEhKXp4KWOjpYIV53W5vcgZxXFiSh+7h6I7NOVZgmIK8zBmgYzy/jfodQQP9
7ZJk2iICwvDnaOxjrOvv/TO2zG8cgn6rh9jXIFE7Z9DYAA6m/3G0zGLnHKDEdpK7
+BrSvrsVywU3HPrBpu6RiUQjepKdPjzTClI5Zf+v+URibfoetAKUltRnyqO5+cag
ZDwK3ky0zzrDAD2umLrhrKkAscBfPl0PuRmE9iaBIBXHed0m3sSpOgrL6WjLwNnm
xceaYB5QvnhLFmrve8rlpfYnuGEK5rFDNTZ2d9xb5K0Rhu+gnMQ5HUhsDAzdnELT
Lp3mH3EV4hEDV1Uc+8zuLyeSl6+aD7s4BzdXNJarRlKhi5gQItyQ29hI38z3VXyq
543TmtYPakvZHPlwDRowGsXE+KJHsNwuL8YmjMyom7fZGYkc5I1QTiwkeR39fPPf
H8vYWauXbEDd5I46oNl49m2/zbGwbHq+iY3mpatsQH1bFiAcDSIjX6x7Jkn4WZMs
H8uKmkv0oNGDB96udUETXvwkZxBf78L267F1GcY2YUhejc+D6HJcE14RxKULIG9F
9Yp6KkRAasv7Pi24KLgpAhtZNpRNn5c2b+PC1uSgdiP6RhF7DGbMgW27+t2ZgvKv
trrQxSJycC9JhGldq39TlYS9DhYQihG3tcHRZd/tK/R5O2RPLFuB2ugcztNWM8zf
YHkrMzWtUDKxG85WU6EDNJaJxbVIOn2pfsmIffOI5+qhYx8NVdrCiO7Q4q9Et0XZ
Co9X9drFPvOaekB31AtTEL0u4A83bhGNXfb56RrYqYM7Hz8Zm0WfnQVPS0PbRmTP
w4x4fpGHa3ihHzyzGmeN6DCFCvIHf9x8Dc9yKAkb/Ps9CIi5S6R7CpQFGpHWnBj0
p1U1SeYmsf1EASPUFb6Liy0GPpPv0AGLN2+UYoCTgsxhu4O92bbBZ8x++m1J8O+q
WJKCEcZqLFVp5CKqC+sGB0AxY0y+s2hxeT/F9S6LzyUbC/BDt+VRdV79zieMTir4
6tcDuIW3NQc1SXiitxNqgE8TmwKgd4SqzVRMF+/MdPPiBHS2GEqb37ykc2DPz7PN
/dOpw4Mze12n603t9Ph0Hz8lxDkUEbcVOsU8VSslQBzRkqS26FLglcSI2BYICuM6
gNqotlooze6Ld24IUjtDBmXtRYocbfMvvA3zQ8TStefDTpRFJ0pYSWGKV38JKxCt
C2OhxUcLR0jJgr7xDym1QliPb9GDmfROFFtfDI11H7nQCl+LMGzqC4+Ch89kKVvh
kCXdHpv73h2Huobijtesru9QBORtQB7KCmrLvNgP+iKhIMbjWeNDev9eJKedPue+
2MH2nDlEtd78fwOT+jrJyipvlykHZG4AOCyT1LunP+GgI4EcXR7kvJm3vThDBInB
onEQ5G3AcTCMEOrweXTR1ZXFGwptiZvqmf7a5kGBWSjX85/njnGeXyJJq5mwxBub
zhwp5yr5jUp4iBDSqGDOYX9NDl0mxOw8BVzbxiiVBsyhTrROJUinxuhWT4o+Hzs1
aDt+YcXPWO3JbiR5KwBo8buCdnhXCx+LDN97YbNZYMTc8Jb4rR6WdjvSWP9Zrwn2
v+IoGk4usrFw9LlhJipHfiTk9a23AGV5R+fjzuNkS0LR7zx3EBtrplnUdggf04AH
YSrBTA+Luj52U8qMlYjvxagyjYCEnMsxMWzOvHbNtgoztl0WH+hCkQg5LV90Cnoz
gM6qYwFwzxJ9y7+QBvoPuPFQoa4cF56ILY1xA4L5aHuznxFjSKg8vD1uE8t13ecG
+9iigNYzLqGW835pinSbTBTOC29wyL/mXz7QlrzShJjmdMGQ3JSvD2I4h3GDeu1v
xQHpBokQGdb2e80KylbxLqaaU61+rrdJBL8+bi59Q7WAZiK7P42TnpIYpdNLcmNj
7MFIvXIC3O+J9Dg6M9p/BnpR4VQqcQk/JVaLPWp6+k0MGdrjxa8DR+yGdreBqf9L
MogfCsWkQs5hPsL9237NhbUtnbOUIrTma5ieAk5yuzV3le1ImWSoKv6P4brQjGLT
FT7K7blDUlNVXVhLUIHAdAPZROQLRm8Y7E654/DyZsKUxYQMdEnjMHoXAy59IHD5
BYBEwSN6REb6JIzDAwvCo/Mp1M57+7TnnIgIVLZNbTLMGP6R6fyOJdUOK21O3uFG
FD6gxiVfLus+6BYoHyDlNCSatSN5XqrTXFIM2lRJQyC5tss9R9QzYMt7VQNuFPzm
4f071vU9yclQXQAal5W1T3Vjxn9GwTKpXRsjoIZM9WbZTYqyE2wrjHli2mzBwEDY
yrFzjzL6a+qw7g+BGDyRd8syUEKs/A9OUZXj5VEeaZtUyzFFa6kZpydrFiuELwiy
piznNXlQzwBqWhXTNLXymv/BbmjrcbCqYcw8SWFkfO61qsNxF4jUgbztiqx3hsnY
1suC4Ut66+9vzfkugTYmLIcRk9xNwTVUyIokcD4qQnD3xUrtsdlVUiDu0DdBmJyK
mJnXQ48rg3kJVw70Lb7/HOVmIkiJ//++qa5QWeUUfKFrq0jJBiewhMXYxkCcEZsE
vxX0GbNNMuWOPDQ3iWwN9hDHGG+TM4nsCHCkCJKj1AjRLKoIDtOLz3LKEOOdqw3s
CUnsbP6ym7WTZxhIR+mzYgCLMz/UcGKT1V1gUZayN/Bz5U84mLVmAkbduAWx3qBH
uCEKyOCs2mq0i8ua54yfXJ71cgQ/fQu+8WdBaUh7UnmydG7Fk4cz1qrJbYEZ2uRO
hu8PevwOOFtRPuJLkhJ7/CZgu/I7FJwXBw8frvoOc2oh98G9rpQ3WRgFo3zqx8aH
hpyPeSqaom4/WFO9xgMhNPOcYmqD9+MsxD6KNZrhAugTn/mtyNFmXMXeVUgIXLUQ
i8Lz5cnDst1O9kiCinMFzzu7CrxcpI6HCuYoEooBVeU89uqXISNGgiKjLo8aMo0c
zvgndL3swCpaHSXezm/qCLph1IO1JnxxSDaytejUiy11kKND0J3vCaEYQb0dmMpt
vHK0Vf8OHCBK7mgMLMwwmzEujVKKINLwlofBXZ3k7VC4kAZ1ia+W7GErgiTPqUtU
sXhm4vutMND39QmPukma8k7AcSWKVNq1Ib2myqTN0HMDFDvz4XOfBmw3qzcZKXM8
ajayNbeAVqh/R77yw1XNieSA0gDFpidWRBEqgjBYZ8yKvTdkZ/Ey1/BpT3DLaZJl
Ot/H7/lwaiB79Zxqs1rWIAwEDv75m+yK342cdM6vRp1jpDL1e0sGX6/W/TTD7oty
R+kO5tvsbzhDVCg9LhdYvwdfC1U/cjfUrJ20iYS3In/J7QuinKBA/vEttfT68Aq+
53R3a4uoE1WLRKUx3NAAQqiirI54swxzcGUSGagVVG+o/w+SCqMvZH+uRWdbfgd/
CsUN+8UVGxmUoWld3xBekVuQyFJnRIEMgY1CxpxC+sQ+VJ6ZDHgaQEG/w83ug6E/
xZqRV8KdmjcJcyqNSHADQcob84YndFPKg86vOpvS+Gl1VwdXmccnwqqxU/P3+qSQ
+amEKwrym17Xqr1O6rR5tjM5/jCxuaJbeiVXWVSe3uFeKcE/AX2RKr7FV7F/dzEZ
460lE9q9hHlsGzgeXMn7PHQKpAdBxD85j1fjks2k0qAU35KmTO7ZRRIAAXc5Pgmk
NOaj9THnBMEXqFXMmmrTCpgj7fo9D+f7DhV1KmZXB1mB+QDJe5pClqPEQFLnOexB
jDOZ09221Fq1ZIhuI1WVmGM+0WKVNcmnjMhIos6N5BBPqyIULbLANfxE9oK13Akj
dGgCS7SJmxS+iLiutirHKfeuzOG6r6HdIwDX8WPHjZQHuzPj2SQ3om/eDAKwTLdG
Rz1aiYt05SvveT+ooCV+O8YfXyI3pAQrocLtHJ2Hf9/Kug8hQdjz+jPCFjo9XmXe
vs9P2i0VPDECPNFebv4C0RiPQM7IzOGVCvU8OwO5edgao8DktT21sdUal/mazfL8
NjAlqVozZmwHJdQFv6NhCOqFUwI7/Ri6Ul3IVYzewrRGULGImKk1m00IN31sI/aN
jmStTW3bgIITos1Nq0LB4FyxwaF3zXas8aWcVo1aZK210ZWFmYpoqnHXZibJYQWB
lA2M6DE/PPOJu2g4p/uH5WXe9jPvV6i5NRgcA0gc9iMA9p+U0lQhS/TYOylShItf
EknNpVnNWiY3aPItDtO9jMWtM6jXtfkqtcxTICKBlYIRzOcKNL/JBJX1V6rWgIhW
mZ/DJJv8s6XwV4flhWe/amB7ZmX0ZFODtIs6L7ZnmrDLPN5DDGba4O5pWiq+84EA
oEVCfohEhFq/v5iXiPA/49Zg6Mrk3l8mXFfIJ4elfMchgS9uOCW+5yFlstc4BC0a
9FOVgqs3EWQ+S1ozeHgLrlUggBf1Dttvacx6vozV+Sm2u/jxHNOxCuEZ2fnsg4IG
JsEELqqPmYEaXqdG/jbTKi/d2YxfOXXTCksxXFE2ZhNpm4cBL+CUGOQE2dZvDkdE
m1PvNs0B8vVLXDyx4RtQCoT8Qj1ZHmtph+VzR/0O14uB3yNB6R18JBh8oXUaJpqs
jA9XMJcO3RqkK0Drx+XllqcSQVRItKvdKv3DEsj8SHqFrSDKSpLGUVZTogEp+jf5
rkmnhAAo0gT66qjf/aqhjalnK4dbxeoYJ+TQ5+uFuLCF5KOUXxgvJ+IHWO/CZvh3
7tNXqKcIbsHADPRevVNz63JtQKWYVfTQOF6u6yfrqgfzSKf7W18tAr8eWC6Nmlhv
736VoP1eAgLn21TFFbqviN1CD/dKASsP6hS6lm/KFi9ImI1DwvMjE+NThPohW5Qy
2PV7YutS0ixrrIV4I8jYfEmIUl/PED5+MWc7lacECUQFoRzwLY8/ROX6uUd9uMBy
Q7eqznrY+iB0QCxEx5twnsjfxkS/mOb8goHqqP3SgPC646NL6E4iVnjFIrFOPs/f
xo1QakxKi8+cJeDMpGvgqYaYWYbWwoIqxK0dDzxUmizwxWG5N1TY/Jt0AGdIUSef
7+PTL+zNMaOAJBAxiCsC/ns87+9Jnha/P1WKw0psb0jSZRJP893976plVY+EIMQI
iqg4WibUzNBO2C2wRsYZ52H4gfOdaDfxD6b4pt4bwi0QnAxW+XtK3jhB9AmbNOXp
wNyzTnp7FTexi32y6psTnAahFFJhlMj2JL6hog71Tg5CjWIsL6V8dW1LKZyf1Hxx
FCNebdj+ilSg7VbpEe4LuavtIR3pg6zHOyy99xZDOh+1tKBdaQKSCiKGE9bgIwCH
hweOYUFqSpSxGj3TDW2m04pluPv5hPDuo/mTKFOnkrP125WxnxoVKaYP8rLzZigd
Msd4mUaiDlbUuTq3IlhU0gLp7gHMz5UDyr+iSjit5Gv12hsG+2ETnfU36u9aTmJR
oYUC+XNhMGKwdaLMNHcJBNKmoVggm3AfpGd9S5NlcbRzrH5/qAClz26WIUaNurHu
ZoLEGZwhuq5ffa5Unrwpo5ehL1Sbrh8rCc5jLhRSmyFhQSRaoeDFNkwWPb43S5G7
ruSRWLIzLjyjfmP3yyAdOYWYMur2bgYKwI1QhidBS9T/aoBEnKKkjej7B4jXIFqP
m+J0qgXE9zI0+QQYqp6hiB+fu/ubXBrLbrEo+VVtCdkph90ljQhj6Gkf65p06Hz4
kBE/s6uEAbkjjKVSnM4kvtEaFSRcx/a94iFvUTRoAe5Z41HntUY0/M9shr7zXTV5
AmA88MvXTc7SlGA5vio0UKtFgdIgRe14TsYHg1JfQPFh0/qZ7apvX5XlXptfG2Wd
0p28h/vm2CZdWl55Iq1sfZDMPg3bYRCOuAeovGIo94hBHkXDzzSgvEhNOKquKdJV
9x3xCr8lJpMVCR+oYuaImRF3o/nF7GfmuWGBinLj915n9DwHgE2wR9Gwcnwd9FRH
E5mOSfe/jnQA4ALe4OM2tneNBEv00Aki+ep35ZbGW5w8lNxOZ+otMgNpKK2UibL8
RGikHnaMQeSb1gVOUfxXM7d/yF8wGhuVdjfJjdr0EGY/gVxU+lxHJkVOaiffiWOa
kBbAF/jzmAQNS0IwXNngLyavVomUtd7svQY/MmoZHn0vArRoojl1y3Bo3fdeDpIq
bjpQZCcB3rcpOUM3jM0OE2sbBfy73dWoo3DneQrtKHm5SU4Sw1ceB7pH9N2dMFPS
DR73mJNfgeSuPAL+zoV7axEMY0STlfQYQZnixtl7BzWYUNidp2GXqEFr6GXVvAE6
PzhMnO8VEcPcIqO96f/VZ0UJXrVmsNyhWWdiSmzYMZIPiglqzc+xUpgmFrQVVm7L
TxqY0D/lftFDKQuNi/bn+9GdBlLJBXd5qBW1dnqeZGHcL7cPKYNdX5VKqI6AguX8
17OCri0CxT5qqhbsJKOrE0VDDehkQBAgfKAwCXSNhf7wMu9KKzkUBLz2O1aGK5nJ
KfsBobgyJAFwPCh6BmtkZVuL+uDwmcXelqm0ywnsSJU78LPHsiXm8r1eJJf5vdWq
teIFi7qTMbY1nIrShQXWHPCtFGh4IsAni0Jfd2kN90Rr3e6hiwIILadI12Gccf54
CDVtkwh2cH7jaEDcRmrWu4VGHqSCSiyxDDU6MhUll8GV6GP3B5OHDsMsuF3MedWk
4a2HZna+yJpN/tZ5727G/ojFocrD+z5uom1vNKHjax1hg1rfs68nVsARESxdMamr
TIyncGQEduRgcCtkg+LxYeRnyTCAYIP55ipqtQJmvHuTl+mfhYu3gWgN8Zwm/l6L
BUbfsOP/BbsuqHJu5mtG6x7M/oh5YpS4qxDKTDF7sFOuN6hzBvA6FFakSD7r9s9N
dnL978H774pH0iAuJRwPRXr29IDexLi71gfC/3XuXMPGucp/XIqGD+WYYDtd87Dv
cLGrLaGYK89wIM3ksaHT7tJTd/C97OpJquhFWOd1oDdmfMFmK5AkULQxoEGQKudo
2P9Jk+yw1bZkSQD3hXvpulw0ORwZBi5ymnnk4Be30k3thdMh0Id3YBvh7PhTILmU
7wqTDy0wnPanv13yQfC39FrrAtKtXYKNXzZ7qbUkCw+EmPhu8dnTq4Vkfi2P4UAZ
RraKeVKSSC3z81HUwLt1lXPi9Q8Pv6WMiegeYDUMLj5eXqJU2/oLpBM2cXLj10mE
cuBeBL/fcV2k0OPXaI4sM9ZUed7+cxgZsYeH9iAkzArW9Ad6hWyLhX7S1MKI3Q5v

--pragma protect end_data_block
--pragma protect digest_block
MuE28aikjikLhFONojMQW96KQwU=
--pragma protect end_digest_block
--pragma protect end_protected
