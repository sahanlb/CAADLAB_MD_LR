-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
y1Vc8nPchqzUXnFXH2u/aMg6pufrh+3iWLC62oY1ZTp3fgMs5/04dcLFcb5Oxfa7
dnfvwWWUB4JOrOBKmK/F/mSi49+9V3syIl3JVQjEL/g1VMzyxQcQ5rrVc/K3mqsO
s94TwGt9dfDMOlZ9KRTL7Nvu4N4RTuc0cyYNCdk5Bqc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13856)
`protect data_block
W0UZz/Z3ggYKOYozYFdiOs4jLGGGS1CRiWuM9AoqtRy3/scRtu3XW34XL/hM77tG
kADxx7d7PymxIAtIHZvih07PU06UVhbYeimR1cFZUyOfxxqufbEsoQkieuulVKEg
e9IQRvBPHbmBxGmffObEfdAv5uk4ml1/2+c74XpO7zsdu7asRryh0rqKR3zBNmJm
H4SWrtnbRAgTOcKMnUyhzA8hGPTqhQ3QkdP4VRhPLts42qiT1z+MuXMWY6YVGm95
yluMxsZaOsZ50buXPGOUA/TBPdCKKsdC1tlSu1CulKo10IjhGh5+zcp5IwLfhCSP
onK2/eqBjUr0XYMwzmj0s3IbqeRvjUrvGXxX2C74D63VME3F4rj934DbVYu0righ
Mj10qfFCeytHhvYUxt9CGgajVxGv7RcexDPCN7IDVcbtciMhYx+a1HhNEFZr283w
I5zMGld6X5HrMeKOZBZFcPS72UpI0mJjZJTxfSFf18AFAzdx0YyFbaDiHIGdI081
qkwwWKZMJ1tONIYKKe/BJ5ipSdUmTpkWEcNKRGtRGVgY04ypxlvPZrFJkm5/U13M
BKsBAwX9J+eMp8kHoqCU48AwOqICbUyE9k5JKK5fsYkj7xRddIGjdxHVdSztXfZ5
Fbc08kFAb2l1TLgOAgr7m1FWCgWrHCx2XlT5/M0Wri4B38tA/ZsLTR52vv9WDe7Q
CWK53Js2LD2Pp46oPNIHfBe3idVP2fmYQrLfEGn7cdblunfjBbIymOgb+jvY5f5C
SzxAl9xCmUCzPWbmlGuCbA39E1HIeSa1lH2sYuyA+YjjcFdz8ZZWoU0pGH0X+gd/
v6zFua6GTAk7qOPyNulV/a0YglLZ1IV7MkAGmp3zouAHIOozE4vvgfuqfUpKQ/AR
MWnnhmEOgs1//oK40wnrHjCte1pqb/+cqUOHHf9aMhmo1gl87zt5SkA5/Bby8btV
Cm57A44u7Tp0PCLOoST5SoVME8QSJFVJ8ttbvuDthMOlvOJkheRY14aWY5seI4nZ
A1S27MxPGN30DR83+0JpvgN/VeaTPv56eMSSA/Kv/h9cs5xGc806SJWLxLr0gGek
eOuAGimiH5ONaY9nZS5thJhC5J9+2jW0Xh/gUM/tV6KT8JTKBF8R8NwwbcSx08fu
EPoyIBsN0VQNNJDmQp/P5wER0A2kYuUakL0KZhhiyz44jgQO9Az095dWjslZG/mw
W8vgIz6hP5/w0jvqsuxlOFxjj7Gw4gkN9ZlpzUnea5u2s9AnEerN/45JTrqO6SuK
op30zxz0Qb8/PZXA0pdsW8gsd3PhKFmxbrZDBRkJWniCR0MUWy+3LGbqs4m39mU2
CVEFeyyVsPEQlJXfJemBEzQ4owjoYTPBzPoRTVptfO7DtwL4ZmUFZu7CZrmOOCEm
xW1B9epsY4ChbBvIFHkQ8evOs3O5+lumvzmE63KRq5AzVnAXJmaoZ9DPXHfX3Qew
BB0C2rwz3/Fm5ZBedBrh25g5sIQJv4ZquK7uZDpi5slTHs9U+OhbROa3Hi1WUGwq
lvkYtMxkmqnV6iME/gWJE6sWfFt+RFrxJ7sO1cYgc/JMippbYRRVk8h5DV0sUPAq
2NzBD2MHnGcAL9t2rg0aaVzTryaTcazFtO4Zjhrxfbdhwg+si82srxeMGtgV1K/f
6txLD/hk3UbXHp8Y/CfzJdDEvZRgN0pwsvnQuxzJWwsZi1DwTiFckn5pUlEm0R5y
IAuvovjuLqAkl/ZaJJGAfBRsAcGt+Icttv9hXussW4+4R4UjZ/gyeuqnuL5ByIJz
j0J/TDJhY8TwYP6k8nTe5kQTTIJ9e7Pa1jbK1UZiwGHhsFc4l0YjxcWBNF3I1Iss
8qwGK2df7U0nAyM+BXUMoLT3ZPXpsLi5/GFooP+8p4ixcVbOuO7lyEolOXTA3FwC
3eVFXw1NJOg3A8bBndZUBpsMLcazPZFLctDQiW+vmTEz6czp9vJwAFjOs85/Vvwa
ACzEndwUYD2rKqlzqnCclP1wpGBomr5wVXoBe+XB2i5gbEHuQbyUWjuBSD/nAKFX
3YoDildhmdIbxwb0Z+O4NazyyVcXTS4vk4YXJqMwJD3m+VVQSOyW4sDZcU6yFs9g
Lxaxhx8K5ZLXcdI/3MsaTcm7z3+b2qs/1Dm3+on87XJ+viVF+vh7S8wXRomT5zbS
Enn3yJBdMLowUR+qHghBRqizZeSV+auUIq7a/Ynmlw2zkeXLEeYwFLLmMhs97f3z
8qnfRPwFFPgUltzs5N1NFBvOUKtvM4+5zPOEk+vq+CpdWWrscUzbqUyx6kRb4bSW
yUTwPjTtFlAu+6Csfo8Xj45lpbEQww6y/RPkKcAKE51aK+nwgZ/0sXrcsNPUH9fk
IvDAWzEs1TG+gkleLJL8zk19UQluY6YkU8KrN7zffkFxLvg7k583bh3Vx/YTD5TI
L7Qwb6rVMUPLbOp6XX0M89azsBE8GK0hKVhW9NCX7uhzil6ijzSWrQ8/0Xss+vx9
kjXmh4dHsDD+Te/EEsabFHX4UitV7dHNqCgNsCuFO4XgJrgLxw3gdmT78IzyfRAW
TAyITKSyk0ZiDcN4AdjgoCLeSW2m9RgRVoPRNlzw46iDE8EJ2gkk97LvUEs4+/Sq
N7cNEgZLiIkGr48Zcnd/adaoEpr4gosexxl2wdN4PIfiYwdES7hNPVRKn4kqiIFB
h/QK0qgrAKkzRjnYvIYX/9nha34Aea+1ku3nS6swj4LbxgXV8r7mVwlTl5dEihqg
kv4mmcCRwfwVfpYm5/ie/dSQmtYAjwa0XgUCPDPoTFaiUpOeaJaGfCi8/PXcymE5
9TVxYvJLjTgOu1IJdSd0awyJp3f0YROOW/i98h4QWNIfb4hOMfWkpopBvsy08ftT
lgnTnqVkieF5ZxNRjNjcy5PA6nL+UsYf7ime4+A+HWUghxHLme+NWbzm7iVZ5wyR
5gQo54zfJOSvqacz7FTrITnf6Slw9r042BPOjHRCcC+CzM7UiOYtD7lZVXjZ9Zgp
iJXoBNZ/692KYWARl2zpO+vAD+3B2oh5HPrR+tAhc+BESrjlWZ+V7TrhDDKxLcCV
sWsQ1Zk3okxGsd1+fAiXEDTgn6TmLZ2+wOoRUXtjmMtdjg9pexXsUjRpsGOqQBks
rxwgQA7s5/QJ0A7D4yLZFLPWTlLNAvs3JBCTgO6R7CDdJBPzlpTtSNbp6a4vElFD
/BlgsDD4gmy9s7tfJ7Y5FnTWKhwHnHEk6GGIakvhFHeydZgesFFzh1x0TSdbha1Y
2cw4FyW00PN71ukSSZM7eqr29GmehJRW8FYI559HO/vAKhHBKR3BnaAI4Vw+l0VK
HFxqDjkTsYXB70dndUDe4RHMCs45ZY5i/nra+TA+TqmrN5A+BUsoEUmFJgVmobcS
EaJe97iXn6Uh3rHE8box0BmUA7zToQoCE/yNfrfabQIJ9pjoZ0v256JSQMMxyPrK
TBOOZiAUhU1RlPboZd3qxOGHL4KSjbTmnoMdYD8Eyvqax3oLjT2gDs9SMs8YA4/2
SBdAAQl2T1Ccj1vKzRsR/YbVQFs69Rn6p8oa4A1Ge7p8IZn6gUUrGPJaAl0wxRFX
DTd5nZiePCwOhbXzWkd9XetbJrfMcPP8v+2T5Hh7hOKw4sO9HylQN4Lxg3wZx5bG
AhXxKlqjD+P0vRLm9kQvZQU5jGdwEkv2aj1cUDIi8jqkF3Y5+hreNpzxTueprQsT
JKT8Ipjm1qut4JYNYusu+GDzeauMxPiJLMc6SSxIsSlXaIGWsgALTHQt9YF8yjtd
KNQKMOWhYNuLnOvyfL4AudBWLj2vqkeLOPYD0/ILbcWkedgBuzKoSLMAiA3CfdZg
vxD6PbrcnQhChrjULXx5jpnKsyLFHn3E5ajgj2oqx7+bGoBu8SvGN13y6T/2OCxG
VH9SS/s3JUotKRq6/zcfhTPKfO7gUqLgXkGcSKyl2wlh0s6sKGt8DAdRmTb9FSdy
ZHraT2RLpqPD6SdnQYyRWSideEhJxtaEf+2PqyskEqcd6euybwqUdPzUT6qTttA0
f/q4wNINpnlnp8hQpZZdzdCEAfnzHKaInfhjT/fpTny0zofQeYfxj/IvAjJN8tae
CtfUZaeeQoYsE55Wgc2g/61aRT3yDc1DgBaGp2RbdfPAyqMUPBxJf2mW9JjCJwiZ
+D06vwD8kyeeSX7BkOx81AXWVPAsFySaLFMQpIcmRU4YEKBr8nw6yk2paloSE27a
r4NEe+LRaCGqbKV6lD9HiIPb5qz15TUhDCIyeZM+pXfObQNeGR1zRf7U0/oXrla4
MLKfb4/QzUYhYt2iA9DZgS1+O4Ss+19swh9Ui0DkXqTxV5tdRqrffi4tVH/WTcIs
sTu/rn/IE+5jhGI+WYoDIBLpkkhO6LZwMTeLE7rfj5+icaEnBAxAW/33iRVkBVZX
7aIFQi4hvqy0L6W/MSnjE9pCWY7Oq6LohIPwVMIlZ5pl//LZD+8c8dianwSFqz4/
zoqD/8FI13ADm2kGNm7nl+UWnvi6mYu0JnFe78CYRfpe9EK7UBSuKbzbMnJYGlOA
zbF+AyBafM0zgYiVe9ezC0EEld6sDMOFDxPZMjyk/SlEFL6RtS7lxe1rWH9Ceg8F
lfIks4S6Xx4OT7W54UKuDZkO8QwS3Ze4M7QCjVR68CzBpNXI091ETd9aw454xWfL
jxV1lqc0tw8g5JJ1Upv+uHgSMqHyalB4sSklRtxv2ZryJX1ZvgJVoRRmTh6HWGQ3
7qakpocOHz/6x5cLf25Y29GlqG+dISoezdwCN+Lg1HdZQTxFTqvINEqMVmzuGw1p
AQsMQOqxhcxnWMw8tJZyCX1tWsCcKL2ZdiCSSSxkHWnwhin5TcRHRqmRi+IDP7aw
HKw1CMzdgWmLyuye/tQFzBSGYLm3FYxlo1hFp+o134Z1ssc+w1HIe9h08eWqxwIO
9/DyochhvtEDWtchc3e78QSnPkC1/9Ebh89GF7QVyqkHGpEObORepGfN+PwqgGiX
b9isgd0UnGIoZBz70HYa3JyVp9mcr45xAZ0WRNMw/ffvK5oTUbBV8s7rV72vp1ui
7+uScHsniDPIXSvDQQtP0+qCtTizdXwkYERss/qGMfmCpRoQrdw5PUiFT+JtmKOi
3Tu1XeYUt1h0XD7lRmSQbowkGiCu5d3lRYri49ixwed4+sK89IoIDZNkpJe9s/vI
CL6lL6APsBstuqVZChNI8TqQeS54MGqWUNjJQ/2t2WQhtTFdg9b+5+50uE2Iu0gQ
e58mJ8MpQCSQhxDrwIpDC3uFMegr8KPOtttAwUk+xRP1G9/c+ui/m0ldpbbCYUyh
uZ65WppJIY5yOdCpOmVomB9NAmJPKsjL+i/uz0d2sOG2mLVt0tb6ZZ460+6Om15Y
xslP7j58zzUEzUCaIdxm7Dk0z29S1W6154BIOiAvy6Q9FT5upFy63VOY4Mh1s1HN
p2l7SoAqpC9CseBMFedpIZmg1aE8IeadDpMlv9onFvISkxAYukZBQBiPsf0RFYqL
b+bmG+AhlMfCKB/+82gck5Rw7FZMFhG2H4z9z2NKTWoZXkMm1c9iSaYUBLK2Nmdj
qt5f2LaX1/P8E9xUnEOnu2HYowPfBWFlzR7v8vRDM17BLvoNAVYnh+oHGZXBwYrH
q3skQCo7+8LGUk2czdgSb7hpZbgXnbsUYNNOk/+tIV4Kz7TgBrDZ66pPx7LSV6LQ
Mrfspv3ni+EhlCdhNYwGzEbJri4oDq1QtU4ttT7AjUr0mFmEyyvlADtiP9wpyF+A
Mq1NSpJ0YDqFsxM87ZdlaAIbNlz7nKd/UrBqeq/YKPyhwgdiCDMlJV0hdicqRzbq
WSX4YPbj7vbzWxU5mIogrItgtds1U21pnBJBCdPf9lSlOsTYJjyIYG3BRd/HZJkh
1zFJoxR7cDNAXSV3lprrPNq/UpfymPvB52U4TRISC/pyxtTOJS7Mgf2Fe0mT1Dfn
oxF03mVBkOd0ufP/jMuk6J1651LcoTZTMhE+gePQT1L/rqtHUNAONCfgLiWWlcrR
M6j7it51Ebzo4qt2ybauooiF9tAIpUWF/CORW9UABN30fZlOxU6QfKX7Vzra4r5l
yp4WnWho9dw4vlheDYyngcf1StL3Gb+nCUPZzBz4YdpacXDm4hu3KJxryhf1Hd7W
1MZaw9zUSQJRQC/Z8Rsh+3yM+T/fc73PTjrZjnhg1CScEutbg7Mp8D5CWObDl1+/
wXyy7/GsBDI2TsRxgk17hULS+bcFfpN0M5w4I9JIsjo1MdHCYH9O7p9pnz69acJT
mH2Cuwk2AutGWCrgT1H65uvxJ4eewRiXU86BcFL601BlHup4KnDx0QLo+h2Z83KW
YZpzIisNEy7mk8TIwXGxl4VKPguXTk8lnQRPAXeOfeRK8gGlP+gcDevUZtSHV/lr
Tm9K0vhyrts9vCb3hzy5aBhAzrhgLZZ63jXd2LJ/kPHqG/xKg84twES2bR/JStif
WTBQ92wawGrf/l80Vhc4ZluKMukWYWqTLYuXqyZF0TJwxPHsoHnV3HyEb4rOJrat
y/bl/y/e4eTy+fjx9RM4HOzdls9BeRL9FgBPLlowqDWtmtd+qL68/l6rmbrVJkaY
lR7qhWFkz63C6e3us8mASeMHo8ZfxAr3CdP6I6qWxMYtLCothww15EdHDyjQsdmX
xbbL6uLj3DlSuEIxyOcZ4phg9dgQkgygZ8jw08t1MrLgSrKr/K023hC8FB195bvu
VSOuvDyNn452m12L8X1w5gjRqSAJ1r48L5CPHPcLyHA+UOcY6c43sQM2pjgw47Co
UpEmo6W9YqbimKEFjmer+hCvgiC3QVea7cwnD9svPNRd5oySgpSfPqzO/uNNDxCe
pYHZ81XBZNq9gSj9pPCfyL7mnPHKv3Eh3qf+cIcIoMiJK+OcIV81mKDULu0FoG11
/z+1Vz3bXJXJVtHJpfRX447n1BtE0twBBtp8GIeIKyPOSd4/7o3uBvE/yAHwK0Hz
Yns7XZleavRG9jAMA61jo0G5mUOaQUQpCfZK5TYqNa+zNtJnPAprfys1Xm2Tz9JF
CTEF9dPP+8iyX9V/Ns8z2KbQgeKdtXcnpT23S8GWwwuWZh7DWelj3Sb92WTR1Xvu
/3tjQNztftSzsDpRO71rhRD5j8JfMewogMDuwL7lBbirtt8vL4HgzrK0UxU1o817
3L004hZkHITDBkqw9l/j3XqTusMdPUuMIMoIBqxcDYDRIcE3Dt3jKB8a05ZjjTHB
Bj6LRt1kiZnCEAKv6GlFuS5Y1pTEUPqfjHoFOAlCi4rVM1F7ZOJxEciLLkEZJ0Dy
sxKaizNVaipisRtDEENTUOkWUYChHwMFFJJEGyUeuXizAX9khqob3Cde2ZaE8Cn2
+dv0bOgGdQH1Fltqm0XVY93UtXMpoOCmZwfT+whZxQYDgyrGGQaQTroYK4jiWZh5
PO9Du+VdIQQ9/U7g3pHw8TyRXc4H5qoGNk2Ig1pDs7XapxC2XKNJTECUIGeQaWo5
hc5SR/bSHB0xRn7wPaSEeDvGSaxG1QhEEu4gHMI2GqGthDkBJjPrcOCNU435p/ew
eQGt2bE4bofDr+rmpNUWweybYQnZ3vKcb13/JJusTNBdgec4zPzTmM8VskyQbWcx
kFmHpkbhED58MFP8SBzt8KuRlIxQTKmtkPvCiJdMd6/KwbPDzNFVaxJnzVWGgVG/
ooFlvpdwwgTtsJhIuThivBRYd3zSpp8Ld/SpW7PuF++UnJDjy/NavzWmOBnpKxjz
9QbILVPMINslIWGV8hDRhrq+INChNKlumhAzW8KvKbwSO5l3XyvC7KaIU17vhIGp
mRmHy49wE2/2NqC7QtiDx+OqfNbHumRCMMvitHEhBh3pO2kp8Q9UU3oV/CuPqUuE
GEd0hVNjHvRvX3hg5nsLVxpkI6BkOCsjzwhhK6FqTRKB0Yv7VSlRbApWcFNr7fr7
gIJ+nMHzF8F3WBEKxcbkbc5/DnJ8kZloH1mTQ2Qxm/j1Ww30HNRBZTr1ZGrro+//
eJJyePtvuJHHCjdbGgf5acfXlIKLsE2s0HB4CZrYx7edne8DS910XqSFZ2kK9SZ8
OHuPM/WrILKkCgzB05n0/5R60nGrA3Zi8YHa+BRXcfRESd3uJMD7todkYZMla3rh
usJCglR8iJM0+G2Y4Cnvt7SRQ02NV+gLRZpWclIIyVRVGU/T+4wFwZzFEUe7f/Iv
HmMaaVf8VSD3gpjyfyJbX8/FOHPFgcYqPO0iI94sn1Cu2wr9jpZJhMkLMTiQWmrk
NqD41TJRqs0DwmVKj6eZPqv0iEkViXnsOyL7hOUQrSgv6gOEpI14eVsktOFmCPY+
Ilu3IgvVINGEDoSPT/z646Q536faqk0JOhJrKIRDhY9EpfARGtSFxpz/q8+g5sTt
oFf0D3hHMy0ycuu4jeEFtaacgMEG4WRW0f9nCAY2ktoHDl83YGMLtGkJCZMXt1+Y
DqRDcnxpum1T2rX6VypNqGbvnPbS4lsty/IQ9O+uafjM0hgDu7BeJ/A8q4LxvJ6q
1/NnZDZxLdw32Qr6uHl4ffSOnfsjywR5vzPizXV/R0N6vVWz/7JNXgOdiSAjCMa9
4ldZbstbFREFiJB8nSnwJAFMtV4MTuiCwH6HH4E9Es6wAaRWckhQVQ5OrkToubt+
rM41SD3PsbLrIhz+vygsIOP1RJf9+cE4U37D1gyoergWmjm77X0wwkhy1DW5CJQq
0bDTdwzHPEtjFDoQt2A7+pnEKTKH3dqpyrbMXBI6qX1NXb8LqeUTamF/Gj7ho2QV
eZ7xZdpwlDKqWeF4DIap17fwR2kqK/inWh+axXdOO1RmiguZFfxJiyOxQ+KvKY1d
96g05kWV+Q20IAZ1ykMe7zHpXWUB4VjaZwg52lHl/7z/VqL6trdl+UXxZjP5e87p
gxp/W8FBvWothkwws6Izzg0sFa2mz2y38dj6n/629WJpyFHYD1R5vuRGGE6/2gvv
sZeP038a4dkjZjQcXkX54/jV4zq7rFiDQhBrFjdNPAVvyFfIJRCs2Q6+2ReaPkG/
e0HNjRu+xzeHFCsBL1kUoCRce6qbWjGErUxejjFJxfagA58VhbShdS8PKA4vJXdQ
UA/3hsxbZOTSkp8bJQdyuYBAET+92CxPNIUOil2v3pSNCCkItvImRcU9IImqvkNd
U3Jj12sqjlHq7zw2UY/QNiGSdKwBzardanNMe62EwCeUw/mshrunD3HDSjhSLI99
3wBSbmkpuFW31TEiuZ+2fPNPQ2psLyRkE64X0s872NDf8MqmyPQ5dS+tEMwSrGQu
MGkMUewWv3F74XzxmD2+hAdGHlpLnWnAQI4DlZLRJcKt+Z0JTGqc+tgH8jrjJnla
r6yw0Gy5gw1n8V584gQNjPoUWEw+a7pXCv+rikLO0q7gWqe6hTqiU10B+7fgMg8J
2DSWE2TNOcmXVBXhJe1FYG44Sbr4R8s3R5EW2huzu14CrXisYsccZElS4PkXz9T1
6rPJA2n5lE/4NEorTq2cEpwLFWpr7QBEFkohQqL/XPtdksIcLcbtcC0/CpwD4C+d
ZNZ56S2FQIXrO4Ur4qiJX3qFHtI2a4V7HYVwCOWAp9hJnvjU5bVW67nJfHAGkj8N
xsyCfBK3xEagVpvnqgm4HIx6UCB4oikzQON/2rnJyERecqgIrcPk0NkWKUWtClMg
dJVEoLiiTozKp8+X95p9t9MVOMYiYrXfl7neFIXP3QqcLCwjsBln57mfUub4VjKx
krFZwMM/i65rSa8MtNgOOu6xJBPiOsbb+frw5hPCHi3wdm1VE/x8YLvfyIjr4QxB
ctbSNRCOJkVdFXErWaHk0NdCHF4iEnlo4J5j8K/GIOk6gaivsjqq89X1OXgnIJaj
0RkQgy25r6+X+b8zYYbI3qie1bgbijL9ayb/xcrRL0X9uzT2WT/pyRRF8NqUQJra
rhaaNQbdascQSX5eJxg8MVKTzJpilidFe3Ifqf6E6UgTUGaCPKzNe35+fNlDYMi5
0xMQ/L7Y3L8OBOpZwtfmmSSKikdwB11j1DhWBvNl4HWbSAFfZrhWxqdOITO8BHKo
HAUBJeBYMVWdSy2z4YtpAmcw6L07Q4YoYRvDvOT5Vf23jQQR78eD4WzXKKI5lEOn
7crwHVI2lam5iHzVm/gZyED88F3vOExX57PHsKeeV23Mf59krXg3dt3bJEvSZLqg
0wgsIAam6kpoVnoEqDyhYeGqg8VWI6MKqLFuPJgZPxvFw3XzYW2XqUSPKVjgPoXG
y2bVWNQvbyjLZaqaWa1u0943UaNVeWgZyXal7uJ3CbGi1cCJuOIz3iQ8S9PQhIFM
wabWWCRY3h9Y3RYotgvbOUC1X7hxGXxujH31TBrXk15WeXdzRHF+mR29xjxeXpkY
DNBoY5zxd0b9JhN0Q7ayYzRykAt5V7fQUhIB52+od/E2Dc7PZVAQp0cU+tYiLt3h
fGUxcSiQbN//rvwX8IFY479C65qmNpuLQ+9oFfV1tSV7d/gMF0d6xg+IVo+mLDzQ
q30SvZsBYxDQzDjFxOQuX/uDQv31BjkRKtF8MqEuyKAqg6wWUrYc17agTb3wY4qv
XO3BnGn5tCYNRbH7LxOtpoNt5Hr+z+d7TffJB6CmBC4jmbGbGfSNhXB3eh45r8Vk
HTLzcpk9b+/STMaV21JjtE+iM+NhcQzLZXClQ7NMJUQDpY5wVOtdo1nO/FWNeF0Y
VgJcXIrDBl065SRnLmstMRmb9a+bHsIQT38VG7N04Ec4gJimHJFf2orECNzgoV1F
QZYaNz8PGyLsAHGxcpx9jBbmfhE4FEYMatB1f7QYRWo+WFiiXDpX8E2gJoBg7HEw
an247xcsg7MnJdJLRwcHSWrLYSiIfRIGA6Xa0qU60lfOit5go7Ircq/AgMlUA66d
md+9AE2ziyODVbFBL67Va1J0WSoImrGFZqH2+YVHoGb5cH6yvGJlh1cA/DyK7l2N
lqfu4yJ0sV/kPUkVtYzi9tfit46nBZlBGoHJe7UOJl6AxvHPDvocCXjKrybg/pHl
icy+Mfa5z6kTpeSGENRFem7t+P9UBT5DrTDTlcsocV4SvFwlzNlkJKP9kOHTSDK3
FAAPd3QJD+fH4Zo+wubHBBlSbbwCFL/hwymfguyhx1LlBES67uIIwPOJbEWr5K9n
BVOzIQTjz+r/zGY15AzApGfoH/z2HRZWbVhP9XBnkNdxksrdVUuT3sbd9cxHWuBm
KDUpodStALIYUXr/073VaQIwvXBQZI00dCh2qg/rB7/irtc6NuC4M007V6YPBv2T
972Jp6AZ5hRa/DGhZDq+evaqEt9YPqrZzLm0mmv7ljfuoW0tuNW7finXgomBaxgG
rJ0N65GZfqyrdW4ZEO0RkIsIbgW2g1qHl7OyyM5B+an14FQGkqCC7J9mEIv5bMcE
I14nx8Nbq5UobM7O39rkIkaBSI1tVw/X5Xz+oXeCrA5qxjRPjDyA+vYxe/Pns6+4
6uaPweL6d2udLAJjCndOTt6+TMCeRQG7lo4AKm2lqMLjEzun6A5Ru0rync+nNURt
R4yx5GSjcvGJul1KNdGw/rTJUUBHvourKVyLK9XxJMPpikUpCj5yj5ZVRooGMQfy
H+9CgyoCUFX3pGKLA3m6gJAWZIABaumYJONnIQuWdXl9+9uot7NQHpWdQyaPyA64
cMkTx+3mRRqEKBTBHGlUcJiczUnGOozECNkpv6LXVVATj1S/l80ElQKCfnIw4aJN
dzpFysZdQUxbbRBRMJhOyQljhI1Pq9ezU/un1fmxY4CbKIVVvGmaND4eTzsFYh4Q
aUaFRCB4E7TatwD1UA899KB+soYezMDyM9YxeFe/s806BvYbdOtMtrexACe4fT7Z
Bq2C2S4XSH64BWh/D9EcYxSCq8QkNGidKfo8SvkJjgTfyLhX4N1QY5sCcG82ochs
6fNG4hFmc2NomMq6926lXhwbYW9NObJDkDv3PzE1BMM5HolB1ZnrzJxRTDHCkreE
gBXbW/aPk+YBOe3wz35VZ6uaEGJFwflo93GhV1GjCgt/9JuhSpyim4uKyp8Tp8AJ
e4IQsEaEip1KRn42XLY+6Yxps6tvSObpNx4c9hchukGfW65xj363o2kKV6WGHW0Z
KmT35lt5P8UV2ZUAoxWf0IMZlXO/VLoECKv5fIp9CS9AB4KbfQ+TN9c/oi8mfTem
QFLgwk8upz3+6rbMMw1TvCn4de3/7LYAxaky8RrYtI0sBZdpJd0g6Fr1Q0NcFa6a
YrYmE08SD2pZksU4QAJPl2UNl2DdLk9LK/UVdI8IFD9zOoybiy1qIv7tTnV8ZG35
EZ5ldm7OcMIwKjp0zVRqrZbUTGnGbSvxJKvtIqyw5EscHuj4M7JT7qzmRF3TiBfL
/Wyj10aCq4SYiWHuR+F7o2dHySTiYeO1K63/+qnw1e/yugsmYt+rieLj9I9lt88R
V7R2zZpGsQBcIKruyB0JZ0hkGRY7SkWrx0CAUS+6kADa1lwKy78cSeSZfmDzixjy
8cW7Hz6THu1GalMsCDj9F7eMeptf+iaaFWPpUXQKJkEB27xDEQfDsk+nNB/OYVq5
9g7cALtufpyOWaBLSzq32io09s7G7lFnI+00b0ACA2n+p2MD/o6xpVhNANzEYteZ
pubAjmIkBBM9vkg/qkp1BBJMP/AOI3hNwZN8z8e3qq65d+d9tEeESMhFR7CsQ9x6
RMx0Q9jhEKZ+eHQtK3lCKt5KoVzwK1mm/hgeUkyRycTS7pfHMzYaStlujl4IrGsm
UwIoAefmxuMjT46YdrtUI/rc6V6WMkPpO7YwGVeJ4HZuy8VbOvtlVXgBqOJQwtaV
54rjShYKyQhnpwdn3VaErttEpjmUHwvkQpHuFYkux6G4h25278aJwhO+4TRaKu4L
2lGQQxvYF+A3lTnhp6gSvPbvG1PS/vQdQg/VBcDPXVzTLpGIwuwpzoMkMPg054Hn
wS77mK/JWb2Ac68uQaUmPYZzFyxIqWbCsU7pEjACmcCMT+Vhopxa2JnNq7zv0dmp
MO4ZYKs9ZfuBSV0KUqdcm1Vc3SyswwbYruifEzzR15z/x8Y/5NMJLNqop3hsPBwD
jLcEldy8/6dloRsU8pQpz4DdP7aFAkyMJQY4JmY3jE4cu4r+gU0yqL5jtdAfO1Td
eK/TW3b8EItj9QK3Hx6LrcCAkL+fBgd6Np+KEKZlFb2X7v59EvpESdVzDMDBm/+r
dg4Dsq8eX+54Eb8hpt9yaR4cojyFL626B5+YORiNcrJIUqMe/FRi1QiIB6u9ZoaE
X5PZdEXufwDXNEGf/Oyq8/R8hF7c79vx7X66ITY87pUQkNN051dVrUxkqQNOiAMr
k3op224UFRuDpP/LpYW/g1kjf4JZSvSYwaMyn+3jCV/tj4T6syJbXWwZzDDlvovC
hXtOaFMWAfORg0TxnkCa93gJ3xQOCmyLIggwMvdHVD7td59+bfT8Cchg7XnNUkVx
mErmnMcZ/7jjuRssvVnOX5m57DzF/Cyxsv9j15xOkr8k/Sf3ujLjZs1Q/RDhNzpV
awcMaMd7NTN4B4nmMS0Dn4Gw9Y+TFg40HkBzO6n73VXGVu1pjgqd5On9HH/9JT8J
7rA3uHYYKj6dx3itJ64D8AnF7jGq3s12isKq3Sk/I2+Ghp3TYq6Zs9ljpFsT+GL0
GgsvIRR8HypXKlsYJVA9KTpLMHZq1ZhFMvridYrWJFDaJIGmTWw4+ljFEhNYaTsF
cTqpCKUs6Nl2RZp0SMI0eaym5r+izlcYuBbg96JnC6/FPsxX9tbTqu9xVyubDCq3
U6J7Pfmbnn/jRuVbW5IVBzvmq2BQV7rcN0UJBY9/y2WXgqIipQ0Ys/V2zEAl2jxx
tH3jYbYcHL1E0TOj2Og4Nk4gjgOEEAZoEuUz02Z93/BM4gRlwFMbPW4blsHYD1Qn
LxzGVeL/XW14VL009al3Ra1XJPclAYZqROHn1ePGnX0nyogZOeN2Ter5hfVgUj7W
5452HJP/tPtDgEABWXp3Fy5TNCKonaNoCeDoGbyV+j7nW8GIi13+Ag+80y4ASrGZ
shtn5ikh1jcdDzNQL0RyaYdX3d2ePWjahF07QVYPmGNVV3CrhMAOzYnV5FDbrfLv
56Nk0hhOZo9tbUclI4FLbx3t2cPdN3Z8a5OkHlSmMzb2Ft4PZIALmu4z8dDYgb+l
rbVGiDu163LIOgT0XWGxL9e5qibKAkDvlaaOQAKYTJxzfHflH92J+857s/5Vt7CH
3oX3z7wJfD3ulhmgQSr5o+JrNrUN/CBIVfN3tp7Icw7/FoRLxGxc2laMsDmXM6AQ
5sW8xeDmh5+3rebSY0KfhUcK4/yyMU7cT8ADyZ6zvYz5ApdElfoWJp5wCL8Ax0kD
F3NwRkj3W1jhmrcXFvwnflGoIST8gGrmrYTtjdcg3zhI2pjNJ8Gmn3ZGnNo4l1l9
t1Q9Xv8FoT9OvQZb6PRiyOwKv6ORCojZHZzCfEGPc9GAnCPDoTld0IjY3wXGFhlg
u6UZDF12p58BpmEBfZRFu6KEZetZTngHMzVHxuziWZe+LjwGW1NhY2VPQH+HXmWs
46lA0nH4NcikOmG2XvVJL5sGzrPCQwUF7g75IIfI3yIJlSZ6uqQ9c64cjF7+sMZe
KHRvQzB7a+Q3mAqDHb0hzaNeamnyThCG6F+B9z8g3dO8YiNq7SOMWaExutYqKfRr
fHQ72hqKPmMu+W9yJPaEqnQMHhyfgyFyeHt/n0PXj60bhHdiidwxfy56qQqnn04u
aqk4WTcQdUO5hUyUUMWLs00JBN+MGGH7dutsOUXxgKc4XKcK/K9QA+7nf05YyZd3
gcnXBtLecnggc7w0N5+NoVzRiazqvamrwes7sel+AHCjDH2uDDNNpb5ZuLWCA5KO
i99oKAt7hOdxlqPfp6gt/kL4O0wiYTRX2L4vas0AcUd4pLl03LxTQ8+/KFZR88eU
xpMxL/g7nbRrWWKHpwlZ6goJpaED63akM/0ZePUS/KZWsC4KOYSpjdNnJigtrBD/
Dg8+7GFHziiIhh6B4h7fAXO6PdEpMQhSP96q8zRgqGPcWbn+ArNYStkMF9YdP0zV
AIVa7j3s6pv57rfWBqF+YGxlGkAcgJhCebz6RGhx+3z3iZe2q41WsUpx4E2Dwn/M
pqxdCrc1+pUq8C0AZbcASEsOkEUyfEqWWYv0wHZXrvsv2lt+7dIGUJlVvTgy/T0G
Nan87rNH2isV2IfHJoFGsTizXmrrqPSOwnQkRBSoYHlxN1MX23vCXc2OvDvfilLo
mDVpVPYNuem97QJ3RJUY6fB5FAaDxSol0j1q81FFNG3kvWnbYOJouCcmcxwW8721
glPysckGIBfoWtpRWerkB5rmysd6oIcKdQDAXzRGx4zB92g8ZQFfcTA4cYxXPegt
Io6jQheIlttAEYnxCufoEOcz+yQcFNL2TF11Of3OAxuvYdJbrGBYjIg/y7mP5jfK
3IydDVvJ0AZlYhPwgf8DwPvSnfjezkkGUSgW1Lz9UXeT5i3EA0CdGK6+IZHrj7hG
pf9UdQm0hveFRXHmaXrwpBZEm7LbY7wZIBE74OLYW8jnqdRc9ZxyjQoVY+NYshPQ
Hll7G298nz0BHBsvQgGzJwrBnEbbtu9zC6Q+HQxMWbbjZYkQOdNgy7y+l75Vx2fL
PDxsaVcnO6huz97Ay92ZWOEUuMGvqvA9ez6tK6mZXlwroz2OUKEhD0nRqIm+Qsuo
05QbTog7WiQ25Ec0s+34LwBH+sM712U2+tFC+jjhRc5Ftbs0AJP78e+hR2puk1JS
cd5Kf7Y9ZKiJ2TY/+TA6x7IQt77XS1TT9piMSUW4xFFiGyuavCgQNQ6jvGg5rjpg
FI4Fe2qc/qIrhsP1NFI0rPVCbBJH9ofXdK76U6B+8+z3KxWscDsi4eAsJ+kxRH93
+qj5m29gfMfJpMwdpXS9cvrFe3u/qeigx9QMGSZ+f+hROAyW/52X1S7ecbBJfoDZ
x+JJAzP1J67V6hkpaCyB9+U6s+xSHdP0+8/kJ7RaLCZmLx4NEiuEWP/xbpktFmY1
Pp2Ppw/jqFJSm1josG1CihXYo02e1+lzmXPSkCa9uWpW50+qj1UpxrroGQqi2mAu
DGU03fDiKNScDhGvNaQ8dsFx6aUq5W31XfTBavXCvedEvFSZ4zf84fwhqIbAUR2I
x3mti7Ql5a4Z0mFZKJeQ+LSY4NM0Iycd5q7KeQOOK8VChzElxHDS81U7b6ogNJ0W
YRiJavgQJBNF1JoWDZy+DKkNFIz4vv3Mi2rMUtZDFksYAE3AGEO+5cNQtDFXbmNp
WnhvjG+eZogKT6BuwZP4DsNJ/ONvkNy71yRCVequEO+8um5yDBPLg/ChKuFMalkP
epAeJZVv1CY7Y6A+mhJ/LjbrkHgII1h3L8pMn05CTpb+iJw56I7o+9SSRxD7eWLC
xKyKwPJg92QfKLVHul9t0b6DaCfzn7E1uWFB36Vkiuq7IsccOSVjdSeHRAb1X6WF
wRLzbyjvaIGB2oPOCJ3+5LRCmqe/W1atWHcf3nUVgHL3sgV42iqbkl/oD1EXD/ym
aNbMfe5BbgsBVKxOR35m7czioNvE9xaZ7QCvplMJmtlwCjYyplAxXbluwvyBXZPY
MjvsrC7hW0JPYUb72q89jqNvOlG1lfegi1MB+IqzbsIcSjuizjQKe906WOvQe4zW
P4LifTUrSfFbnk8FnuzMVb5UscbwO3tXGrXE+4E8JsFMyXMMcsgHwylyjHMMOyZo
lSsFu186Ll3ka1a+yF11fXXOREbV/TLl5i9QGhrxSdEBvcKPR2HYkWMwCtD5Jr61
u1E0InkwHmcBtf4MDIcmcbkiu++ggjlCHzcU7nz8WTTzaMi790bkmu9zTXmJ4dJw
iEkIAvYkPatEDEcAQXH2gsSxNfc1Ayf6dzwgi7Qsz+TneLITqaK9HGbLKi0fN2Nc
mZRJxu3Bm6kTeK75MBWKzqvvNdsB+RGsNNATZo/TBRmkqoOlSN4V0q+py7toj23X
ZCYQlcMC7FUm6QypDMLihcjj2zRkCWmIIfvVZ0uiBD8trTnKL6MR77DTdIcLiSGW
L9LIN721D3W4WMr5Llb/I/ZlrpT7j7rnZEfhZk6h8KWkAZyWz5+JBoPBDpmWoNwj
nZWnR1gFcpui08rGBCiTYFiePebrntjvhnS3LEwRm0bmag4RRvaPt0FlLfT5CtRh
8bwpnKu+XO6Fqy12QgFUVP9uHwROKYO1wWhrcfzNytJRzAjTeW3VyWJ0b4RNJrhR
mK9E30Uy1bFAD9EhhyQ+QdoeDj0Evuyh0/Z7OJAaXI5Obc3lqH1fLNFv0DVqQo4M
wI8F8FXUIYKZCh7BrxGZreHsXC1mswwUfblGqh9V/G+LOAavzTVcleU8VCP4YcIO
uQ6/BlFs6Y7Rcq5acIVkeezdl49/itG2+KRxsEv2XdcKJx7eqAoZ8vQ7iMGJ5AWE
Dsy2cQD7LvzSBjC21HjnTAQujFN9gYMBqk9CV5lEUcKnvFg4yoPqYE+fsQ15/S8x
Jsq7tJ2CPKy1e4mpbh6eUm2kB7ZAEJDW28EKcHMVx4gkHXc4+WdRxRNkOmjHdIHE
Cr+aaA/pe2E9iau96OqRF+SuD2tUcZxJLPOu2hdI+J0WVi35VUVJIInPZ6/f+rj9
R68PngF6h8l6ig7dc1lUIHW2ur5CxCelwE1bDUvS3f9MEzvAPAoQkIPFYldizgaW
R735WxJyhxAZG3bOBpT9O+UJ1j7bRfXqnExFaQ/IpWHPbCWFXcvUg9cpWZFvt5zV
wdWq/UlS/1oUm4B2ciQwrdd3lmYrZrDJBzoSDTXh6Vag1lnHW3OjZkYGqQTND5DO
nGpkRLqcvR3HSIo8fyhQ/0ET/I1AVxMgAd9dFSzPBiC/b37eKAD8CqlhN3JKka/W
axDuWQxHVRnsSk4ITTovVeXhCggjCV7shlXMbDGa95DEHUrFsQB4nOXYWMjcQNTF
VANLqJn7CmFyuqu5Cy+KU591NTvJ9Hp2tn7ajxxUi4NcsZvocUDJ6e+Is5Gy14l/
0hcr8GCd2Of4kFRscRFInGSz5SXXXlfzTS4WYQYi5Zg7n0ddZrF69tm+A5hUqhaW
XZsAmmPIL5cNmPrl+JyTxQBE7rN02zyBxDqLrWQ/wba5dQ4R54mblc0G/Ejpu4fm
uy4jYON59oHbz3VlRNhrNMYrpNnj4pLGJiMuLabu7p8e1X0GwLsYYyynAZF2OYQY
tTBw+ewgaWmgqLxl0MYMUyK8M8dk/x5LoA5WVhX9KvvBM1c9xULdBhNkGav9Yuwm
QL6NhkCiKUv6bLsfx06r33IWc2qyqiCyY/tJPnmhWJsB9VHmH8u50xMaUox27BpF
YhkZh5eMyzf7G/PRCeWDqAOGf8CG5BElshN+s6askLS1KjFJTOBB75DcAJBlQRP7
xXXiuf1MkcVtf+sZ9DaC8EIBoh8YDIh1xN1YhNbpr5iWUTfNrWv4XfxJyOmhRSEY
2RBRt4PxG86BkiAHZZjGNWpINwZRQka+3nqKYj+c/bE=
`protect end_protected
