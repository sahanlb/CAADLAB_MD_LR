-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fOZSShno6oDfyoogdyJCpXpMJVasVBRZsUAO0IR6AWDYusYe399YyWOB8W7XmAYmrRWv9nmX88tF
Tkcqc2aecN/3jMwizaaunEAproHcd0NVEVwLMpgpunBeItDsUM73zEsmipmgScH1cBUbKcbmgYVa
fEG37amlT+BNCuNC8e7s6JXIJ2UtvKTWKEbzKKl/ARPDbhXUGvqrOzaP5Z0YMQtlK1Y68ulVmalO
kssWJ8iTuHyhjeIiKNIDIwMhuXWGsZHNrTIHNpFrXGjdky5F6fdNCJCrj988EDMoWe+nV6IjkWy2
4dDB9zVGWamopOy8NruMLWpYQP2StJ74jrq0kw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6000)
`protect data_block
UOmqCmmMmYmNeamRF+U0Y91bYFbjfq6O4bsytjFyqegpVvaCt/PbXbYTIuRim5adad6hd3PPTTfU
HWthSCQ+8KrA8Sqw4Ifyva5AwlmozaBe0qaQZ5CVHoZbhy5B+wcha3dzQWKCqpoxmDgPDdNc7wbf
886atryAw4iAX7IBOCuP9PXwvancieBTDrXMYn21CAVJ242Snv1f2+aXmfg8HQfJWAU2UyAnhRAT
E8sT3NqMpD6O1Ek736K/4dDy0F8m4zc6Lv4/FrJSmcHSXgxOYJGENq2KhWMYbFemYX2J7hTy3Dll
AB4M12GodglM7KgDJ39cSfI9GjetC7jbLwo4qxqRIR6GLcdRijh97pdMecpLjk9YxiXl8KxTlIXd
rwuBR1j2FBNGocr+7R7CYuJ3I+YA+M5gFtEeZZXhR4kxTMMT9FzrlI6aKe1tSemEWqss34rN7NFP
fniEUXs/fHAKWSNDujecc3Cl1x+GIoKK8xWMXf39D/8+bSs40UDl/4KgrKGpTHup5Yye5LnSWykh
B/K1Ag9WPaktgYassOs0tQQ7sL3rfZOAfFzyPoEpXOjofnyktinx6li3IoxIeTbRmweYopLyRlbR
sAB5KeSpXFe+dlIte2a02kHDjLbdFvNWW4oBlfnubPeVL2WzJRpfqyXOePO/7MDuskDwX+wJEwth
05yfi2CyBsihe9dZjV92TiqwyGWHHSdPycTwU1nBlR81/YJjPQLotk2znDdTVDnQwYyp6xUj5j3H
47FhZ7+SX0nZklbf8wAZMCqqOoD/vbh758G7ILzseTCVPbukvvAM6HTEtqDjfsV5r0YlYM7qTmnc
bNAisFMDTtB8Rt3r1CjOdVXCrVkcltQKVlbjC05EysD7xfX59K5URfyVhrCjxiRyAs+Q1RZ7wLs8
ia0pp+H5BcB30wHCvJu+xtb1D6e8WWXV5/6Nd7I1U7D2QdUUbeCMlPOPAl0dAvQ6uZUDmgZFs/hQ
wAoY1nEvUZ6c+Y5DlvKEhkzbDNbyS2xQ91cJe5wdcs8rljAt+sjzKv19wcldeDs5+xfzlpRHH56J
HsOhbm7hDQ3BxlOTi11MrhvPdJcsXaitBAbH3n4vEQdWubKXYPwWVxWDwtXtRu+JcaQR2eLnVewk
GeZs7+zVGRgzTCixjNvhsKzm/8oyzGW1HzEH5O89Jvo9p31ETYJym1Si62eyqVsCl51lcQC2R1kb
T/H3qtoJ37F8Yz2y6o/4pDFHKOn5gVJ4o3nDi++F2ZPkcjbroPnDrI2moTmBrZc0cxzwKF00fwwl
BN+LFi9Rkg/8JM5UjV01Kh/UU8is6pK6fgbAVhzFOIFihz0k6Bi8MeQXm8ItdSn/wx6NLDSzhfLm
F42TfFR90YC7usIUhrJQcnRAZG0UXXyhXT0LwrgD0Ucylm16dGWTdvN2bp0Zn1lBbwQEDGhbIQWR
vZSxFwAGSH2tDOLhjgJq6bFGwN6uPnHWE+pMw1rRaOuTcsZ7KWPKbkEkH3daQyO5EWAgoN+x4rUz
uIitu2r96jFIYbwZ5PFHnBG5TIeGeW1/7eAkwUUDgnZgQkWJd601h/G0P+wSBeLDhoCuCuI23uqN
ra2nN9V6/K06ro8PvgWUdyvJueyG3DkZzjRxyKTucjf+SvkFoNTNeMA5+Glys3lCCWC06VtqrTg/
pWsjpOcYouzDePwiSoZxjBWLIkCKs5unqZxsZTURG+B2xDK9FuhBvEAgh8RbF3xurC4UHsbKmeEZ
dmKmwFma5r+v/vLV6Lz3iY9fiinyvsl0Gf4a6UoiFDsOW9SaWQKgnGVx+4zwzKyNm3yNuUib1y6/
8X7sBx0awbkZ9QgCLrgKZ9IN5QIJIO/05pDoyUUDogA1nCceajPfFzn4htUa0iy3ifSL40bGEOqT
bchQnp0Zs6Prs0cULAosbtsfUpfH/IgnV0dIiYkV/OqnMYxyR1BzByC+z0HlOQE2N5crloNMmHJ7
E3xvVe7Glo6SW9CNdvFdFMqg6aOvy/ouDt4V42Tle1fsfq3d8FnTRUNbYj75yBV3BZ7i6lNybQa2
2lcgA51Hqh/F1sInSAQjfcee7bumfywnrREdv1055DnPENJKo7Tn+FzSYG6O+WhE3VIcUmL5fx13
0ZWMYTL68v+JsoxI6uJ58WW9wX/wAuD5K+SAaJF9hk/mAzr0TiGQyPEjwYVPvYNDOOtcWlTEKWWR
VGm/ADW8yWYEARq4kKOJ5mcb+QEBJY8Iyf/y5M7o+QVorfMyp6UbgXLq8IrvB+pD9Fq6ugzwvzwm
MJRGQUA3zPu5H9KIjXcdudpCRZJvbWRhd6drYuvDliRG8S/U5Ss0Q9cCjK/H3YZsgcdUVFj9z8Ht
LVlCjL9VCfCkaN5+QgnfFBquHJsJB+7SOFx2dEryZQpPEimKRPtC8rW10w/h4SFiM3g2E1mQkyu2
cfepN3SkZ8mjBe8CNFJ6s+YLcvNmTKtaawk1Xue0k/O7/CAeQgOqjLk8i40rNWcsMRYa7QAQH5cf
qinJn6J9X8HAYutgqOyRT+uzQFSRZSVVyj4p/mPDQmEfC5NOd/0HiG9CGUH/quaYHIcURbRDZyz6
OfcOmdP7zLpGD9QYiLH/PTpNerVbHEhLCTejc3eJvSX5Pbl+5slj6Jbl0oOebc+pdDnbiStmSz68
grey6FAhXBRK68p1cdoBzHNcPla5DCwCJMYAhXqhr6DHbMqRInhb3378d+pAJ1EWKTBgXTVNJjLm
jUy1I1DtgMZayORvkXYZpRMc0JNH5sWTgk9DuOuWZFVBnnycbgAuS5LOmgh7YRZKVgdhZgja0c4I
/9980sPKVOPONHrLog9v+xKQr02+skW1mKoRdz3IXeJN1TLnOa1QPre/+OCe9GiIJyAwQOPL1MI2
sU6W7QSKhOVKDTrnSIbd5SMmyeRfbFvAQ61GDa/qsqCL49bCDAksZP5nsIwLo6KOcS/M1IzKsMTA
4xDxBTtxX6eprVgbIpbYq+sUc+kaBDLCANFZCVSKH27vkvtDUA1uPQuoihgQ5lIPbxJgNYR5lq5u
U6oxOPAUUJYcUiH0VIN9YdUj1Ei/bpkGpTvMaTuRHmHH6XuIpc2sOia37GJP4w7g8Mrk3C/bf+/x
lHQUxV2j+CkfnwoU85C1fJnOSO2edKdV0JixViqp7t7OlJasNUVC4vuDZMpVjLb585XbWvBvrhfh
UBYRoFEP+xJ1e2l5IsAzme7haU6GKZCCTZ0doRuWBfOwSHJxBjLbEUOVeSwDT04Nkbub/GGImeeB
Qhy3u/Bj9MiDN4Zk4pIPCH+rWxRPS/sqoEWsBmsclcI4IJc8urp7AqMGrRWp4HDPK+74rF+oaNlW
0oMxxlReHok4GKynTpV4KnffCzVGLoQDZ/yLdIZNpefTRvGzaS0W67sJpjR4hC3MfUG5Dsr/PHvT
f9tAcJrNKPJc5N6ObBg2cjCdYgIXC3cvIE8Y+yAyrpaPse5BkQo62GB2uYhSUnRvntw2gbJ2OeVJ
c3tFQrif7+O3iE27YZrr+X3LbQaJsQAOvwxJDJJSxnORkQQ0ghiYTO4XrNtZ4LXglkbyfXbnF7os
IfQB8N82Cn3M7gvGMEZGfgyqK0JUI6VhheH2IsSKDLmmZn4Rz+H/rDUrojxryJSafwzpM/qdgtt2
QyiYgq/qnaCSaoEJHpln2CbeuRaQWIqcxAG45NqsVqyVnhTusCgDg5zHn1fJPKgVipqfsBgYVVmb
s4Rexw8SRfGnySTPxJxBCLP7lPDG2BYRZZHWZYWUTmiSnM7VMGS+ZrFiSPeQKPGsHW8nsJnUyNZK
wj16jI/ATOzMHX8rNWgHVbEQnP8oeWbAEbtx6NAni/fgZ4VUHRkD0J+lelvgmBuFCtgxfobMJH9z
1cUgcOmQuVnz6q9PHEJ5ofKYIyuZqqX4uKFEtQsW4sqMZVBg6yOFUSBFH1AA1Gjru8/akh47VETP
Llavoqp4NNllwLh37bfLr5GPBSPxrZF1TWbekmVIBZ+LVhUHT/t4MKuaxcuc/wv8GcHqg9qSKGpD
XNsQsQ5Qd0AnOwojb543FKUaCk/bk1JhooWyNUz+ZI2SNnPmSdudUJg7s81PJW7r+jveFKdth/G4
Z65RDy3Zk9QEFB2//CWiMk7eXzBkcx/uiaBKh15mZwp0WxNEHsVOr+tYoKNa0d84ElsCPjO7WsvR
99AOdvmSmAuQve1OShAyhJUVDuSCbeIw4uuHYSKMADv079F+rGCeTXaY9mR3UICvE8yuvjTmS/n2
iCEsnv0N78DrElC61uh6J+iRwKxgHI8KDwaMlDd706nCmbckDXU74VnNT1R25qwFSI/hFXJCmFjW
163dS/KSk4pu4ADjL1s2fqFmvs2GZL216SEMcKWM4rxlUmSADHPHOj0empSQE5Q7W9mFblNZMgWH
dTR9RdT05FAfzxDiZ0jEZDnhWrDAaJlDKB539Ho1uSML9zQCq5KJ47Qz7yDSLWULQySsJxt1eHrm
HIM2/ColJ9GVhFNACxKYSOiNwNESgm25YxKfVUT3Gh0cknEmnVypXYCxB9BxmyJjB3bO7YIDK/uV
fBneUzxwN7xeT6m7G8z4bK0B5usGQdvb7AuCFueh2sV3/1JxKYIq4jeJItWaeCp59usQGGNwVXlW
Z8WEXd5+FZ2wV4QXPvIeQ1yhGgWO7z6a/UvHm8cfQwlhulqHoR9U9/LRXsHVZmB7bYf/7HFjINDz
uPudmP1cYT+617t0M64WEjuKl/KsxgYCn8AyZo2idMGn9lr7zXgLPY0/1lFBxijTCABabU1Ro0zH
1C5+ypfXGkhgle78tf8nBaPGsrR8lDh4EWAOx1MFOcwcsRByrtLZTyi6oPvRLQlTkb3ShM3ULcD1
vKN7m/bosuVjO8PIiqkMWEE/QY5LuHgdInFZhVSFv8mZUv6PWh3OnMzRgACWrEVjmK7HM2wXou39
TSxUqg9KWUz/IYFoBrOVRlyuRbfdRp7KYl8m6z5hQmDFnFQl6QbT06H/lsbpNF70TJhEJQtLvAq/
9mS3DW2BOKNqxKXG21BjX2cPpXLTw2U2DOKZzk4kTuv2ba7LoEYPx0ksX0ua6oNgBdZZWyOsPc8S
G0KKauavi1njbC+YcJqK34VWJTZ5gNdcXe7raUZinBciwlcwq9c1O+5Lj3Zf+SXsiNnWdnekFcOc
1/WXhIx9cDaSWhwkn3iccLkN4vdlOFqkfvN96r+lGt/Pc1rDgI4ZPJDqIVU7DuYRew7or+PJDk+g
H6+Pr2GN9H8Pnb6uwFGAcU1d6t/J4f5RjziX8BJPvOgN5GNEGhWQOe6leXgFuIor6FV1eHNKxrWI
kFRwAwalP46awPIse4FPbPLCcPFD6JcGUgZaq+corffdBLMWLfCdsDPfRxvEc8Q78eYSTqVjm0uk
7yxLFHNnD2TjifNS7yYuF9CXkJw+W4GCoXbiS6DFkEg0pyBzQyITwAGjvh/VkuDP/gD0qbqvzpRD
XN2Gbcx1sKnIpyCDu0/lSboR4NI0VdNiIaiNvOhlJrKN8J5WlCR6LJPL6WsrBTpxISW7hT6/I2cN
4+KPpLiMJI106U/U1weredMJHHb6cty82JyPaahQMsVeRipBOFvVJxaeHn5h1rBBLwoXOz4rzp9u
4B/E57Y5znO53sp8+Bmd9wxVYz57+zktExJ/W7nULAXCfu7YRDEbtOxqQJYP2/i1/rp8lOK21B7B
iupV4CrRdV5r/R9j7l96UvAuNKNv+d9fwQu/Ic+3ndNgyQwM8+d6twT2Qstsd7pm10PJiJTNHR3W
NYjgUZGx+5uaZAnL/1g5LErQmWquUfsrUiTJSqzGd3HunR+Av+UujHBeEPlfkCJL9Kt8+hGLomjE
EzRWryH2W/Z5byvz7R5fjpwlGutD2Icibl9uBOG1ZsumgoZdNRrUWSBiAJbZJ4r59TncNq42d4+y
HUu6eN6YAPkNohewKNZ9L+J0NJwv2oYCFfy0uIteV499LQpGzvRIRK4KzPWYCFgwTPfVl80mkF+k
f643lNRZYvM4QL0z0py+piKVW8rZqv8Z5Vix5hLKJhBM3cfwgBnMMhGrwWPaV2uxpm3DuqH/9i1M
XI+t/E5iFDhQaMiUpyqmd3zQ6Cyn1bofEgjYaXhL8ohL6zlDXJxfs94MqI60AML/yfCsuoBpweg1
qJiuXGeXbZnWKKbbqkzjbPKQIyw34QWDwEG/lOR7llzTVOERIxBpiL/1TstUj22cWfscXxyb7zmj
/hG/v0CBd1GHux8Ut5je9PZedk2po7tUB5c/TEUTkrDeMMetpVdygPIb9D5lZHFitGraRLlQCCuG
g7Ff2FyaPEuyMYozYH9m7dip1gG2ALeSWUYlu/P/XdJfGMtPFrZgITZm+1I3BHe2mW/kgSmZnbbK
XOIMMprvhoybDG7paKi2yDM++B8ddhXzkcAbN/Z7KXCK6fTQYSTTB8Jq1y7DaVpCiuUaBPOUR3Hc
G/+KvMf6TO1VBCZlFTLXSWLoYFT8hvkiC9qU8q4N0BcYFbyJ3eXqIChlj/SV54rZb3WkjZHA6V7J
N95kg7NIS5zEwshsgqVaAQeGBfTUX43+Ilm4RqqsMMSJEzUSvnR+XioKo9AfIZNn6s6k3SfZxFlN
O20yyoqRWRU+puA+ZWGoZQW0rF8hAFHuGBg48KMJwuPCiPN4Gpu7Eu0OWx8EK1szmcRufIZO59Fd
4cI/GddYe5lWVTZTrer6L0UErsV4ffusTILU6BqMXGaU2yvAg8KZaVw7NgFS9wJNzTS9LM/v6XcY
pwcilyR/Gkcot5+NCUJtVk1fMeaXXFkER8xcc8WMNi3WmTU5CIoYhsKXy3c9Jar7L+++QtoXk2qc
cOrqw2pZjBEArObwCrltVuZeWYIMT1VmuqJ9pdIKUBUxFtzKyjJYmiWF1WtFicS5lH/1AxhbKrqe
CSCZDoXPw0s692XzV18+xCuS5zyeVtByaHoFPSmtpgAR8/gPoWSEsH6L/ipcNmvm/8ZRY3AGpZ0D
mRt20RCWkD8BKZuSRlGXLRxTeV5lmq/+htC5H6nC23dHdpAh+rJs8YBBphoi3FHSqpYzEEX6OHSk
XvSY0Ao9XKWJBEml1ixE+u7MtXv1h5PYrV6WyEe3WkrYLKasQ3LSU7+4XjXWqU8CiaiVWVzUVMtK
9k1NFESwZRMw9SB08LmZkbECyBFLuP4NmSEThqLhYO5/6xqWfOdJtAmU16gnzfuDgMtnweMvD8qj
YSRngaTKdjFrkJ/Ph8/w5IDgg/D3FLxRSe/krZDyvGcVakrS8JgPLoPKz7GB+XSYZhA5PozN2o/A
PzP5XA5qG1DLhRvJp2AaYaHgWisnA6vGFDwOjHtQJiAV8X8T2UQM7O4DxYZlvlnsC0FExlnjTP6x
1jqFkDdMLxbt5pJTORRkgDHOh/ztIHgxZt412ZFgA2lKhIzryOvejlCvQfsq1ycPpBADcbFCux2q
o/DYie8+E12A9IgBYyd5QZvJcT/SNnBnVh7sESz9xp4g3n7Gtc0A7f26ngnwt537J4DS3tGlWnJk
NZDyqI0V5m7qRvzqjG/DGDgEVHhDYqaCeAz3W8Hzh53sZVfK4JcCf28Rj0SQf9U/jzpldE9SkCvF
OP2ePZrnnfm5pYUGWbLRWX3Z/jKr0ZFvfjDYAcC233SSH4mItLUydQ44aOkIHVfKo1f0DzyAws3o
28D9MjpXyoKH/x2IVO+s8VnBUeCLOUK+zFw956/V01vorMJTqqhIjlybs2TIhO65xpRxAoDw+KJ0
vodF1zeXKAzDQ5ULo51l4O2U54BbOQX7jX/8/uQJPGWuMbZVbdlOaQLhxv+fjSxBnrbC3cYAby8B
/PL/ex/QeWQAnoY6aqNv3qqkBqxkZPInkZewAqDMIup9MI3Zl6eWbYER9uuERzSrwdye+WFSaHWr
gEJNvOC8XgXsBxm5uzOvJitIFIdR6tSi94hk6L6cDrSwrBQdnQSxUJzE7IvO/3JpPtvIuoa7X1YK
Ut1qSUqQuForTBeKxj4v
`protect end_protected
