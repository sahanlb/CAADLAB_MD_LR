-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
RLHT28U8doyPJ14ybVI4/70IQoFaO3V8oESpHSj7JPSBbGrtzBzzIlVUW0aqRroY
FspHpq8k7DG2k06Lh43homYQV2L6nGwCasfRWtokt5Y3kDuUGj+b5y8HZG9NhzFo
vS8MZNkihCnnoV0TJJJMQiMq8QD5d6Fk8g9070f1dJ7tVcgV7tH1HA==
--pragma protect end_key_block
--pragma protect digest_block
a5fswlvf3LsJiAH7dsTUv0nYaG0=
--pragma protect end_digest_block
--pragma protect data_block
M7KVRCKqKlr/f0MJWcFUI9f89NuKZafjW8xRiQTRJ07SUazQKfC7+IFGDXaZTxTa
Yni4iBYnbkXiZQR+H3Uhj7WIUvjAsNqrldM5AsL8qeM8ao9u8OWlahtqH/rmDHAN
aW9Cdf+gV6jVXOPzg+sECH5mdr24vDvmik2seJXL5DAwPzPnJGx4EjE5MvyDvkay
ZFfGaG+aueJvF0b3dv49bcpiHOJIAHd/5Ldmrn7RarBxBvXvGDs13U5I/Lq6kdNx
kGS9WjIPX/zlrNMAqThPGvT79Ns0JH8osp/8IxwL9LXOzrO3p/kbKvAhwFARXXIe
sBOKwG6B6YC5KPlsMkYWRH8d/QbSI8L6265hRYkVLfKmJ2FsyB951vJhHTgxqxr+
UcZf63n3lLQfRtQar/2aSnxrVkxiWcMmxeBB31eU3bcVfG2P35WUQXQmYcOJe+Sb
LQY8O0MEXOyJTT7Kknql/iGrhftn/6NkMUSi2Jol0AmRN2PkrKjiAGy0/q4wLJby
eDO+Es6ydCnDkfpaMc1YlsHJ0lHJy2Tg9Lz8xkc6yZqJvTy9OAYD6O4+nvasfzMz
d50DdsGIP+Shma7Y9v3t+DnfyqBg0+3EKYk2/YxKI3WTokURc41SsVLcJFoiB53z
X2maA2nwCm0VaH6lfOO1HjHGxDv6YiXdqheQX/yIPAdmY4prQSAl+ctfytnCYl3h
1V9Rj6HFVppMPz/nn4In7Vp6PHsiTOP82tBBfZOnvRks9hsZDHGmI5KbRRenGFAc
cA15uFaKibQhhZYGXBiB2ydprRQRvO9Ck5WjQMzbbs6FWzbrYv0Jgft/mTkjuxA+
npvcRMR65zO4Hqe1KIA+6gX3L0fe6tjDXksKyYmz17VHA8ECH1aYtaris3iMTUgA
8cMFuZ9NdqpaWvU9WWWyLWuGxvQd4y4jo1FBV5JHfUuVdjvITeWN6L88/cgevsZS
EucNsoNgFEqoacpX7Im8h3wR4Lgniz+hAD2P+3tbCO4BZF1zadMWcMs2GrTbqJJQ
fMQYfMAGeRWfsQuw+jZ6TfHO3XuHomFSGdbzl2NDbLN9QRBHRzakO+gS71vqhYkW
F1ey2DVPJnkhd10Cm7nbJsGlSxWvwbYXgp4aME1gwTS2aOz2vDuXWooWHODXb2X2
1Il6KZ0VtyiIFlgMHULkgsr8RxbNlAoSPo8mqEGjjSTD2yhCAwUrVcI9l3p1ks7y
mwyVJX+K6MHKWH0eV/xNhHD6nwGCMvpQ24A0Gqg2ok23dhEkGK1EQ2znRR8Rt6z1
6hm0N+TEylO5KQJff5bHx/5H+aYhK8BjnumMs2KmYjdT29op/tbFkUzrT5ZUSNgx
sdDJPk5Dp3jpu38GWMpKW+3DTh5vwlXRujUY/4e5I9yKpiWereUgkStSsZPYOtFE
RapAPpyYo+vtZVWh2L8Z7i6EekMDpbahs8pMBQilK/m9w4LCBks+61HeO4BXsdV2
iDHAUV/ALJEm7MR1OEKePXJn+B/E+y83Yw6tEo6R0ZR5j4X82GZN/gSpVIYh4Dcz
luwpjDK1DHjgBLGc+PKwDZFOaPkgv5wa5yvoSHBvPgVKXVYRio1+V6ts+XXQAP5h
R+4Av+IN9BJNzlV4RaVega3wSD7syqbpj/mF9y1Ct411fitMxq3q1TwqZ8CjZtZ0
IqtCG6wJq2i0QyG0Vmb7sRGG+wfqxFJ/vM+ZZVxW/K9irygWnTpL+hr5VRUV9q5d
hKwCIUBe/BFuthDeMhhYEWDJBCJDLXTBfvJXcNMTEpQT2Ol9xTDRnOkWRQkAXo+B
shCStgXHhcl1dmK0cb4FYDOE2GXZ0PwSYoFcmqzoujyOTh6Gepg1YBLvHk0BDq4M
oe6DERnnDfVok52MFntHqcvV5OHxJsLq+oXV7Vg59EzXUXlHmNGvmmQFyaeiCwsP
2CHxpCrWajRCr9tC10QH2Iq2b9R4BboVgvuj8DCC0aYz5F7TqnIltrVt1mOKqTSd
E2h7yxerYQcRUuLf8lS7FAfcaG2KDSVvAnY6EjZUT29E3Wl/nCRxWmze0RjVBLoh
QPtEXT9eP039WaaVqQF7/F5PWvONndLGE7ZZibt6HveWLAEOkRNH4ug4+hcfP6/g
0cxN6oL5dA5GYtpT2Q/wpOZsJmvHj7ZUbIVfuvrgaJ8z4AaxmobjdSRBmwly9KTx
3KoN2epw7LpNWFlBqlQF2o7CXOLgmZe3lqvn8Mdg730hkJKCqBrGOt2W/Em8e1iT
wxNXRRDIPnwzPB3ZDQSNuCeNf220x6jmApuENapc390y3Uv+HX4jNU369qKQ5g1X
Gq7C00MMeI9aa7J9xKoQr0RdwQTVik69+vJNt7HRvYZJVkaL6K5TI3h7tkogmjGh
VInHuA56AhH6Z2K+GaoCIG7Tz+VzXUec5DuXYj3rMq+6zrHyd/zhAwJ6f7esaZFV
wlEeYXF1zEOb2TiNzEaO62WjX2lgaRD33h00R2J+XMu9A+vkNSuKvnpFXwQQlJTR
RhWmTgaq1B/0l5xn0q74rZrKB6nGGX6YgRLXG+2iycD5rTngNE92vrCqMJ9B5ai7
uegmmTIuR2tt9sutdhiKxcCxxG6dAdpdcAZyOu3GJNT/283UrQqkwbFkW3tE2qOc
fGtlFGw1ZkFNj1XdQHDsVU+Y9BkPcHuBY4gDUHAOTt65Wprg07fIcUD4xeJJOkgi
5sxv9d3pwWWAMIDqZWuFDm+dFDu0CX3aB4Z/MozsgVxrkGsyMPqpbznBkRjz51nX
YMnJJ8eS7fA3RipFz6gl8i1gN8utaYwm7gDdVDvnaiTq1VbvZXK2WsKf7rybLwmu
qN+1sQbQuliKgIFLwdfGVrmT6Q3Dk/sK1P10IxJ3cSzPPJ2FYsZbuosq/UXWoOIv
umbW7S1ZeMyvD3mMaLWTZ6tvQyZVaR+jO4TH7ZEwHrvHglftQCHV3ngzEBrLssfC
9NKaWRcPjITrYAF7dOBbW0aPrLN5Hgj0kQUwjICOTyPhFYTuytOUo/HF/h+07HL4
Xk5hFeeN21kyaTIfT0uv/HM7Qs0xRzaHqVEDv6cfGcsmTKFwVSj/ZKTvfTNUnkFx
9q+BpTb6hssBUcmbZO37lKIY/FQL4r+/RyggbM2+dK5wXZ14WBwROpeMfdjATUrh
CXzUPBCk5etRRTWKlryO7p+DKW58U3JHjBEtLwJ4Kjydzp7RdioZQf4fF8OuZJ4A
9i0ZNIZz65JxVAqHfmKqP47ZeyQ49YVBz8nYwjrYxKYBKtzkTrw4xlrSLrcoCgzZ
sfBUIngXIKefitYuLpMspxc2n81vL/7SORfxD0PkbByKKqh4m70UNQYD5/HngKQC
XiPb2c3BqhJ8wlNrJL/GF8u8fKb0/F9VjFGvHavYuzpOzFsPipMjrr+cWJdSb4Kz
Sgl67VtzE9fHrJlj853a/817LkC3J6+WDY1XTtBy0JXTejjOr2NNithm3TE6aj8+
ECw4pIDGN2UWav4x9wQ+pg234Lsq8UyiWAUpMZAGeL4AwaJ7TcSQ85dAfG7o9ScP
evQP6ucJ7ipiSZ2670CbzcJHtVyn+C/LPr3LtCewrHrp1/UNU8VcWDDwP71/GuPL
GzhHTsBDyua0j3Eqa641M/WSP/VbQih1Rdi8bVxyLJ0HcYCiGvAA1/8eimGFJtlC
8xi9qKwvMeIBb+Ly/qTeQSc9wWE2CTdhFoK3+fQwQ+79TY33FffVvi1BUKRfkz9D
eMqhWKM+Msl/cMl+Pk8zqmuSJqcFBuDrmZ+LVJVOzskRlMMtNvs9kxvx2GvZyCgl
xopdN0PbjoCJZNMfzkCynrFtTIvvjI0cGuKd/FdRNGJqnlQRoaISMAHs4i8spJxK
mqAyHMjrPo3lUp5edOQDVx5n2u2k/XJ+MQmfoarUk/l/sJkEJ4g0L4LcN96jo/e2
qhQ+9d5jCmF8H8eZszVDWUt8tJnx1jENguZ7quba8lgoRcks9aSl0KNNuer5kSVE
k1yvF0SasfreCM5ARmUMJdXfD2PBq/P2cFYNCRgmBJl7/oMNKn0n6i9rAQBGK73a
N7KGJkXRCr+hYSw20uJprS8Xc2aX7GuZBYUai6s1mdyN1zj2YKmbWqT7H6cmQHeU
QbcQB/vtFbi8jxjT6H52UuN118BDDCMafBC23dtb7/hsilkiSX/6MU/hoOevYzeK
/BjwOSCIdD1Mb8fikZTmOVhCrif0iPXnfy5Ng5a4NQ1Nl0HPW5QDCZtmzuGNq1gP
yb8fv5XYifdRHYcGSq8iFHBr84PpvrY112iRq3r+m1ay0AOPojoLlu9GrNlwJWcG
kukEp5XUeyWOqWIT0n3Qsqr6qUpU7DkcQbZ4uZO7NyQhQiphVLOsG9OSOuoO5GcK
UhMTKGn/6mOxoprdaLl2LFiF0YUFx85/U1ufIzNnvE5TV2/F4SWpP0Fk79YSwxp1
og3evPgJfarXI/QJhZ17xczosyfUOwuvSMkqoKqDpSWPyTVD+TWFk8A2MVC1OG84
R8mWYN/kUl2WAcGXbFTdXWJH+n0Zl/UoEFVTcDhJrfvB3FDTuTEsl8rqrbWY4zh5
kVCV+5MlVq3pRUywYPtF3AY4JZTcEEC1+d5Kyu+kvQyRfwryHTXfcFDXrSqWPwyh
l1PQzqWjVzMGl888vrmn/khKGo4zCM91jzSw8ND2hCv0mPQjXtvtHRama4dD/Sue
0QTro3282H0mItXG1IUJLYcr8weLfKMAv85Cz8RGKtoi0pMbdso8q7a6pXepNl8O
ZOXOWqj0soPG0Myh81R59If4Qz1X7fj8wivmNdylj7bVHwUM3/+57tlObJmkkkTQ
fpPwJREssVel6mTUwlgTAP4HZx4z/vAmeDEp4/HjWdk6232uq50BNKqW37Rcnsgb
WEq0xnvxg/dzkreH3Gs/ghZnrofZpnqr0lHZVwDZ6OGUYL/iUWL6jjvKSewaxqAD
fHVj2bw0/TiOdQg5lt4vF+6+RSU5QhGzhmBMIHPlTz1uilUYEhWpKEhrY408yYUA
QRgRCYZOuzQleoY7UQgpLKeeXcUoqwbiHAt4Tvc0in5RPtiPnlEE3otEtPGjC+dA
XQGS9SoI5RkWZJHW+UM6i/AM8iILfkjIxaMLShhPwjN/yG0VomKsbNlSRZkRaDwv
VILDVMuws10gjKNQ1yu5Mmc5yJp8QtU4anJrWGxvzWMtNfni3D632gqXkJwXAUDc
uwTKu3Pq/7K3ihHGhQjSjMfYySKnuK/8wtYn4/Ig8ZSPXKFayLsxmcwgTEo4dk/9
TscJi8Et0o827jylq4OR/GYAOvWCjCRXcVV5J9YFDKxm7o5zzbFDxK3IFDPHqRl0
1YQYbyoppyaNvQV4e+1Zk+uqxjofpcRECQyK6JaTRTcPJteIedgcC+Yjq/F92EfN
YrMX60srknNr9NYZZTIeV4rGhHAcF9oBsukGDW+XBtMUukKr8oIjhB5/Ff3WelgB
xQQg2y5GLdDG5vriRH0cNajzgJcvAcVszmP/ygkwplxzanNyslaTGR++mIvN3zWM
ZY19J8eM5l7KbsdUdMWvrL91fljAUGAgdyqEDwOIl2yaCq4gG/wFDUHC4yF1n9r7
odEDpM5Ng+Pn/AvGeuqlj4qoxhw5Gz3sPHNvuvl6aCh5Bq92Umv16bVnpK32bahR
dkXmp4T27G6IMVnjD1+FA10YtfigJTuKeWSiMySJ7hP6/OVxpVxFxC6qN8003M34
MJTBpRCZ5ZILtRftHS8Snw1teHpdZQGEyUz3O3BS00iKKxJhFBSLKY4B/HpKsiAT
dbLzrRC06jMD3fHDqAiva7g7NunoLPw43MU3Qiu/GJiUyXO/iVMSD3GIZOQtazU1
KaQgQTQqO53nIPuhKF44Fv5nKb8WcdsB9R6MEhXNni0NaQZMlNKkMe9p8XHTEEeZ
ulO1rd3stoz0xVJquKl7gt+s5RRGOi2tMOQZoqZBNyfshwojWBUVBaEOSLP0jbOm
9R6u8LJWVIiDVNxXmlahrNd9ZLq4g82rQkwTBflwiZkP7o3IgiEyTpMr9T0wj2zl
hbgFQh0N68uDDk8Mn0brTVswvTwMJagvdDbaPlnHIIKSDDtcUrb3mpZoqfa9yDl5
krllhm1kz4MhtVs7cS71JD+QsFeHZgjpOim8E2GmBrlT1Zwlf1hpziHocSQM2SzK
gI6qyB+DiFDu4Rf2UAGs+vUON9ooHoJXWS1qCm33owjvqiKYakt2AFprU69GbnVR
ZWX1F0iQtXgvT6CU8QamlbbLB3KBiO0kRgNFUmhrpIiIJXXaDhhAO+gY9tf1vxGu
kmTJT6DDY4SRV3wX2SZbVe7FHkcXAU+WE8H8oR+ILG4KBOvIMMyvHMwWBfuIYNiP
8ixX0WjJnzAFe4/Fo164YMZNxd8j+n6SmR1yKqrAfARojpzbXlDRnrpJFxk1WI7d
B0ViSnO0tXMCVQvj9nES9RgxsgeX4qHxh0ROcQiql/znY5om6RAkb3m9Z7kLV3YW
7bjxhLhRz7SIpTwI2Ah/isi54qMVXGuuhCV36C+fe528LQeMr9CFtzYY6TON02Xp
Ivp5JigjrwOJbHcE6H1sz0e1hKeze3YII+9OR4VH7ticIbVP9iThwGcbg4+3FPnu
R6/wtsp3U5oDm9GcQ/VWV90QJTOrYkre9QPozbYyhshK7ituWlHOUKG9GqbjoCyj
0l7ERdzV09IIVYOcyDpQhEr+D3BuSjQQiUwUv/Q3gcQ98Z/s/bY9t1cqjl+tNod1
kSC2PEwYMzAr2oJZ0L/pcZRbKo300GrB/Ms5+i7XMQ6wcJdz8YEqxOwEUw6rupGn
Wi0y1kSKXun6bV8Vstk1xvK6BWqZLtt4EEgmO5XP9FIhh5fsjY3blmBc4qN7h5J2
+JOmQr1vTX2GrB7sLj6+SZVNap/ZRcpo7F5qGiLRDo7WA6Sz3pdY6psT2EiPCAog
ldFjq7uUAovaG7IHVjjRatevk9SV/uz75NokYnpJPc6ytY/eqxQnqwRmhMLsyHcH
vvgDEvWN5I54m6fOrSH2vQMMHYPAlw//7re5Kh1z07nHtcjRGYDsWkmRDVPknQf6
afDQyZfMqz5Ez7x8h3ngBrM+dGYDPgIfjJYWU6yJyvtszNMNKyS9dpe5D1GY731u
SuLgMB2BBx4zlfSrhwgdeUnWXsK/nUJV2vNrxPkG1IPeXQ4nzzsVXYYCBSSk3jgu
c5QQCyZ/bVF7VbOwhHZzlwAJ+mZMecgp2jSgScVBjs6GOswbR1PgMnf244y0gYlQ
F+PXFZHT5rrJ9M2Jc7drtFwjGJe0gNaiPtd4MO4gWiby21FwwpSPWdVzeAi9UfGw
8lm1urve9kWZ/t1XjjA8CEHzWoMEquitTBg0gyaE8iw5dpF60eVa2G9Dr7S6uwNx
3zdCe1j554RxCzjmYkFZHQYpB4/LuORGjn/UbkS80ENuWwNQ6pjLKF752S+oXlvB
HNHqcN6SH6bqdDnUGVfjqsWvjaShpEPUF38fFiS9n6m0K6RT62OprQfT6bH0L18W
54EYH9P9b8y7K0KHA4VXPHPWvAvWOvHUyYL/8V7obWerFtweA+kpsuX1s3sYDDkP
FQuNPsdtshNuNAIOWkw+5GMEUNOo2lxG3c7q+04gW2loFgp9T41a/yef6CCyoiIy
NG8893qLKAJTm/gkMKkSADhoK4H4Fu+2UT+UTVY23VOe3dwV9RAwS/5zEGWOLkfa
YH38QJM0MPu2GqQIErDQp0/lmZSE5I4BgT3dvCNAZSIb95JMpFKdE93v2isGeEUZ
Lx1ZToxwfnBThp3v3H3vpwjdsbnMBDJFVSf5tkTyM5ahk9ft8eS+V8gXPP+8T5Kp
5DGC9AF0nZvf+240fNejma1NOvn+vnkjmu6/CrZ87KiwMzSBWcjxClmDHZUwJdDI
1MWcYC4UVK33LkSk+P0HaPvlcGfWBMXohhFpYEztxWXIOHg31y0LBfsLJsx7uBbf
uHpGOZ6Ln15PK7qduJUNuedmVrTBAC/+8yDoimCjQr5QR3vh6XNsV6eMBk7l9uD4
VS9Iy9OywRxq8aFMVZd0fcaLiWadhJXO8T3OR4qwSIWpNSWCCxlBN+CG6E/u0lTo
+WeXl7uTiG3RzfTS4R4cf6lLn41P33jk1WxhvLT/5taRonBb8tET89W5EuadhrMJ
ax3Po6QbAq8jVDrcjTwujbrSgL/oKqtD0jRfaIqda+FmaYX9QjNpOkfQBHT+sv6j
LNGuP1YGS4jNUJk2LGXyKqc9amE4s7Z9CWbxSRXYdOIMge9vznaa3NafknFM7jAM
nkRPlxt3AxsaEOD5Fk8WiNPPthFWJb53QxZmNNcPmjz3DQtOrWw1FQTXJGatbeLM
O5rwLl/KzcPBl3vm87BjkR5jQ6ENjogQFNzCOd6/c1a6ioQTJ/qotQ3WaQhLCQ4W
AJrt3LwQZw0O1iex7/ccVFL87NQ2xeBSofjPOwMb+VkNAjMhDl0PqdQMG300bgx/
XBTmIT5AtC2/TGx0pXxAiADlBAFZ5FwgHLZ97zZ7SZCYTczfK98nJe8sX18Lty8+
yAGk5qRrYzxC0w+5HVjNfIRJ5pZmPCg5phBtyfLtS1IGsmOPGd94Zy6eGEqBXbx0
CocoJqSeWTcnyMMADBWlxgfQHcFtLtzHlpxMphSVX4nLQD+KIpa4OMK1dDAGuGSs
nHiceRtGKdiiEXU5XPoCezjz7t+gyKiLM+0q7zPYD3AmPf6aSJW3KZAdoVM/OeKd
MZ/RAu4TtibNLsfQo8hmcJ+Jt7VShqQnpOXMdEFS+k3ncaW4FQAimy+bxYeqDK5n
lRMuykz177RjN/yYpfxj/0rlkT+zoutMgSHDoM9gF62mvlzJNLsBNxzrK5LlUlYT
FTn+DXyOXIjyJhSpQlTqeR87OT+XezBaGayzvvJUJoNWwmL67nlWPZyPH7aVo4eB
NCuqni4fYq67DQl3iZ8Kpoa9qSFXd1lN693zUdIGvejERM1+Z+bvcYrlFfNC5FFA
PmJyzM783ORnKnth11vPSAyX1UU6+llMPHgohAGQHPiCGaMRemNpmu4qAnN4g9tz
l+vW5aMe1wuB6ns43G2P+t7IGnjPofSmEmI5K0qbDNRzpDR6axD4XezJfV5oWrhJ
7RbnYXdQsZJ4hKH61JhfZ0FtPDh5+qK/NpMXQ1h1LMIPIlodL/7ljrIG0dP1waOD
v8tk/8+6bzF/iaMsrDbSEhCgvf+V0fvvQS31V9um9o+ROJH9QnvHJcHrV72i5NnO
g/a44hrY2tMIQpTULXJ8jftSdTlIWaVqslEK3PCmfTmygwQ9wAHWGMDfHfNKzByw
Oy5kB0eDoUU29LVbH4i3EOllbADQbX6yPcWR6lLZnzoUzsW7B1++hWuF2W0MRV0q
Hdn5zd4v9fX25sLZQFs1eQuSQkLDAf+KB2ol0EMrLeUXRuy9hEM1HOFUbDqKotxu
S8+Fq5x4fgr3YyNeOWMqac8aNaj8QwrBeB86QTTEXRDRoSGSR96gd+HAGLh9lQ1Z
Kh/PQZM4frUM7+WffqLCeDywm1KeL5BMzuNLWYWnNCBcTeIf2r4bDKrw5fCeRB28
QcnMP/Y8BTcFdgyWSc9KcNp3rF4Su9NbzipbCCO6IY4VMeYvWPH96h+19E/nlovU
tpa8/Fu4KP3UTNMuf4brYHHP3tbN+Q45m3EGdrYdgiDhcEHhPVnTRDrMdpex+cwm
jAgV4cQJ+qgLEFXGiU9ms4fim4ylDGEBqzhZh8NQ7Uj497gnhHbuxI+rHZnSBjfC
j+tggCicLujvA68xYJMPY3mGK11GmVSAQHkZw1wJbW5BqJJ8yHR6xV9tA+Zp3uy3
4ZgwKDxdv50wUOBYjLQqgNxJrk3m8W3IVgr1RizivWKjI6x/ayu1GC9+x0WQmrqd
EShYpOOpc/Vv3Ves5D+7Ciog/r/NRW7loZMPg5wSG33fbVIPgKYEbxbbzpD1ulPG
oGlenzXmV7ylSe7El5YpKSCJivEvI48kgMQpuDd23S262hjMIJ4U8pYHUZTdjcgc
898YTANoedCo4hPtyVRE6AaKxQm4vpgLJbVMqyLgWwGPHbpKIJ00HGEO7Fu5WKiM
Boi66wXqwW28E8shsQlf5pWz4pibD6IefRUTUb0BVBIGfuKjOcdBKwNLaP70Tg8s
iui7nuE2PYdNAf0CDI1bzif4A4TGj9tsul4C0VPE332Iun8vItok0civ+q1LxA0T
6tOdOe2WttBA7Gx7wKBk+XQ2TsMwe7aFhf4K9xP+dy6ihXwhYfGAJgth/oPk2hOj
lF8Rrk5QFXlYQQh/UbLuKa8+1AT++fCVHDbqXe23rOiz3wvYuIcFOewVojxTQr+P
GIVEdHn8WvMc9UZ8Q0rN/ua35/ub3vBnz69F9zjtKhfGu7FjGmI/g3HZ2XKPmfXK
pxQa9iJk1E5Sf+38SqpbEoPeaD5eXsIQE84VxQavzBpTKXqWyf6O7nVp2KhO0Uky
mLbNk8OjIlhW0ZFXv6ZHh4uB2Vy/hB+hyAazE3mnPZvCwsIoLviN/mlsmCxNbdZ7
yshUoaNrPpS3ccTjiTqOa6A3Rd35lRvrpWa3L90hR0TsfZQwbByfZW1rykcxZv68
QjhC7vteYXIefCcLQEflyuUPofSzNkkAb31CbQ/ZQDpOIc8INo2+eA5UVvwuu/Od
EPZ3Y9Et+dLCHcQAK8CvGxxujj4UXemG2g1us3Keg71WL78whlnGTta+A2T5P1BG
swjoj7vL2b8MAtatEYS2OUReCSs7Oj8an/UhqWETOGBAbv8Rsw/I8tqM5Mvcqzxq
hlA7XAW/6en+8ZdWOaES1F3RJsM5JAjnf2IdIQGb3/QSbabRFgwrCc0tQEEWrZ7q
7g+c9dMiNebS8VGydDzHf+FEzdSTgWyuuB+a2kHHm1STKUsxCxzu2hU4JF9lLtwi
9jcJbQ/Ud7Nx3eV3lG6t0b78gf8pNxqOAjNEFUAac6CX2PDJ4zzdPYjYtaMuE16Z
BtbTT7w44HqCTStkJXa3PYqe87jkEx3aW/M2U02VNX6PEVT/PTDcLPnORJy8zsCv
yXZw+VUB/KBLjpqsMVogudqzw8f0NJoDQu1t5GUN3kWSm74FLFsPT4aivj1nq0Mn
YvYIyNLohown3UPBbw3g8+L56Z1Yo64K5NvlytJ8TvmNsksmSOmbc6Ngqh2HlWHI
Cel2pTZZrUHXUuxQ0neFVP3SxwRFNiTyDymXu1x/LsNN2j+HuTD2YEYcEuNk1kjQ
b8rNtwj5dFgF0DAzDpGUk5Qhj8SMU970bMqhgWfpCsJ5Be6M4bfZvmivXqF+sru0
iO3h0n+VPQMfiBbMn294qE5falPVnH9bGHzVLrNYYwROTKJ4uzbTthstcn4vtyVR
qcU322GL2gOg+UEN/YYKS8qOZUIr6nU9CiL/zU9A+1kJH+FuJ48RoVYtn49YhDgX
kFQQZnlhC036bSu5qTA2ChqaBhE5GMy6x5nJasH4BhUu+2pmuV9RjxqFa7LUXXql
aTgXPsgUsCexCDa20iCv/iHxxcFq1shSFjpy2grhweQ/ytnhlZZWkGV0Od33b7KB
5vbvhhb9FsT5DB1fcvyFoS77/4bbqzhePiLqZB0tjnZgpJgCb5DnAke8dQ+Cs42B
3MIjaawwIrIMmn+ymFr7ATvrgnVUMbO9w4RVAr/hAAiPGq9VEuDTHU5XcZmL5ti+
eemro9+22Gc0hmPW19fw+JWSF8rUzzWdy+bLYy047Y8UQzLrkE7Si0mD//l7FbAH
K9BidfMHcSPwRhoF88WJkarx2NLqjJ7EeOI6USHxOnzuDVmC31aLi0wZMdaGsN1J
5l/fm+SYlsWOBf0dR1tbCPbloGil0ZswrqfbVXfrCvj5LzvG0NrfYlL/nJkUZHT2
RCGyJOMOOCITeEqBfJKQESJv0nfz4ywIw1I+cew+SmkQiyQkd/kn917uafXKggl0
00aajhy1Jv5uEx+2Vfu8B9rrjkXNhpy0YCaulKZRjdPNjIMyeSQZqUUKGeUbxWYG
LdqWABhp98LnaUPEl1V7YODVRPoq8Y9wgkzyAOKySegHZbMZv6Lzoq+Ie6pEyQVS
kvGV/X7XuQIQGeDB9kLSTczhDKzON3qwAeu0oF5Y+HssL9Gt/dEPZerp0aERV4Ac
lEXNic3PQyjdXbRijz6OCW8zavs1WdFyoMgqavZ/5KVIWTs+QxQNzEHZwC3XXiWV
xPMoltl6RQT8RA8NaurxkUJFJZvOPkY4Iyxna/j6lohbwiZTddkGOH7d6T36a841
VxBjJKYWmFC1IP9dRSjZ3/pRL6OKxFk6MI83V0mecF4XrBwrmOD6PVBIWPvPyVkP
K/Llilpoa8iQr8F14cvqH91v44wWSkubRr/QPVtEZIiMvoarCCaR4tILKvS7Is49
J9ElmexVB3SBNZaXuXZYertARXNflBn2gnwP2ObnUcQlSnNm5jcNHujaTdzlBTbq
Yyap/WGk3u2h9DzNz4WE/41kLNXVPfyscLEubVwC+lzOGibMy863Oxt2aUl8/AK+
xfbJNtYTPQIGsS94ZH3M4XdstGzpau69Mc6X+nR/CfGy+jbOfRsVKyZ7M9Qx/cJA
kUoOb1utMmRSLrMxePYNB1/mjMfYjw6gWN1LitDMXkGAeeGDQhxTOl8wYaFEOv1y
z8vr1N3niEjJ27U0ZF2t3MFQyldpMwWup+G9Ia28+Zo4GZKZnzaojs652G+kIGmA
nDW9XbMR+9YsltfLHPZJRZX7T6FHLdUrI7G99IsHNxYpWXVbedv1UxJ574iwIVZZ
7Mp99OcpCZtOrJtn1rLwjuxaM3EKxFOyzSINuU1a4X4jj9HLd3evslk80+99ycRS
sjr/2wXC2hE3VzIuQPcTNpqtzyk7Qo8gHXAKHG34z4CoM1BGdju52bGuHkcE8Jpd
/Yb4j3pn6Cpn4APPWeOQhC2zZd4pMIT4liFrIkiEyf46ruB2QtHbvriVfHdS/MEO
l/dl/+dvSXu92+umj45h7Lsu9EPYxjvHAx1Z1suzMSyLROxUARDW6W4cCwlDCaX9
ZKzqPqSE+5lhWvO9+qPD4zAzri0IYet7cvYGMU4OenaQwUz9uFFuTBN9ETJAmWEL
FUmO8FMP4FXSMjcFxIYWCVKqAHtni9L1Ruxe7ElkIx625vA/6yvszXKytpeM6vxV
ae8KIEaMEXp/xnIB/CIuEPAs/RWmuVejZprNOFnaY+gid0cfytQbNrQ6pw3zG/7z
Vh0p5M7alHfWJpisQvLZC2mjPJKzy65iGlFmbJdnlHIqHemKREOessS9/TbWOhd5
OycusNjY53zYgCdQ4TM8nIStltBY9zfkOiqVHj+nlxqmkFVSPYTNNqa13lKUkhX5
PbCM1U6J2S+TFrIWWBc5Q7y1mJbmQLymnjuEDkJ7bzznobEvQOM+D+hBi5IhlBHF
D6twSzGNdrqmE6JqqakYNourkMXBG0ivW0RA/yIgSHdKNef8qsC7dNUQh1OMf7E4
hVzggMvXNHlrhI+TkQtEQSf0XtqaORR0cLGmK9WBkwB2Ule4UefJl6B3jew1BWmt
AjgoRcRajWybMsEYG1IgHOefheEl5fGc9GnbBZbos19lGijqsTItb7GdeldmI/q6
TpHR5tqxt70K/Smm/eas58Xf+Wmstfv7IB8q4NP5Vb6k9I8SM4HIQTDG4laZuJUM
GTXH6wadGAjvfoCqpAjkROGdnEJROCm/soWP+xO0bck84TtKHbCBJayo4ZVl8j4j
JCtBzI7JZCwodthtMsxUiD05GqtdlZ2w+7cN5FAqE+EXKsXCYrwqH/jTW89yx8Qa
uXv7It9yse/wCxWzgJEpaEA+cGIY6snAk8rD/FUBFe3SC/irerfRrZhCiv0P/AIy
THN3bkYawoSA5kBySH9tjIs/CKSPgInN4ERhyqO3ni7vBmIfRALnUYFyoOrQENRQ
MuNANzNpY6eWG+x1tDY8MCvuC+74I2wQ8E5xP53MoP83legv2loIlpwWjVSgJM5U
d8hR6x2BXyQDLah5BF9Iuz2Ajmc5wZe+Y9DUVfEdRvEZE7hJE0jvz3bN1FChudbK
Y4MdxpWJrQbBCtyZM0lbLoRP54q3oD+1NsodovxtiS+/V3L/C3L4UJEakN4Awb5T
K71ySs4Q5hsuzB+FGidqOLIRYv1MxP/V8wtd4w4v7b5yuO627O9mRpfhltSgG1x4
LiNHTqUoX58mFGvq6QliBRhlg0vLG2IxqYEVyiOyTrHCEIWSHNIOFyzFACh1pZJZ
T+IUEd3WqkbtYddomaL1kM16kBqkZH8wM6A8zYwr9z6gOKZyyvEBPfGL7wGDSBpG
HpeSvaDwpFFsu5jrsLYl88ZkaVXtTuUvDzipTZKEwmvlF1GhUsOkOUZpUappI5N/
NFDk59iBq6bBb6AV/5lwPkSXVttTTRQeF9vVYFaKhdecSaEIfTpQ95+nsz6rYtVO
27Q46QMIDoZYzFwde/B0It3KxZ0ypLspIF87SQA/bc4nzNxOlz6b2GfkkbtWeLmj
oDo3aVXd+fJwT52wPdJ0ZKYIs00z3HOGbjnkPh8n/RYeCx20o8njUxSTF0RphJpP
y3hD2K2DeE/7dkC2TALRMDZCzMQ5CjM5zwDGDRaftPqvoYt5jFoEARHb+4WnUsBK
51whY+0cYFHmRNa9CcmD0QB0l2ugt8viSenmGQRTh61nOBh5KktTHXOdyFRwbuhg
ag0FDvqUIWlW+DaIPDpaspa+oGiSj/V+c2NNMzNtuv86lncwpTbqCJy7OjSwpBhM
djTwz0Qo448/+6er0ZEMPHHZrKwNw58P1PblD2B/g0jqB/Qw4cCF1PC5WKjXZ38T
g9J3QKGC6ClIgEjaiNPamnUmEZO1SBVLymhj8DaaaEnQ5akHP62IlLlBJBo8gDA8
zMMfOt4xZKVBXg/0V00UZ8eBaOEyQ9QuRZ7c92YuY5Difb2V7rYdtST7WevEoEhr
64t8PPKw0lG/mpb3+zZdEyWFIjvUhoCg06P8t1uRTxazXB6zmHnrhmHV3KWih9RT
FD5HZiic43GeY0Aaw6XiEbQYQBSCoxsbt92ocURxFvvdpVbUpR6zMc8e3bW4Bb13
FLsSmfsGdeYp6MPmfxY0KDBHBSHrTtVQG4cfMfbLaJcrWzlbZkI6AseijWx/FX9C
zErCd5+koQuDxKpLEwKDIZbzBi4D5r+kbAG7YgcmWaYuEmlk5zMq8uR6I0p/jG4w
ZsXk05oIBQ0jCatux28PQbFGsl0fsVxlau4FwSs3BCj8hzzsaHUnaUq0EF/zaRvu
oNxoGo3Bj9wwx93Lpksc0UxctJkz220OboT0KWfUDCQ/0i1Uy1YAQVM9d3MJi+RR
ZTQvEbP16sx1wADg64fDnDgzoJ4EMjAnjTVOJi76vCv4E44KWvha7sjojm4Lzi7X
zMYmR65gSp18p0HnJ2Q0KRpCkAOxfFJjBDzXb6hjxgcHiiXlctMMHXNhuebBpS++
iRN7QbvsJ5gWh039sp6q86LXYjsW2oOL3Tm3sC+GPtHsBulgiCRk0ZAwlZqIIfTX
fEo8zLiRsJj8FwFcQ6LFCYbuykfXI9n/76IKfCZCJ6nfhrS/BmLlIu4JrOQRlqBQ
sEls9/q/kn7rpJ+d+LJ0fBt/8q9ZkWkOjrRAmH5D1zbCjP5iLNUg3S99S23laPXQ
8YrV5vrlUVgo5QGQu3Y1u93PiTBl5vJtRkhW58Ytc/kasGye6vktVw4gjX4uiv0g
jFb+WzPG03lQRYOVGduTCwHUMmwAPoteeToJet1MCEVh2Pxi1nU3lYFY5dPCDonL
lNsnJGrwpOe21pv1YvTGGpe212y2yxuKam1oaMoZY90bQI4wd1M3J65HUcmwMwdT
OQC33r8X7fjjsWA3ZeVq/ROOF0ksDKyij2Xv3jL/ITWxo8GKK6pnbOJUvgLUae9G
/Y6J/KVJiY4rGoat0BUdFzo4pMm/3x0MuzxeOYFWukkdqg+mvoSkdpkVBWio5rPW
ZmFocWTbZFDWwKMycjbtGAdqO7FKOV3JWoFBv92mgWUXK5jVr9ogZ45ID17MB9tO
57ByKrzqvoiGmzKKCPE7OAxC6t3HGW1g45WLduOsst2Nd2NKbG/Z1H9rGjk7eXxg
YbquuaGyE0OXQ25MVzf7/nFN3gvEI0sJyKuHyG7tivVh0Mht6Fo51Aqm9KcE65yt
i+Y6N4OJHiPR5iK1OcBrFh9BSh298ei0axXUsF81aTZmypvG8ysWMwPeIGD6FPZy
0SbnK5tY6oFxO0V6zimvtBzIKgBtF0e/HPLl6fYaer4saDy8q9c6y3bzR4Q6B0+h
vjOzm/ycWta7RP4HI52ImvpIZABTjfaprj06o+hSRCCMBe4rCqt9cog1AVnvcUX2
Czvvbe76IOlvHJbqcZo61ZMwzCyiX1uRYJRuucF1LhCZ3E++RyNcTodU5lggOg4d
QTF++V5p/saJGCFVi9kXvw5sPh2M0p3boy/IdKZgZcVfC/KVFTGiwKBAhhzmTRk1
HuymKNRJBn/f8xpN7/+wvpnc1i2gUUBwHDSHF1SBs07m7JGhL1tXJW0QtMqIpHoO
uhrZ96DB69QaNe3eTZ17EULJ3uAjLozWZjxE2QKAQR1SCW2Myy+UijKBInPHpDgH
4YbP/7cBbBuyIYQXbat6hK4CVJvlihzDhHq75Mz6OmZNPWUyVxfVbM3mEyQuwUYV
DXFhakSiyIaXRM0gfmcd+mFrb3DkUGfgNTIOL3oHucsblN1bXCYf3yEW7lmCTG4U
dD5aRfAU0BUfSYUiyTNolGQAWhxsT1WtHco0SpB34T4nN2gwFEZe/fPAwz9gNA4f
GlKxcNrNzL2QBzkZsWBq14lgoQfqTTMwfLRWlJBtHjk28YUfktN42LjaE0sKv1WG
d5pbK6stas/OMaLuzSpQzNo498Ja5sSHjYx/3ucgfCLMZR+gULEiH/INNUhJt21p
ZxGrexwrJL3WSoPUzsNJRxK14M8556Ee76DRwne69eTIm8eC27JVziyhkSaWweIW
qyp11xaTJ7ClOW/FPUvKWxpxUodKWEGbL4jzgQevLHzF3XDgmQcvZkS5Hm1vEkPO
skwV9JYv6YH/jHG9ukMvH1rR/OrhQ8XUQkKQ2eqwpaQNyzbX/TsaPItAnnrPo9CJ
A5VtxXYXDYVzIw6xdFYVKQvEkvK4DHcbxdwDpQxkTo4uAzH7+z7hJV2Jxv/pLbdP
KNzZ6tXPHCH/1cvClbrb+bBxu2fvPOsHyY7YPuTPj9jphlooDfO08qkRnn55rmxx
Z/jq7/b6xiCnR8rSP2QJzoJJyJFjNNGFi/BHuYbK5tFVgpEa1fb2rIadanBcU41e
Wn2WIXsD8v+gAJI+h2swozmvbp6BnLES/Wf6bdJac92moFXuAbseqmBM7heV/HeV
NC51lICRZOv0UAKt1eERB1dk8k1LkQ+7kvR0zY1gk1g5EtqMjLT+gvV4cRyePkbD
HycWuVfvsZgl7l0dgMYdk+zQmF/qPNPxWRASf3TJnRqkpCyvlgiB6qg6ibt6Hw+a
hFIsgRWgKmQvOdltUDLEE/bLmD2H2/s8IgUDZlQwSXv8UERZIDw6syX48DzY+bi2
oVZSl25QQDiPWCYYQJafkQ71RDSrBkTacdPe6Z25cFqOdkAyhfqCMbMAmztjrgIA
+9yyAszgP2gHTlLcSsR4iOel5DzvSM8z5J/oVJqAkS58rpku2/KQXXpcZ6RL0/2W
e79UlPooI6Ws3CnbXZeQpHLomAhBobSvoRPxlmL1zj2ZVme995ZWgnAZ5GJkquXF
wqT98n0NHTt1cUcy+sQ9+ugIDuX9edVfsWhdvOabIbCIFxjpdJt7xhba/1TYiJML
1AWD1F19HQDaaLIIDzQ9XNgeI0WAEtpvtDnwAxeFPCzoN5PxDmjo4eH79nFyNCvL
6wSKQwAwTCtju2AWjJ9VLiPxqdRElDB3lqrKpEAtH4otk/OI6VyqQL/sxrNn0QTo
cnG4+KzqE4ipV9b+FDlh815XjuZQQN66GzwNoaGNjShHwIdMEAnNURsL3NXIt3F3
3glVZsnSJgDwsjuyPSf0lpCqXrOUST6IW5bRFGyU5IqxZWMmoB9K5HXfHns+cwoz
HEsSAQ7FLbv6r8YsuX2Dg5iL1B9jCbIcLPGhBRuXRamoUFC3gBYwlREcntq+AqKq
DdmYkCAAnY4xq8xh33fpQaMi4f/QXzVWbNa5/Wr4a6EcdSR4hrWweLY9VSAFw0/B
7ccpRyeVhujXIjTSUi0+v/U7B4ndi1JZKrAGExO4cP7jVS6aPirMZ7OkrGTpus0j
imdiw93Rcq1hcpDZMWoesYWXzy2p7HBZzoFdSfYS507J4mQ/qsshH9pPCnCtDhVY
Xq3VqAHY+9xZNhsRkLQJop5KvaFKP/mcErObC9g/iPqJwGgTg4VpOYv6QcR3mIAs
FcQmDNcVrMgYG8q9lvqoB3McSjz/n4meowc436bdCNjR3bDVyJdMRiTpL8Eq4O6s
gXi232CjFrvcpYTCffIzjbD5NeF7nKHo97vcMUZMILXKTA1dWC97EoSinjyMu53D
b3SF4OBRt5VDDITdpzefKzIrKHj+LJm+OIvf+MrZvK7UVkibJuvTirLICg29ZIMp
ieqV3hJMrwh7zvpyxLNvOWxcfZV85zrhUK9EdUI+MB8Kb+JPqYeS/29mCXhnVjiq
990tXmk3QN2I49J8fgHjSpAjuH9umjx3tmtVc7eYIuvGmRDIOExYTz0vyS0OsDR7
BR78U0+3xsDJcybwIXr3R49qpa/EY0FXF4WIG7zfRi/xqPGIgmzx98KMuuxIu7iw
1LHsrbNyDCNGVeuCXuywZA==
--pragma protect end_data_block
--pragma protect digest_block
Q/ojGW0xyK9awVjtTkrlSJ72v+Q=
--pragma protect end_digest_block
--pragma protect end_protected
