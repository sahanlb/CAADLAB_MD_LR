-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
oiX1mKxW98Q4If4geBAt/dFaylzw3Pf3GSBBddY0f/ui4Eam8jGDmhPcglyLyHHE
5x784TYL59W+RRLto+TGfDaXV/jT2cd0NdlSWbFKuAoybn8qXG1ulh7mTxsNZAbp
oYOi8wKdB20dXWsYoaRHMfIOOYSFI8TYvH0BFr9Ez2xVIVWq8nEv7A==
--pragma protect end_key_block
--pragma protect digest_block
EvwFnX+jZO43iUnV0luJ2L9xnFA=
--pragma protect end_digest_block
--pragma protect data_block
yfb0cc8UEW7G9U35gPNce+HZef2q24aZyM8nsrCjBd+fp2w8NWL8aB2NxBExY1Gj
yzROWrPgo7FrMNftHN2yv6k2VcD7G1fDkcpNae4cShjyl5wZH+vrz6cn4mFkSzJo
XbqTecUD2jVmIS1TP+fdBsBO7a6bL601w4OHwTOHgXPGMIlwmWeDx1otmqnZLlQZ
E2PcekTzMwr8E0K34yzGSByHlVV9ZZkcFCTSku0pI4RYSzYrCf3w4+VABj8UpFWJ
W1wD8OuUmfC7GrlXOcE0RoqC2UjQ7A1GRbzaEmXarfVBjfQGqrgwoKy3qANoaqRw
nDk9y22aU+UNl6oD/s6dDmkzcCt5hw2b8OjAgEnW66DV9NJ6RixltCEvK5Ucwf2U
SOhK3q0lHl29Mn5VI9aZNMpe5gM+kgMzVPWiPSAFYxHta6+Rdbba+BtB6QptISzC
ynVBr5WNQzVFlqDLx2dxF2Z5RKGHstRUwyUbGmbtKoLCoRxRYX5gUayJBerKT4lI
aW1IvfD+uBu/O27f0mWo4B6rj15PCOuulk4p5cpQku/C3Xt08DG2NU6cGTmgM97f
UbPkUTm5WyWBQi12xtXw45MWyHBoNON3msRCzM+PXbSLw3cWGvXCYIJUBXPzyQ7c
twyqDA3ov2nByLRXC9ZKX/JwHSl7FC8sD9Fn6tITpue9tt3WfwYc8BwcQhr4Bk2g
1K92Kc9fcZZ5XahmeDoXAwUKFlFPDQcKzHKvI7UwIB7LEqMYRMS6UEVr6mDf4f6n
OP3oTWQ0gM9R2HhdceN+IaRfRPIptYI34P8LiXyxJKIK1Oa+qHnUgUjyMaQfOYyc
vnU+QIZtooveHkSm3zaCc4J5JcZzLU9PF8XT82bLhUXkEvbWqhkj1Vv3uJ7Y6XHW
XY3wX+rFSUSTrHXLxaIm36ukKWXL/Nx9c0r1L3OnGnEGTggcA64ZyvPCXIBnyViN
nb7C+fuU6rEQnMOzlUtcEuIH72M/1PQSpnKIWQKPjhsl4Crd+Y0dFZzl4V7fO/Ig
mwReJsKPGlSpkyWHIz7U4w+CR+h9tzKYbXkgKxmsZVDcGh4mjNs1F5+mII/+FBtd
Y4oJbB/DEWh0uyGwFkopWlmGVGL2WYvC8Pscw07zTXYEg8Kz0f4wC8nr8FRyXgk6
c/QY0RzE/u4CyLBwf8M/YsEFbDG1u7vAwbmKHjqWzqlBAhiICt9UafBSGymeAQLV
EA/+Nfv0XptFIUKvShJH3Rm+r2n50gee3Muhn2u0QIMhOSn0bsY7AHcqgepAMTMD
XeFRdkksdWFJa2nHmoSQR/aXdU99XqT6Kc7qdYLMGVn1PNukXtxmT3tmY71LXEYr
8HetqPf9ZCfuNzMMlJN2fZxg/BzMaymNxcxpuDR5URqNUAUxKgI7CxsG0teQhA3S
D4+RVljZJzBFqAQ8PoE9IDTZuQJGHJMaAouLjb6OZSaBBZrEulHMmVqdRaY82ZNQ
ePQN3wY+xkc24MW8SjD3gyOYtQyG63FHvhcNZ+ltJ7g+5n6XgKxlMpGiJFDwDTFU
Kf4ye2XPFYsvrJIAR4sfAG/0h5kPISfgVgYa/7oKU2FN2E6OI5SJ3RiLrY5sN5cn
OJVdDwTt3J1e2cOb+8oP3nkjfviIqLKxluaEsCfRgyJ4fMdmcT+LAcfF5F/kgMpu
MYp5dC2hT4p2VRqscaelzocld2KBjatxfWAXt1wnUSiKcgsbmfkGGZcrR6FGy2jN
ew5Wlsf3YncLCrNpUtz3qffw3hcN1upAyidG+ToiOFyJF7nyLp1rmbiEH9aMYtbc
UvkGmpRwbPKA4X9DBHrU3R3o6saE9/YWaz1+k5M7JAFQ3Mc7XZ592Dhs027/KXzV
pc6TjdJnjyy5Rn8wO7xyfy+wOl73lR8Pbq3qXGgF6aWUfIf9ROwP93hshQEEO56P
9rT48XREGW39KUnb1SljkgBNhSjLXPgavbdZC/SJSMmcCz8rMV/aoY0BL2wCbi1a
VBjrZJ+7gSB84qxA1+B2sMjX/q7np8p5TmanpQLzPqx8HKLwi5j2T/ud6yBD5doG
+J72lVfjeNb2f9zEnjjXTZxpTMKVmZRsangtNKkD7aSmJ8BNIEIefTxWusi0rkUz
s5yIDU8l5pfFg/9qAIEJqXKos84atEiSgYN/hbyfeZcWos9dUI0rziBKHwlZkBJP
6vaKWEZaadkapcZmFe2eCuIBEVl/DiQyqc1W1Fv9Rxne5h6MH/azdQqZETBwawpi
SWwxZvoB65VdIzYIunNFXpDz+NMTjL6cgkteCbCjUltCLL5WCKVqpztpJhEEpmVv
yStXy6Rm1dv0dIr7I2/to11FRa9Hs4xJKBa0qmPOXKMGBfRXa5Ramv6vF+GrYOE0
JJD7ssR9lW8K23Ga2/DOpfehJ8t4qXW9WQ8BkyWJnSLXPvdunomCZtiLGk2p6Snt
HDL3OgBPTDw2QzSXqiQq4Jr2E5SbS3EgbTATr/P0z3WsAbz0hy2MIxmd05MVX8nk
jBEvFcvmOM3XwI5nJmvupM5nLhpSzaLdFIc4WEBVozQt8s1aIbV4dweupbNjvp8E
ltCC9s7qJ6q/iJEjIGJ2H4xM7PoggiMqItf7aPrg+qYZDO3Cw3HlUG+K+xtuGvU5
H3MSJucOoslQEf8Dpkm+QW+V6S4tBPgXeNZ/fAV4kYNXJluvjWzzdiPsBLT9OHNg
r4aJKwAGojnQBm4xXtW2MiVJ4cMQ0Xoub55AMkcMNMdrYgXqC0tWb6cwM1RGb37V
GfPfU70XhR59TAaaOO1pyvQtOx0ukouddFa3oSDQHDijNNqKurbNt+n2ue5eX+09
IzHnJ9prEbDa6Pp3wbQd6y0j0e6sWFv1/X0fkybGP4r8NsEn4SsXrl8o6l1e1O1t
Dv/flK3sAv7+TcrnJLngbD7NyroL5bVuQZ3fNPsPpnWHJTJecoBaftudwplMwvyo
05+nMBqxN67QpsjW69qvGpOoAEtv1SaxG9Ym0pwx6C2m/QWW41l0wdQqVTTL1EAj
gIIKx+UW3hTKghmGQuDlW0gORdAT2CO5C6gpfDPROR4Quq5FXMApvu0nTk+Bjj4O
dhzNRtK2Sqw+u7xiKfZDbhvpxIYTsbWUpFLNn7mkyFKKk2lKqHJQcKIksXbRVnE5
7FX5pJKyO80SFrB5ldTZDvqt0fLQoYz6dC71W/BJ2N43zND0Cbex/AO2kobEwbQW
LVjcKWKxIFdiXmerbKuCc900ZWZhqW2KaiNHIJN2p0BJXGOaWCfuEc1b4roYowan
+Z/bzZGaFeFXZO4NFxCnI0FW0e/z+QLR1H33gItCmUzAxc2uTQqndpbd0nn0uWoB
3kneFJnzl6lVRBbVbmPjaB3HpmTVqxqU5YyT547aCwy1Jg38gheTKAHK+wFrrURM
vcVPi8sot8YARbItLD/4tX5NWFBb4/TdgDChsTS7IAIt83DVjb/Fw8aXMzxg6QRc
l2CXxgGuVuoXZMLadnk3HfNZgroLeaJtvx68G9At7M8zR6PN0zaS5Mot+DT+neU/
Xo5wxWbcItzsMRtmYpAdA7/2BNxns1LnlPFm0twd4xqw7gJSEK/ZNwtZNX83LnCA
5Pmxs26xqj34SU3TD5HG/LOA+vS3wUb9cJXP1sQfOD5dQR9On1cVfEjg+VVzw4oU
aerB+eZkYd+Uto3VtnGCir+DixUJdHakZk8U/G94XL7s3yxcRbcW6RSsdCztd55j
Wt9Eu/OF88BFA3XRSs8b1E8sUFey74z7QdHXOSVvttmU0t3+zOpDHHrjUt5wNK/W
HGpxP/GdASVqb8/Nw8PZXH4YQax3b5X6td9646yJmAKsjKpxN8Cpf9tzaDB2H/En
JnrSPtsNpZ64uUBRQpg6QaUdrFkLL5lZrkT9xKdLr8D7p/gbg8Dh64hCIEN1+XWq
j9QtUMFL519pnpJmSQdVFBjPzzIkDYnAVZBXNo33FSg+qBiQTV555M569R7LPeNG
Mmpw/AxpLsQt5QjOBbhhGZykJQXgmIDYLV/gZwhk2Rfp8m1CEx+7UmiRRkmQ8qvX
bkg65oPsKcvFcYZGSgzXvAPWdDYpCIxor8NXoMXEnw3Ewr2bfiyZAAwZN6s+UmYb
IuEfU0IgOwjGTqOpMCFrkHv4doyXUvFIjM89qpXgGNjG1QsY35QTARozLPbCgq85
PhbofkZLDD7h4Eqs7kn/he+Hlk7MkpYR3e6c0WCWSbfPhlfzHRFg0Z07TTbyEZPo
KXciRMB3gyiHabNPF3KH+abCKZBRv8bSX79X/3nK4mayJ7PPNrarn5hyiwEiWGw7
t6zSmjjxy4QYrmrySk6ribvitn+ijX2UCQYhHmd5mAwZvLQ40GKNGnIjOFARdQnt
8Q1V6f6ETi9dGM5xQIUwlZ2hmD85Uiv3Cf9dH/GoKucJM0GscK9yypv5mbOrpVed
NVobMgGQSmrp5gyoUV/7MsSPY1z4J1j3NrodNbgeT4igAlqKHtIcURHst1Ou42wg
zvzuM7VEs3pqcNkIQVYQjM4Tc2l91YB4bE5nqLy/vrnVgUMswajKM3EYAoN69Vrf
4c4Xc/Skw7PLDuVzk4f9NV3k8FLfJ0HIkUD7Rg0xYpfB39u5b486uVbPexRcyZjM
C1zUZ17SUAmLuWSjQClq2B1xY5x79sQ7mtkB/Eg5MW5d1RhJclh3AK2il56Gmok0
MNBnXy51813G+8OkWyv35K6sr7aGxQmVZENOh894d/GSWB7n3kNRyMTTb6yl8+EN
Xtikjarjq/opw0F3FVl5z4AD0flps7HzN8PQupt9eSp8M3sZj8Sh+ZB7o+hh13TE
gfDCD2pnGziDEnTgkdYS18saR81wQVcuVcmn/0tVR4fIAb0Sx90S2TmJOiZD/OX6
HnQ6UE30MnJI0y96TR3oAXOZlxs2BLbzcb71UtjQa+DYbSY2rWWIItAtquMv4e/d
1I2rdwwbioNJJIUjmWB4GkCcebG7FFSqiTXMpixT2K4I7oqdc1Qt4WEOArxpGwMX
ucYTddKM3FdPLztAL8VwDb3J4PvG3ZfJlusdQEA3aJaaHgBP6A/7acg6T3D8zcH8
Y8dtRAz90RiQECMdpfts0pe8fVtmt7OyQfPgTKlN1isKL+JYnXqp8BsRojn6C2Zw
fLC6hBdoYbb3yOtA3QjY237E4CcJkXWIEzZH3Wz40qErsvcD2maW18DzLRL3XPuV
nDQJEiAYVKOJzkTklTxe/cF6n5ayNT3TuwpFZr6ptTO8PPvlpZ3OlCW9/cx6y1YO
ItY1DkcfpKKFxxvCunpLyos5t8sCvrM5pbuyNSvhYh7p7bacrGqGVZ1pMgxQ4zwK
3uhMF6snEmGdHJqdKeMLgeYTktEyhIyvmAh4kLHUKlWONeK4aOhyuqPUbXyDv+LK
d5Xu+PqnLi8j2Wv3XuuqcDxS0wQL0KBQCqMoMEt9AanHH0K2ofUA/iLuV7erkpp1
0Odal/rinzLbgM9t+eMMBX86iLUPc1knKYqah20wpUltQVtHjkV2rBqhTED0zZgz
e4NIpo+e723wmOe5/ZPw91R4GDzavfTSBPu85yxeRx83B8rGrEXpyeYumRj8299H
H7EjuMw+nFnK3Zp2S2Us5YgKpS2YQjYcqkNp2z02zX4RUODxahRw8P8mxSpRDIjs
0COTtJCEzuSjoitF90QD6btnwecT1/b8ci/teqiyJ0wGRaVsb0S+sz/j3eZPWVN4
HVL7oQzAcRvu09fcc5MpFtfKkW6USapdRM43UBnxFXTJBElgEMeiFzgInL4ha9td
ST0Ns6IK4jglMPo4YtBnDdL6i0Db4LBjJddntkG/rjxgKQ0rs3RIRujypRZQYAW+
A9gSU7A+wNBUg/3F0iRD5JRlLd7P2+E4jRpIefZZBz3HerqYc0Y6u7bqAuGOfOjw
YLl+uFSC2A3YkNSzquGiFtM+Xd38LBVeeC879wViOpcV1/Bw5iKGEKzGnPnXLP5z
hKgR9MAK2BV7XgYfpbmZvXxfYrxFiuGLwmMtrvNFss6LW7NmysHeEmh2YNBSbfVV
1cbT3c39m+aBo/JV7680mW3Hjyo+Hvqb+pTpGxDoiu0DqkciCojoEHLhASXMPKTh
T7PKkA6wNfJ6y5CrhSBwPvwYc4zqGinHoIdNMcaoC1FGCcUtlu1BIrRQqljuY1YB
ZIC7KH4I425qTSjPz/AzzLWCP2PgUHsqD5Kaxw3qzjq4zCfwRXOe8d799lsLF3QF
fCgTA1tFcbyYCYx4l7oxHhTXL2UcnX2d8+CGzwjS68VLyA5YldJl8OJhJN3ZO8Ya
jSWonC4T6e39mAV8yQtfpjXe/F8FPLFLg9bbTvyGJRuCpD04rS6nkdFrPItLOszl
CMMuNw+gQCTy5k7JNVXZTP9TFMLddLDclLfpEPNxRyrl2MIwS4ZXhiUb627BBF2M
m66rCq8os1ZVaZR9xlXfarat12QD/zNL25ndffw/hfhDwT5RKp8rnc8WFvOTzbPt
zcESvvTRPr7tiPX9KlgI2jsZtW7WO+T0PBrcGXG6kk91G8w5UYzvdJ/WQ1V5Fot1
lk0wdL4F/XkTsvvZa1dFUzs3NmxMwDXab+wO3it10bLvRzp1Lhwuv0FhlS8DaAoZ
nA6Y48OLZN5hmIQ+xR4GXiYir2JjHSsmH0bynL54dIJpmYkfhZj+i6zvOiJOX8eP
0K7iZULPW78OfbEGiDCChrG0FsmAgMdqbUL3yi6RBeUUuw0ZMv27dP64f1QyURwg
M0+2iCQaVUcV+N+NlllLhzOhISLNJSwOd8RW+H4IDeNTrJqb69UzfzDWL5DylZMa
y009R0aiF0PuT9hYn+L+P4EvTa/62eSxur4g/1nVM8v7TV/uQNn0B9z41G98IszD
wpt8Gn9yZwPe2yTae1naHvkLff4Vkifco5Ata4QIsbXpndaE9lMM0v1jq5Xx77y8
2sYMnRXcHHJQoq0CjjIzqKfKjBM3jXkArp3hAVqWPHCODNL1wp2TX08HDHwFRDQx
7Ar3vQdgDKeniQA3jzzFoXfCpKNUmNLYGbEyWnMUvTe3SvSx4sVR8roxwsPX4kdI
Yj2c31Co3SknY1/FsPASGk4dzxafX0vrmcQnQB/3NQrFcmj9hZc8H4gpfd7+1DdA
a9XnSSQwCg7cKnJjmiUHx8FBt+XLDGI5pKElIF31O5POCxg6Nr9vpQIhXOESJuKt
sTpmUYLduxjmpyiVVbtkLRoXNHpkDEPTgwNp/JekNkLSHBIqPrBKDL6HzysTNUQF
BjWINTlhXyjZy53Ds7Q1V3zIuwR94imG09surjRhKf+AWtJHv3pma/ixXw7ZG/ua
inqDzEBTkqZ9oO+on8ngO+xs0A4MqcUS2lEcoIaJlXHX/7fvMwwRzZhhhB1Dcb+f
s+i48CvongyB7GUeIwhMsySgVDCgAvmIvc7/+FGkxNfmKK0DpbQPhzzdJj6vHhMb
MecQvCm2yDbznzEK4FfxvqV4DRujk0+CElzqOLX6cDxdoxhwe9ggwxxtT+dy401t
nHEe09djzQb5gM6PE75YEnJ6rpBihT8awOoQQPIKI0Hm6Z/UgSTddkCfjt+WnW/L
axBa8tf3eJaXw72VRJv5XpTiH8SiGIxFnen2TQ7i99a0rhtI1nB7Mx/kE84o1O9E
aNKNKUlul+tMHPS2/NCaQwb1KyU/4OreKGg5maZt3Djidrmftlm1MqHQCUPOeruo
0j8leuYA9wAXR6iLAUGhY0d1Z6LFgVcS5A8GscMr/BhLXco8mkBSiH19kwt8zOFY
UXKMNATeyb5fcLp2usALy1adXCUhAB3b/7PaL/ZT9Y+bRWeRQaLboQBm3E5RJo56
rfw6OIIqW4pEBMI3IBaZl08pID7StTwNTNfbplaxwk+kLCPOU+EZroK/iLozZuyj
SIfUKTpf504ypal4mpZWFSPYsL+h7/eURR7mVCag/TWGMin/gkKlXIxmm2jwSHKM
iM9xAcnb4z8vGeFnKJhxrGLkUzppGJYpazum6c/osst88zNqwdwRmt43lmCvNhDB
LGINtcXUsmxJZjjj/zf0avTP3I20sNpWdhXLlOcBTFyJ/E4V4KiQlHW1Ac/15Uy3
HqtaBbJ4WIjjsQGvMFrwHwC+WYmQKib5lknUH5+4ff6c9YLFO0vAfpaw6I0WBmdD
PZ6YIVJXxZfASugxfr4v06L+Ybckm5UonMvMz6cmbKhXRjxoJ+9SUGf0TLlP4UDd
HrF39KdsIXgKVeuvKfMfOIQiuCp/dxUdLsg8y22xYHhoiAFf1djUKnjqre3qI/fM
37CwgYFXt0T04g0UfQm9ee0hkQ0rtlsryAZAsP6hC+jmvPlwGeRxIQzIbJzm6qCB
JZqi/vdUnh9f9pW3tqsnvo+BjpLLoJr01HXS4TDG/IYhrs+T1H+naCTyx6xIC6cP
+ovDGHoBxDV/VRs0Su0VHbFJW0+Km/Ro3xl9N27hDcwDZOnoCJFeZqO0Cj36RZmY
wZ9xJHz3xLPB6iIK4gjnhGQ2PRpmYUcrpeH9liQ0AmczRYYEu38l0bbgkRmDGlmh
kvkGj90way2S/x8t4lDV0XxGXv0ghp8lO7kCYhLWs6JuDQvIq98fED4qSEPLUmSl
TnC905vSegPzuGMR+2E1mFvopMh5XReBT7IPZflM8A4/REmm1QpdEhjCw3oJ8pcw
OsRiLBovBXFXuSbSET/EU8kmTXDpTtv9HXoEEFZ+GO6lyqkRyzTUSQ5TI6j9WuLS
xYFeSdyjI/5mWvkJqiHJ4C2MN3S4j+wqzXKCH1imZTe6o0mZK5cJTq8NJnKJZC6A
GEi0ruvYhOPpRgdCwYAsr2kiCVxe5x8uADP889fvckMYLN4E+Xv7n1BHxYmuFQ91
CKGXeA93nDr9mW/FR9Q8C+AyVv0vOWF/oI4v0yVZ4o7JwVSLfZE/+wJLgDlbIdBu
+u4FG13zeRetKFRUZtedHGeeKupfIlIzwuWKCj0i4qWEFx5E0RYoaVGBr/neu8ay
XmWZ+LfO/gGEQoEN2dz5lD4G4+GHMw+WxQiM1bveB0fbCDERDsSTVbbssYifBrD6
r+xCrw0VwGeTU8/kuljUmP4S1URF7LSqo4sCJ7JsMyA1YaT9z/b+UIw3/dgX0o9j
ktDkiWhZ992DzOVd/K8ZzPUihc5dQMuvSwhuAG+L9bSpe84Cz4fRuUxzTYsYl7IM
I5hDVzIfg8uWqmgID4KUJ5v1x7DJ/65pZQMhHBsQ3t+LEBIPYaEvQMNtKU+ETN8L
rUCgHsAWLvXznq4IIuUG0cJmJGDHLfA9+u0ZiVR2afeEg8RTm9w/5480oqQXYr2l
3jiHfC7VRHsG4qICYkuTudQE7Wh1hgtJYUv+M5wJVxJD2nY+BLkiRCL7Tfm5LMVT
IEDQijz8byAr/uJ6zmvyrb+8UJZIw0El3wyDJWfUgx6Wm6cUw9+beKKWRo/MkOrh
S1aWcLE3myAHP2SkeLYsWTIfCfO8I8jnKh1oV5WMFdW+NVegC3iM9BYNuMgNykv1
DqKWy165tO6AvbxywMfK01sY0euWwgHuA8SGvgNB0tgeN+uQJTgqh0dpAd+FtnCb
mczPmJjudJGROqLjJzLQQ3IAyQcxq5soltGWgG5rH08142gSCdajxxmFRzJEogQ2
tvVwl+gV7ALFNzWQTYsQp8LBcUznIQk8P9viBN5DymXlJ+2AZrBkG1M7Pqxlsstz
Hs2ltQZXW8nnaS57oSYYewOcNtc9sGNTySOGgQ2C/CzU6hOoqwkQ2/6fvE6atmE1
wJIA0thB1QV/VYnANGeeEsZc0C4Xd7529CVGOKJHk3gWE/a1Idx7DO2pwRz7p4w1
rYJT47r/pRrdfl+Qlm8M8366nkxx9l+ma3SYRVfIgIYS0NyNhGXt+MT+u4SRTsPe
Yg3bRaVHaRD85fTGGSMm+RK6z7E7uY9njZsS1+3ZV71fpCw3T/slJp5geEWkGet1
/V8+XANj4dJmJocCQTdermdWwvbZt7Cz+Xo9VVarT2CkTuiFwKYalqKiSWduBfj0
LMFYMmq38dDeSoTIv+lzRPeneURuMOOsLqCvnM4PPTDo9A6v5mVDLmH2Uedg4GMA
H+dam5fpZWqkr7igwpV1qvbhjUZ79uJzkYgC8jixMRtd9XUyp+k4qmJgWtmef8Rx
zEN83kXTLZwn+ttezOYskpkoLOW3TOAXU7UEho7Ti3QFcK+q0fR4rTw7YHRlPTwz
rPdDD4J6TlBS2giiEMs8fP3pO+BWlucF3UIFGAUqXgkdSyUOcLAhoCrt4igSXR5d
xOHqjJxskd+1QbUsR83V5Lkj7jAlZVYWylkLFyS9B5ofa21QDqjmxin4LLiarhWL
K9WoQWOciLvfrHvSUffxaHX2+HJa1bwxYWy/uszDqYziAXq7/E3yi6XYG8zTQeZ/
jSy2l09Z3XB0O8pJDed+mW/HiZFmvj8xCYUY74xOlfaamaP/OS3WfBa8p6PyQzb0
VOtgJH3yMnIVHtRUJ9qMvR+b+XxU42fW6qn7x1rn73/4E1ZLt4zg7lRN+h53aNFR
yyO/N2TbX398myojnVTsQRf1vu7L5LjatP0oKNqXsX7uY6skqQ3sRjvn/1nPPl88
xGRrjiTUzaigk2MY6jYkNix+KCHLKBiNLl+NmLzgOPvq7WfFHrc1BO3oVxv9OwoQ
8O+hlzAEiGcEFZAtFhD8FyMJCbkFDbb6Lsh94UfhGulrT3SBaYQVUimCzRH6dVYo
17eR+lnJ+eR0xh43Vvs1X3km7ospj3+MKdjCPd5aWJKRBsn6nhCXZ50RG3QJepVb
bFJfrzYwNUl4LynqhCRSaMRgjGFO6a1fNZC/3eNEQCLoDwz614OMMiOnQDk6J3kG
dG6Xabc1uTbf/fpmyNMGRbyJOYB7bA2v2m6ErUgOA1lmaTz+MICwx7vHfCBql8YX
IUJ4pGsCmjnb+7tk9poiB3oYH7mT7vOi0MTrj439P10+TPmVxe0PnQtZIgi7UwEV
hIlZaaCSwR3/I6ri+BH3Sm+1+qml7FF7uUQ0B54RGiaw88q5ihuueHClWhhn8xRY
xwP6RMn8LHYvgo5C1W4vLoYACGxq6hnCNc51z1Oaf5wbPiv9Zv4GkW0IFt8813a5
7EMDpGyAPWfvIUFANEqI7l6bEfYLJwuAZw5JxCT+ZHM5WNBQbWTVMlGWf6P9ZCvG
CBs88AX3dZ39UK0/LOLHODyZh1TQ0fP0B6ksN2Q3wnQMiXsc8pLSpEN5yqtMjghV
ZiLkv7kJYArTqpdl0rler42eASjozLGhF0fle2k+D24vSnM3L9ef3fTk5V6VaU6y
P0AsQh2Ykb5nMEmeZFZYzjbNtl6dfkE6kPYrEwRnwNutbPd/T5XW2iErbXzlHutB
85826uO3OIQyqSolVoxKF5LVKYvPRNkkSvjW17djw7ZN8ByJXT8oCs9NSlUjOPfv
/Ta8OJ9F81/B4tQMlUOkgidA27ScjOR6ip1uTFxUjdQe6kFJXSoDoMZZPCsQ/OM9
xvG5eCaP9KXu6JOAy92ItF1VWQj5aINxOU3KGDzn1CEugYXmMz9dOs8oPqF73CUh
tAAxU7xJ/f8N14ga1vND+9FYJsN7HY55E3EPNXhzJS9faEIvL9egno4juxEjOzCr
ZBwQq3qirMmLumxbTa6P55w0pTUvlhnxtkKOr0cVmNEmhOKX9Wv0MvcLzLAq/w4T
LzRkY+5dvxmea4/7VrciN+6pqTaMH6UUcYFPjl4bFf+qXRnmWEfgU1QAwMNXopKq
s+4UezbeurFS6ta+r/lO6ujM5ONMQjKwVki/87F1c7zCKlZqydXgpFIoVKJkKrz7
BOc193zEuMLbINIQtJzzqRJHTvhwgNmEFDg37J56IK3DVl27DA5+ZVddz5semXYV
OL7y6TPezPAQ+bNNd/FfhbobFmyMaZN8kmRYZyAQyTtlcciWSoZINxn3SOfI9OPE
PlTC9XsVO1wBA4QQH/2Kr5FhNbCPPECjKDa/TaPTY42onyHviVIzn/ohPjQM/Hkq
xEGU9/I4MTzJ/UxgX/BqWmrtDa2XtFLPAQedO2Ezl1zzxcydB7SP1hg6G0FfVsDJ
PQYCEf+fQeGlUsf/6IC6wvJ9+Lxrct2QtxnV6Y4fdQ6SqAHiuKSLoJcsI5nVH0uy
rxU89M3EZd9q9HriwTX2nI+kK3C798YbPcTGfJ216+50cYY1+skIFytEXcNZiMi8
CScuFEy9ib9GxxOwtB6dRJ+LBq2ri3XFVbVyRtwFIGFNSfDrqWWhiwvwhsy4XEJ+
s+MdbkRMJYVs9/a/RTNWDk9PjZpsnJq7Mzbdam1kXLTPNG9e0d5mxHmJRwaPbYLl
CcPUNQxX1eHnKv4FM1do0bnvbEfjEsxL5c8/Bf32M1yn/KcFKzyx1OMw/cwZaNmM
jUTiAdNzMAWUELY/teilk5OqZRThJ4HAFzCcoWND7mMbhUHVUz3eceqa7gJur+Y5
jpXMA6KLjrYwClV5Xg8yl70NNSP/NdrykKOBwFfXZg+eIuwZ1qQ6vpBRNR93V8bk
QvhQI+e+5snu6mRDpEJS8GYZJWSmkMIG2NbVHbq7W1nFL4lxcOxkofchj8TM6+yf
loeGGFT7/e5qq63eOHjm4QnyEIcnEMfYPtdtTiVq+gY9A5LLVx4vuR5rscwjUMdk
9h+UCG0l+17NuSOVT0iEQFu3KQQkhYQYREUAeuyMNrDzMAVlq+9uMifNRB8o8je0
UZzM4bxhkQV0WCLCLE0YRzBF9J449gcI+yktnsL0LNWhZLj6OYLVOvAbja+EC11V
YDOUSlGrRl73FjYxt9n530vf0t3965OMbpW1tawxTq8U4ugTuOtNZ63ieyx9q8a9
QHfo8BAU4chPNZLu/zxlpphDFhImWNPkcA3IEDjukLkFW9ZOPO5QrjkRO82WKuaG
3thn/qnv7Y9ZQ81gDfIfevX0fUVN3fMc3UzUMwaqtX0cscYkiLSWsvkS4VkO+A8S
bZdPzAQxldjl9d0NWL8MD0wP4vxCq71FNEhYWlo7/oSjNsvx0dMtuH+zRHHRMgR6
bXHel5F8CTQGcJvATCN7Fqjvo9akNCasM1OXrb8lspzf9F2cbumgBSQGZ+/7iN88
QAjFT+nOaKsG0UroozXJH04T0iKEPqPdhg/LP/GNhcQWGd/rnFn2C8A3lofyAB9w
5VOqq+XrLuv2Rt7kO9Her3q4lWHHd29kjpI10yBIJ31fMabBCaJQDjg28X1aBz8R
tUjEVIljO5+tIT2Nuqu3OjrV825jHKD2aoJI+RpVJzXrblkin0+VIwOYOjQ7UxdU
y22i8W+7Ua5SyetKzmOizMzmfGyWiydASi/lzFnJWfrNACtF5jKgba61aHGlsWNW
XbahK4kvmOE0s0m0YFKATZZ6JDBOoclQfEdFZQICcCyCrx2n4l3gEnW3QvzAxDAJ
Q+cy4c36l1npdYP8TXJCLIAcPJM4nJRF7Ff7fxU6VwXZmBA6fzr/1kH//JgERH3c
IMbFPToQMDQZxfboEI6yqtZDBUY43BZviDd7omOVQLm1MJfCxmsOL3PKjvDICWvv
TXwvVlG1iue2OqwY5by3tsay9Eg2+bimH0SVEYdJ95T2JyquLHzZWPku3bBi/SUC
uzNhvtP1rvjRgGBKgMVP/hdIt1DZ3EkbhPYz77ZCOhHWtnP9BDAmboFZ28o45wy+
VfurQqjHPcZ6EuFvDQAnMd38U90S1GPFMKrMuv7M2FVIhMdaD0VC4kcZjMhk0k/C
VH9bwamuEZYUencDEf/vBZaUm1Tg8bxRZlF79xT/0tKUglbFgu6rfYqPmnamYO6f
I8q7BAWCH78fFkdX7JQRKYkyiDnFNlrxf9X1BMv5VSnPyt76CMVU7bFU5DwHTXIy
dh843apXxHBNcdVWsSFBOIMFMAjkXfq5aTKyP54qFTklJeUuGrVrtFO3ei6cNhKy
5PGJIefA53tbBvDb7EbsjiiIIvN1eWv0gzFGkzQP2xpGUtEOcOmr/dHFSpKbxj3j
jCTFR6ioC/XWaU/ET7uaLBXftlTSamfnTlWI1ObWcIVeZZsW7xEFXBI5XopnTIGZ
W1Xlva6/JOoLvi2YQ/wOdcIBlwF6lwcyVmBVbf0G4K+IGkLozgNOfvOue7NJBBTf
3XpQTAVkWgUGezvAFN2fZ+YqXwNZVqIh5O6LQRIq9Wv3KMsae8lOCU+EHD/S7ufM
jk9pGdCvbc/f6wCxCn/7ejKQntQBo0zUf74evvErhUBlc7WfOXBcc2MnMqmt9Oam
s7i/osahYLRZN7c2dyxh2DEl5I+vxUqkc5V3PzHXlVgaFM5S9cgvyzE6ZmoHM6/U
6Mqz3Pm6I0d8MDDk75AmBvPKQ7gRHUpT1vh+IK/8II3oov+u7jXHnHhMhGcOjtvF
KcQBwUoi+x4Xx/KkCPyJQUnhBT+afsvKB4rk6KcMP28eFUhxEbqaQk8Us1Iui64X
pMNqw9zAMbHy8tksKp0ophlzbkHHNfthq2K9C9pd8oKgziaW0C4EUEOyxEUyK8p/
C0cfwIOOSDN0hjRPjRvalMgM8UpHvt2NAieWBQZGlKbKo3iTudUaOt86o5PShbea
V9andVA18heaA1GWYFB8OWEs0B3iqOLUZOv9gJ8SWn1x11NUz/UKG0PsapKTDi0o
vNr9XjkCGFNidV6JDr2SMwwrT/D4XMm94CITpGF4bR2g6CeVW9AhWaQbRq7asy9l
GmCf6tVAvColIryJNL+AXsCHHqra+Q3UIDFI1BtMgezvP9rJeZBkPsHo/SUxG42k
DNKR4nzYEmvNQJfVu7b+GUv5T3BXGEofP+/T7YXYiRBc9pV3n92LBiRik+23yhh3
Bt2CGIiG1ObRIo/Km6YJZV6v0Z1iTGX7BRIe/4ISa+cltBP787MJOlcXeGz9E0Ow
J08z3G1W7w0W46bfDzyQ8gfGAVnH4bf8sQ5qalhE89uGyhF/Nokn0MLcdCAH6XgP
OnqhTKgmwaSulcaA//V/z3tIz/yewR6iqBOozbE41Qwj9zl6col50Vkvwpdqj3WL
Yn0OqO+Myez8WDpwJDLvjfzbW80TB9QCpe8CG8bTykhROPz3G/Hhp0+ySKLluafj
zPiyiZ0IZcM6AnsgVEwYag5Lm4c4+OCMONXnAd2huuFBVzV4FrfacWLDgHuRGz+4
12rGL20yJFSlgHaEJx3LRiF72UMvxL3UC/VBPbVfvmrmIxZs41/twZuRx9DiGmRC
IW+S9DipitP0L3gy6AC9WuS53CpA9pPztn3i4DEx5rJp5L4E8e/ibDHmS5i1vvIk
DY+sRio0aIJ24h4dVIylspYCHKr3PPVSz4IbsQjijucxXfA52uYoRKH1qbgTh95d
S2unaEpV1wfuTHe2MdHTAvI2QChMbQS74Ccfdum8YUS5h3V+59JSvV6rsOtoORrN
wBpFbrEzAB1rBkTBtchDBmTWAZ2hi6QpZoTu/s0ycxTXw0mg3U9fBuCcSKOwo+db
vv/GvcoZ7upRl+N967R/0NWecM0mmwWB2OUkeeww+hR8PpnJRQjEbyDndrXLV0Q2
pUJPHc92Roe+eIWXdGTgMi8CoH+6geWq3/MgtUqBy9zDT1y/7bSHHQFVzSj7SNDE
2P1Ly4FYDIzDxpdAHvbU/rijCwDjiKapo2IGDcjYjN8uIk/VvsL3jrWMyk+s0CjJ
Pcm+jWXJPduF6Wt7IxD8rgtPsiqibLnB95AqoP9JSP07FiwvjAiYsiuVFCZheXJn
grcQi7cwCtVv6fLCWKwI4pdrg3jVEtZSl6ROA8sycITrCyHGgr/cqINa8mWRrCym
NhLEfr8PXcYSxV+6Kqe+FqjKtWh4ebY5pG50qk7NjkMkPg8+AHTo3/pRYawCjxTY
h6vJvJrXmLugjvAMCu/BAZSHeudOAx+vamDe/pgEce8t1wqrTEI+EaVpzIVxewRy
P04obvIONUDLMc+SMpRTRME9eWoyDnlDlFc+Yy/YnE7G5Cnw3INb5VkCjHVdcMQX
Gd1hVXO35KRCqHtkYjNMIR5As3aHV8BebzLSU4DV6dzGv64e+ZMNUgwPmxy6xPCS
l4AMiSPO/7/1KcBpg40u5/lhS4wYOd0m6q2nKxyaqmsfDjwVYfkd6/8l7EErSYpj
5XlKYUxpzOc8GhaHm+zSfr7pxPncszr/UL4mtu8EOmQU7/umlMbLMSL/HCRfA6r7
AqulZHnhLjXZO9VatpN/pFLbmAE7DB9smNb7GcZpIzV36MuD9pTtgv2Y+SshCdcR
dmOwqdgwELdNFx9T4qhZ1ODahw2S9cTg115jWW2krzllVasooG7gWV+tHHmQfwWb
7j6YLyiuFbon+HFD0Ba+Qi1Bjpq9952Qjs7VESdWlDH3ZPpRYcynNeTMo5bJpMlJ
UxhK5dQKR6HC4vWdXG55QBECynAKCA/Zwlj9usJ9GsVXqkozJPCwNB/KU7jpn3As
kadD9nvj/Vi8vtOjYTQFY6GHrBgoY5xe3gtHarA7VYPnuwMlFuLw2jBLbwEKytlg
DtXjnMnYiAFYFNwwn/A+qIBu2VoIFR0heXrkITYJ4Ss4ZQgGnrxt/FHiSeD7HZ8o
BvfgpecxBgb9/VH3l3U3poQC+rRRVLSB+NhUqdC/g1MXjWqTJ3hN5Fu9AKUkcC5P
ji7TMtVGwVxl9mVeP67cFIGGZj+bLPOVpMilQv+xTi8A1tWRw3s+wcmIG/t5fAB7
DOoOFKL++Hs6ugx3ZrxqMcvz0jXZHMaOnyFZ4v9LciAQlG+SCOalnRwwc65ceCYf
uSQitRsEfetuV2PrvwgLAA2f3h5Yis2RGnWo1/Qnrbh9WrFVCiQDiR9zeeCca1f9
9w57cPSLAno/ZRB3hJJbBiOPRDlHpi/nlmeY1Y1j4F7SrdLv7UiBHFp8GckFcM7W
5hjFRWOcP5haBtayLLDlIuckrW7SgU95+d295VZ2KGEew9N79pQ57xZxRw0ffRTZ
EPTo99Nu3/3rlWXZvdYZmXiqeeDJd1zMIgUs7ZO7TdSt1CuJmcPQef9PiPM3pDrI
HfSKiiuAfBpbey+Hzo+0Bqqzy34RHWoMsPhHUF3OY856qcm5p1QBZUXaOATogBrN
ZATomvRxdorvOBOEwDmERjM02tiNDpSW/eDAX/DeFtU+h6tWBH3+Veeiolbdbf12
JOKDQHjcFDpw7uC6kc35YasUr0vMnHsG2pVArkWh09xUlZLtI2A3EIwgmOoBvL/9
e7ErfT50UOAUSyeeMCdXLuM20fIWxKVQvx5MuCFuqquxJtVQmTEX18LYp8swByyM
Djg1VDhb8RoahKkFUraGPoPGfGRxByK9JpMVT9ENMYfrvuzGL22yai+D1GC6YaaZ
a8BxgkjkxWAJOs0cvdR14uKyjBJXUEz4i7NNnG7y3+fvQMM2tdYlRyZDX2kK/qhV
siSIPE3U0yLo+dJf1Nw+nf+OwhfHc4a+KHgIXId8kiDFZJs/cIihaw8zfCOrmGmG
CRqjLZQ9Fzt7mQTJSmOltvZLoHTlpvK2Im1Fa5Pih10yMtGRl37aPY+g1sBu+14Y
oMEot/yai8zn9Gi6SI7mmhx1Ea7BRTgCu4HyCqYheBnwiEyR3dzTl2WrbD7xbVAz
WVVtUzrCe39VukMGI6JI6TZMEpvQV2vsk80WgRVPf0NvJa+kuZalkcQcH5HjCMJa
4vudk+4bD+cM9b3f9W6o58Gp0VKUZzLfZqeWL4V1/BAxuP4LuwUfwWnHVrXEfz7V
DJIO94BEswwK8UD2HQ2lCtGF+vlPUoF5C+hnGItCONfPlyqo0J8QkYrc6s9ADYme
COGzNeVnJLkzxbvWgjO36wPx7m9IC+VUCy6uXRa2rRJjC5GJCnXLlVBYDVn7+AHv
IgOf+HGulbAgFyCCXMwPSvkGDfUG968Z6sOqkXwDx59Lwihx4edOVemdiEBTjP3V
o8ksjJa7wFz6PcMu8rdkHikEmTvto9olmsJWn+NCJVxfHfLsj7S8f1WPOTw8thZz
xWkWoKA94YAbqETuFVeEnoD/cZuOYuex0cEoHmvJoWI37b3uZ1+wRAIP0LUuUCI3
sMwuOJOc/HdoNOQbZml4xSDwEpHrV8dQGur1AcrSqqAtwCQK+aMwt5CSvFQYYCfm
Wyxby3p6YnNhj2wV6ZZE8RrFngkdDWT4m5oaAdMBqHlHq1/8T3utszN1HgZWoAa8
ni2R92dKLlVPlrIUmABU2HuL19RwSVA0F2DCqJ9OEFzKmQ0GvwJabU5yIVDwTUxg
19kpbs3WI9vNewl/7AXvtxaZDJ5oUZg8+kLdt+NPMr9iXXSsx9Q1/JZxapU9S/3T
UwyA9Qm4n1ieBg0Oy8VwJkP6rG3qnYNH+vdR5cdxLZ760b8COvj9COFtUJMfEcEt
1tr5mDzugHSau/dajHvXYa/0aLksAb4s2sN0bY1c/chIsaDdbvHTgSY3oMKHVJOW
Zt5PapMVEKLnzDdcDViqNDtY65lMlWogO3lZxmBNXdI+m7MUfEUIRkpfFS23p6CG
p7+AoDGraD+cuXdN+3ZBtbS6hC3FbvqLsEnfC6Z+X2tDgDD3LoCY91RapWHBx/Os
nwRd/aYomcLdvkfM80jezjj4NBVOiYbKWyV30lKkCabS4g9HV6XcUwLbInqeJwkE
+4fiP7Kt1ztQqbMOOBnLpTjUiVqhyEztrZq8pLNDiQqZtwhZDkfsk4u9zCDDZW6f
o2RrBfoHRbmSj5znfPcU+OkXTkNaC+N6Fjacw7pMh9x5QzCMmAlSoWrypCklF7zu
TrvMnQmMIwUT2itQwrXgRaVnT05krl/ErW+olqtEgCTI+xtBobG14wEY/1zovdMc
yWDu+nKHj61KUOFNQKqCk7bEcAVNzmU/1bHgG8YVCyImMnmyPvm3P/VvUr7mDljW
LRlR6A9nKj9F0B8AXOZepBsZzvNZj5nvvUQhLee93xJ63N3Hxbxb7kuB1Gkw51PH
ZN93OeZ6x0H1P2Mt2LcF9zIX5K6lGqVSx/Ygo6TdmxSbtGv2pjAE68whi97iKeEA
4qqdkRjSbqYouBNlVqAD2kkk7ZcX0U5mcwvSPYW+IRkjxZZezQZETlGLCR4dHdpj
gvb0t3KwZ44As1rJwztSVe8Z/TB4Z853Ul6FU1aGAT14TZPK4i7YuH1ktKxHbXyC
fJMu4ad+Et0z5rxAqPUokUyuTZQ/BbueNsCFroLFbUa1mQa3x2OtD+qLXMROKF53
Lz+j3ToOS92R5SicCYzDVdvbNNATWFvyl/KXfgx2OHDURIxzrLsDv1iiY5k0pQ54
vf1lUVLhgfyPRlFK0nXl72pt4F8O/wnjnSoJ+vEa1ZBVRwZhypdeOcUY9833AeQt
RRFaoxaPBZBSF4zuTJTd/YHELvVCLbVu+FeQO7qNZu+bUBujPWTE1NZuRaGrSC7Q
6J6Tpo38AiUdM+5TygV+40uIoFmxE7Z/02YogjKZRUkgEbRcY5qpmcZcebqCLYLw
cf6kEG5kOoxvo6Nl5ftEaW8EngCsKdh34vR5ymnYY8jLSuV+zntMqfeLpsDodcGO
rxMysqSuJrTRhYLAtmC/XnJwG975h59IUQiwpgLPCS1RG0xrsHiQkKcqbf92uKyP
o2/q9uuq+dLyhR51kuVEuCIBk28K+fV8hSlWi1r4ve6zD+AHUQjQV67PGZbEWmnr
iBZ0YtCracNJtt5FmVHTtC/hJIvv0ae7xbwnHZpu06rGXu2XZTGS9VtWao5RlT9q
4RQK032heZlb8bf3bzo2c20afcvZGuoSPzrrrGVZ4lQn2/aSgOnpi093fZcNWY0M
BFIzSCPPYHPXZ8HJN9HpyuwYm2vVBfi2pI72cOkcQID+fQNzEEYHRFn6ftO2XL3I
8G5AwfpHFr99kfJkIZPuR1DmR5lXyxm5NXcXgP/8+pZny5zREAaYRKMijfc5XI46
BQq/OMmajvv1V608ETKL4qxdjuQ1WMs6N9BmMo5yxJUl36CEG1u0AQr7fZ/MAxDO
cFCuQHFFvcDPdSh+iciebwsPJ71RoQIVmXXwvE15EzRIiawBKl9G5yyWyAUgKk6u
KQes4mluj4VxSz6EiYqpufNTJBsYEuUK7l3cwvLbT0m01LCS0TyCuRmnHyk7Uh2j
ScJQAbj8nr8T7184x4+rf/E8YxiIvoYXNqL6Ns4y9YlPb8kXlLdjiB7EM9WBPdyk
f+ejtqOLn5PNd4BqZZnVnjnSGtKwE8epr12oxFit7U9YSysQ4HUZLu5KAEbfhy+L
oYrhpudGS0FHc637+jhWsJ2cKPfab/WZQmn74UwYMUVVzUkE+gHAfKMFG9h2/GXi
2zbVKCB3jetmfszaOEBvhDuajnA8HfOupkj7WejdL9EyAtxZZpR+gVlXIPkLuIo8
BUk9mDsuwt05U76I4/pxze4oRqFqrM0Zyf+ap7WC7Kaj0feCbRhweNG4p27/xrao
1GC4X5KQwaIMskII8O8b5BEIRkZzSSIelVg1bmTxT/P2hzaqxAPOM0FLZp5AUi3F
5IQ5OhqHquMakqX7koyesFpWE23Zb/IhNbMNNE0Opnj6BKxszTos+i7I1Cm/Cmu0
RbqEL0gitbaU4Z0KeIymR+M0ElRSHeQDEUaDJqmd6Vu0OlX68hFvNfhAwW0G0fmD
cKoZxwGiAFhr7BIzVzyRkRknlDbNio8vzbRm5g6+R+cc6Yiz+9BNJrZFFXKA60dV
/l8+b10ww9krtVhpwGRupPaR41rT5vjT5nBPZoxKRlEWNc8cpIA8Smdibx7Q46+F
Fm3rbdtqARexz2/pzIS16d93ifttjNg8pY/MqXkjO2DSziP7DaSASPP1t3bNslfH
cbEWvspp67nDI4+ucLeoAC/aQvtJ6N2wqTLnsJTTAFLf3bfp4MxcYxY48SqvxfaA
YKxfyjvXL4YoHwz8qiCAIRhtNvzUIvTgfy7n5/mISKHI1dZCOibboOiKFs5Sicr+
eXNtsFmbSHAlAkKqfAobgpos1H/5I8KT5M3h3tPa3Tfb1zpnT4+koQzKWtYHeKIe
oqwCpzVRExq/8aZDqaY0Y7uz7VUpAldZCnLIltJZTwBMYBCxkPYgZC7xCme6r6tF
KbGfNezTmDvM7COrB3Y/NklpvaCuTP7xZHZDLn2spiLd8OA7xiP7fZ8SUHxINpY1
UVkznhGTMGjEbZYluPpSFQHncZpNScck6EROphxT/4/1p9FoNbQyn1BR10FftIHk
l2/CHt7sq0weLfuSuOwpwLpvASiM/+agwGnvXghqhcjC2TRJIO1jA7wMF3rgfwBW
cSj1yLXHdQymdbNMVgv3F2TXCv7OpkyqveTKUzIZe3EHqgoxjIK4zjDFQF+OSgs5
nivh4zXD+WEbBVAmgU0Z4KQhI3f0OZWGdVVhUl0jg61KHyzn7MW5MViVuhV38VNi
PmrxuZPXC7bWeXq0wZa63yHweFoGdwUowNoYjrKbMMZ/GVJw4/byx2yHSJ5LM4aw
gAykA8aiucJlkfcOoKwO8CSvalc/pPQ3fCteV6hvwhAMst0CmSNkAZNDUhqJE1Q2
J9GavQ4mUZDxoV1y7QQw36oajSFltuWWkwXpX+aO5buniHfZnNZYr9LFiI3l3CFS
x7EEaiz8otK12LsBbbzgxs6Jsv7skUlfU+grxKs7cA9A2Wgna27n/mi21EjcpqwG
WXNLsa6JJ4fzIHp3zr10W7MMIGaCL9nnJq4F6t2FwKfcLJBRZ+4vj80shwArGyAQ
x/3v3FF7SjAHGa73olGLRfjBIV/FG6pyF8SZa2RDRpsbYItWQFD0KDIs5Cmn2ZoY
mFlU5g76b5RFn2pkaZltDqapX02lCplTULneSmDi/NLlpziV1UuPnOVzTOVVzQYT
wgc2lKOLBzCR92+Rb7foBbVWzL6F9TXHhSncq/gmXR/eEIiaI64CaRvAyvTEimjB
3L1YRtehcgZQ5n4hoEAUrfZ5XyoSP6UllTxZ/KSpRH+D5bWdnMRkKmH6Bt8S0SI1
bzZ6bsDC1JWfz8xnfRQ68pkC9pyaBgv0C3bu0ABJMeV/HiIdGI7NzuJ7ljvT/Eet
9z0fyvtAE/WYlMnNn87lPdL1tzrv7gH+q+dPf7lsJf5RhzkWk54ptVsQn2DRYpB0
uPbzkiZrKNOjGUIXqNPChIK7XKj2qpKs9p3u3o0dIMlj2RJk/ouSgmdGuaJQP5Ke
BNi91t4D3FpUuYcvPeUATqIuMgIm4hPsiaUwVmvyMA5KTdO/TdT7QN/6t3PGNVPw
q9CncEmGoVyzlm5pDNuZrfC88GWsuufJqEibJMD50td3WB1o+1hk5SSxkdd3BcFi
y0Qm1e7eveluIx0S3gK1BetZt30lYjqhKrPe8M81gr96zbZbP9RKoJtVIRRDjg7S
YscW6399gR71siZZmhOr1Jj5B0Ce6XXl/gQSZt/1T8aJQ6f9QBr4QTOsxK6DgC2p
aM6dfxWEbx67JnhoWzWvlmPptg2nUtPeJjraGA5AbcG7wIMue0jlhVDBE91/HSCp
baEOfHgY+hyc9ISnxZQo3V0/9XFDLbFYZm/EgGcHt5/6WfRTipxOczVRcv+UEUnD
ylegpo9ovIQaMjIZACIkt4BkEVDI6UDvdTvvPv1mdOEEXrFx/Yc8MxAYekdFB4yb
yJpVRCFFCdyINN1U7rxfVWIbE7iLq7Uvv9HI2l1wFGwR29CG94JX+j+EiQ6UqP5H
eRNEVX2kpkEwzm+x1afBWFaan5bBV7v2/Di1ko17ITqnmsoRXYWhV74EN4kEb37I
B8wMV3j8QJlXIax/o0T9aXTXTxFHCyJuv41+6sCkK0gxegWVUjJ5FfxWCpsIex2U
Qvxo2Pxm1Ph8uA1NBGTAiSp3Co3f+3PBlT0xCyyR18rGZJRiXgTgM3mp+/XMnUkm
SpTxuPcSA/47PsbsCsdQhw4ayBSen1ihsfrIzcsOQWdhJjy71lQT/WSWJtmjxD3s
Z0aXyekXHPFM/5HzVGpRb3uBs6ghiLGFfBa8BBSw6hSDDpHL4I0Fad3ECajpyTK9
awKnJEVqpFVVPcthsYMCgl8Rjhlqyy2xSGocIwzxplnV/bLzR7aEA04jfSIuYpOj
KM5VLDOaAWQhIwufYFGsBfoAnTn9DeSDyyAam7urayVi17X1H955TADqNYOzjGOK
X4NuJREF9C3sxduwLJV1Dl8RFLaoTaLdtzFCfhufquSyI1EqbOwy28BK2ATGdq2I
W2VhV/Zo1dkz9Cz36v0UOhzp12bw++fe6NrDnQ9IBn55Uqs/kcFIJz0c8/r2rs/z
IFNnnCVP55stDvgZcyXgv0oyYvdo3ZM4+C9F4G1OOuDz6uiRmyQFHY8nkKWhxkDy
uRXPEzKfdj7tqbozzd2AtJv7cGB1ff7fEz5CMCkU8T8R3B3OzKvEEucnZ4JGOc/x
eO3Ldzk9x64Kk77xYAURJc+ncdzj1upeVJ1c3yiuh9vnvdTsGD4ZLjvvvEQcrFW5
0dgeP5nW/CsMtx2/UeF5IHYnAeTYW+7vZaCVNq44AvvVwZpyHilLqdM/BswqtedO
rxyTCBzv3w1/C3rhkVDt6rPTIBapzDPvN+iKaHPtrbEhB6Dx0lB5HtuN/RhUiP3e
H3Biqshe4G1SvXvKipQC28jcnopprZiF9kMb5d9ZtgDXIAiEYTUGjNhD10E8jcO6
l4VBTvGJAfrYlH+lJeKXJae076yhfHBcQzkkkPpu17HDkHwNH3XPV/ZvZJUo6sjg
Fer/f0b/sbwEX+HClLq4As8Cb5GBDzeN5epLaH0EXD9CCZ/nSSNBrrKYGQ205C2y
hCvNIk6QEN9io8bz/btcKxRmQv9I4sRTvATdidGtyjXCkBWKiy45qOIkq3x93MWy
vMxqiPV3sPXF+R4oVdR4pT3wHwx8BXVICmxTRJGLQ/hOBdail3Mkz3DcWW57KTyO
3/agih0szUSGibxYBaiXgSJc9eiGKqzF4unQOBuz3ia4wo6kfMrTxwzFbM4iDPit
kALaxW/ufAqZTArpmJdGS+ZvQYaXHRdqXX5Hc6HmpO1PZ5xrbwYQ/dUmSIQWFQQn
utgbtqOYMUg7fKoFYzlSSpYH+3CA8yCdg1FtGiX3auwN8ue86V+fv2F66FnoHYSo
4rsEIrsrxcVZzIQLfNnR2PdDNqYTpejBfhDrksAeN5mCBGZiil2BTJB+vOCQQLff
SvRd7wgZB772Sn0wA5LzrQV/4Pf9j/8bQmv1xv7DC6zZjFeUdvfFfnSH98Ws1I2U
DpAAM7h1KZemTQLbyqlSUZ1wbadsDpK2HlNIsCTV+lyinPVKpZlCG9uA3DHGPm0M
zaNAF3Tf/jrCSYwXJXGOVMWbYWClFsvvlER8rcOMXQ0EopAC57CkQw1C0ddJ0R2h
TBmvtHwsqY0Q7+simox4iUtMNEmbGFoPDnD6YP2TwFepSCavicX1cBIz1SrCCvJv
lc86sGY9pWvlY7+rSQDY6mX3BCT0Q6Vs0tpNjjsJw18ftHpWAhddsQitQipOa+FT
ToztsrqFFjJycZBoqMYSjpU+mB/eJXLFtKXqAEyvo1b6cosWMe1NBKcinljn0FCp
p37jqGIqKMao6sqihM2bBmTykJTcjPvKxrhBy7OfLg64Wg++DCCrWtWBO1zbSz8h
L+tOr4dm9jk7dqS0ZM42zHwbAt0AfkcYYKSKSv1AjcmiAPOyohHUzDVXFfpRJBaL
gj6JQpjCBYkEVGmcEf3msTVvJ/rKAbSk9Tfg7WCx8AFhkduEWKMB0JaM/34CrXJ6
LnfN95+IPlpsI0A+5zQAdUbu5BgGICfdK5KXxTyZVmY14CvhqyN58HNcsQGnabdT
qDnjzFwuyDeR13TeM4kAhaxx1Yn+Ul3cOAuCQuFZ5pVKjImJAF4NJTt5HZRz/st7
qxuddmQwvIJifr0jpzxNm8YCWJODbvrNZXpjhv6BINBdVLCCYYz1hsWj+cv+p9lI
WoLS29BrMn7NqwB0N+66/viN2DnPV9WdXR04hQtjPeHLku6uQzCkDxhs2XzsyqAZ
wbMkS9DdXZRLXoewAIwXZ0VX1JEJ2haox34s8DBiBH1WZZubb10hn+/9UJOcgkAf
VjJ6DS1lxTVxC0wjvmKJ6aQ5GlnP1FOdfx98F4IsaaDW4iGul5eaw4wJKORLKSxt
i8l3DT9HR/KtmbUtevJVdPIh7VE8ppzQV7L6J9AKx6wm2YS82ALBhN/dmRwgBhAt
tJD1g7CE1zWOua79jnELRlfYAARcqPUSU854EijpWmnpYARwmQY4rTmQ97KaJUrs
WA0aVRwbCsVI5fGAlL+qUmb5pX1C4jqTovjeH5aC/c0VOcbOPrLyoYZdZ7s1M2nU
8YZkEGpZOwLJOT1R4f/csxyeYKarjeLy/c3d2DCxR8QKx2SBf+2h2SDKcS6E1o/I
bWYtyCoLu1mjqW5bXmDtv77O4y2/+T+1x5SQZldwOxxiJogLY3XJTWqBpwsW78n1
ARhtEJUZvs1YjOzXhg3NLZboqRtfnZRFGR0dvIpaMtNUd4GehQLmjn0eOo+MZrjq
jg5yPjKbBdNdmLDXG4C2dJyq+kRg+InpxhABl+EHxwPnoZEgcrocY4qvBTq2P4wt
ui56R12nkljW0HkEMEvq82ngXFfB0Bp4iK8z9BkcM0dtBfmQHkMhKhaA9cUpfa1X
aUzzPliYbDaS3XFXPyWkdZIHri347eL9zyyK3g9h+0QqEKs2YoHJlposk+ZRo9yN
TAL5waA5Extp6QjqRipssqKslQcG0hsOr+JDJ2dvLzwaYpBak0ZsSO+rIrgQlafA
6RF2XhHILCIR0yxUDsDD75OIAMpnQXYLttATz9K5XN0P9tqRL/L6eU4HJGCMK2kP
jvmpzkGxIQ4YAL9Hg3o2ZapvFqgw2i96OsP4cjuU/YJ6NiGgOAy5ouAYyf0GbqMh
dP6V1wos8fw755tUmArrC4Y1U3TX+yYslebfKWSwi86VNtFYRfkh+yv7gYGF+ePB
DQMEonyH+kASjOh6BTKFhBEqehLOxNzp1K5DseHvMvddwLnQfTKJ9Nq/LVJn7H5k
wfk7qaMwHEgOwKDqdQIiVV3TBFEFP7/RnKJjzCGUyAD9BK3sozMUemq7dE/MZN2Z
OpMSGIBsZdriHn7BaiJ87Wa0uNXDjw+TSmMWV+21/X0nuaTWg0x4Fk1elyFrVC+X
BUc7Bl6EhJhn2AUAHJdRG8iC9N0wQRtNX9vtQlOLRRW1clJlzSmvoprsF4Es87Q1
inVLs/yWXZZWBD2EH0cZZUOaGbObf3rGXSeF+8cmLHeD3GEQmiUNfUZHUq2TG0Wo
3yGiYKNu50lZSFCVZ4QY29wRipMa+nkWLgBUp3aZuN+oZhmf0AoMt1uMr1apmIPp
i2i6YKr5Dn9sj/n2EqsXdywPKD1joYndbUlC3KAEIMRfmEEgBZms8WP3G42gKOdq
69XkdEHFYHtb8NiE5Qv2fEqMF7zJCauhNNrfS6WGg6/xLGrsn6plsbQ+byzYsmiu
gK+JC7FtIYy0zIoZE7LFFnAdY0eWCzxjDi/KSqI9mRVdEMh/B1TOdRQ7SQoOYr+Q
ZWDBQTv9UKSnqsW66uEmr8OB4BfTMfMDe4bV1vfzSs85LU4iotLkkW/ElMsSIyH/
Ad9EeHgc2YxLo89j1gR/dHKvBMw12WZFeN2wbl7DW6y/fR/6NMH1Feq49mxZT0uM
LGPD9KJvyVmj182nmio5gslYZ7WPlfkU4f+I/YW53UL4+/EUwzazd8wy95kUXS1w
VYOan7VIDPasl2wMgVVD/vXQozndd120aU3deSAru48Q28wM1CXcdZNgjJ71Pvqo
Gy7E8Y79kWQ+vd1SPxDZWcKVZ7JTYZ5sPUyfFDTaqJIWKjc3/hPaVc4FVr3XaecP
3t/F3WUdvwTvOnjhPu2SFK8l+SP93xY8p7Mo7hNBcroyMfRq14uaIbI1CDaC8nr6
TuAw4n9U2uE0Wxe02XlTCXRq/kjH6/KgeLVeBdMBp63fgaLEanAHTeeVAcp9YPft
SDcZQ4LSP7iBdkm98wnHFVbPSTqvgBtwHNfiVWbDuw4Fp0n5l24+ghn433rt7m5q
XiXMvNcwu4v3b0nCOTpdJkZshvHsORjxu6GKojVAzuYIIGNwSBGGZzuBvjyxG9Y2
dX5qXyoDgsTfna806CynOp9K2QJGks+e0To50p+N5OXrJQJBHY0snQYo2fOG1kCL
ZZrPdgvzU7UO807lIkDuM1YfkjE07DFjoOsEB6E5hBmSOr9KjkfjjD60RKM+wy0x
Uo4K9Mm8kupqgIVWyo5vkIZymdb+wqliBYSYHdwwpHvyEnLoxAaaj5+oFnOyGzY+
DdoSayo5GmwSJfi8VXibxb4wkQGmbkCGWcmMQEG2YRtVhTvxZrePIqJyuOC5ffzV
4JYQ11HbgGADLBnte7CU7vePo9AKHYmIlB2JQqgaqUG90B0YvXlIjG0oWc1l8vkZ
cuuzMrXHIDZ3QOK8v6oQDGyyF617r1L362rUiZaSR1U56iSdX4aqTlWjaazPZDtB
2J/ZCJ+E3XS6uHfWwMcDkb3DhKbQyBcTdl8AuZ+RQzPJsAPuVfnbgaTQGF+ZBAFg
kiT+TwMLzhIC8z4UROhguliHHJI2lODrU4MSMEXSXUpRw6gUoYEArI08dvMMiXTE
PdOCbCMiAL43XP9J/VYWYtPu0AjcfMfAlBrFfQMZn75iiKR4VRQB3bwtxLzfvL+n
IViGSx0bWMzIHR+oabGnGXAr9df7a3NMq0fOGqvD77r2dWjIt78fcWLU2mXI6HTL
9pcgA0JV7gozyj79G4FsGoHBrTVmPcpBTZINnY62YSTEeSEHk+8TT6zyXHsUboe3
guG8WW6APfJjY+V4tJSmfzTdXRlFhRVs+mp1z+TVoinHaUgYnVEDGxXZGxbRHz+C
G/fSnW5A9sDMmuHqde5+7rB/UQlCKlXpotkvMoT1uvjekdjBPDuvHmaQrbqwDskI
sUmfylA1LxI3CDwAoGwj0OA+wlIFB3RHcUwDH7OqZKQ8I3s7NyqQicll0HGLWKj+
Rt+4oxd3HHxQHcMPpyAAjLfUvXU1giNVJxuDyH7oaBNxMhiUgbH23oEUlIk5xAQ+
qRVyyVzqLrSWUbxCeZxdS9nKUiHYSmlkAGKiIea6VS/GjOuqYYwkaJIYiM6yc7D+
uMhDEJnN/sRwbz1Z+Z4TE3Q9akTdO1si4pczPdVSfwu0MBvNpGq43btMfR1wxr0N
1gKGC6gT/DNGwGutLFYdtKofVhA3PDykrX6WjNDXaGcu2sMLyrV3ert5ajPTXMeM
Ru5epcnJzhoeXww79+/OqXzpjTqh0DU/IIvt3ArullXte9ve2Ru6S+6Y3x4f5SxM
2M1f0NomlhXJuo/oDY4HEeYFhR5b4DkLYSOG9e4gbP5Gi9EEXKwcRS3BX02pUlHW
GdVYAHhUwzesGC+NUs8zTJ/Rf2PG/G1pZIFMihs9Ub/nZ0o4PpcU1wT5DfESkIhu
sfbiP4Bt3O+5RzvTRzjy6LqiHwsnVA/KHmB8gWJ6bIuBtOJ4KvcP2C37uWLNXcnC
yNDDELIXp5GbhScWIgitZsa81OvR0SxK6a3/0eebQHZta7AGF/aVvN5AjlUbQiBN
En5hLAIQH9Jq5Cn4WuG7Z6bMA7oywEAa6YSc23rrFukchKCUoqDraBAIxI6/EnAY
8iZ7vI81NSJXcPBrxZV85ORAe+1BBYOD6e1kRD1uL4r6qjlG5uzKuH3punrZjoB7
W8C0rtSh/HZgobiDKdrHIT0EZRN6BI9oI9i2PlVIfEOJpHppdzQoxs6Jwb3Ot33Z
ctw4pQjW/B6uB2Dhv65yc7/UXFq3AIbxNoiWVSk9JDpUR1TBSQClwDz80v9dUj2t
Jns/+xLYp/maBnzOJ5hH5GDIA/Oj00a+rj6l7YOMIdkw2k0pB9QHzNrOztLtXHo0
g07RxJhGKiB/OMP9xh+jnDSxg8jfLUl2XhzlyFEeV85xP+JBFMUiPIZ8eL0TQzeF
cFc99J9pRjuPsHr0E86ZTWpM/vYPipmwRRnEc0klLw3fTnbOlgaa5s0uKH/c5xYu
WnB1vBD4vMNCN9qKouH+nry7QlNQT5XhlidzuioiQIhfDAnUxndHdfK8TBy9exhE
+OG3+siOfPajEKgDIA+cobUvLmvpLdhXhZeLiHDS/cWTRNs/p7CjtjzjnJo3W2m3
jXD7smuHIRBjCP/G4FglgWUsN+JiH+7joH40fFHw7l0NhHrh7ImpzNj1GMqMbb7M
p3bP6HMwCJTeAgbhQ4SwRzQrnE4KGVrzh/3C4nhObXWfFhTLwed+HTyi0k32ESxS
3TlzjHucUc4oOl1/gjp1fLBcHKMCl99+PbEmvaDrt+VQ/flFlF055TmMPPglHLVT
rXuOcCuGl2OX5FP+7sR41TpWNyAIejQnFDRsMa3hkIzbotBdBfkAen8M4hFI8viW
Y9gqJuCemmaTywPi0P5gsTrIg2K2/pb0rYVD+QXsD9cb1EAzfHqcFG8jfaEiF6jU
LRI/PvV0MZxaShrUxpKbEn4boS45rkwf92h3PkCcsokyvfAyNnvPNspArv6ueazK
10xmeEK29R+gy3q+Pbs5LhhH9Zf1xGxLQAWPq5yeb76Bdlr4cXlgE5tppEnhGXXY
OovUhixY69PBvxi3kISSGe9x3ynR6Dw/XjA93VHR4011Czc1TOFug5ctxMqU9eq6
hSgqsIXv8q1tG5d5InZaxq/7aNTou/tSggGUl9A7ug8nAEr/jIDlkVVc96Xz7i9J
08IUiyt707KPjG4itX1ol2diVW2oNqPXd5ekcPRMYgKmOaMysLhsJTJVlNfd6qlT
rnOjbfjjZKOerSBYBA8ALarcKrQ6HaPW9TQTFGS3WPKsjqmw3eUQcdRRIRASoSSW
rZoDMuIOXfU/SOq8hjZCtHEPTbt8mma7gXryTRJTtE0xNfCc31xgRm75XdzEroHL
I7JkL5cvGU70tWXXHnTHNhh0EyMJyj71p4RHxGQq79YO6LS7YHlAwOOcfSVBmNRX
TUe/HkpaEGWhE2KTD8hzdIbEH/UTWw+sTKWFlXeoaDpmo6G11xaSjaKu0ogXLoyK
o6MGLKtb1SA52EvhVupRkbww/NOwgtYUwbiUEclKpou74ZOqP3U2T9Adua+bZAv9
mED/UATakFIqp1CWgsWELTEtRaIyMAO/Wrga979gNUNqiWQhICLNPXqnSqVEY0nt
GEOAT0HjXGcCdGqHZvIYo7Qpp96CUerHoR3HVmw0KhqCj5yj4o+eXc1sbYCYrceZ
Ih+OwAwC6wH1Sgp5Jy7qQq+MuEKRKMsuTtnWmzMB7/nEt45woL7AedOfN0Un4OsL
l1R7tjOaTYV70RlTm05RK/k2Bxam6b8f3rrIYYsMgZCvaFmeRlmkbx++e/Swwzt1
S49xI2t+wyVKA+XPjOopx2p2MsmU6jiz+KYWm9sPhZDjhB5DiXrQeLbdysa6wOj6
nRJrAsJCkKMMA3uU3hU1dpHyqWHpGuCvRAXEEnC0REkKSsb1LoiNmLg75obEOWDD
IQ6fc8mCF+g0ypMc5Je8ikSZ62xiKr3dV8oAd0FggvorTEMXBq+NHr2xzd4YbY+e
J29XDOPZRJiYl3DeWpo6DejNUhb7rfYEYEgcizeopA0a6LoPJgedBD6IyPBCs8qi
GzepTAfWGPYfCbO4mR1kruLhHYTKGBfRXWlF3ZD2zxphtZj6/tpJwePbATX33VJf
7QZ0Ym5nfVuMG9bEha6D6kRY329cirqPRdclCUykhN2oOS5vif58Btewi7iTz6PC
SUn35UpgZamKN22yJwByfx5JVcTyASwyiRWOj3YP3n9efBeogBABnU2ucAgR8v5g
ZCnMS7u5vdOL7qrl+TL0D9GB3Vo8uqC/tW4zHezJafa7LPxz99DTUV/K8FUVW0jU
wI85jpOGTVDYiqtS79OjXQywvl3N5MImYYBCCAWduqgQyYOPn0UgEtmLiSh0Jvry
Z6pdQXg+r2xlVheJdGoMJCm8bs2TRiPn8n9Ol80SviMURDxSS7qzsBm/UY5AuaEI
J4hQme9vxPTR2VQ66ZsA7tpsXOMx3jPQVxFe0LBtCMkEsSP8/nXC3pDC2pGgXMao
7WInmlc3trL+egLYlMtJc0mOu3KQf9dLWXUKo5Z5q+zNEcHLLrl0YmvTWhRb4rty
uPyICX5loAVOFNwISuzPMCLamyRoZrHo+PKqNGbzStkDJCwYTAVCb8US8fQm2l4w
PsrSkA2R50gFdDB22Fg1TA/a0lJfp8QyzFkoC2+kZ4DxtLBMT/GvvV7Go6b35wqc
mxL8Fq0jkyWsDh+9YWHlbX4kTEKWiATqAwropTl4CG3S5F522o66xMl50p9bPoT8
uPhG30kZdanl3wiEgl/POfvkaSolusB2czm8MJFDRLkMFfE+y5d9CCvkgTTrtxoM
jImLHF2necOFlrjLpUPqITpyQlHQ5MnsdHyL45o9HuyqwAd8Q1AmV/44zG2jmIee
QpGMOWW1Y8uoGC/laHHQvQ==
--pragma protect end_data_block
--pragma protect digest_block
3ZVpX654kyWEgDOGypZV7wOddeU=
--pragma protect end_digest_block
--pragma protect end_protected
