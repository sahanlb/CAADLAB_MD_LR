-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
hqQuwBNF7zhyTX94+zMBXbZHD7J9InUrxhE9VAITWDKF0OWXkae07QnFu9QnW22v
NMs3AWh+snHlD6hPnDlpJDzUgn6TcASAYmsesLDOhbewLluymdA43IhyKTPLjMUI
KXHqsBMmew7cF1L4SsqpAa0FV38djwKMxAsg5sQ9UMk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10668)

`protect DATA_BLOCK
iHTZ2DHnydvaLxxXh9bxjtXyiqFy7qNcmDMLHslXy0bO193FMmj/4LGr12A6nUp4
vHcMM1hTedxsB5yC6Fg148FDmeQyGM9ZPOjX91LhiJfW9etVafH/idslcwrME+Wl
PNNoajQOWu7ifI0Ij8t0x5IBwxUwKLxlsEj9kOf+t8A5o6eUV1s50nYBlKNBM0FI
pHtD2w0ndImSJ9YzzeQl0jVq6rYYnaWY9TZH7y8bTL2JSjNLNt6o91UD2vaVt9aN
CZsu+7LTgsTmjjpVjKMmaOH5L69/irtW8L8dQGlrWY3I0QaalPyrSusYd3bXmzWG
Bnv703xDBOKfFjzuuE9mQYF6JML2d7h6P4Mj8wivGg15j0df8j9rGrDfkJbeK00C
zya/ZQyDwq9N+I4AKYxYLQ/1EmEZg+SlclLs7Q+PArCMGjcdh3MCGfSvfJ3vDILq
8i4Y5msFMcYTxHeiBEHKNDV7tv0kNKeLrquGCI1GbGQyLk+XD3zg6O/0gw3Qr0E2
wYQpHBRjZSU+E8fqzRyAohGslmBAlOoD0WaFMy9RSbveEaHU3Dfxz0axcOItRtZu
q4M23gXN9Oj+PfYN5Kz3K+v/YnlP/86IWhGMf+QdF3UqZAoLIk6PJiegTIU/eFGB
pT4FDrxjVn2F+9ncE415LztELmAuL2b/OD51djmgoCnsaDx2HInhV1Orge6+5Aoj
LhDb21l4/SD6m0oUfrTWak3rRuoxrXZoN0zwDMPUAUZIfH3w3whEE3OVN9VtZM0g
iPEZQ993mizQhWk7U6RVKeBxq53tIOMH/+r3rBFpiq8Vr6fBcbRL+srpwWzOT+GG
hbjxYcgIgyY3HWdKvLdwIR7S0LEmzjtv2l90iVCQzrVSgaUNwrv8GYscLwAkiqW7
eaoviUo8PzkUSrRH+xWwBgnFZYoEN+mTk5kgW6q0WseUsptWZ8/oZwivQqpL3f5x
mj28qEEEgY5DqE4HddwY/3agwhFpDjKZDS3db9W6s9CkxIDc/yDKZn/i2t6gSDHu
NBXxx6vj1icHhKaTK3w8pktMXausUlqGTM+yzu9/rK0zxiqMjTLQg5TbKOw9Np0f
KUJxDDOpHK7GDXAna8kAVveOuVbzEKHYkxIXoYpkxs4Ak9l2GISrzLvlGF/GXCQx
RPEyztKXN7fy0csPw/V3yGL3RrPkZam9yVICCRq30Qfw3CBaC7wpXb2/eSM/fMtP
jlJjMlIdk4aATbamuWQaOPQGBtbWMVbuVQtXINz2na1tJrHcYsogyoQSBUPVVpVV
lRzsnX1Mjiop1BAwapPsmTQuTvKEsF4qxLMi9d6XUxyGHq62/jOpasDEjzzr7njN
9g7mpzf3h/D6zI9OJ572bgMP4WnDLDRklhbxMgMWkvBW3l+6X0cP3Dgl5mA+57i9
g5ccGn0w0XbUfD3yl9wv5ogiLP4GrsdK8llTkmtpg0b8kvoPt/ZbtWXjX+vcbtF4
N6QKJoi0njI42r8yLSuCtgsRyNy/Mn5EPZl7pkSWrRan+Pr5MR7Qw22SYw/DICx0
k1/oldnS5nc+51yVIQn5AuEderENXCQi/eFgqoaFuj0d/SLanlQpnzL/UxiClLRz
rEThUvinWy5ldCKuYil39VObTg/EW9DlT2zTvDbLVk89uoouK7QEOrKkzduZGC7t
t46HsOVsRFuojxaNRqnXJr3y+968hQ7ipXBINyqdqgBZhx4etdJN6mDW6Wyw0Ogl
ZhKBqkCDfGGSAnR1lD/Ma5HDdOajKNOKSGA48hO6/mfyU5hs3YIp5kYCUsyK5zQ3
dVryrjYS7YxWl5OF0fEPuiOK3ysuohCAO5orYkp2YPP0Zy4gqcU0l43W/3GOVIgu
yP2b2mTIB/JQ58PNpFsLVXrnfHxC2bAdMG15xvGC5Cg/rwEQ5ASqa4LiyofBYmXU
aeN219/2vq9hf9TXtXJHp7Vyz/XeMZ0TnDhPztft5vHugB/3gSvXGwE6+OZEa7lR
rrvHDANsqemMPRliSPm2qkF4vv60r3Vtvo4xR5Zoe9zsbelPfFLjY2Ikyx+0Ko7q
9jPCEzTQLm+KIbYVQ3aHVP7TcDQr9LNLF22fuuoZo41Xo+URr8QgDzSmdixc8BH7
0K7dzI9F32AD1EOOcS1P00loo/N5cWRj/3EeSVNk9AOokFfUMLG/zE4WCmeSVYfK
ckym2GagH9ITDKCKq2xWB8/FvoJiGw2MHj6Vc65s2hMtWREmjS0WyQh/MRMaNEIw
uY6iMWsTXlIONzS07PW51kUihZTwgSfDvZA+RY0WU7KRvq3rbE+eHkmMyQalxNhZ
mNytIuJ9Q+fBFArI+7UczfHEszJ3zt16Rc06lW/qTZ3+fBazo6VARoGEXAaecjwm
JJFVsSGtCKi8afiBctpOsT9bOQtUkjK9RRFN8oN4TyKRyKTemhPEAfxakdjF4tI4
+ryMB6caVl8v1wcYx2OsuArZqaxhdA6jsQdZSQK9vzlMw4ONpY5BHn7yB6H7tku1
+QYrFcQcBL0qb30iv2XegwRE2mOdwRTbgY0ULThAA6yj+r0qxLynwzhvM7oOiL3k
LjPuewaIsjAX+WZs4UfxWpPQfkItyp7uoMgKxEi7ulKQdhq/eaBaGFyZr7Q4T65W
Hgkbg1QSjAqeRCfYDn7/nnfVQ4UbSiBE2smmhnhgS48Zxhc4KkW5stboiaeoKEdb
sSDhOWi5HM/eo0Matmjdqeh1CCrlBy6yiCK2bFq6dvloq9kYnActfrFfznQsO4AG
ZF3slh+l2ypmLjS3N7Wp0Ztv1z9FNgNhzjeGdOtQIM+kaWp53rPkZibfHYGVIijI
F+81piqrMH10Aa0rAFbIa1hkCzzwO/kX2YAorSptiineWSsbz/TskyFxzdNBu4o0
ZGRXCF6N/0Ex9+ZKsnzWew8MabxmnHWbmDN8hzZN3aQW7rwnTOqbUR0TvRJTjWRR
tkiYexvq819igpSfZxS0xeE2Hmnok2ExNLmLteyf8nGX9RNumP0EUKk60/k+baDb
ELjg9jvIzMHvpG+8ZfkOlF5r6hfxRtXaTnw8xTeHqkCDCU0Bi4PqEQ2tgJk9iyGl
Rhuwmy6q01gpcYJlWsIocIblMet3y7NnKO73ltZNrvuGPSPXb+ZlOF8nJUOb8w6B
BNHr/3kOIWan1MRBYoj/szGJ3I2R3GL9covgh54flwWFg2rndfu6ByKU/e23sDXp
VGQad5xFmjXN3HJgJbJ+KodomS6xV/AN4VaimzdtEYreUnDikuz7zT3fD4Ts6mYB
DOfBzGNONd9ClL+bCwrNSqQp5q5iYAJn9tKaMQr4qJgKbWSyrm2J1UHu/+iq0SLu
kNPG31hYYhAknoiMTmKqK5iMabgV/Ab1h1E1SZewhylsvAqXEh3ctR8tR2jidzlX
pBZyCDuKsMaAqw5BN3xRHhknRMq7CWxJADijQdK2I17PqFQM7LJ/BlUzeJyJwcDJ
ZMy6PE+atFPd2K+739PS2zIDRsik5ICQRGKEgDMUQ4uLZ8qEe/u8xWl6Z2eD5F0K
JcYEBG7Z/qMtn980mVPWhcJ+f/1slihylE7MTTU7jrWy2VCULc8nC7zEAXvvwtKk
onlruVKbmBvVJFWH1y/z+l8Ij8OKdRVb4Z9VaCFtp9Qzzz565K8yEfSr3FvYfhE7
GvVvQkKLVu6u78qtWUAOoaSvjH8CdpTRACgoZ9ENYuA8l462JZLQJyG8jYdClFds
3pqITiWsqPkDLSC2Kjg5w55CmJZx0PMvo6g4Jfx2elsnXQAlI8cQ7lcOIOCKNq92
+0+RTWb1xCTrV+zdW5+tmjBuuQmIVxMoe+xE2ltaiy9FfwKnI8U07SZdkfmQ33+a
YqGC4aeYKQJV7PB6/KjvFdYwtg6ugEpxoHdjnhUdaI1nvm/MRdeTFJLswq4xreMp
J/PI4hQFbemdIpajEs1es9gB3tOJzPV3cqaTGgqv4L24KjrhV/2mlG7Z9stT4w3E
CEQUusQP4Mc/lRHvi1vQWISGb/dlBVOdZ8bKuQHeIeZbWPsSIYnWblxDaC+sLc5E
OjkWIvr/rLj1BcwvlGetDAu9lr/V9G0bLirpEzo/KlVnmABnMMkrdX/0BJup08LJ
F00SBgqr0jfG6K0GcAgrZ5L2VaOLG849x9XmJQEG8+McR7U56FeTn6ttpH+E8sn/
9QtTP592QlrMAQDSi3z8nNE2SYnIPXGZyhOL+WB0Wv38TQR9YSllUnJAnrsJEpXp
XHGKYMQ3fuuasGNs+ShAKKuaZ1jZLUhVwL2qsFKnvzhTScMYw7m6VcNj1xrs0B+f
hJ1DFe6e5ktkDKXnl3YqlxkEoWKAOnZWtVPZMJ4a7CPw2kldzfRzUJG7lrlfUBLD
pqfqGfqlbUNxGDWzofPkFTdTA3xq82xVracEUrjA3CJuofO49DQY+R9N1imKmY0M
Wp/ceGOc93tybbzD32GPq2Emt6wJvhvJqK2y4SdTODN3UGB3wyFdwbrmiPbK/U3l
iw9RZf4M8++/7fPELOm6tosjPxq+Hut12bkolOePXmQqqlS11p76Wm9HAXc9pgAl
8SyV06M60X/Y05+X053Jn7A0+J/sRexrp7DQlB2hR9d12V7n2/aceiiAxrkNWXIk
Ipv4ivBLVeUsw4wJa2Pl6886uxGosCsz2byvIF9NPoSOfOJEwizGCAMMBo1wndAr
6m86oiQpoFy7a2TzaG8UeTjXWON2ikLjIocC9UV3gOr/XozW5lBvca/HZ5yx5le+
v0L1ORQr8uQc53VF81oHiDXz7SFQs29MWMHiqjqhkspC4XrNxqRUh9ISqLwIYyW4
9M2AoS84hWAR+pJbH79kNrgU0wrJF5IagXJaEKZEQ/O7rsjnBq5egwOmPsaWQyRj
7QsIilCtvbisQazsWbIhwnCwXYa2JcCDUs8BBxWoW1v2m1Hw/Mp1KjdA5YANo9dh
MeownyWiChqJV40oDc2nMjD6bt/7/Xtv/Lz7FVpCrKuDnN5VTTZX1H4sxNvOmyGI
LSCFs8tHN0u8JUKoZeuIHzcX0VYz/aBX9qURl0TWJkGws9n99eo5frAuFYJTN2kc
EJ1OR+ChZnueiYsRRWusSz/YmBSV1I4b5BoRzV9EUcm2j2NTAcjtqCStxsQ/HRlk
qlhv42NIN0xzaBlCW0/QUgHSkw8JAE3NGcaKoldHaYLHtvbMs2ASmm7vGSJ/LPyu
wGLsCPZ9SyNIMCyQ6NKtkDh9DupSNa0LFkFe5A95ySYmsD3b/knpdSrCJh+35pje
pp3BBCEBHjw04L2/j9KFi+OzwsBoKxDiqJCFe7llvMh/BhDDRp4FuBDgW31kqg5x
JeGzhA42/RiOw6FgMWMO7U8/LR6WXtWRfRlamPsvrgCwl4qjva9j+8O4QmoqZAXB
uYCJA7RHZWCiZ1zdPJOwBUxdWzj6kXNx0KBHjQjKzx8RyFGHmiiyfrlkv9YhZWLA
4aHxEIwdE/+TJFu6WmJzyH63cXmy0KECn2i6V+yz6pvWUATRn68C9glhm6LYU//1
90oSXuqo3+jlUV1QwKfmeWdvlE4kOl1hRtZIoZRwErgiDLpeiLZUDZcATS62ivVl
pbKUvswaOznggDuLw4BaxLRQjlhZD3wGDRSO1tlsZlX9LBxWRpj8XF5je0xHFa1o
7S2rGp3VlPkGm1ImBRybvjvsQv9WIJmuCy9DUWyU+VfziWTn95OF+mu2ipurntwR
u/pCYzh+3bfIj/6Pt01TxkYgT9f24XAsguTGC++TLEhWiYt3nki6lEll587dYhUm
+8IIJiWU4PcyOFZgNSfJWiQdyJGodjdT1VFNXLZ8puvX/UsYL6jXIxC6raTMH97/
tQm3M/D5dlAMGiHDDEzuO49W/VJq4SR/YaLXy/NMXHcNiQT84Us7Veoc1PoAPlPW
zPrimnp8qCgNRUKQssBBj8WPEsgMGhoT3k8WHJmbJuFymppOqAOtp34dvyEaJrKE
dCBvaPDXxmPzHuBZWxTg/3TWp7I3cPzJ9PMHKXcVcr2b2DqCY5xGj4YTnGpgWA00
Ts2h/s+Ag4IRypWlY6YBPzRvmohRiAKZFEBoYxiCnpI8GKIP0DIlcQp91b8hqbfd
karhw1FTYaIczq5LFSJLJaYpD22pc84/23wp/3JO3gQ9rw3zbikQMc/13Z00abgE
LNb/zdNB5I2FEHUu+ppqilncACntwH+WX7DWLBhgfuRd6UDVVId+1wiNWmdDr3VU
1m1rN+bIvdaLOu9DeY8OL8V2A+3ct6XTTOGm3KwDFBRNCKmrNhxI4M9W47KCz4We
LL1M5Gm2gslIGPm1WwVBOy9QUFiDPHNmeM+iLhxQOp1nfaV12VHJstFiqySefYR4
P1OYqsMWnreskX5YbX4kQYROgFNhJ6Q1lGqvkw8QjNBdKMw0qLw6orI5JksQdg9t
r0DdNSuAmiSwpV/UQe6rEonK+IRwxDY8/oWS5JoQkhgASrxWUNVhDpaDlLeUOtoC
kt8sToGrrOyrNWF4GBYP2ilaobAnK4pI7VA+tjx+/gBRc+Oq6vK5/zrnrU4c6M6H
7sgA+PhqFfqryV79YxwDxJHjZxNTZYRrsO3+eHQiCP1bAWaGOrprAsio8FCfWBCc
GI6uNtv95ubnMU9grGTPqqiWsdh6p5Tn2E0Xcm4oZ/6sjJYVFUefjastZUkWbK/Z
WJpqR+6ArZZ//ZM/7flIcB8mNFtqCcjUOvwm+qSXrASwReLFJ2xPFcRQ8x5blJDD
vRiUfYnTSAkvpBGjdn5lb+5ONaLEEpFDBeO/EJDVcjL02mrm0oO1uzkkFkZ7xR93
6VA1G4ORQMSnzyiD3i5qjbdsAIpUOlsLB12ZqFvO+sCK46gB8/DLtjJlFTu1pJQq
NBIOaG1i1oQ4aD+PkePrcaLPK7CrHgvcFeSp4PbLvkx3j6J/Q4TPz8t19Rba+WjW
rzV/iN3rI4kT5c669myeNafn+aRX4aelDQ9IEp9yujzEWbofnXQyAy57RSBjkjg7
67ngNGdAf+aZGL+FT7WeKAL/xc5a9zkjZR7qIstDuypIM1osYpAcUQtSESQvXu3h
oTS5bI+8JSB9cqE9D8K5SiGlRihOISEp+HPylFaxOa5xg/c/MHZDVaaqO+vRfKTC
4wKKRM0pIcH/eS8ocnPHtArJbXmXWsB5+sb9vC02kjTANsS9X7RxGD1LmDxdr7Yn
nbJx1q0r+lT8OfEen/HaUiuQMxR36RmTNCuHGzAMDOPoWukkEHq1tnKoNNHTzWRp
2FfrSnk6oLwNlU8jqIEFLbtr6SOc8iEeQvUEcAbNa9//qmrCNZ25DHmymhaWqaEA
n5OkdjJ6r9dl1ZlxgZwKv5Oy+fjn1+rrsxgtSrk47efbhkthgtcXKD61rNP7WHe7
/5/nyim9lnH9jPrTQKl1gumnLk6I/njh1bLENCT3NpNFBgOD3rMfTiY0gpijEowZ
j6JM+GpNONf6JT92FN9LMUsy1XDNeXyI4ZCdjuxlHHD0IHW2UO8vZ904OAAEy94p
92zgvYb+P0zuYH/pf4PHxJlUn2Uvc4LtscF6GG/ILRESlCqp2P5YzJK5rsP7f0Bc
unF7QFmM6PMmRw4gnB7+TJp/MjiC4jm1CEx+wnXwVcO6uMQRvmd7FONCzh8TLPMB
FKO5FYNRtx0HdgxWrP+hvtQaP/vdLpb/k/3e21PjQLcd6ymrusbZ/RwW9bbUZdlu
BN3NP1hIe2jiSuHK+P3jAhXpyAQg0rmY57o9rlKSdoPomAUED/wc7Y80SzjM3opO
w6XYeVAAi8RYUEp1OiiJI+byet08a00CUMWlPSY/rykEbbmBHunYDoYSeFqsCZdq
7ujs/BZcWFQ0UTOfistpwSnK7kxCplm432VFK/EU6Ex1ni6dFAh7Hu80VzsjVnuw
m7mXeZQdLnNrMO+kcc/Wy3zX//mkQJ3O7CgCK74dNrVF1uB/1O38Qow7EDAEXE7V
YIQrCpA5WBNXY34Vu0zWqKF+Br5Aitl5Hk0jCdSNdnXUuhE5w4raz7WBKkVBGLER
p4sTIE9m0q4cfUdNQ4H11CVjKNRyJno6PNJ37AdAuXy4/BNDUAyLnwuAX+crvwKK
mFN8QXesWj+GOM4K2b/U03tTyHiCBHKq2+6WFKybiyLasz4ZKanQed3ZFByaX4d3
C7SSJu9PdrxZStLPg/ZcUax4sRTjeJ41nKFXavFqBLONpOp5CXCC/Sfhm5fRWu4X
WYfeZkvcnzV1qch2oImh9R+X5UyPRjArXnV3OpGYAga4MdxEH4aVckQQ5mxDIKaQ
24VWLHol7eHUQhaohEAPoBV4JpPCZKO+o7wSVbHKqNk0i0Xu65f11Q9IfnCMlPZ0
BvmPL17j37D3+UpMY5HNpo5fsMqg6vEz1sDh5ZqaUtFUOW9ie2HcQEZSbQ9Yk+eT
Bwxr81n1TvrL9RE0fDrxl9Byqtkh5K8T/F9HFTOS4OP+sicSOH7zRTqwSYMhOOPA
P94/5JtJtzf6T4IO4xY/qw2fpYAFo5A/MCk428hGA5cdaQ0k/cEXnv7alj/lJKuf
hTU7zryYcN2ubG0NPEwee1G474GzE3q4t0HyYMYZA54X+/Y1TMGqZoOGOLbg2DRy
7OOt8WQCB7VXEGX5ojVbqTTIbeiBHj9oIPGg5CxX35GCotie+4eS5vBXrnjYSF+p
50RiFDQ1z3Fa20HSLd5F0rgHZKcO2F8OIOxhB4QhCmMd1lXl+pQS1yAHGqQ4r9zU
IBY3QMoZ3y06xk7TIfAi4A9baIFmAlUKvNZXAPERe/hq2214Gdbyy5lZ4mDz9wc2
s9+jsn8WlDTD7uSiFePOm4ag67B8vuRMLWx+qy6MzM6fdeeHWIapU5SXKCNDJXyA
Gh9xK/ldV8Bwa/m3tsqe79S9n0lFzUgNEVLBNfSEYknBpzjDNkC0ILyR+UTUdR8/
sYAFIqn4HsOPRLqtal0/BNHT/sqLa+3hwLj6fLaUb4ckYWdOnXibIkK5xibhU3XV
9hSyM8+Vj5OOg7CM4JL5SNhdVFSnzReRRddSgACXM/TbxNMy8q+mheM9WKY2OlA0
inbQ17jWBeqEPhsJ2SZMPBE3k5uBEbwH36rkYSGaJuhhNG02S6MuWdnqO1hbvt6r
e9wAniP8STHhubO8Dgv4prZ4PnJW6LHTMHINGlmuBGWGF6LuIebWIiDbBXXPZq4f
f8ys4g7ZUVnNWiWUwoD/6ppvWF1Q4F8/YSJJv5NQ9OSdX9AJ7k4JZoCGRfJW8WOS
Mn+ANyqN4LYsViJEEHBPlgEHcPjHStMCmrv8EUI/cjzXNbaVWTS8Q5UBdnhCIamE
PPMxuZCb18z9O28iUmXpb7O8/gsCFs6IvSDqhZusK+NQ/qgRh3d8F3Hm7Ti+NkQU
vrGVYPlBHdO/WaGlo1b0O+WUMMiukoHXFu5wV0/gR/6n4ZgPT3JjK8T5rh9Hu8do
YiprHOrU3ZCkXMgLW8zmAfuZjtam9XsDOcP418Qs0S4iHf90QCuMOlmwDlkR+K1+
jYj8mu/meYuIOSyZIZuSuOWVR2xxo2l7IEeEU4VoBYjbADktnSQZadyvogVpEshB
WM3ndFqplwxHPyjMnLGUWsmRf7j8Bk/No51zBhwKE38JL5GoF5R2l+hRghk44/5/
T1C0imMBTvPVS++vF+GoGfiAe8n3o+qijl08LuKxUQrN2zi+P7WvwkTJQs61vrfS
TjdsP6REOlrXvh8aRzD/YyY7aKRJVXZFO88wR+GMr6QZm67c49RZiC9KRLxxrFAF
0FQMEDCaU2vVzxbWCKXVT353xS34n/vE5rUZCMtJIAcgaK8LYvTJZJWokzvvZ+GO
xHId2FliWJdHAPDGihejC0QJpp8vSl67F0G/kWNrXd3ogMgHwIAzDnGfTXe0xIoW
ecYT15hsE9CUrun45FobCK3XO1PGh2BYzWeQg3giMBOqBsnGFWeohJltwAVX3CZM
RchZeUXtmg5Xg9/QfInxle5MbOHAwjGueM8kBYze6gP5TinQkemFZZzS7/2qZCPu
pIjisB7kEh5Aj4Tznl44bAP8JsdqGvgXCEL6ACIuNhjiYVULigWw8nz79icJsXCM
lUPDPgQNagSJyuUSjXXwxKJABEEREEF8+kCfdSzPRIdqRYC/FxvvgnojkoWvlIWl
YdkqasWv8T9Xeq/GdesX7Ro2kY4yVOONe5GJGiN/pBPu1Cwq+jPt/hsL9sl8W0lQ
+9OMMdpZGJ8Pz30G+1yIFIpkhyikEVJlZaFat47Lzy3ccpx+NKYPh6R4FZhReipj
1HtSFNPUV45O7qXy0B/WKAyBcHAZd3CEuRclyBoYzdeotBnlRhUTiWuIV2KTnm6j
o3CYMbh+cHVo1xofs8kj35BP+SVgazZamVO5fnu+uhEoyD7sUtthSn0G41fIOrLG
Tn4DKPXtGYX8KkQX03czbDNd8eTL9YGg2Psmq+aPnSOSS5TJ0f/wnIBwCz3VAsaP
BX5DKPYSzDp0Dz+/7iDoMCLc0Gs4qLNf3nO1LrD/7MSoiQX6S0AhsT08Zhiy8lll
oO06cF+xqhykCjf9bW1ufDDP2N3/7pfZURKql2hAiOeej+b9ZoAB7EqbOdE3tqmo
gTZqGPVW0tpK+2IbNbCnibp0EeVztFwsXc/7bDI3SSjYIOO0S/sJOfR2AQZIYLAd
BAqp7UaYpFZcMrcU66OgogrQTKsOq6NsNz9ihMwdHGlkGx5I+vmWOu/GhXKbvKQO
YuI5MKb/S1DdW7sRhwyilfV5zZ+q8cvFxZcUrCCGoP5KdMmJBGucdRUiu8zVZxOs
XtZOZ1BEUiZ/2Q4ImnzUV7bhmInutFkvdLcQwfUqQiwhWtdKZB/F2Y7qFXImxpGU
GGmyw37NZoKOFtntKBFPyiz+XQ56/t3WYTFMatevhFggAJwysFmE5eAcN9pxec6D
G387+mTXZOQtXTyDFMwjPFf0W8pAazS+9jG2bC9WEgJLlpWuXc6ieSy60E1LqspO
hzFSk71lvZJNYkDklpnV7RhXJ1gTGAaFBuBonxDXqlelZ/LhD4s3LRsgM1urCK3E
faZ4g8a8C17HR5435dZMT+Ea1dlsUenyEoN93+rnbdWWiuNRq+BOR4z1Il6kA1eR
29n/eyUo/x+esMA4Je8QlGu+061PW6CMR69/De4GL0LnT3HMYqUgpeLapBi7Y7Oh
7koTM+BRIJA4Wnzv5yCI/AKSwFYtIL/49MUDxniVGr3OjFQNLEruv2s7TJpbGdfO
6sgfQ+5+lwspc7dpOeBsndsgCjqqcRs45CDu4MrWaiF5wLS7/IyJle7zsXIie6xU
dsCMMywolZYsYG3j8dlk7MidU6O6nXLQXulFlT+wZlU7/ZCceu+Ajv85kM7pQRtJ
qvw4l/GDvcUVqj2zg+oHRQNUXGw8EHZCiktzk4cqEckMHyLV/MR+g0ZG1YiSi21y
W/96gRu/kq6Dj+N2xntOuKBVxDeFYGfEWhgGhjkgp4RE76DggpKfTRel2J8m4+Cl
DGfxce88f1wJmxBqu/akr3tK3u9ubT+YkBlz4+hI1k1gdXB9r2HH5GZj1yON9pgF
bSWqf8Vvsop0p2UncQ0cQM4i9gJy5mkeLQn3BR2AZ0AyGdDI5/l/yHJZjQKLViKO
V0AsW3XJ9tqohRVZR/s7WOZmf/A7O1LiMOMe7hD5LLF1FlnwNC5AowNxVolXiLVJ
bE9eJsT8TYE0YMg7e7pB0ukPn+7nLHUG9IF/FKKl4pq/x4TR6eULCxooYMmAybdF
rOvodgANBLx/IM5CvkJUuZU4qUHH3dkZRpDJRkUKSmm6LbUGhRtyDHONuR2/cnQP
uPu3/ijsGdFx/gYq+xu0lTXQMHMuDifFUY1USTc7eTtUcssFF5M07PgYAhvmICnU
pXWXZbP30Y9982XuJX0c1/JVPVAiQElnQ+ogOfHdB0ugcKEsEn6yMUE2SS4qWTeA
oZbP2FtrEYdvjoi1wJRFyrK/UkOcyPZXbBIRR/ew9abQGdHgYBHfSOxk5peTLPfD
4Yic9b+ME7d5L47UNZ9Lqjtz2na4hXJlllpQi2AnXozFSR531ntY9gI/Rr7Cgvr4
UL1oto9Z3y0BapuV11pUr3oqlXqLhPRjihQ9W2fT1ER9iLWHJ9YpJn2E/LhaULcv
jWVM9nQ2jfI2NDt9U9HCjM4mHoBxvvdlLE2K7AorsivKqh0/CzOPe7ecCkqulauK
XqfWKCYZJ10rsOtsSL+38j8GICgNSfLYbTwLAsjwRBZdfcitMXA/Sny/key5aWMp
xDPCNKs8v7Pcz/ysHp0e400xm53qYtLW8IIiCg3mNOLCV0cZWi2iiEKDSaf2mXVn
TAkVLeFIci1h9nGdz/gr88ubKFzT2uw3HdDr8V7GnWrIn8ri0sKbm3f5TLDitKml
sqb/VgX9j87ZnBZhCDRl1xOS6TvgxrqZ4B49gb4bo3akVLGHjhdJlUIFcygGSrrB
YLFgdmRmXkrE2ORk5uIPVz1ReRNXgO+nPiGQkBRb60sdCZCr3HfRrjHVdP5tYTDb
MpszbEfroOOUsA/jdEFJQZ2ohzctAagorohZz9Z7TUEtHktPfG7u8PSgcWb6q060
RofnFNuSi40f0X9Ep/8K8yjmqsH5K0FA7zlSopy3BVuTwTKo3nZ2TM2L4khD3pZd
/b7mAy46rMSSzXh+cTXLlz5UTXj6xctNF68+DibDIYV9b6zqpPmGBENKSDC03VBh
y1Lpac6BDWcMV7T8h84E1vATmQI8uH0kKzj4lxZbDSMfHGAKNvrq8sgZxGNTwCaP
XhDwYOI+/0WInSYiuHl39hFpPBRjsaiZ3/iqbS92LTiM8uHYmSzK/eqgEBdlcrpy
WJ1QwjyFDCLkkI4BdrHo1RR17MQFUFG8z/mDbU3+rCFbOA9yMCBRXDS+epT9CT26
2tk20BSAdszLT5UuF0BiXVy01RaB6gf1adzXXetITeGvNX8+Y3olAgSy7cKHIHAn
Cd+EmyQdkpk5Rf1IR7m/9f+Ou7MxGjkMTx3sfRKBPSrv1W4/Askp277tq7yK7UAw
tK8n+G7S8CyemSdIn8+C6RV6jBKu7W6FP9VvvlbR/5aWraMJOJXnxFjoHD12Dy5Q
6X0URuYspT3kXlK8OgDNRYDT5dJNRLdvjow3+Hb2N9cT+tXvcTMPTSMPv9HWWNLE
nZ48bTqgqoFnmDfzT52x4itJqZfahLm6yzPMNLya8ERbIgQYkDSl8c/jSG3zXDiW
9dNc0llPH6F8Yyob4m4ehwmNJ0KLFI2I5oV9FBHi9qm/r7+tLyyh48MkYAnnPiUh
LNQ1ruhudvOHGH9P9PkebDNKHqoJ834QohURzQwuxOi3/hN99KCa/cxu6AiMO+X/
hLMujdSrVmMYxEhU6wllP+kGtbX4JAPxMVJ0OAdfpURZ0V//uf1fK1t8gBH4I3fH
iiiykE9hG8zSpXHAj5cmYhXtUsKwOt1l4r3LcYTYCC8s+JM3A9AVu22UqWlwAVOO
nT7f1cdqjNcLTj0aadcMOz1UOZMwqTpQ2VOXcZuBjHCnsFu6MI26nsAeQnT3GoBT
COkGESEKWgiQqZw1WY/EFt2gadu0IPnuyn5CXA0R5MxzGPl9OQ7tjGUfmSWQtNHu
+mYSmUEHSRVUmpdYNOuZi7J+xDpZvGo3EJkdPG0bYPIrTHMVzpdRon/ScCuvw9o3
eEx3s2no1Z3/4Mk9qCU5QlbDcYQ8GKtjdO5durvwTxYc0mMpD5QIJf/JlzcJW1XL
MCrhrBL/ZlfMNUS/sao707ctIBf+mGxPJDHxchE1fDheQk+9My9a2mUaYikn9pcL
Zkl97eEfNHGq0ArNo0nyN1x7hLmrhM3oMZwHd39ZnSU4ZvulVLonYltgIrY5qnZ2
lJnkNf2Gz3Dp8Uq5EGCwDxvFj2b/kR82GOrRrae5hqRLfH9q1ESnRvfK5YeEl98T
Jqs/hYf9s6txuaWi8IucHnwjgmuODcvCV8oXGuzrJWo+nThwaN5Z0PXGd2c82EKI
mCFYJeDJUMBVIupXq1GvEsgMriDpnyrQMdHSgxAMBWLYfkTfc8CaCHaIi3/kGrti
h6lMlxVO/UzeeTcy3Wss19uY8J2cbOcfBL3Au7x7kPAOjmoyrJCoHgWW4Bpfj/GD
VJ0RI8+YkiyRIS4R4GI4lyOd6TUsuA7lZDV5938HIySLZ/PqWS70teZf4yLI0AjF
ePceKAgcKF9uqAzK85MPVZapz4dJX1kyvNG8OZrHUPcPHdMjBJLqRnTLxkvzthlZ
s/8GLNweKYehFvfxWmbfjjdQKzMBm3MGW9gOWJqcfvk=
`protect END_PROTECTED