-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
IDWtstlgxmH77jq5WJOucUsOpmjn3YavxCWpoQmEDfrpPK7YoLr8gbwcWPIlzOl/
9Pn86h6g9fSU+spJfeQCEt3rwaW9U3lUv84SDTelmauev7AwKGBWslWA2Xsa9Ksy
u+rV5UqjmJ7Vx2dtG8dDQ24EvCQa/8hc8NM8ji3wJjc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5392)
`protect data_block
psocJTU2e4lKvmQtQSq9oopRy3NYNlG56kSXngCJa2JBSFEeVx/DFIARMORxVEE7
1cUf10aIN7TPq4xMcdB8T1/oEqHvRtvnn6wgAV/JTjF3jRbLLldhaa5XefcgTa/B
IQ6xt84bwnYo1FJZuiTsvsphjjd1L4CJ7/xMOlCCQfXZ/I4KbOOMlZ2e5yA51EI5
YcR59D0TkhivrfJhxYT0UzcFwNNoppJU9ftoNj7ThTxEia9cu8ECrzOjXRStWCXO
EfEGpk5+pwFoI6yf5a0MfXZDdHnxOztpkdZxEYGtTeuaU5tjyHyu4y6COAZT1AHY
5Cx07Rbd7WHROlYVNQrNzpO91DDNkPaW4X4ii9U2dm++/ULcm2nOwaMAMIpeMz1k
kOcnEpL2c+2EMgPFAwPuquCE2Ou0gYd/bl1xTGJQ6fQ0JYw2ICGG567GTGQ8Kh4q
kV1k/rtft3jUkWV8GtL2xUpV3ZMEQLvM7jt9MYRn18CRW5FqOm1XCfG2CKzGKD2l
RBlunsVzMdRIZyBeYZYzTDEcfCXbcadXGrfgbQEMcZWJWcc/V/lKop9BpqRQ30tJ
ajUxjmNVfwQTZnATX7kVMQhDBWqxpvo3QaKfL8Aspg2+GiyWX02O/Sl/5qoXNiVr
SqMhBUT2ooTscq20zpGwEcKgwjyutASgcKRAI6/SSZC7kfosVgxMgSs30pgDQMqY
UMcPWwVet5cNZdr3Dq5nmHnXDJxWwqit1SaPgEe8BWWXw0qOurJ8wVdro2VTkfaP
0b5+9Jh4nsKFBLi2WByv4FCJquoFCL9VAI4YYRTGDPfi4LFZNQW1C6ibHqNRZDfa
qjLPZT1o8pZCS+mMRHcx/M1V7CdbeShjDIkOTOLUKk3u2WfI7bDSYtLiKHa8+WBh
yChRC81oZdEj8OAoG80BYu0XSBlD9rz0eThhKMnYaPvyVgu6JVYgijKJEvvr10FF
dHEb41Xd0vJN+Qj0EJiUgmPi4ON5n1jVkH32Tkh7oHeAxiTolQZsPGoVzWy4TF5e
u45rBbKiiOvCrdNZ/UV0VJiCXNmMNC5bplBJtfvxBxYaY627xMAsLk2VqNIXsEHg
y0MQR1rZMvysZZkYxOS7IpmfeUr/zNlj+PXxIRlY9Op0jBOkUtqQr7B1iuoUnD3N
RyjIDhMbXwBWiiUdRDjnVPnT/Z+2oLiyLvxPLWCsvXD+OpGLkKgFnv94u+3GN7qp
QvFtinLmWQz7lF2jt5XF2bBoTnwy4jIcEq3uc5LAMhiGUt/3grLh0RaNmsBZ1Sey
+mvzIfjgt+2M6cUj5M866bdJFgTQuml6V0pAq+1lJ3Lks54wZ8FDEW/NEKt8xhBe
geH9+2ZEcOFo7wOS+rmCWYzBUZf1cBaJxR7P1sPKbuY6tTddlGte9OwMGI7bWg3C
q3R0Ne/wJ20AxTK/s9HJtrHebufEOuhRMiRM8zzYCUTHH+LoCXVseRFB4eWJcPhD
bi5fM7vMP0NiJshlVU90UIsjxvLw11g/SQsK7U7G9USHLCQOyc4LIWiSPD2PdgdL
oUKIFqcYayiZJNX/8lEimdA9voFVWdDysPZRifutxjvuEJc8+tT/oZrtoR4PQSAy
OBIhd8PcJ//yZk9mhRNC2qnJB30hYr3VdlhXY2PfhEjcniqUi6RTnzUsNc0xZorc
qTOs2uFcCD2JqXju2r9I6rvXpLqm5wGCaFZwTeGOaypR8Oga+YmZNmnP2tx2ZwFP
XGGoIYxsaxHRphOF6HLQUSyqXAvCULfc65obtMjQiYf9KZAUaWgAuirAabeuakT9
ImAtAfBhEPadiguquAcIcuyx54td2eOLfZ4y7sfczAwm/GQO9zyuo276Kq2VnDL4
QoYV+/rfd0ya1a5TAqZHXjcqvnigqM0F+th6ZKYB8pZr1e1GQFqHjykTUGrWYoN1
q0py+lCxsI5xXMPh76Ka8FyDFhIxCMa+rx1mBRsZLhTx3SwO/p9BCmjNZKW78G2D
SrU9eisoi5Shp3ZEk+/qXM0A8YKv+wrOPFABxnsUP2hzXcNKmECmHBdV0GD6JD3j
9JXsEbd+sj7ys/YJ9j66HmbIuxmyALgmCWKJitxauDj6lddUkzuRfkcUMOX1psKU
sU58bphp5F4FyADvZ+sP7FXgc/ex3D7I9+JbtFPCv/+Z1/Uijbg7KDNjrM95iO9Q
51anht3sWljLdogq9aSjIYzCiT3XAVxkLLt9hQfaNtOhBehs1uM2qGQFuxQ6PfVG
x0uM5hSxNktzZt94KPmiQKy8932XTqCJIEbklBcVCVxftcQtPAPUj+ydqUondSxX
YFNE/zsjXW2LIwmcX+3cKCVTjFIFEEp1Kk8/2jvdIYM6QMwIKD2kK9VKxAFFeCKw
Uqy1bHn07F6kk6NkE75eqKalLGCPBFGfHqkekkzxgesxww1hmgZ55FhJFrloFHAk
gq33D6HzehyOTxuH+td7MievCTjDnFKWtguYm9vU1KYvZb98m8ywhWOrv6vqGfd9
oY0MAOHUu7Gd+9vM722T8JD2SK040PFLVLj9uq5RjZutaU/9kPqFyafHrLS5Myau
sEGZ6UB2PHJLCx7quisfru7Hc7IYi35E8xqE3UHagwaQFCVdainM4Qcq397c7r5R
TlPAsWc3cw+ayWVv6X4zSemH7Tp8r5iOrkB4MpVEuwpPg12eTzsPat4EVisIfMFY
s2/ml1Zn7yzuLRZOcpqHaeGtG7RuxZGOsTigIjnFUMoWMzKNkLMX5KhKDDavHmaD
arV6FAtGaEa7rd35U6nbsIdRnxqu8BaGBUQzGXpYVBtV49yB5WUI4vN3mgrEKBXF
cmLtzKl6GZ6l8epJPKVh7FGmJO/xGwjHDqtqPgBG1ousyfVSlRUHLwA55IDR2H+F
JKP7Kdh2ycPCAqfGXfFk4h9yW7E+JtITIPEfEjTr0OcdvblcIUDE2RkSxhfFnMfU
G8b3EqKbsusoK6R2kAznAhVv3KUrb9eOC0sWOrbXAZYyuun0F3UqvH0zmyFc6c81
4fgkCHWv4uSRa2YSYgHiEzAiqwWsR3maKsaqkoo0BN4frT62+o38nIMthjZ1MZTQ
5JTqA9EdWCRWQi2LwAlrtRvpWkS1NlwEeT8LK/3EJpwy0HSnRzA1fi/Wz6cIxFxC
QrPF5JtigrOqQFQUMarcsETnUig9bZ6paNFQznw9f7nlkFDkni+r4txdMInlLHSz
hbssoZtMYIxlQUnknCDJyb55qwBS4JmmRE9DjmR37o4UKke8cn3R12zFQPRKVlHy
aQpzpa077EWA9lZLpfOzQws1iuyY6dggHqkUC8OaSX6RVbckOBlDupmLND2kK/Jg
yPRYlKEeSdzLABPoOsuNCXUR+os8cXCrWReOEKqaxDniwPSRPk+ruhri3vQF1EIs
7/TOzy7xWvziBCSxIvdla/dDK6uVVjRgFG09PBv91Uv7U3STERlO1l8SNR951YYq
BHraVAGHUJ1Q7FF2WEt32Q29XRIioWnAz7qdUNuVZxpxv32pleEmflJZPL2HPB2O
mmUyU61pIuFG5kQDb6fTBQF56C9OsuKTDbx+mCH9+CatTI9aGFWmKtexADTu5brE
jiA17PnFRGcfwrBxTIt/1AU3CM0VItbiZ5HHu1aMYNGsr4a64gbQ2jUvM+lczxaq
KhacUcQNAoB8uI6ICkE/EolhBysYZCUtyV8cA1bNTGX/sZv40+7R8Rye9NKVtZuF
zIyarZoS8jeEB1E4nmlLs4LqM1zmqd26d9Rp9NkjG0m3MpbcVBJZMdpRn1kFRkz2
fOq4kTU0Xm4LHiEs2Ti9igWTeeEAFJDyrQHqdbTE/ckzKbUKa0vEYDJyBLu0kDc+
VlS/qAEwxiw7kuLDPOWaWUmNYUAHuO3lQJdsHB9Umvj40tvNuRQj3y3MZutOEdzd
P/foAktTasM3zbB/W5GeXFMO4GlrbbaHjgOA5S4qljLnaqFGjOQErwhBfeu3nyXp
OXQRa+bMBN2LIt6j2nMk6/RUiAJg5qUYuICc5UAsjqruIUIx4XyhrHrBGEWW6cJ0
YqL8e+emjwOfdrFw18Fri/VuWSAMxidurbo7ogVrW1ijInrnJixA8HQJhrAE/lCA
6jFF/XRD8lLcYTRY4Pf+RLWFmE5yShHM2YVQb7G5qCr8bzluzkk9mcYrDWwQnGX3
+e120Ch39g6+pyGNHcy+pUjMrI+Hxmmqth4idKsFQxKEZHVjlLoZdevww+OEWTHf
qepiXdEzbZXjOITZR9R5VfpkPSd89jhAYeyDUeFHIPlbaCx22EPn7bnN7UEZRtgT
j5gQr8pkdWFtYPBUy/2Ma/wEsLViNVMEW5tHflUbpZX1zr6sPA27SE28K/XnzLb+
ihY2vnYalArpJ2Fbg4tUPE6WyasX5EZo4Cp4rFloN+ZVL01q91MYt9hJj7Qn/MJU
H5PsRRiQ/Ms95SlowpBQlUmctQBjupwZD5eYkpA1njysr/4kcGJpnhsuKKBdews1
Odj4GEwEFZQxD7WqghyGj3mRN6hM1tc6EBumDQ+0Iu4LM7tmrTFi/E+CkToMFTJC
/XoOpNKSU/GV1zWs7Atoy1GFTXiGS7w7zBARtvt76rE0rAVK2jNxoaOEOxfPYI3L
GoFdaaOvbYiOI89Vq6a7ph1CpQDhOGeFKXjXNTQrWZJ3IhV78qN5ODyyaEC/oaWq
32PjwwQCvYFuD2MoTzxwtk0RGHbEnR8XjD/EGpAoZpPoGGerzdf0DKcd8jsk1wI4
LioqQfXmhgIuoNlVIfWOQrWy/8hsQvdOPIwO7A9RdFdgHAfg+CCPea2zVTl3OWQR
usMJ0SSUePM6oAzvIVOJtM/INpmfKFjNy4ytDoTOCI4NJ/0PR0LcdgmP2QD2fxQe
Sx93ag/W6sDvkKY5bqzi1fe6tuq7K1ApGtVQPBJ4XJ/chvzY2J4DH6M9Ex4xDYMj
bTP9nQY7eMZd46LxXlKfEIO+xn/R1IBf+OZfLxkVAeKM35NrxWD5mcrj26k9M+Qv
Zoy65t2Te2nldPbtAPNrrkZOx071pEfTtSz9wcAK3GXebLeXHi2Tx4i4+4CShK/d
UlM0PkVR/EuPGkrRQkNATOnDm/w5F8CwG0ljtRENvsgGHMdU9GbfNHaMY2LSr/wm
oUXDXzO8PLrvIVdFuRpdfRPM4dZYwIcA+ulOyuU7XlgOU3u5dX6SUTTnHqG9FKke
p6iYqkbPRDaz5N6T1vThCeN8kbczGylPmPFEBauZqJj+6N+XPjEbJ926G+BzvXy8
Ar42NK3DaY7ez8IZl+uuKcgV7+OyXK0qYpTKndmEjnhI2xmelkOCWHJ9RK3gjymg
863TNYMfw2i8l6dU8h5oKj/McZqIxtlumh7oTV5JMVXyXyshDW1+ivtx2OAGPtdB
VvNL1jPdayS9ejfwk339cDJFpVw1Pv5pMM5dv6osthuSYAxfWflJbIu+HgvpDOuI
oyiTmjj6NTd6iBSIDwbqVRii3j9pQvWqz2aYfGKv3V/Jywl8bi+hCP0tFuqr8Bf+
BWa+r4S1GAtQ7j+RUqNsxNMbtn5cphC3CLKeueXPRWUR6GSOzCPdAUI21s6mMBrX
z2hVIFgGH6GRhRszh5OyF0/jS1DxA3+IVoqfbO2xhD6xMlfoo+x0WtthQI7F+0qY
26gwagDhYY7J+zeZjBeFJE7zplmuHL6TUmtE0AlUjNIKMtlBNEtVPyUaWmam6ICo
U5ZEyRSvKqkoDSrvhM05CukhtIAcrubXQ+506pQaZS6BC/vMqgaPqLEkHyfuyxzn
UCtATvjoU4ICzAxrjFl+YUYElxSmor0AkHH5qfXkUxoKGAiW3FLdDbRVeH6K1X9K
RZq/fJ3uCTn+m4e0cC+U8rQGq1CeixcB9lFpjmp1/ueRo066wL/U9dSXaEi3d11j
eeMiDWEsPR+qBL4MB/AgEAJGyfAuRPR3b5sYCqaHU01mM3BzmdqV17ZlBbnWE8Wh
iu/UmBhDoPRfTzgexkX5Xh4qDReXOWRARhO4dKMLKiLLYi5zOswK64V2pzDy3F7L
/UY6tV02OSZaJ2Vr+CWV5CGFejNDZWjK2BiDAxBx3RGgF3vo1KRrQAO5frIpTO4H
DlMdQOo/8aWbK6sz9JvZbuHyYw047guzazjT3H3MFwE1gE41p9SzYgmR+I1PmOXa
w4JF1hSaAmqKIov6vEJeWcgmF0artV4T2CV0uv78GlWhaQGO3q4Lj1g09fz6+ih3
ih4mCdiJvJLv0BYk4WnWF77+BR/vVjHYlgpACuBkfG3XFIz2pBtEYl9Yxt2gSkZw
iLmj4oTo5Id4GMpg4YSMSylj1/l4cX4dMd7wijDAUC6lVVR0hocZQkK/ZLmZPBAP
LpqbCqwkmXje7xvwAErTOJfbqCTMcJru0zE2u86suQLoYEXIIRuQJIx7Hh3FmZdE
M2/ydhHgwktvJ+w2sTr0wJFqOVESX/ufMKyMMwxjg5w+ZimGEjBahHiGTrlL97JB
4RYMVTumW1GgyiLH+NX2JIvry3Y9O1hWDTJvyrtK+y9K9EBzWPZHsHCPjAbx6wBE
SJ0DAEwpzJDNwD6oZQD9gACxCE27R+2pJKoMHo5dPxgomGQs/k9BuWnXVxZVIvTW
zjmKv2LwEu7z/eUqS0Pj/r9R2eiuS435RwVzV7ZkARRmpp3tsmCuol8LspD1+twA
o8UDHlEgtPGBEPAUhS+DJUzKw/KmYLdepPIefcvkxPvUmVZDncl2P95Zdc6GXiXn
yLCOSQk/RY6y8T1DyNmQwZ70H9JqbNM4yc9HWwsASrZQz2ghI+n30JMi5HBmFmj9
T3UGdFLq3ApDhw3GzdJ0gd6qh6JKZNW8vGK0xBVJWhV8ZkVRycUBCoZSVi2F0uW4
UeZTuB718G76XQ+wSJmteCnnAOMIHlPN56nhb94qqOkfStiXqNb+3rkYhem/okwZ
u7v3O+zH+X6Ezw41CsQUuYJo7B/nsV1iYP/E566E7BAnQgRvPeGO4hYfJMkIQfKL
yuJF/xcJIysjG4InFqbyNvcOoqv8GFMozsqLmbGF10gEqdaftsYVmLJNuvZG0kwa
7aLX6SHsvUC3Mvh3FPLp72RsnyHIUAq19UemwL6QGOWfbQTfyil0fWQp+SpnGAj3
9fcv1cFxQCEfct2m19WejkrSh/XNDbRxWmOTVBUbP6qyEz1DpnRYklpvT11gCpgK
B25b0VirduoAyCuI9XQUNA==
`protect end_protected
