-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WAtgRtu40fHzZaiaqDIJd9vdZSaEhHqFYRuXeMPDP9IphP8aZm5e8ENGyveUZnTs4t93yTwzblOo
mlvoDfv/r0g68S7pPyfr91UCi1BEyB9Rj7qeuiMKEnjkHklI7egMR7fJGjkHj8lttMAxXG2khR0H
xTwsuJ3CUcxwaKjCi6LnVfOsnSiIFisvBSigYPMhw220q+a2gus/TnBKH5CuV5+dTaCtGH+05aDr
85r9+pwFD/AkqOUn/a/NMCUj3xX3ZRp5PDbnC8ORz7QK93rsxRSUn9pz2sUI6/NzUGxE6igHpneV
rj1FxMxrod08CEj5BqEw7pmPZlxuFOPzPw6QKQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10688)
`protect data_block
Z1cJ7wTR75/zQzennkhMB0sbgFVHCv8mF/ar7ngHLiwmBw2ooWCV5twzb9ZGiSOlo9U72RWIRisi
LOnTS06RaFp11gHVbGw9rQhXK67kusT/4I5M4IdroYN5c/T6JQhB3030vcF5+BqQnP1EcCCC2Ljw
mrqdROXxDfglwVyMAnDPb0PLljPwt7AcGm08oKnwprlGq717rx15QKInXD3g6J0nCCSoiQxLtewE
yoV7c0BK8CB0lsrZzHrxlXi2+Qjw6ncJKGNJiWOwHduRDRQK06NzGFt8AZ8SY71jnQUj5w0a5p4R
WLMasASYWSBJBmHoDWgD31GCejhiavzD1luZwFEjC2H3OwmbIhYpKQaWCiAALxW/9gX6izr9R/I9
TgF4ULjKetxHIfVMxm+SjqzPoD/fRHzGcYk+RgPjjPNcDhvO2CrYb7HaxV7xCfDdJXpOd2aVw5v4
Ay2F2Dh+AFaq4gSlL/icDs3cfjhVnph26U4bFgHcbyrdu2LblzboMBm/BmYjb7yTJEFuiCFQ6wNV
VAE9KcNV1PmwnwJ8h2PkNREHkAdhUMwwi6WSXuC/+FbwYbGtvWp/tzgCFwTalAJ5rYJ7Tn5mASBU
9eOMOumAqv5tohCfQ+1LD45IRZCPJS2tuUw5Do9SU6vlc2j77DA43AkgPr3bh6L2rNv41o3PlKtG
MhuOL5fA2abpAQ6Vinhw2hKru83CgQ16wTmCgTxfDQ1gQIttL2OgqJAehCU0A+AwAsyPsOa++61e
mg/FzeCBX1QpTbSBNlwYa2P/LztkLg/6k5TPhTfw+EoLGecrBBvGFtYR19RM9g1U0HdaZXiF76L3
LpKAeCYmn3f9YOds7SL/CtnBGTJcSfEEFhzANNNBbG+VgOWI8EKKQNVZaN+CtRaDIG6oyTFWNiDk
4WpHXPMuBbmiU9lHzr1QjCzP2Wqt/crgY/lTgvIS2fhplg1sM33fa3Ukxm8giG9ZgA3YzgcmCehV
arYqUGsN4CkuQk4FkMUBaTySjlhSp7iGtYxO5+1DaFI6DXpaoPr5kumaIP4r816L3K5KkNFWEIPo
GAuyLSifo6Z4HEuKfN5vDERWWfBIckRa25nOytPvgdUrlvtLkkul8t9s6Xj37VVlwlefVOettAnG
nM6BbsM/AtPALTdIVXTyOaWICCeucU6yrx6YbkvUzlw3j5wU7thc7mH0JyqRB3Z4q7vMd2PQLo0G
ISQ1TTu9pivXGrz7j+yzc4wkzIcD6aRRV65naE1s9Fu1/w0XoW3m8HBKJEB8VpQuaBHpdVqUqiJl
jP8BFnvUmpbfEdpMwUrl1+A2K62Nk5yBvh6HQzqVyNEBEjas6Ix7+XU2CaGrQ9OpJuBukWJuVa0t
4P1SBTMqNJMy+e54x5mVn4xfatAORlUENJghBg7kE4XOoVS7metUm2BGAegvvg/4DE9Ner0EBmj+
AHAxEBeykGtrXKvbpzp/mGHi/HPdi4nJ4PR/ADdW3N+oPD4LdX77YApdllfeROmdqpE6TeEpiCll
H26GN5ku5tUauMlZ2fRpQ5BIdwfc84JpHgGmXjRxf+jR5Z8EtuBV2RYsc6UOXm49mDnZOcuQHBYP
A0MLeAhfWl/FlatafvQ/a9GUh+gs0AtHLIlDfUBXHkBoLqO3l3a2FT4YJf6xfRNRsR03xwHLBNuH
aMn3VqGpOEEglmnch5SOa+VPdZIiR5QMcx1RRP3ysSTJg1vVrLMqXZK8lVQ5mIUcWYQq7KW2UtGk
Vm6Zaoh183cRrw5RsxnwllLZSt2t913gdA2Avtj2qyS0GYoWvS1rDMsVt9ubSKTWnVim37Y9oPzx
Lv9QyG51wKTzjzUi0E3/fL5H3drbNfLM1jGh2EYwpgEK4Gq0RxTmQO3KE7O74WZFn4GOucvbQ5na
ESf9kGtUU2aaxRwQN04vD+GyvWgu5xFcrLTi1UQpXJRXNJMgUOdkh9zy2/+V9bBiVWQzabeDtj9J
mDZp/I8Z8R6nPH0HIftagqWJJwkAKDuFG6M4Zuc3p57hOg172jkpjizKljTZ+gdTdspY5t7BgC9d
j2YzrZ/T+7xNGQVP06DUh8fEk08L/5fhWg0oyrNAS9hTXhyCzN/d6Kj/C29ncHzBRIfab+Sbh+4g
sadMmb5Z/RukvH92l907btpw8z3yp3R5pMqTQo3qGz9ucnL6FkBnmjlgdKAapI5PzFmUcPGDKrLR
jCDmoieG4TVlddobVUSSfhF/qq+0Ko06QSTgtYx1wOelzXgjozCt9fKfsNdFAb0Ldhp/NO3iUYts
iklsFPrTR/JzDkyR9L3bv7R+aCM59PyoaxK7mluvXQkmlSxZPuOubnH0OZ+9cWi1ZSGqAn1hOEvV
jMKn8ux2UthDND0LCK/eCfEvXA3QvWnx7/XnLI9TfGZDXY1SsYTedmbAKtEs1V3jMFqx7pXpc5Zv
7D55OQf2TUTas3xsPTCTohpT/aksHOJ5/tQS/Jtjs4/lQEe+pbRzucZAyGsdrXPUFxtrH9KJ2cK+
c97xVFHMrmu06r5atLlQDDV5xUqHj/ZWDkIO8iBTW1NlMX/v1CCl3i4gujYPDQFzXATpfRpWvKyO
S+MwbYPApqGrBRg9125oE0xguLqfQmu8ighL5hfdL2x9oxdmp3teO859cX/qes6BxsiLwfsSZhSC
VcSQlXXRRKTfbjk04Yk1cfBz5cl8TtYZPVRGN7aaV1DuvCeOWw1BirRxMozBSx74WH/d/TN5+m63
2Fq6SQHSoKvulP7HZtOvuVLxopHcxOojq7pzsmQqPr+5IEpPES7oHnfQCFErOPC0w0vqFrrhyXCs
5j+Ku4HocsqzxeYgL4ddgDj6QEJ47BC9EZoUMinlHGuAprjn0rK8GbKXVOU0uc7KUVKHGQwBOfSr
ssDVNlEv7FRlihtbvPRsvR5l4Y6cwIm/U3Ig2RvWgXgEBFv0bV9uLwtVTD1wAk7Ms2fHh8PZTcsN
p4+bEpTjG5kx5a+Ale9QIYe8+637EA8CKUPKCrw8MdagJk6W93l8Xc76jXP1vodd2pHl55TyrMyN
1hS0QEVq2PxwEEeSF1RQsY7qOaH4dABi8K46UqVP0WOUAlB4CQpOekKROrvUe8NE1nqy+hfA7AiH
1gyLQ6wRExWb/akt3UWCOoKwc3123O+/sEiXzELfTvVfjmeP1es9jfQ/Zpf1ReP4fF33jFObcY1p
M9WvvWsTMamkBElLZF3Fa1ofHivoSn4UuJOjfUYb+g7/0yb8593dxz5KIp0JLUOS94oHISMm6UDs
lM6HNZmOswbuCjxgEPxF8Xscpt+KWGNFwHIuBPhEIhBTcrJF8V1rSG3XyRwiFpHxx+5C158X6Y4d
T2mAF6Bis7BVpmafxo3u9+lM6P1poK5aHIug3KT/lcxYCrZAmVA/nkBlKvxsMxg7KxrABspfqPNP
3qQEGR9jAl6BfBYcpY16QwMeOSDfEFFd+zP3i+rDJlGCRNGES0yZAUDBAcB+BWbwJT2g3cUt1iDv
dBc7gi2sZe8Ov3+TQAFZJVIYixkWh5psWlp5bAxHGKOfTbVeL5rxzpdKRgXL3kd45E/SAAbXaqjf
n+mgrmi2JLXmgnJHyj7KmqW6kDiVm57hqbozQJJrXi+Vag3yb4mCjl7e0rLOQCXAglVLrh7F88pw
5C7bs0sZ6cjiAjXR8+t5w/WFpk5jDndJoojEUoYIq/odH5vMjYhNR/umpFU/cmc+e+vq1494GFKG
gXwEm89rc3deQxx+zCy5r1Ro8gPfkfOMtIfVZiw3mdXipT3Bc18lHeikPPDCxmQyvtUhn8+tbLa+
lxdLnPUgFGeRkb8GlhKesI5Nm+zEDwhHs8QUqfMFhLnAos5Y9QQQO0AwRP+s/L+gu5jiEvuRCOz0
D4x1PjQkKVO3Esk6XpzhAi4r1UpEIhHKdiimFG8a1xwgwHbQB3VK3a3irWsJfvYmaGYFk0kcJnso
4jl7hRhZlvTTRAL/Ki0MQyCdOHxye2HT7pfZ/z3tczzj7Wpnvf6QlDYD9pjtKanp2+f0+hJiTp5l
daAchyKddCAs6gySfvSdPxHKlnw08cvF1a6/H3apvhxBMdGA1sgglGuUV11pnpNHrdfeX/fI2llj
VdSLzMbhMh3gjFQkbu3tNJUyke94OlDswXVMnuVTOJXbeI1ZTLrFgizmD6rEb3+R003JdkD4DZ4x
Q0BVLwvaBij9ivSfJ9pn3HMOblU9YS1KOsZEfXCGdXvPxP54/0mhP8fkUNrYqAXAPI16RL0mZRky
cxs9bRiEHVUmVWns7ErL0rl2a35W2+kHoYvnJoM7aGrS395ZeaQucbUyW8irKuZVtmBUm9hkw7pg
ZUoQPJSHVFell4fQ0PbORUmpkVS6k8wo8ZpSIFV3qoH3QiDc1dcMVOwIsyVifKSOVTlVP1MpUddp
U4i78mRd3MOzoYZUhdi6ki7Nv5s8+7l2G6c09GqoJfvklmM+UprvUf5gq9ZgWXQQfEQhvTFke96Z
LHU7fS3I/2Pamd7P/tHZy6BaIf64Rj+ylD+26hRx0X4r3s41C5UiPpb/+wvq9p0TRYMBzhUceFZT
UzJWaDU47d+7hdb/ZDeejwXGYO35u6qswryimrvvWopFoSMRpTQCsyU+GvJcoXK+SFuUHC9HrLVq
Qvj0lc6r9qS5k1LHiBI9GylWU+ei4TghDyCdbWCheTUQYtP2tPdBkjjyQoGXyJRo2ZiXA/rLhMaF
wW/ycwKnJ96xJ7WFSzFBMUs7lAxNHUzLZlZ5No1fazIeuQtsFqqtAbynpSrQs7SKhujyumbfQrAR
PiRJV1w85hPPSNo45U/YvbByoqzuaDJS7FwSGlenxtkgP01Ui15fg+XdPll5zVDtm5Bgo4hj5L9u
Zrpfc2zPzCF6jJLD+2RJgcAGrXfjGzWMyPqKP5eu/cw3noE3BmcQ7k6Pm04vCMakfVfXGaeFcfb7
emFBBftYCoaLw69GnthTpNx5Mg1BJBISAmPaQEeIFgLWZ5zBBy7CHDVxIJ/PRjmjfUoCSLTNkyof
y02CyYABUUxYeH3/svABdPgb+RHSu3WuqqusOFOnaOUfq0ODRZLJiFsAXVrf8lWJANicfid+Dumm
tGRNl90RW6aRDQrjE8VNw5QythhADbtF3t5Ncql1ohoo+Hr28CkfR2lbBbqFhfo5akrNmFdRZnKV
pq0fVcwsE4IlowVqY3uVKelx5cDZLE6oIG28FX12PDTs2BMKmB3Yis0LGn4+iYVTGrzeAU1i7Vjc
SxP50lg67lSE5hrI41fh/NrAwBLvg4VrGHJmKNF03K94mYkFSySFU4OeX57E1ZuzNmMtgV8Q7ADo
quQVngpe0ltj4UBHchXSGybPRPRMxcCzql/3oonKDgQASn9s3vBeJOeeTegtZAj2AthcLYUisLo/
rN1m5ByiQ4xkeGm79GIk3jhIAtwFUwjJwGGTnBC/aOfQi5NIPFTLj5JYmBJ1Vtx+8g89shS1C77K
pfWorW32jW1sVSxMw2tGW+reg8JCJV6Jp1TemAaxcX8KPeqqGTpu54eUSa1+a8D3pXaAoOg5XHie
a84c+QwRSebzUoNKQmYHKSNxQdIhVVxvXmzCim8+ZSZIoFduyw2veAk9s5ma97WRKYRZ0/18yvJb
34EMPE1ayiRqblM0kG/bHRyw2dvpeorOhWU94ZrfZkUsEFii746UfLXSxTFbwjAcjHmMRD0otiVi
wBKCjBOfu9NGtcYiea/ZV1fvrUNbgILam5xU76m0qp4YqG1Xp2ALFaF3F3Mphs0d3HtnbbWn3U41
bm8WXrYDoJqvdZvzM2Km0PD+6r3manSw/XL4F+kkn2xF7zCUprWht01HWCLtvRrfAm2rc5ATwNDV
87YijLtkc1neqoq0oQE0D3k5oeHBDDtgjUBf6yck0UAMjhHlxDPnxTKgmUa0XUEQMdEN2jHqAuTR
SEe0DwvMa6wMGnGvIcUY3wqrmr+S+58tN2nISOngkwWluW6TZ8nfCfpEb1Kfvx57Y8wVfsLNNK3v
HV3e0Ieim3q74FReA+HFcshh0z9YOphQYPYyTS2bxeUAh73hij524Z2XhYDT3et5pfZRSn1/ZhvC
1Au9qNhpr8Lb+3zczg0EDJXXmdIbJ8GP0tOtgVKzpzqtSjM2mB3C8acdIcBbStQAfLNHCApT1qRq
vEmxra7RCyt3iGYQri+89PX0ckRzEU+TK72dz+TFhresgmxB0AuVtor6UpI8aKS90LSL+HdKaDSD
ydlyReaxVESoMXU0pO9VEnOethd+fOZUGZsgDqmNxHh3Fm3P2+MQIq+gQ0AxJgoGsCLYxYAli43o
DaZMAWvC0p4eTF4Ygd108Xdi3i8hRKfgZEYP4BhZHf9BJX+sXNGbJ350vNnXce8l1vn6aFXZmMql
Dhn1GdrojzBiHnci7XcN95bHxJCtg8Mc9ZXNSpceivbvU4LJboLWowhQNTXo5rnVj+UoKIguSSHh
ARZqnMmqdCdpeGpuw89YxgQQbGRzR9RDsCDHlbL/O/tl4H9Lb3S0ZxcfREwfEApZoqXlInBE3laX
gQPaNiQ0VqS7+U8gB0dRRcFFa2tGKoiJXxs7US0gjC/siBpGAzBVLKvjCQaMhmxhqB/mBdOB9U2Q
Io5KZ4il9bulPJNCYjM26UP3LMUrLtGl1lxSr3bF4szOm37EeLD+CodMOdvUC4kai/U1Ya+kp8HB
9fDHL7JOv0zfq6io3Fyo59x/BUvDH+O5JPdudE/nr1RBqIUGPEwCfsBIcQwS7jp/q+1zmHVz0PL9
SgTXCwZeqEsC0B6bzJ3P4AvFPD/Z3exlF93gCNeTiJsVViz8DxzkVXObeiCD3dN5Ja85G6S2w6y1
Ei1YxaYt1EZAWMSXenLbTksGODISl9UpDkVXlgINU0o/rxeDnlEFw55zscnthAdo3BtILTRO76O9
gI6PJE/M5OC3CBjpPNlu3OnQpZRfK3LbL5teuzVfKULRjtTyFjgtvHUT0+Hg039O5pn2pTMHMN1n
hcPXOpRUNP6AOwfagoIQSWqDxTGGZbkEZdw/ysJatizjXWyZfjyciLKHDTNiNzUjR0Sgg3HO0MLr
r9D77bjZwP8Aa+/2luSDA9Iz4Esmxa0uD9y0exhRIdf+LKys0ZTm+M++hckVUZw24knTX7wgJAiG
vzrDVGnoOgpD+jBtuxzqpCjp0oJjyom+WNlazlWwbSO1jHRfgIfuiT+AN7Yp4XqzACaG2MBRZ4Dv
9puewht7pKv4242RnmnwvACXdRE/MjE9juYlECoY0orS9j/9YeXZtSrmEhyny0EqpF8n+afYxuiH
ylsU5dyyqjebKlKDbBmCFbWUvZ3KVCZ5DZqgFpBbUHD/obrXpaeMQj+B6vXBshFFZU/UIECJU2g0
spC2m0B5mNMgRQtBGEfdLnOxU9SlQ7kRXUo4YO29naHvkIZO+sFoUOgXWRbWnMLx7V7sMU9cLEIM
QRZIo3WGAhSQzij7DRIdu0fnD0faoGcquLwPVnAW0Cw5KDQod+6gswl1deyN4bFne8XKROBBHERB
9E2gLShAQSD/s6V96lyBxGK5M9FJs+7rE9KHZeNSsTY9n2s9+7Yy6PckPfEnXnslceKS4WCWkl/J
PmwD6Werg/hxCfO9DpxQxSK+aMyZeUEKVjXd3l9eRVhtP4IiRm7lJcUh99ZG+n3/fxie+NapCgZb
i+vantrwPue+b/G5toqZdODG/GqXt9oy5qyOl4mnhUpLVBuzkoYxs2CKu81SAmdTTDaoyGmUFoUa
FLCZyPcIyst7OF33Q/N2cHXyUSnNU/sXPmgBmd+gnAC2h/Tcxyo7oFjtkrMzreVpFnjF4BLELiXX
TGX5phYGtUkMshs8HFtN1lvxBxcxZPcnOiRqP6y0Vvna11LMiTt2QbPx1m33IqksK04O71ASxbeO
27RyEVbanWQ6c0jBERdbLJy8yKZr46rWnUb3borSbZEYkv5cs/HCEzIICQ6kUG293IWa2yupOsk0
8i4BfoCKG8hLmKuzQ1HJPa9ak/pYEoKh9y5D211kvABUXsIE4LtECqoIztSdY2aGzufRSViR13pF
fkNS+1wkKmKB6FU2ah0s0pVK8YbwLHYlk8e3pIiYvYBD1fnI0iJa4WPzw+JLQx0V8B8jBKdR0RVd
B4APBfujcXuBJPMQZLiX8FT6oV2GhLJw1PZy3BHTGq8CVDMgFKwA6kXdi4ULR2aVtNmfGltim2bO
pyiVmmOPN+3mN/dR3z5kI7cKa6er6L8k53IsHnVPKmEarzjhF1N88SDSb447HjgHUxmTewk2i0T9
97PYrCMKOAanLnK2qF5BJ70NHHKWcq7pi8NXho6gAqCGWkXGaZPBtJsu1HU4W+5kljka0223RBle
rxOMEMZE2nmJv8rJ8tDVJIjaQ3Ivumys9ZDN48wvIONoLR466hfpW7HCEbJAo4zAJcnpBrhKgQnf
nLYTAy0HLaAgRihj8ZCcj5zCwo6SwRkj53Wp4oXpazXe6cC0I+c6J81gMzmktmvP1NIFvzXssLp/
9vAEclaigvEaGR5r2LhBS4gVSnb87WPxwYiaIXbC6E6KBas9R+CM5DgdaGM4EHXWIbfG3Prn9lGx
hcLnrPfTNSKCAdJHpZLGUC8XcoaMHi5VRssh7Jvy6hCgbK4dAKpY6M3YxHEpgrrqwAwFarxvNgp2
L2COMSmssDHMB6lsXJ5XvdY5F1z6pAi1ePJB9MgT1qtlSqAJZNUxGZxrb0NbZbgLf56U7l3JEGVa
ueuUjIwbUsUJ7XnT0L0t93d1dVe086NFPz4coLouxMULTw2LRCunon/D3Kl6f0x17Ww8gTQXSh0R
DqSQ7wkMmPABv97FYHGr6aFzguoJDf/XktsXhAb9ztYq+Tixz/AwtRLqiV7DMC9Eo2xS263AUaWh
nvJ+HebbD8C3wF7y/Rlb6ngwhkRAjTwMHD9/JykE6RPMmBNMYb1g3alhpQ+nH5x4C+VskB56IlmZ
tF/dDUZzgXwjcLWkRBpXxJZhDQS4dJ5R1B312yezYmVvWMIcVSHMrea7zxI+XhGX8OAJ8+KTdiej
basuYhu8gMKacIuzyuK10LW/guxV/xm9+GlJkg3+rhuczt/sAi3FZkr1BsTR+Ck1cKlxo1Y24jK5
xzNDHkvwedGNqNeSx+XMQyUt4gHMrIVGCAa6bUie9TC79XdmDLqiHv0fHG8e4wFEJgC4EDV3wDJs
CMP2HqTvgxKJdEHjWrc3nePggzFiU0OPdZe2Ifnw1EymQYGNUkvF/xrZjvgz0xWLy0g648x9lqBQ
N+H5pwHrDc9ug1VpILB1turWxYWU+z8QDJXfjKLArl9goyaanY1JATu5sxWkVr38Ddn7aGCT9i0X
uYmHeeFvHLXc1xyxxThAPGDcnAbt2HhNeQf+OJyyULWLYgmOGH3pEDytovBpV3eZyDcOkagbwneI
bhbuqAa7iMPyqcH/193U0+n//lRxbddju9ImAG1xenY5teXUd6hQGAahD1868Z/0L5RUWdO44NCQ
qGVVRYqPEPXqNxaKrQPl3v5bgz43CXxI9j2FUAyGH6bwDz/vCBAbBFUGsjmhFtX6Es5F1IETY7rK
uLSnc50LKY8I7wDZkQVhbRJo8vVT4I6K14VmYzfLW9EJKnA3SLVSQvBTmgt98paWtNCfbaUO3esJ
Odlm8VImk7ol6n1eLOKK01x0x4KhDD1lF62Us1zx67fpngbboC1HEUp3Hc22ISOAOeHwSWqrUn3N
z03mwilpCO+htKe9aUOZH2VIci6//cJWURfOpjKAn9nqvwpsJ18NUOAITIaxWhqO70V0d6RwwchB
lUugZd/tnU1rmcMS5HT8DaexwNSKdNNtzLGeodea9CeXRtjik64wMB2EjJ+e/USJjqY0U+QhhfFK
EcrcdTkr2uqYjUW7TRjMHdGDIxHL4oWc3+3dc3NeooxLKJu5ayL+Ne8XDiPUgrlVXLubU/KeXkpd
ZCdEAUQUlbLG/e1lPKvODRA9TGeIs9itRTUnH0D5+JVGaAuFQIvics3Da6SkgiOAktGlQUrdpyrw
vkTf2741XqlDN5bzGrZ1KqxDVsSPsB14YmQRvRZ2YcaymzgBwIL2+oXE5hv8K4DxyL2LjKLl2Twi
AzTK+KwCggMb2vAEsQZ+pxlBw1oR4sXW69E/Gvt5JZ3E7H8Ln66YJcTPq8mo4H/UxJmYnQzdeFNG
I2ydulMbKO+RjCrBm0N8uAopFrbpQPOmexG+8UvuYWb0aEBlBolznPbw1P7qfCgPF1jJPpaNOlwQ
bir7aS6QwkdccwOdgAxR9O4GUIrIO0sNPht36RCge4DHYzeT9zYU/SJR8clz/Hqe/6zYX4SQJmR6
viCL1oqOG5XNun2aoEgl9/ZAaBt3QgZLHBOaurROgNRKYGFrmQ37GQCfjzsE2tFdaogI3wWQQsEH
WJRpA+9Y3uxeigChkQ1qSt/n3Q0NdxheZ/3rtI4gyOABAYOYVEAjFJe2mBsw4yzX1O4gnzRhjOQB
my3yrCRf8SKfdwsZLLRtGEwMqRaS/mbwrz6gNpReHIbgmOw2rC75lOIuDu9af1uA7DrPD8ZeQVp3
wovWBeFXkko/iYFA3XN7PJ6ku4/6MF0fiwOlwiE3D1UHzcKgTaYpCT1SCt4/UyZg0MjmcQ/K19KA
acIcPbU5+keI35koZJDdNdgA3STD/Og5279TAuwb24RxyX6zNGLdN/kmANp7f0RdM/Is2ZHvxQqo
tHwES5F58/T4py3OT2oBMj1uUVojVJVlkYbrT7LGmOMJPy1JxnYMd5KjlIQi/KwbdTREGYn18uHt
PxMknXJF/w/7fHrvGpZCvR7J78eaQeYSWbxuC/IlGIM2/FvT/ANb+sPoPcZ5iz9TYBHuEkS5Blus
Hg5P8c9BwgXikwNHA96b/vKdpQCGss6f+1U6XK84vokqyF1pvkjg3+g6QbY1NeRoreLMmBuWpIMR
h67m7/9T4FeUgLY4oe/VJQ+/351H2SpMPg259TsXdalwNHx+JTdxIlXiDas/i1dlEgLdu3+COfXf
uHWgeE/R3nccDSA3nbuxOQuPDTkx+6isO8rLmTUXVvY0INncYy2e5PA9Wr3kKDrK3lLd6A+Mcyv8
T/8YJiqbnVp/lQY6MXjlu18KHE9mWralDb2jbK1tJE1nA2rSmVb/suRAx6sup4QQwzJHurnngI0W
JiT8YfAbGUxl8YCzqlYnQHXc6g6UlcIMAVgLByCm52PzScNDsITbLYV0ksiZlCbVQNaLaGjiL7yN
mveMdhU/lNSFYTXPMPA42H7gua1tm0mS4iu81UoZ2SpuVE0iWW+9eoP6Na1zr3Bev0sDJ0MwWcBR
+m86+EtH02rFUkB5HYxi46HXuvVsuEqDJz1Vo9pBR7DOUxRBucTHMCN1USSssM6C2jHI1rQ7vWOn
7J63/4JOSy9AO6WobYafUFDDgBhipqUkaqCfDGZEHtxUa/JK6Mi3WdZTuMAWGRnakzRlHddE+ecQ
drZR+wQqB4zKCLOO1y/d2BXQifpRw3uhQWlxtRPQRs7uuxWDJvt2cVFMIXL9EqfIvHFR8b9s/cGC
Ce7RE5GYffmfWM8Lm1U+OvGmpWJCRbfSKSmkYtOJX1VZfVTGWnX5jsWU/T0D5JmCiWLN1rfDQCJ2
OiNC/bzk+JhNVIFqRHn/LkKd/P26aEzidZ+7j+CJqNhVIe5zENyFp2LDXMntlcKWu874XyoUDFFv
SsHb4Z4DWZaCr4gFHcFJE51+no8SneZM52n9HWcVSX/emDRBbPiiujgJQYIfTk+LRWohU3N66Vh+
1oCNH3dOkPCH1dwbGkYlK924zZnWPxCo/gkImelAY1DU1Gh1O6YFhJWAo6jAD8uik2EJZX34bYMN
BcoQxTYJ1+XntNoQXoTXifvSdEE+L49pAAsvPtvEAUYRBwTOVP8/C4IgGT/rF/ZxxFuuDqTjqzTl
P8Oy54YbWFjlRd2InmpLKWeyaKgKSUIMV+9II+y9c4zOwnrQVDhpihkHOZcfch2IS1W6k0/S29jM
f3VDFzvOdI5cnwMohGoraNd7ibfK2iXZJcIG9bC+DG3v031g/FcJJGR+0OJOOAPmhQsEa7xseyhT
ta4/XqjrTRC4xL2MKMpSwONrlq9FuuSU29uneKeX/q+clMrC5NVF6jZhMSIxNO8VRBeOU07MeuLQ
fzV8XbBY/hqUqp1SQptDSncSCG0y5g9d+NJsHn9jhDUDVpjzM8Ov2he4mIhH9Z320T7FPh/wrH4i
rirY76Dt4G43LOhe6t0+LFL0XYCfLU2hWBbGfw/KCDB70tQP0oyy0ocpIw9Bg+yEO7W/mqas/05p
CqP7IeBzmZ1TSv8/Vk6O8yTns0Ze7kOkyx3zJfvR8y5hgjmZv8sSDbrdq8rim7aFNWzLOu9jNf4X
0YsVmRj/nM7qsohcZi4E+PsIfEyWWZKxf/CW1YIilM874JiDCJdBVOuxAOv3AGr/jBwKxG+SpRiG
evd6lFgpQB3qhrQ5lgtD3X64qP7o77m2CDfdU/cMgPfujHM18sItNN7KfLy12TW7aWf41uyvdM5O
t8vQOEw0QlpnuS9zZ5qcNm6yiOvGDE/8xS9lJASgSUFN7Om28qO11il+yQxndOPlosAKUbl7k9du
UdT0J0C6F6P/OcZqF8RmLrAioKbM8JSL2yqiqUIRuWC+zxjKOzQCRIT5zAL/4oX6NJvctRnauvvB
rpb4XhY0MT5MVHTly2nWmx1G1E8hXu3E8G+XE3UC7MeUrNQ9a7K0c/T0flm9dh2dru/DOIEQH7Tr
tFHkfZ5vrcvqK+oN+DPA5MIatBs8A+ASYAcmMJCMbg4Yvj7z91xdmj2CVkpqenfsDuAMT8YFKcvK
2UsrEao4zdvDNAzyWUUW7nQ2zTtQIMOG+I3l+fkjVybE7MM4aIHlbALP13sGvcuCtHAGLAYxn3H4
68B1/jnrFVZtqZXrEL189YrNE6lfDWtLcwrFVIsU+5OdnsO6Y3gfj5lyFAJvD90fmr11SDlRHrgF
7tf/95lP1FntG82c2ff4yXzajmM8UqPsvq3iP4IpeOrsMV3lkTbMwG4W+RqbsfYxKV6AmA8tFGoG
qP7Dx4mZGeLB7GNGm50KQujXCQJwxbkwKPdZ82KX+dKJ61nVcjKI+wNkWptWtzA/qxrXZJgBksKN
qYXr+vVdtgFxV89gp6KmsDz/S+9S5aa3MNVrFEQkespw+le0yJRhqYYp8aJnBKstuBa9HkE1tiGF
1oWjvSRPy7j6Cn9PWwAIXtX8HX2EzcvRxrj3MWohyJazlrUgIqWWLarG2aqSdEW3jGkSzVpZ7MSa
6g+bBitSI87BmjEiwwcwmLZmDgMXFI577lL/2/jGGOoqG1hXpIb0HIDAroDbqXK0sqV5aa6E5k0l
y1MoFX8ipqjWbfr2gfVcAsWbyEbj4JX0ZH/d7YMl1PoHCqUuHsBT902RLNqPi6pNJ4uyBBLtUsiq
8XLfugG2TCedB3CcAmuhaQ5+CXR2QpioGPjhbhBSkKM/X3g0jG7K95nwowwFGKg22nXyTObZBEAg
RE+LjkQnhyoS6z3h694DEc3Ur2fujN8KpmRkKBoR4XDspARwJk3GJi0u6zVTa2kkixQ+YBit4gUz
ASr6nmKyN/IycXXoPoGG5Ebh37rJIKel149rrBhhwoULhYREDMK8r4OeQVMSBuPfo3KXaQ3laZNA
uZ5RZKwezTAr4EzQmePpwELR15F/9kMa0VRNTgztkO63xlEFnCVRT9nqDF5yismXV/l5Y5ULbdNX
LgM72sn1dhkA+/IF3QuYi4X4a15CMCoolx4qWi5mh/Ose5ugE5deRiYBb/MnxTe5/U4GchZm/T0R
wp3+m1drR0lKvngZxZ66RQ8drSOkCT4MxeQDxQHKGlEVmE4eNZeAy//a7xMzxuySKK0ABmEw5WlI
l9OKMToSI/B+AtLy9QM/PKu7k7gzpV1p4RzE58JXqDgJL03m3cAbuw+2ZDdqDx7aI2aD7mtJjXZn
F6b9r6DT1MIWY9Eg4KredGO1+jPnSofJTOurMn0LnTxXAnbtuAePBUlV3iaMf5Fz2D4bPt3q0Dik
pW5JD9sqajwDWTHYcBJtgPnt34k3CylmXKsrmOCO4zsW636OxZA+Zdxjpsrq2ydqcIxtjw+U65nW
DXV186YMV5z1qY5YL7Jvdj5W5zgqakSGJba4J9KztVgARxrTbmv7+Cp1kDt4zNpKvRLMST0QLKp1
FA1OvI0PN7H0pR5FhENpocDwmLmwXKL3pS0V7sQ=
`protect end_protected
