localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTX_CHK = {
  {32'hbddce957, 32'hbfd03ae4} /* (15, 15, 15) {real, imag} */,
  {32'hbf42cbd1, 32'hbf144999} /* (15, 15, 14) {real, imag} */,
  {32'hbe5b6e19, 32'h3f02a37a} /* (15, 15, 13) {real, imag} */,
  {32'hbd860cf0, 32'hbee06bd9} /* (15, 15, 12) {real, imag} */,
  {32'h3d31f09c, 32'hbe413c9f} /* (15, 15, 11) {real, imag} */,
  {32'hbdcb8f34, 32'h3fd6470c} /* (15, 15, 10) {real, imag} */,
  {32'hbe5fd664, 32'h3fea310e} /* (15, 15, 9) {real, imag} */,
  {32'h3fc865f2, 32'h402e56dc} /* (15, 15, 8) {real, imag} */,
  {32'h3f85fb02, 32'h3f06d42b} /* (15, 15, 7) {real, imag} */,
  {32'hbe8c1c14, 32'h3e0e0b54} /* (15, 15, 6) {real, imag} */,
  {32'hbf64c87c, 32'h3db61c14} /* (15, 15, 5) {real, imag} */,
  {32'h3de3c068, 32'hbfa165aa} /* (15, 15, 4) {real, imag} */,
  {32'hbdddb576, 32'hbf9e336e} /* (15, 15, 3) {real, imag} */,
  {32'hbe893456, 32'hbf4f3cec} /* (15, 15, 2) {real, imag} */,
  {32'hbf8afe46, 32'hbdd4a2dc} /* (15, 15, 1) {real, imag} */,
  {32'hbf5d92f6, 32'hbeeb98ec} /* (15, 15, 0) {real, imag} */,
  {32'hbe413a1a, 32'hbf975b16} /* (15, 14, 15) {real, imag} */,
  {32'hc009584c, 32'hbfe3bf25} /* (15, 14, 14) {real, imag} */,
  {32'hbfde3372, 32'hbfe39f05} /* (15, 14, 13) {real, imag} */,
  {32'hbf45b899, 32'hbe2c5798} /* (15, 14, 12) {real, imag} */,
  {32'h3f724c80, 32'h3e4476e6} /* (15, 14, 11) {real, imag} */,
  {32'h3f9a23d8, 32'h3f4494f5} /* (15, 14, 10) {real, imag} */,
  {32'hbe4266f2, 32'h3d4efc00} /* (15, 14, 9) {real, imag} */,
  {32'h3fd34c82, 32'h4010338a} /* (15, 14, 8) {real, imag} */,
  {32'h3f7564ca, 32'hbf6b1f93} /* (15, 14, 7) {real, imag} */,
  {32'hbf69e52e, 32'hbf86a9e4} /* (15, 14, 6) {real, imag} */,
  {32'hc0183169, 32'hbf0e3f5a} /* (15, 14, 5) {real, imag} */,
  {32'h3f89f6f7, 32'hbf721139} /* (15, 14, 4) {real, imag} */,
  {32'h3f059cb4, 32'hbecb36dc} /* (15, 14, 3) {real, imag} */,
  {32'hbda9c35a, 32'hbd2108f8} /* (15, 14, 2) {real, imag} */,
  {32'hbeb38c7f, 32'h3fa24976} /* (15, 14, 1) {real, imag} */,
  {32'hbe0f180d, 32'h3fdf6edc} /* (15, 14, 0) {real, imag} */,
  {32'h3fbcd73e, 32'hbf48610e} /* (15, 13, 15) {real, imag} */,
  {32'hbf673ff8, 32'hc03da6f0} /* (15, 13, 14) {real, imag} */,
  {32'hbf944b2a, 32'hbf81d694} /* (15, 13, 13) {real, imag} */,
  {32'hbeee4a5a, 32'h3fe96f10} /* (15, 13, 12) {real, imag} */,
  {32'h3e1be196, 32'hbddd8f3a} /* (15, 13, 11) {real, imag} */,
  {32'hbed04fa6, 32'hbf50ec2c} /* (15, 13, 10) {real, imag} */,
  {32'hbfffae79, 32'hc009005b} /* (15, 13, 9) {real, imag} */,
  {32'h3e8d7b95, 32'h3f351512} /* (15, 13, 8) {real, imag} */,
  {32'hbea223e5, 32'h3d989158} /* (15, 13, 7) {real, imag} */,
  {32'hbfa7b48b, 32'hbef0f244} /* (15, 13, 6) {real, imag} */,
  {32'hbf1ea63c, 32'hbee19af9} /* (15, 13, 5) {real, imag} */,
  {32'h3f07de0a, 32'hbfd333a6} /* (15, 13, 4) {real, imag} */,
  {32'h3fa1fc63, 32'h3f93e868} /* (15, 13, 3) {real, imag} */,
  {32'hbdd46489, 32'h3f247e6e} /* (15, 13, 2) {real, imag} */,
  {32'h3e9fbdae, 32'hbf22a5fc} /* (15, 13, 1) {real, imag} */,
  {32'h3fc57d38, 32'h3eb18521} /* (15, 13, 0) {real, imag} */,
  {32'h3ea33948, 32'hbf88287c} /* (15, 12, 15) {real, imag} */,
  {32'h3e55eb90, 32'hbdc5c570} /* (15, 12, 14) {real, imag} */,
  {32'h3facad40, 32'h403f3e93} /* (15, 12, 13) {real, imag} */,
  {32'h3fb24a14, 32'h3f1113ce} /* (15, 12, 12) {real, imag} */,
  {32'hbf632b24, 32'hbf983af8} /* (15, 12, 11) {real, imag} */,
  {32'hbf7bcb4e, 32'hbfcb01c0} /* (15, 12, 10) {real, imag} */,
  {32'hc00c5c1d, 32'hc01c9bdd} /* (15, 12, 9) {real, imag} */,
  {32'hbfd9ee9e, 32'hbea9e262} /* (15, 12, 8) {real, imag} */,
  {32'hbfdaaaaf, 32'h3ea987bd} /* (15, 12, 7) {real, imag} */,
  {32'hbef3a57c, 32'h3f69c163} /* (15, 12, 6) {real, imag} */,
  {32'h3fa75c05, 32'h3fa0d6ee} /* (15, 12, 5) {real, imag} */,
  {32'hbf2a2c50, 32'hbf8d57b0} /* (15, 12, 4) {real, imag} */,
  {32'h3d4934d0, 32'h3f1e695c} /* (15, 12, 3) {real, imag} */,
  {32'h3f057ba2, 32'h3fb98222} /* (15, 12, 2) {real, imag} */,
  {32'h3f9c89ff, 32'hbf8acefe} /* (15, 12, 1) {real, imag} */,
  {32'h3ea02d2b, 32'hbf80fc2e} /* (15, 12, 0) {real, imag} */,
  {32'hbf28f806, 32'h3f2b9774} /* (15, 11, 15) {real, imag} */,
  {32'hbcef92ac, 32'h3edca1e1} /* (15, 11, 14) {real, imag} */,
  {32'h4021334c, 32'h3f56f80e} /* (15, 11, 13) {real, imag} */,
  {32'h40445e15, 32'hbe36d53c} /* (15, 11, 12) {real, imag} */,
  {32'h3fb7bedc, 32'hbfad558d} /* (15, 11, 11) {real, imag} */,
  {32'hbec4ce80, 32'hbf8f9a9a} /* (15, 11, 10) {real, imag} */,
  {32'hbf678232, 32'hc023a585} /* (15, 11, 9) {real, imag} */,
  {32'h3f920e18, 32'hbff3a9f5} /* (15, 11, 8) {real, imag} */,
  {32'hbefc6f68, 32'hbfc325e1} /* (15, 11, 7) {real, imag} */,
  {32'hbf60988e, 32'h3f0b4873} /* (15, 11, 6) {real, imag} */,
  {32'hbf01274e, 32'h3fc29ebe} /* (15, 11, 5) {real, imag} */,
  {32'hbf8d43c9, 32'h3e54f306} /* (15, 11, 4) {real, imag} */,
  {32'hbfe6e698, 32'h3f0afcb5} /* (15, 11, 3) {real, imag} */,
  {32'hbf9ccab5, 32'hbe6296e8} /* (15, 11, 2) {real, imag} */,
  {32'hbdcae7a0, 32'hbf90697c} /* (15, 11, 1) {real, imag} */,
  {32'h3d887886, 32'h3d57f890} /* (15, 11, 0) {real, imag} */,
  {32'h3efdb21c, 32'h3ebfe6ec} /* (15, 10, 15) {real, imag} */,
  {32'h3f160f74, 32'hbfb1aa8a} /* (15, 10, 14) {real, imag} */,
  {32'h3ea1c956, 32'hbf38f50d} /* (15, 10, 13) {real, imag} */,
  {32'h3feeabf2, 32'hbf171a3a} /* (15, 10, 12) {real, imag} */,
  {32'h4011acb6, 32'hbe7b563c} /* (15, 10, 11) {real, imag} */,
  {32'h3f926d24, 32'h3f8e3fe7} /* (15, 10, 10) {real, imag} */,
  {32'hbfe7e2c0, 32'hbea324e6} /* (15, 10, 9) {real, imag} */,
  {32'hbfb08e42, 32'hbfad3dec} /* (15, 10, 8) {real, imag} */,
  {32'hbf41c3f2, 32'hc04bb998} /* (15, 10, 7) {real, imag} */,
  {32'hbecd34bb, 32'hbf6132b2} /* (15, 10, 6) {real, imag} */,
  {32'hbff47b57, 32'h3f9501bc} /* (15, 10, 5) {real, imag} */,
  {32'hc02550fc, 32'h3f356682} /* (15, 10, 4) {real, imag} */,
  {32'hc0292071, 32'hbe0c7555} /* (15, 10, 3) {real, imag} */,
  {32'hc059132c, 32'hbf6fefbd} /* (15, 10, 2) {real, imag} */,
  {32'hc001f86e, 32'hbf980441} /* (15, 10, 1) {real, imag} */,
  {32'h3ef0e84e, 32'hbe8e62aa} /* (15, 10, 0) {real, imag} */,
  {32'h3f0986c6, 32'h3e3553a3} /* (15, 9, 15) {real, imag} */,
  {32'hbdf71211, 32'hbeee68df} /* (15, 9, 14) {real, imag} */,
  {32'h3e130b15, 32'h3eb82619} /* (15, 9, 13) {real, imag} */,
  {32'h3fd90d1e, 32'hbfb3a6f6} /* (15, 9, 12) {real, imag} */,
  {32'h3e75f1a6, 32'hbfd489ab} /* (15, 9, 11) {real, imag} */,
  {32'h3fe993f5, 32'h3f4423af} /* (15, 9, 10) {real, imag} */,
  {32'hbfc23180, 32'h400062c8} /* (15, 9, 9) {real, imag} */,
  {32'hc013fada, 32'h3faeb4b2} /* (15, 9, 8) {real, imag} */,
  {32'hbe643e80, 32'h3f0e7f22} /* (15, 9, 7) {real, imag} */,
  {32'h3f564217, 32'h3f983905} /* (15, 9, 6) {real, imag} */,
  {32'h3e3a3768, 32'h401bb2e6} /* (15, 9, 5) {real, imag} */,
  {32'h3d878de8, 32'h3fc198d9} /* (15, 9, 4) {real, imag} */,
  {32'h3eb3be7e, 32'h3e43688d} /* (15, 9, 3) {real, imag} */,
  {32'hbf7900fb, 32'hbf91dd0c} /* (15, 9, 2) {real, imag} */,
  {32'hbfda3832, 32'hbf0459ee} /* (15, 9, 1) {real, imag} */,
  {32'h3f780130, 32'hbf0033da} /* (15, 9, 0) {real, imag} */,
  {32'hbf00f561, 32'h4005a3cc} /* (15, 8, 15) {real, imag} */,
  {32'hbee9ee98, 32'h3f90ecf0} /* (15, 8, 14) {real, imag} */,
  {32'hbf232305, 32'hbecaad65} /* (15, 8, 13) {real, imag} */,
  {32'hbe18a1f4, 32'hbec48946} /* (15, 8, 12) {real, imag} */,
  {32'hbb1c6980, 32'hbfaed098} /* (15, 8, 11) {real, imag} */,
  {32'h3fce115a, 32'h3f14bf69} /* (15, 8, 10) {real, imag} */,
  {32'h3ebfd930, 32'h3f49e5ee} /* (15, 8, 9) {real, imag} */,
  {32'hbf741c0a, 32'hbe077018} /* (15, 8, 8) {real, imag} */,
  {32'hbfa6229a, 32'h3fe779c6} /* (15, 8, 7) {real, imag} */,
  {32'hbf4c3313, 32'h404e4f34} /* (15, 8, 6) {real, imag} */,
  {32'h3e41dda8, 32'h40524e34} /* (15, 8, 5) {real, imag} */,
  {32'h402f61ae, 32'h3fd7767d} /* (15, 8, 4) {real, imag} */,
  {32'h401040dc, 32'h3faf4004} /* (15, 8, 3) {real, imag} */,
  {32'h3f7493df, 32'hbf4378d3} /* (15, 8, 2) {real, imag} */,
  {32'hbf5d1100, 32'hbeedafa0} /* (15, 8, 1) {real, imag} */,
  {32'h3e953955, 32'h3fd3b40c} /* (15, 8, 0) {real, imag} */,
  {32'hbf5a8342, 32'h3fcd61ba} /* (15, 7, 15) {real, imag} */,
  {32'hbf9726e0, 32'h3f7d712d} /* (15, 7, 14) {real, imag} */,
  {32'hbefa222c, 32'h3f9111ca} /* (15, 7, 13) {real, imag} */,
  {32'hbf9d9d2e, 32'hbfbbbbe6} /* (15, 7, 12) {real, imag} */,
  {32'hbe7bc3c4, 32'hc03a34b8} /* (15, 7, 11) {real, imag} */,
  {32'h3f407460, 32'h3d91f768} /* (15, 7, 10) {real, imag} */,
  {32'h3f78b51e, 32'h3f033e1c} /* (15, 7, 9) {real, imag} */,
  {32'h3f480d34, 32'hbe9a843a} /* (15, 7, 8) {real, imag} */,
  {32'hbeadd4ee, 32'hbf056ec6} /* (15, 7, 7) {real, imag} */,
  {32'hbfc6ffc1, 32'hbee97d58} /* (15, 7, 6) {real, imag} */,
  {32'hbe774fb4, 32'h3ddadee8} /* (15, 7, 5) {real, imag} */,
  {32'h3fa7a2a0, 32'hbf009a3e} /* (15, 7, 4) {real, imag} */,
  {32'hbc2232c0, 32'hbf3a411f} /* (15, 7, 3) {real, imag} */,
  {32'hbf0520bd, 32'hbfa25111} /* (15, 7, 2) {real, imag} */,
  {32'h3f9a9836, 32'h3ee835b3} /* (15, 7, 1) {real, imag} */,
  {32'h3fce3dee, 32'h3fda9158} /* (15, 7, 0) {real, imag} */,
  {32'hbea186a0, 32'h3f37d958} /* (15, 6, 15) {real, imag} */,
  {32'hbf8d372a, 32'hbf8ef550} /* (15, 6, 14) {real, imag} */,
  {32'hbe9b78da, 32'hbfb28eda} /* (15, 6, 13) {real, imag} */,
  {32'h3f807bd7, 32'hc0001b78} /* (15, 6, 12) {real, imag} */,
  {32'h3df818dc, 32'hbfdacce6} /* (15, 6, 11) {real, imag} */,
  {32'h3fca218c, 32'hbf173a58} /* (15, 6, 10) {real, imag} */,
  {32'h3e984551, 32'hc0245570} /* (15, 6, 9) {real, imag} */,
  {32'h3ed972ea, 32'hbf012477} /* (15, 6, 8) {real, imag} */,
  {32'h3ff149b7, 32'hc0187c10} /* (15, 6, 7) {real, imag} */,
  {32'hbf9832c5, 32'hbf947108} /* (15, 6, 6) {real, imag} */,
  {32'hc015bb08, 32'hbfc0a27f} /* (15, 6, 5) {real, imag} */,
  {32'hbf2c0256, 32'hbf87b2b8} /* (15, 6, 4) {real, imag} */,
  {32'h3ed012a6, 32'hbfdde004} /* (15, 6, 3) {real, imag} */,
  {32'hbf86cdec, 32'hbfc31053} /* (15, 6, 2) {real, imag} */,
  {32'h3ee5d73a, 32'h3fc7646c} /* (15, 6, 1) {real, imag} */,
  {32'h3f9d8e4e, 32'h3ee7885e} /* (15, 6, 0) {real, imag} */,
  {32'hbebd6383, 32'hbfc82aca} /* (15, 5, 15) {real, imag} */,
  {32'hbfb1667b, 32'hc0166ccc} /* (15, 5, 14) {real, imag} */,
  {32'hbee2d63a, 32'hbe8ee6ca} /* (15, 5, 13) {real, imag} */,
  {32'h3f346c24, 32'h3de16b68} /* (15, 5, 12) {real, imag} */,
  {32'h3f4dc4a0, 32'h3f194376} /* (15, 5, 11) {real, imag} */,
  {32'h3ff97554, 32'h3f35ddf3} /* (15, 5, 10) {real, imag} */,
  {32'hbf81171e, 32'hbf7ea2ca} /* (15, 5, 9) {real, imag} */,
  {32'h3f630c40, 32'h3fa3e505} /* (15, 5, 8) {real, imag} */,
  {32'h3e57178f, 32'hbed6344c} /* (15, 5, 7) {real, imag} */,
  {32'hc0189f20, 32'h3c81ccf0} /* (15, 5, 6) {real, imag} */,
  {32'hc0778c04, 32'hbf3b23da} /* (15, 5, 5) {real, imag} */,
  {32'hbfda30be, 32'hbfc649f7} /* (15, 5, 4) {real, imag} */,
  {32'h3fad6898, 32'hc01504a8} /* (15, 5, 3) {real, imag} */,
  {32'h4006c8a8, 32'hc007990e} /* (15, 5, 2) {real, imag} */,
  {32'h4064966f, 32'h3eaa8a0b} /* (15, 5, 1) {real, imag} */,
  {32'h3f84cfe6, 32'h3e65fafc} /* (15, 5, 0) {real, imag} */,
  {32'hbf47728c, 32'hbfb9d202} /* (15, 4, 15) {real, imag} */,
  {32'hc0247742, 32'hbf62b116} /* (15, 4, 14) {real, imag} */,
  {32'hbfaaea25, 32'h3eb32e60} /* (15, 4, 13) {real, imag} */,
  {32'h3d900a16, 32'hbeb86dd2} /* (15, 4, 12) {real, imag} */,
  {32'h3e29486b, 32'h40031728} /* (15, 4, 11) {real, imag} */,
  {32'h401f367e, 32'h403ae798} /* (15, 4, 10) {real, imag} */,
  {32'hbfa5d034, 32'h3fbaac40} /* (15, 4, 9) {real, imag} */,
  {32'h3fa91b54, 32'hbf1dfd8b} /* (15, 4, 8) {real, imag} */,
  {32'h3f4a4a37, 32'hbfe1efb7} /* (15, 4, 7) {real, imag} */,
  {32'hc03a096c, 32'hbf430522} /* (15, 4, 6) {real, imag} */,
  {32'hc0706b1a, 32'h3ff08703} /* (15, 4, 5) {real, imag} */,
  {32'hc01ea482, 32'hbf6a4456} /* (15, 4, 4) {real, imag} */,
  {32'h3e982c5e, 32'hc069e406} /* (15, 4, 3) {real, imag} */,
  {32'h3fd1edfa, 32'hbfe8379d} /* (15, 4, 2) {real, imag} */,
  {32'h3fd0d09d, 32'hbf3de33e} /* (15, 4, 1) {real, imag} */,
  {32'hbd61b45c, 32'hbf1b1cb8} /* (15, 4, 0) {real, imag} */,
  {32'h3de90ae0, 32'hbf05f7a9} /* (15, 3, 15) {real, imag} */,
  {32'hbeba578e, 32'h3f49f18c} /* (15, 3, 14) {real, imag} */,
  {32'h3fae5c3a, 32'h3c39f850} /* (15, 3, 13) {real, imag} */,
  {32'h3fd82592, 32'hbf99ad40} /* (15, 3, 12) {real, imag} */,
  {32'h3e50e37a, 32'h3fd98e87} /* (15, 3, 11) {real, imag} */,
  {32'h3fe03dfd, 32'h3f83d670} /* (15, 3, 10) {real, imag} */,
  {32'h3f4055d2, 32'h3f35c02a} /* (15, 3, 9) {real, imag} */,
  {32'h3f2f355d, 32'hbfb5d758} /* (15, 3, 8) {real, imag} */,
  {32'h3eb5d4bf, 32'hbfb424e2} /* (15, 3, 7) {real, imag} */,
  {32'hc01022d8, 32'hbf9c29c1} /* (15, 3, 6) {real, imag} */,
  {32'hc04e5738, 32'h3f6aeb24} /* (15, 3, 5) {real, imag} */,
  {32'h3d08533c, 32'hbfb2841b} /* (15, 3, 4) {real, imag} */,
  {32'h3f8d607c, 32'hc05a6f42} /* (15, 3, 3) {real, imag} */,
  {32'h3d2e2468, 32'hbed456b4} /* (15, 3, 2) {real, imag} */,
  {32'hbf4401e8, 32'hbe9aa051} /* (15, 3, 1) {real, imag} */,
  {32'h3f33a094, 32'hbee9fe71} /* (15, 3, 0) {real, imag} */,
  {32'h3f110423, 32'hbfe7ae2e} /* (15, 2, 15) {real, imag} */,
  {32'h3fdf0243, 32'hbeb6c472} /* (15, 2, 14) {real, imag} */,
  {32'h4036c0f5, 32'h3e5f7911} /* (15, 2, 13) {real, imag} */,
  {32'h400d7868, 32'h3e4d36d9} /* (15, 2, 12) {real, imag} */,
  {32'h3f7995ae, 32'h3e36e6c6} /* (15, 2, 11) {real, imag} */,
  {32'h3fcf91e6, 32'hbff6da95} /* (15, 2, 10) {real, imag} */,
  {32'h3fc5c834, 32'h3e445d59} /* (15, 2, 9) {real, imag} */,
  {32'h3f872a9a, 32'hbdae501e} /* (15, 2, 8) {real, imag} */,
  {32'h3ecc2a27, 32'hbd517e6c} /* (15, 2, 7) {real, imag} */,
  {32'hc01745b6, 32'h3f9dab3c} /* (15, 2, 6) {real, imag} */,
  {32'hbfdaf8fb, 32'h401ddeba} /* (15, 2, 5) {real, imag} */,
  {32'hbf95475a, 32'h3e43aebe} /* (15, 2, 4) {real, imag} */,
  {32'hbed527d8, 32'hbf39d1ae} /* (15, 2, 3) {real, imag} */,
  {32'hbf0d90be, 32'hbe5c9612} /* (15, 2, 2) {real, imag} */,
  {32'hbee66807, 32'hbf8d5e84} /* (15, 2, 1) {real, imag} */,
  {32'h3f986950, 32'hbf1f3f7e} /* (15, 2, 0) {real, imag} */,
  {32'hbf38f11a, 32'hbfc6b26b} /* (15, 1, 15) {real, imag} */,
  {32'hbf7cf252, 32'hbecfadd8} /* (15, 1, 14) {real, imag} */,
  {32'h3f6c896d, 32'h3edec9c8} /* (15, 1, 13) {real, imag} */,
  {32'h3fa3a264, 32'h3f23b86b} /* (15, 1, 12) {real, imag} */,
  {32'h3f1c720b, 32'hbf3d991f} /* (15, 1, 11) {real, imag} */,
  {32'hbe6f99fe, 32'hbf98758c} /* (15, 1, 10) {real, imag} */,
  {32'h3d42d0d0, 32'hbf801163} /* (15, 1, 9) {real, imag} */,
  {32'h3e547750, 32'hbfb80e2a} /* (15, 1, 8) {real, imag} */,
  {32'hbf76c161, 32'hbf2260a9} /* (15, 1, 7) {real, imag} */,
  {32'hbfa8e45e, 32'h3ff96ef7} /* (15, 1, 6) {real, imag} */,
  {32'hbf6145fc, 32'h40330d92} /* (15, 1, 5) {real, imag} */,
  {32'hc084ce48, 32'h3e0d8c36} /* (15, 1, 4) {real, imag} */,
  {32'hbfec5327, 32'h3ef0697c} /* (15, 1, 3) {real, imag} */,
  {32'h3f795920, 32'h3eb53774} /* (15, 1, 2) {real, imag} */,
  {32'h3f4bc28c, 32'hbf61eccc} /* (15, 1, 1) {real, imag} */,
  {32'h3e13638d, 32'hbf625a7a} /* (15, 1, 0) {real, imag} */,
  {32'hbeedf410, 32'hbf842654} /* (15, 0, 15) {real, imag} */,
  {32'hbdd92efc, 32'h3d7a9a00} /* (15, 0, 14) {real, imag} */,
  {32'h3f187760, 32'h3f0a8f11} /* (15, 0, 13) {real, imag} */,
  {32'h3f9d39df, 32'hbeaa4ace} /* (15, 0, 12) {real, imag} */,
  {32'h3e0e545a, 32'hbf2a52ac} /* (15, 0, 11) {real, imag} */,
  {32'hbfad071a, 32'hbe6ae869} /* (15, 0, 10) {real, imag} */,
  {32'hbf8cb960, 32'hbe99a2a2} /* (15, 0, 9) {real, imag} */,
  {32'hbeccabf4, 32'hbdd05aea} /* (15, 0, 8) {real, imag} */,
  {32'hbf73290e, 32'hbebf1209} /* (15, 0, 7) {real, imag} */,
  {32'hbe137076, 32'h3fada07c} /* (15, 0, 6) {real, imag} */,
  {32'hbece395c, 32'h3ffb62ea} /* (15, 0, 5) {real, imag} */,
  {32'hbf7a0334, 32'hbe8742fe} /* (15, 0, 4) {real, imag} */,
  {32'hbdf7fe7e, 32'hbf16ce5a} /* (15, 0, 3) {real, imag} */,
  {32'h3f46f216, 32'hbde21ece} /* (15, 0, 2) {real, imag} */,
  {32'h3eeb609f, 32'hbe281bb3} /* (15, 0, 1) {real, imag} */,
  {32'hbf0a98bd, 32'hbf30228c} /* (15, 0, 0) {real, imag} */,
  {32'h3f3d3f60, 32'h3e8a8b26} /* (14, 15, 15) {real, imag} */,
  {32'h3f6ef991, 32'h3f145b34} /* (14, 15, 14) {real, imag} */,
  {32'h3dc94b89, 32'h3f1f0ebc} /* (14, 15, 13) {real, imag} */,
  {32'hbdf470ff, 32'h3f628f20} /* (14, 15, 12) {real, imag} */,
  {32'h3f2590b0, 32'h3f8f7e46} /* (14, 15, 11) {real, imag} */,
  {32'h3faa1e0e, 32'h3fde5ae0} /* (14, 15, 10) {real, imag} */,
  {32'h3e7d3989, 32'h3ee177a4} /* (14, 15, 9) {real, imag} */,
  {32'h3ea92fee, 32'hbebab11a} /* (14, 15, 8) {real, imag} */,
  {32'h3e78e48e, 32'h3f5bff3a} /* (14, 15, 7) {real, imag} */,
  {32'h3e7f0ffa, 32'h3ebafdaf} /* (14, 15, 6) {real, imag} */,
  {32'hbf7f840b, 32'h3cef8758} /* (14, 15, 5) {real, imag} */,
  {32'hc025ba54, 32'h3ec73604} /* (14, 15, 4) {real, imag} */,
  {32'hc0112e82, 32'hbec73788} /* (14, 15, 3) {real, imag} */,
  {32'hbedc6fe4, 32'h3f129bde} /* (14, 15, 2) {real, imag} */,
  {32'h3c2e4990, 32'h3ec59b69} /* (14, 15, 1) {real, imag} */,
  {32'hbf37a027, 32'hbfa0d8aa} /* (14, 15, 0) {real, imag} */,
  {32'h3f0d505c, 32'h3f8f6d78} /* (14, 14, 15) {real, imag} */,
  {32'h40048b71, 32'h402db0d8} /* (14, 14, 14) {real, imag} */,
  {32'h3fbc6230, 32'h40227609} /* (14, 14, 13) {real, imag} */,
  {32'h3fc34ba6, 32'h40098e1a} /* (14, 14, 12) {real, imag} */,
  {32'h3f93f600, 32'h3f984dba} /* (14, 14, 11) {real, imag} */,
  {32'h40078a26, 32'h3f81e78c} /* (14, 14, 10) {real, imag} */,
  {32'h3fc29478, 32'h3e064484} /* (14, 14, 9) {real, imag} */,
  {32'h3f6429b0, 32'h3e2f6e50} /* (14, 14, 8) {real, imag} */,
  {32'hbf8bf688, 32'h3f381db6} /* (14, 14, 7) {real, imag} */,
  {32'h3f091530, 32'h3f54c23e} /* (14, 14, 6) {real, imag} */,
  {32'h3f35e1bc, 32'h402aba28} /* (14, 14, 5) {real, imag} */,
  {32'hc00d4802, 32'h3fa89d2a} /* (14, 14, 4) {real, imag} */,
  {32'hc000ddc4, 32'hbea7fea1} /* (14, 14, 3) {real, imag} */,
  {32'h3e729850, 32'hbe97c36e} /* (14, 14, 2) {real, imag} */,
  {32'h3e233c81, 32'hbe1c3930} /* (14, 14, 1) {real, imag} */,
  {32'hbf7e4662, 32'hbf50b3c4} /* (14, 14, 0) {real, imag} */,
  {32'hbef6b7e4, 32'h3e8a1b22} /* (14, 13, 15) {real, imag} */,
  {32'h3ee14698, 32'h3f56c201} /* (14, 13, 14) {real, imag} */,
  {32'h3ed56290, 32'h3fa8b14a} /* (14, 13, 13) {real, imag} */,
  {32'h3fcf76b8, 32'h4028eef5} /* (14, 13, 12) {real, imag} */,
  {32'h3f875d68, 32'h3f9ea0dc} /* (14, 13, 11) {real, imag} */,
  {32'h3eb371be, 32'hbf5ff8b3} /* (14, 13, 10) {real, imag} */,
  {32'h3fd99c98, 32'hbf8b886b} /* (14, 13, 9) {real, imag} */,
  {32'h3f29283c, 32'h3f5ab86c} /* (14, 13, 8) {real, imag} */,
  {32'hbfc801f3, 32'h3fefb1af} /* (14, 13, 7) {real, imag} */,
  {32'h3f536e92, 32'hbdcb5b80} /* (14, 13, 6) {real, imag} */,
  {32'h3fa95842, 32'h3fe576e8} /* (14, 13, 5) {real, imag} */,
  {32'hbf23c9dd, 32'h3fdcd4ee} /* (14, 13, 4) {real, imag} */,
  {32'hbfddcb14, 32'h3f0222cb} /* (14, 13, 3) {real, imag} */,
  {32'h3f2c5611, 32'hbf3a5486} /* (14, 13, 2) {real, imag} */,
  {32'h3fbbe7c4, 32'h3f99bb2b} /* (14, 13, 1) {real, imag} */,
  {32'h3f69e73c, 32'h3faf0255} /* (14, 13, 0) {real, imag} */,
  {32'hbe0e9a2e, 32'hbf2f9bc4} /* (14, 12, 15) {real, imag} */,
  {32'h3e0728bc, 32'hbfe52eb8} /* (14, 12, 14) {real, imag} */,
  {32'hbec8f80b, 32'hbef4cec5} /* (14, 12, 13) {real, imag} */,
  {32'hbf42e1ec, 32'h3fecf978} /* (14, 12, 12) {real, imag} */,
  {32'hbe79631a, 32'h3fb73436} /* (14, 12, 11) {real, imag} */,
  {32'h3e095c25, 32'h3ec63502} /* (14, 12, 10) {real, imag} */,
  {32'h3f4aa780, 32'h3f03fe1c} /* (14, 12, 9) {real, imag} */,
  {32'hbe980317, 32'h3f473203} /* (14, 12, 8) {real, imag} */,
  {32'hbf1d424a, 32'h3fea0e9e} /* (14, 12, 7) {real, imag} */,
  {32'hbf462cb2, 32'h3fcc4615} /* (14, 12, 6) {real, imag} */,
  {32'hbff4d480, 32'h3ff7dfdb} /* (14, 12, 5) {real, imag} */,
  {32'hbe4e183f, 32'h3fb6dff7} /* (14, 12, 4) {real, imag} */,
  {32'h3f834706, 32'h3cb46ef0} /* (14, 12, 3) {real, imag} */,
  {32'h4010b3d2, 32'h3e04970c} /* (14, 12, 2) {real, imag} */,
  {32'h3fa1ed3a, 32'h3fd49f45} /* (14, 12, 1) {real, imag} */,
  {32'h3f5060d0, 32'h3fc10a5e} /* (14, 12, 0) {real, imag} */,
  {32'h3f6ae236, 32'hbfb58516} /* (14, 11, 15) {real, imag} */,
  {32'h40286cf4, 32'hbf7a4dd9} /* (14, 11, 14) {real, imag} */,
  {32'h3f8a763c, 32'h3ff775ff} /* (14, 11, 13) {real, imag} */,
  {32'hbfecc81f, 32'h3f89432a} /* (14, 11, 12) {real, imag} */,
  {32'hbfeea524, 32'h3f732857} /* (14, 11, 11) {real, imag} */,
  {32'h3fa6155d, 32'h40040c58} /* (14, 11, 10) {real, imag} */,
  {32'h3fcf8b4f, 32'h40288662} /* (14, 11, 9) {real, imag} */,
  {32'hbbd18320, 32'h3f4b8170} /* (14, 11, 8) {real, imag} */,
  {32'hbf85e5c1, 32'h3e8757d3} /* (14, 11, 7) {real, imag} */,
  {32'hbf714c1a, 32'h3fa0fbf2} /* (14, 11, 6) {real, imag} */,
  {32'hbfb586cd, 32'h400be4a1} /* (14, 11, 5) {real, imag} */,
  {32'h3e553541, 32'h3f88468c} /* (14, 11, 4) {real, imag} */,
  {32'h3e8877b9, 32'hbf5fb92e} /* (14, 11, 3) {real, imag} */,
  {32'h3dd56074, 32'h3f353296} /* (14, 11, 2) {real, imag} */,
  {32'h3e9e09de, 32'h3f77e47f} /* (14, 11, 1) {real, imag} */,
  {32'hbebe7297, 32'h3f8dd525} /* (14, 11, 0) {real, imag} */,
  {32'h3eaccbbf, 32'h3ed91ff7} /* (14, 10, 15) {real, imag} */,
  {32'h401a7c18, 32'h3f85ad02} /* (14, 10, 14) {real, imag} */,
  {32'h3f812054, 32'h3f01648d} /* (14, 10, 13) {real, imag} */,
  {32'hbfc6ec4c, 32'h3f588a7d} /* (14, 10, 12) {real, imag} */,
  {32'hbf7dd158, 32'hbd6be6ac} /* (14, 10, 11) {real, imag} */,
  {32'h3e96b178, 32'h3ec99397} /* (14, 10, 10) {real, imag} */,
  {32'h40133a16, 32'h3fb60bf4} /* (14, 10, 9) {real, imag} */,
  {32'h3fbcb976, 32'h3f2ac954} /* (14, 10, 8) {real, imag} */,
  {32'hbf4fd2b6, 32'h3f39288c} /* (14, 10, 7) {real, imag} */,
  {32'h3e993e79, 32'h3e5fc5e4} /* (14, 10, 6) {real, imag} */,
  {32'hbf10f41e, 32'hbe858718} /* (14, 10, 5) {real, imag} */,
  {32'hbe912ae7, 32'hbf4cd5f6} /* (14, 10, 4) {real, imag} */,
  {32'h3f409e34, 32'hc007ce2e} /* (14, 10, 3) {real, imag} */,
  {32'h3f5f8a4f, 32'h3eef4d36} /* (14, 10, 2) {real, imag} */,
  {32'hbea63d6c, 32'h3f2a2b19} /* (14, 10, 1) {real, imag} */,
  {32'hbf917a51, 32'h3d761fec} /* (14, 10, 0) {real, imag} */,
  {32'hbf46059e, 32'h3ea74cf4} /* (14, 9, 15) {real, imag} */,
  {32'hbf6900bf, 32'h3ff2d218} /* (14, 9, 14) {real, imag} */,
  {32'hbf289c12, 32'h3f1cf427} /* (14, 9, 13) {real, imag} */,
  {32'h3df7d729, 32'hbf450d27} /* (14, 9, 12) {real, imag} */,
  {32'h3ec5a4de, 32'hbf957fd2} /* (14, 9, 11) {real, imag} */,
  {32'hbe9ab212, 32'hbec05bc5} /* (14, 9, 10) {real, imag} */,
  {32'h3e9598de, 32'h3fb70dd0} /* (14, 9, 9) {real, imag} */,
  {32'h3eff1f64, 32'h3f265eda} /* (14, 9, 8) {real, imag} */,
  {32'hbef37d1a, 32'h4008eb2a} /* (14, 9, 7) {real, imag} */,
  {32'h4018cb4a, 32'h3ea2d115} /* (14, 9, 6) {real, imag} */,
  {32'h4011ff64, 32'hbf8cb800} /* (14, 9, 5) {real, imag} */,
  {32'h3fde547b, 32'h3effbbe3} /* (14, 9, 4) {real, imag} */,
  {32'h3ffec19e, 32'h3f4d79a7} /* (14, 9, 3) {real, imag} */,
  {32'h3f885b3c, 32'h3eb69803} /* (14, 9, 2) {real, imag} */,
  {32'h3f09c4bc, 32'h3ffd1862} /* (14, 9, 1) {real, imag} */,
  {32'h3e2585fc, 32'h3f95d05a} /* (14, 9, 0) {real, imag} */,
  {32'hbfb1f350, 32'h3fb2d16e} /* (14, 8, 15) {real, imag} */,
  {32'hbfac85ca, 32'h40870c9d} /* (14, 8, 14) {real, imag} */,
  {32'h3f413e62, 32'h40182bdb} /* (14, 8, 13) {real, imag} */,
  {32'h4021128c, 32'h3ea86ec4} /* (14, 8, 12) {real, imag} */,
  {32'h3ed6b492, 32'h3e409882} /* (14, 8, 11) {real, imag} */,
  {32'hbeba6832, 32'hbf4e3da2} /* (14, 8, 10) {real, imag} */,
  {32'hbfe2d90e, 32'h3f3720f5} /* (14, 8, 9) {real, imag} */,
  {32'hbf46e04c, 32'h3ed68e1e} /* (14, 8, 8) {real, imag} */,
  {32'h3e809c6b, 32'h3f9b42ca} /* (14, 8, 7) {real, imag} */,
  {32'h3d15a0bb, 32'hbdc31738} /* (14, 8, 6) {real, imag} */,
  {32'h3f78eb60, 32'hbf23274a} /* (14, 8, 5) {real, imag} */,
  {32'h3f392ac9, 32'hbd3c83b2} /* (14, 8, 4) {real, imag} */,
  {32'h401e75e8, 32'hbee30210} /* (14, 8, 3) {real, imag} */,
  {32'h3ff3e60b, 32'hbfb26bdc} /* (14, 8, 2) {real, imag} */,
  {32'h3f26ec78, 32'hbe9d6058} /* (14, 8, 1) {real, imag} */,
  {32'h3ef8bc20, 32'h3f1b7d36} /* (14, 8, 0) {real, imag} */,
  {32'h3f1f692a, 32'h3fbb9f74} /* (14, 7, 15) {real, imag} */,
  {32'h3f0d925f, 32'h4059a264} /* (14, 7, 14) {real, imag} */,
  {32'h40069c06, 32'h4058a4b0} /* (14, 7, 13) {real, imag} */,
  {32'h402d99bc, 32'h40306e87} /* (14, 7, 12) {real, imag} */,
  {32'h3eb0cc24, 32'h3f770c30} /* (14, 7, 11) {real, imag} */,
  {32'hbef48374, 32'hc006fa80} /* (14, 7, 10) {real, imag} */,
  {32'hc005b92b, 32'hbf425a5d} /* (14, 7, 9) {real, imag} */,
  {32'hbf82e0b3, 32'h3f3362e6} /* (14, 7, 8) {real, imag} */,
  {32'h3e6c2620, 32'h3f23d7b2} /* (14, 7, 7) {real, imag} */,
  {32'hbf1a3437, 32'hc024c82e} /* (14, 7, 6) {real, imag} */,
  {32'hbee19b92, 32'hbfbf8aec} /* (14, 7, 5) {real, imag} */,
  {32'h3ef52a89, 32'h3ec5b72f} /* (14, 7, 4) {real, imag} */,
  {32'hbde93da2, 32'h3ddd4f61} /* (14, 7, 3) {real, imag} */,
  {32'hbd99d33d, 32'hbf5f8432} /* (14, 7, 2) {real, imag} */,
  {32'h3ea9e26d, 32'hbf8c21da} /* (14, 7, 1) {real, imag} */,
  {32'h3fcdc39c, 32'h3fab2b62} /* (14, 7, 0) {real, imag} */,
  {32'h3f44c8a1, 32'h3f8e2ee0} /* (14, 6, 15) {real, imag} */,
  {32'h3f28578d, 32'h3e5da825} /* (14, 6, 14) {real, imag} */,
  {32'h3f8bbdc4, 32'h402541fd} /* (14, 6, 13) {real, imag} */,
  {32'h4000d2be, 32'h406361d2} /* (14, 6, 12) {real, imag} */,
  {32'h3f9af807, 32'hbf1c287f} /* (14, 6, 11) {real, imag} */,
  {32'hbec2d341, 32'hc017d23f} /* (14, 6, 10) {real, imag} */,
  {32'hbfa9e33e, 32'hbf236b35} /* (14, 6, 9) {real, imag} */,
  {32'hbf440dac, 32'hbf223124} /* (14, 6, 8) {real, imag} */,
  {32'hc028ed73, 32'hbeae78b2} /* (14, 6, 7) {real, imag} */,
  {32'hbf9dbccf, 32'hbed2f949} /* (14, 6, 6) {real, imag} */,
  {32'hbe93d0b8, 32'hbe9cec2e} /* (14, 6, 5) {real, imag} */,
  {32'h3f2f6d9a, 32'h3f12a707} /* (14, 6, 4) {real, imag} */,
  {32'hbff1759d, 32'hbd63dd04} /* (14, 6, 3) {real, imag} */,
  {32'hbe9d5050, 32'hbfaaf2a0} /* (14, 6, 2) {real, imag} */,
  {32'h403f1a3d, 32'hbec50a56} /* (14, 6, 1) {real, imag} */,
  {32'h3fcc95dc, 32'h3f3b00c9} /* (14, 6, 0) {real, imag} */,
  {32'h3df14941, 32'h3e91418e} /* (14, 5, 15) {real, imag} */,
  {32'hbcdf6df0, 32'hbf96d0ee} /* (14, 5, 14) {real, imag} */,
  {32'h3f725218, 32'h3f383c20} /* (14, 5, 13) {real, imag} */,
  {32'h3fc3ad85, 32'h3fd70cfc} /* (14, 5, 12) {real, imag} */,
  {32'h3fdc424e, 32'hbcf508a8} /* (14, 5, 11) {real, imag} */,
  {32'h3e0810d2, 32'hbef23159} /* (14, 5, 10) {real, imag} */,
  {32'hbf9d4798, 32'hbe8f3f60} /* (14, 5, 9) {real, imag} */,
  {32'hbf0f971d, 32'h3eb76ee0} /* (14, 5, 8) {real, imag} */,
  {32'hbffb019a, 32'h3f0115a2} /* (14, 5, 7) {real, imag} */,
  {32'hbf0a8384, 32'h3deadf84} /* (14, 5, 6) {real, imag} */,
  {32'h3f5e098f, 32'h3e9fab19} /* (14, 5, 5) {real, imag} */,
  {32'h3e45b1c8, 32'h3e384f5a} /* (14, 5, 4) {real, imag} */,
  {32'hbfb153e6, 32'hbe6e4c4f} /* (14, 5, 3) {real, imag} */,
  {32'h3e38bab2, 32'hbe6ce9df} /* (14, 5, 2) {real, imag} */,
  {32'h3fa77666, 32'h3fac91e4} /* (14, 5, 1) {real, imag} */,
  {32'h3f296bfe, 32'h3f85f914} /* (14, 5, 0) {real, imag} */,
  {32'hbfa9faa2, 32'hbf56bb23} /* (14, 4, 15) {real, imag} */,
  {32'h3f11c595, 32'hbfbf3b90} /* (14, 4, 14) {real, imag} */,
  {32'h3ff5cf3a, 32'h3e7815b9} /* (14, 4, 13) {real, imag} */,
  {32'hbe11da34, 32'hbf985e42} /* (14, 4, 12) {real, imag} */,
  {32'hbead7831, 32'h3d8499e2} /* (14, 4, 11) {real, imag} */,
  {32'hbf749106, 32'hbf1cb7ec} /* (14, 4, 10) {real, imag} */,
  {32'hbecbc41f, 32'hc01c2963} /* (14, 4, 9) {real, imag} */,
  {32'hbf4b81ea, 32'hbf230090} /* (14, 4, 8) {real, imag} */,
  {32'h3e878916, 32'h3d2d91c4} /* (14, 4, 7) {real, imag} */,
  {32'h3f63f21e, 32'hbf7830da} /* (14, 4, 6) {real, imag} */,
  {32'hbed9b872, 32'hbf3cc040} /* (14, 4, 5) {real, imag} */,
  {32'h3f851c6b, 32'hbadab3f9} /* (14, 4, 4) {real, imag} */,
  {32'h3eda8ba0, 32'h4009c653} /* (14, 4, 3) {real, imag} */,
  {32'h3e85a62f, 32'h3ff059ca} /* (14, 4, 2) {real, imag} */,
  {32'hbe903222, 32'h3f804332} /* (14, 4, 1) {real, imag} */,
  {32'hbeb9a2bd, 32'h3f29b50e} /* (14, 4, 0) {real, imag} */,
  {32'hbe03fac0, 32'hbf428171} /* (14, 3, 15) {real, imag} */,
  {32'h3ff3efbb, 32'hc01ebee9} /* (14, 3, 14) {real, imag} */,
  {32'h3ed10b3a, 32'hc052e44b} /* (14, 3, 13) {real, imag} */,
  {32'hbfba5476, 32'hc0343ae1} /* (14, 3, 12) {real, imag} */,
  {32'hbf510ee0, 32'hbfb8c11e} /* (14, 3, 11) {real, imag} */,
  {32'hbeb2ca7e, 32'hbf236644} /* (14, 3, 10) {real, imag} */,
  {32'h3f264b74, 32'hbe192775} /* (14, 3, 9) {real, imag} */,
  {32'h3dca34a8, 32'h3ec5c395} /* (14, 3, 8) {real, imag} */,
  {32'h3ebbd6d7, 32'h3e5f40e0} /* (14, 3, 7) {real, imag} */,
  {32'h3f46a5ec, 32'hbf80071e} /* (14, 3, 6) {real, imag} */,
  {32'h3e93a8a4, 32'hbfaa38c8} /* (14, 3, 5) {real, imag} */,
  {32'h3fb343fe, 32'h3fb97e9e} /* (14, 3, 4) {real, imag} */,
  {32'hbeaacdfa, 32'h3f9f895e} /* (14, 3, 3) {real, imag} */,
  {32'h3eb8ed89, 32'h3f73c216} /* (14, 3, 2) {real, imag} */,
  {32'hbe9aee6a, 32'h3f5665eb} /* (14, 3, 1) {real, imag} */,
  {32'hbec5ecc9, 32'hbec3248e} /* (14, 3, 0) {real, imag} */,
  {32'h3f3c76c5, 32'hbf876e09} /* (14, 2, 15) {real, imag} */,
  {32'h3f4b402a, 32'hc007078a} /* (14, 2, 14) {real, imag} */,
  {32'hbff22585, 32'hc042dabe} /* (14, 2, 13) {real, imag} */,
  {32'hbfd737cf, 32'hbfc2adb5} /* (14, 2, 12) {real, imag} */,
  {32'hbe8c1f38, 32'h400c0ea4} /* (14, 2, 11) {real, imag} */,
  {32'h3f9bc1d2, 32'h3fe12394} /* (14, 2, 10) {real, imag} */,
  {32'h3f5a7c9e, 32'hbef0b2ee} /* (14, 2, 9) {real, imag} */,
  {32'h3eca07f6, 32'h3fa21018} /* (14, 2, 8) {real, imag} */,
  {32'hbd1629bf, 32'h3ff28989} /* (14, 2, 7) {real, imag} */,
  {32'h3f3e5946, 32'h3f87ad3c} /* (14, 2, 6) {real, imag} */,
  {32'h400b5d49, 32'h3e119d78} /* (14, 2, 5) {real, imag} */,
  {32'h4027d2f3, 32'hbdc053b0} /* (14, 2, 4) {real, imag} */,
  {32'h3f1bfe87, 32'hbf4eb04d} /* (14, 2, 3) {real, imag} */,
  {32'hbd1e4ea0, 32'hbf422a73} /* (14, 2, 2) {real, imag} */,
  {32'hbf73c6d8, 32'h3f8c1656} /* (14, 2, 1) {real, imag} */,
  {32'h3e00abe8, 32'h3f576d2c} /* (14, 2, 0) {real, imag} */,
  {32'hbdd1f7cc, 32'hbf1f91fa} /* (14, 1, 15) {real, imag} */,
  {32'hbfcb949e, 32'hbfe20bc6} /* (14, 1, 14) {real, imag} */,
  {32'hc04617fd, 32'hbf831d86} /* (14, 1, 13) {real, imag} */,
  {32'h3ea3b0f7, 32'h3d5c40a8} /* (14, 1, 12) {real, imag} */,
  {32'hbcff2f90, 32'h407d11e2} /* (14, 1, 11) {real, imag} */,
  {32'hbf90ac0e, 32'h3fa9e774} /* (14, 1, 10) {real, imag} */,
  {32'h3e88e8a8, 32'hc017ba9e} /* (14, 1, 9) {real, imag} */,
  {32'hbd953b05, 32'hbde5af88} /* (14, 1, 8) {real, imag} */,
  {32'h3f7bc2c2, 32'h40568383} /* (14, 1, 7) {real, imag} */,
  {32'h3f8a3fc2, 32'h40414c94} /* (14, 1, 6) {real, imag} */,
  {32'h3ed018e8, 32'h3f1dd222} /* (14, 1, 5) {real, imag} */,
  {32'h3fc48ba7, 32'h3f5199ed} /* (14, 1, 4) {real, imag} */,
  {32'h3f5f87fa, 32'h3f3f418f} /* (14, 1, 3) {real, imag} */,
  {32'hbf6642b3, 32'hbd23cdae} /* (14, 1, 2) {real, imag} */,
  {32'h3db04f13, 32'h401c7438} /* (14, 1, 1) {real, imag} */,
  {32'h3e40d054, 32'h4009df71} /* (14, 1, 0) {real, imag} */,
  {32'hbdba27ea, 32'h3de48640} /* (14, 0, 15) {real, imag} */,
  {32'hbf3ad4d4, 32'hbebeed98} /* (14, 0, 14) {real, imag} */,
  {32'hbfaa3c5c, 32'h3e51540d} /* (14, 0, 13) {real, imag} */,
  {32'h3fab45ce, 32'h3f4c18ca} /* (14, 0, 12) {real, imag} */,
  {32'h3fa752e8, 32'h3fce99c8} /* (14, 0, 11) {real, imag} */,
  {32'hbe834a94, 32'h3fa70f20} /* (14, 0, 10) {real, imag} */,
  {32'hbed9a0ba, 32'hbfa3f402} /* (14, 0, 9) {real, imag} */,
  {32'hbf5fdc2a, 32'hbff2771c} /* (14, 0, 8) {real, imag} */,
  {32'h3f47fd20, 32'h3fa66fcf} /* (14, 0, 7) {real, imag} */,
  {32'h3f74ed57, 32'h3f570731} /* (14, 0, 6) {real, imag} */,
  {32'hbf10af66, 32'hbfaaa620} /* (14, 0, 5) {real, imag} */,
  {32'hbf95dc2f, 32'h3e47519d} /* (14, 0, 4) {real, imag} */,
  {32'hbf3ef01a, 32'h3d13c91c} /* (14, 0, 3) {real, imag} */,
  {32'hbf091c06, 32'h3ed15047} /* (14, 0, 2) {real, imag} */,
  {32'hbeb1d168, 32'h3f90b1e0} /* (14, 0, 1) {real, imag} */,
  {32'hbf1aca4c, 32'h3e7eb2b3} /* (14, 0, 0) {real, imag} */,
  {32'hbe8ab3fa, 32'h3f33eb10} /* (13, 15, 15) {real, imag} */,
  {32'h3eaf2c72, 32'h3f08622a} /* (13, 15, 14) {real, imag} */,
  {32'hbe28b414, 32'hbfa5a8c9} /* (13, 15, 13) {real, imag} */,
  {32'hbe42ee9a, 32'hbfb44e04} /* (13, 15, 12) {real, imag} */,
  {32'hbf3ecc43, 32'hbdc8f06a} /* (13, 15, 11) {real, imag} */,
  {32'h3ddb94c8, 32'hbf30bf62} /* (13, 15, 10) {real, imag} */,
  {32'hbe76f8fc, 32'h3e18c184} /* (13, 15, 9) {real, imag} */,
  {32'hbf29d2d5, 32'h3f2bc001} /* (13, 15, 8) {real, imag} */,
  {32'hbe5046a6, 32'h3f4a2994} /* (13, 15, 7) {real, imag} */,
  {32'h3ea1b065, 32'h3e138a16} /* (13, 15, 6) {real, imag} */,
  {32'hbe3bca3c, 32'hbf9a121b} /* (13, 15, 5) {real, imag} */,
  {32'h3f9fba21, 32'hbf1cd670} /* (13, 15, 4) {real, imag} */,
  {32'h3ec76719, 32'h3e92de88} /* (13, 15, 3) {real, imag} */,
  {32'hbf6bc195, 32'hbe26862a} /* (13, 15, 2) {real, imag} */,
  {32'h3e9e7976, 32'h3ece91c2} /* (13, 15, 1) {real, imag} */,
  {32'h3dd2daac, 32'h3dd6d910} /* (13, 15, 0) {real, imag} */,
  {32'hbe6ee96a, 32'h3f9d9972} /* (13, 14, 15) {real, imag} */,
  {32'h3f693a0b, 32'h3e745450} /* (13, 14, 14) {real, imag} */,
  {32'h3f463444, 32'hc01480dc} /* (13, 14, 13) {real, imag} */,
  {32'hbefa795c, 32'hc02308d6} /* (13, 14, 12) {real, imag} */,
  {32'h3e29ceca, 32'hbf1bffd5} /* (13, 14, 11) {real, imag} */,
  {32'h3fb7ee7a, 32'hbfaacbe2} /* (13, 14, 10) {real, imag} */,
  {32'h3f6b1dc2, 32'h3e103184} /* (13, 14, 9) {real, imag} */,
  {32'hbf4575a6, 32'h3f3db862} /* (13, 14, 8) {real, imag} */,
  {32'h3f332d1a, 32'h3f328fe9} /* (13, 14, 7) {real, imag} */,
  {32'h3f89f4ee, 32'h3f3f1460} /* (13, 14, 6) {real, imag} */,
  {32'h3da30ae4, 32'hbf632043} /* (13, 14, 5) {real, imag} */,
  {32'h3fa54301, 32'hbe9b018c} /* (13, 14, 4) {real, imag} */,
  {32'h3eaa4eb5, 32'h3f84a748} /* (13, 14, 3) {real, imag} */,
  {32'hbeb8432b, 32'h3f176d9c} /* (13, 14, 2) {real, imag} */,
  {32'h3fde22ba, 32'h3cb5e870} /* (13, 14, 1) {real, imag} */,
  {32'h3eac49a6, 32'hbe86cdef} /* (13, 14, 0) {real, imag} */,
  {32'hbe88df6c, 32'h3f1ac332} /* (13, 13, 15) {real, imag} */,
  {32'h40248dba, 32'hbecfd29f} /* (13, 13, 14) {real, imag} */,
  {32'h3f4d79d9, 32'hbf85c04e} /* (13, 13, 13) {real, imag} */,
  {32'hbf9c24b9, 32'hbf0a40ca} /* (13, 13, 12) {real, imag} */,
  {32'h3f6d72b2, 32'h3f58b756} /* (13, 13, 11) {real, imag} */,
  {32'h3fb604e0, 32'h3f2b9e4c} /* (13, 13, 10) {real, imag} */,
  {32'hbf0f685a, 32'h3fa8673e} /* (13, 13, 9) {real, imag} */,
  {32'hbeb2540f, 32'hbda7e1f6} /* (13, 13, 8) {real, imag} */,
  {32'h400696f5, 32'hbf3208fe} /* (13, 13, 7) {real, imag} */,
  {32'hbf1a521a, 32'hbe6d4d90} /* (13, 13, 6) {real, imag} */,
  {32'hbfc71aa6, 32'hbe75dbe1} /* (13, 13, 5) {real, imag} */,
  {32'hbf085865, 32'h3ee62132} /* (13, 13, 4) {real, imag} */,
  {32'h3f44fdaa, 32'h3d10f910} /* (13, 13, 3) {real, imag} */,
  {32'h3f0f92fc, 32'hbe099704} /* (13, 13, 2) {real, imag} */,
  {32'h3f5feb97, 32'hbf404bb8} /* (13, 13, 1) {real, imag} */,
  {32'hbf0f5639, 32'hbeaef546} /* (13, 13, 0) {real, imag} */,
  {32'hbeb2d7dc, 32'h3f0a0869} /* (13, 12, 15) {real, imag} */,
  {32'h3eba97a7, 32'hbe2def36} /* (13, 12, 14) {real, imag} */,
  {32'hbf57ca84, 32'h3ea97e67} /* (13, 12, 13) {real, imag} */,
  {32'hbf627d58, 32'h3f8a4c2d} /* (13, 12, 12) {real, imag} */,
  {32'h3faaa4c6, 32'h3f93f3dc} /* (13, 12, 11) {real, imag} */,
  {32'hbf31f822, 32'h3f1bf634} /* (13, 12, 10) {real, imag} */,
  {32'hc025dcd2, 32'h3ef4ff7c} /* (13, 12, 9) {real, imag} */,
  {32'hbf885a9b, 32'hbf37a20a} /* (13, 12, 8) {real, imag} */,
  {32'h3f898306, 32'hbfd575e5} /* (13, 12, 7) {real, imag} */,
  {32'h3e6b88f8, 32'hc00796d0} /* (13, 12, 6) {real, imag} */,
  {32'hbf7206e8, 32'hbfadf80a} /* (13, 12, 5) {real, imag} */,
  {32'h3e9e3926, 32'h3f0c766e} /* (13, 12, 4) {real, imag} */,
  {32'h3fc6b56a, 32'h3f9b5b71} /* (13, 12, 3) {real, imag} */,
  {32'h3fd9d638, 32'h3d8ea3a8} /* (13, 12, 2) {real, imag} */,
  {32'h3f81d7a0, 32'hbf524b23} /* (13, 12, 1) {real, imag} */,
  {32'h3f18590f, 32'h3e89f79f} /* (13, 12, 0) {real, imag} */,
  {32'h3e5f3fb4, 32'h3ee6c7f6} /* (13, 11, 15) {real, imag} */,
  {32'hbdd84353, 32'h3f101f09} /* (13, 11, 14) {real, imag} */,
  {32'hbfc6d120, 32'h3fd61516} /* (13, 11, 13) {real, imag} */,
  {32'h3f3805c2, 32'h3ff8c328} /* (13, 11, 12) {real, imag} */,
  {32'h3e9b33eb, 32'h3fa30f52} /* (13, 11, 11) {real, imag} */,
  {32'hbf09fc4f, 32'h3ea3e6f8} /* (13, 11, 10) {real, imag} */,
  {32'hbfb8c620, 32'hbe4d61ca} /* (13, 11, 9) {real, imag} */,
  {32'hbf99774b, 32'h3f4b5ab9} /* (13, 11, 8) {real, imag} */,
  {32'h3fc3737a, 32'hbf16b924} /* (13, 11, 7) {real, imag} */,
  {32'h404890c1, 32'hc0192b50} /* (13, 11, 6) {real, imag} */,
  {32'h3fa7488d, 32'hc003bc2a} /* (13, 11, 5) {real, imag} */,
  {32'hbe48f41e, 32'hbfb26456} /* (13, 11, 4) {real, imag} */,
  {32'h3de31b9c, 32'hbe020175} /* (13, 11, 3) {real, imag} */,
  {32'h3f663014, 32'hbf4217f8} /* (13, 11, 2) {real, imag} */,
  {32'h3f93d43c, 32'hbe891de8} /* (13, 11, 1) {real, imag} */,
  {32'h3efb30de, 32'h3ea5890a} /* (13, 11, 0) {real, imag} */,
  {32'h3ef52c31, 32'h3f3da638} /* (13, 10, 15) {real, imag} */,
  {32'h3f76cb93, 32'h3db0b498} /* (13, 10, 14) {real, imag} */,
  {32'hbf3af132, 32'h3f43ace2} /* (13, 10, 13) {real, imag} */,
  {32'h3e106aa8, 32'h3fe86621} /* (13, 10, 12) {real, imag} */,
  {32'hbdaf5fcf, 32'h3fd18d78} /* (13, 10, 11) {real, imag} */,
  {32'h3e86a026, 32'h3fd472e6} /* (13, 10, 10) {real, imag} */,
  {32'h3ec97cda, 32'h3fa13028} /* (13, 10, 9) {real, imag} */,
  {32'h3f3cd786, 32'h3e835b6a} /* (13, 10, 8) {real, imag} */,
  {32'h3fda06b8, 32'hbec9e9e5} /* (13, 10, 7) {real, imag} */,
  {32'h3f6fe303, 32'h3e5b90a3} /* (13, 10, 6) {real, imag} */,
  {32'h3f8f8136, 32'hbeb98274} /* (13, 10, 5) {real, imag} */,
  {32'h3f708ece, 32'hbf2b358c} /* (13, 10, 4) {real, imag} */,
  {32'h3f1d5f10, 32'h3efb579e} /* (13, 10, 3) {real, imag} */,
  {32'h3f8f02a8, 32'hbe21b98c} /* (13, 10, 2) {real, imag} */,
  {32'h3f5f7551, 32'hbedd083c} /* (13, 10, 1) {real, imag} */,
  {32'hbe9594de, 32'hbef770bf} /* (13, 10, 0) {real, imag} */,
  {32'h3ed035cc, 32'h3fbac715} /* (13, 9, 15) {real, imag} */,
  {32'hbf5d5292, 32'h3f3728f6} /* (13, 9, 14) {real, imag} */,
  {32'hbf6c6445, 32'hbc28d420} /* (13, 9, 13) {real, imag} */,
  {32'hbf134b6b, 32'h401bf926} /* (13, 9, 12) {real, imag} */,
  {32'h3f027c18, 32'h400b64b9} /* (13, 9, 11) {real, imag} */,
  {32'h3fd042f8, 32'h3fe4d605} /* (13, 9, 10) {real, imag} */,
  {32'h40052cf4, 32'h400df8cf} /* (13, 9, 9) {real, imag} */,
  {32'h3f73eb8a, 32'hbec430f7} /* (13, 9, 8) {real, imag} */,
  {32'h3fac0153, 32'hbed4bd3a} /* (13, 9, 7) {real, imag} */,
  {32'hbf383f96, 32'h3fba9a10} /* (13, 9, 6) {real, imag} */,
  {32'hbfd17e04, 32'h3fd2395e} /* (13, 9, 5) {real, imag} */,
  {32'hbf02fcca, 32'h3f892e6c} /* (13, 9, 4) {real, imag} */,
  {32'hbdf84e6c, 32'h3eabf526} /* (13, 9, 3) {real, imag} */,
  {32'h3fb7de8d, 32'h3ebf957e} /* (13, 9, 2) {real, imag} */,
  {32'h3f96a043, 32'h3f06e0df} /* (13, 9, 1) {real, imag} */,
  {32'h3d8f95eb, 32'hbf56c565} /* (13, 9, 0) {real, imag} */,
  {32'h3fd51aaf, 32'h3dff28e2} /* (13, 8, 15) {real, imag} */,
  {32'hbdd0749f, 32'h3f45090e} /* (13, 8, 14) {real, imag} */,
  {32'hc0086eca, 32'h3df0b494} /* (13, 8, 13) {real, imag} */,
  {32'hc000ed25, 32'h3f9bc008} /* (13, 8, 12) {real, imag} */,
  {32'hbf31b9e4, 32'h3f671a49} /* (13, 8, 11) {real, imag} */,
  {32'h3f7e6ac4, 32'h3e8f54cc} /* (13, 8, 10) {real, imag} */,
  {32'h3f8858b8, 32'h3f55987d} /* (13, 8, 9) {real, imag} */,
  {32'hbf4e905c, 32'h3f3705ce} /* (13, 8, 8) {real, imag} */,
  {32'h3d871ce8, 32'h3e9e52fd} /* (13, 8, 7) {real, imag} */,
  {32'hbfd66200, 32'hbec0c640} /* (13, 8, 6) {real, imag} */,
  {32'hbf6f0bcc, 32'hbf2f8feb} /* (13, 8, 5) {real, imag} */,
  {32'h3ebe4f7e, 32'h3e8d69f4} /* (13, 8, 4) {real, imag} */,
  {32'h3f2b17f4, 32'h3f8ccb3d} /* (13, 8, 3) {real, imag} */,
  {32'h3fd7bdce, 32'h3ececd90} /* (13, 8, 2) {real, imag} */,
  {32'h3f88d2ac, 32'hbed8f95c} /* (13, 8, 1) {real, imag} */,
  {32'h3f68b058, 32'hbe97b013} /* (13, 8, 0) {real, imag} */,
  {32'h3fa870ea, 32'hbffcde20} /* (13, 7, 15) {real, imag} */,
  {32'h3f9522f4, 32'hc020f5a4} /* (13, 7, 14) {real, imag} */,
  {32'hc0008905, 32'hbf477280} /* (13, 7, 13) {real, imag} */,
  {32'hc04e711e, 32'h3f40247a} /* (13, 7, 12) {real, imag} */,
  {32'hc00ad2c0, 32'h401f2ee8} /* (13, 7, 11) {real, imag} */,
  {32'hbea66ac6, 32'h3f4594f9} /* (13, 7, 10) {real, imag} */,
  {32'hbfa82638, 32'hbfa7813a} /* (13, 7, 9) {real, imag} */,
  {32'hbfaee6a9, 32'h3e500d72} /* (13, 7, 8) {real, imag} */,
  {32'h3dd1b060, 32'h3e9d15f0} /* (13, 7, 7) {real, imag} */,
  {32'hbf95d224, 32'hbf99a5da} /* (13, 7, 6) {real, imag} */,
  {32'hbd6eef2c, 32'hc000ab89} /* (13, 7, 5) {real, imag} */,
  {32'h3fa16720, 32'hbf0ad65c} /* (13, 7, 4) {real, imag} */,
  {32'h3fd6320b, 32'h3f71cbab} /* (13, 7, 3) {real, imag} */,
  {32'h3fdc104e, 32'h3f65edc4} /* (13, 7, 2) {real, imag} */,
  {32'h3fdb1d92, 32'h3f8318ea} /* (13, 7, 1) {real, imag} */,
  {32'h3fdaa221, 32'h3f9a446c} /* (13, 7, 0) {real, imag} */,
  {32'h3e93aa27, 32'hbfec3b6b} /* (13, 6, 15) {real, imag} */,
  {32'h3f73a43c, 32'hbfe29afa} /* (13, 6, 14) {real, imag} */,
  {32'hbbae8f80, 32'h3e99916f} /* (13, 6, 13) {real, imag} */,
  {32'hbfba2bef, 32'h3e0e5454} /* (13, 6, 12) {real, imag} */,
  {32'hbf4099f4, 32'h3fbd3074} /* (13, 6, 11) {real, imag} */,
  {32'hbd2d0f88, 32'h3f363cbb} /* (13, 6, 10) {real, imag} */,
  {32'hbf19a4f7, 32'hbf06f904} /* (13, 6, 9) {real, imag} */,
  {32'h3f0b8b91, 32'h3f66abe7} /* (13, 6, 8) {real, imag} */,
  {32'h3f63ccf2, 32'h3fa87c34} /* (13, 6, 7) {real, imag} */,
  {32'hbf0c54eb, 32'hbf3ff70d} /* (13, 6, 6) {real, imag} */,
  {32'hbf14fdc1, 32'hbf1768a0} /* (13, 6, 5) {real, imag} */,
  {32'h3ebd6aef, 32'h3e433508} /* (13, 6, 4) {real, imag} */,
  {32'h3ea21a5d, 32'h3da658a6} /* (13, 6, 3) {real, imag} */,
  {32'hbea6803e, 32'h3f48ad38} /* (13, 6, 2) {real, imag} */,
  {32'hbf7c5ddd, 32'h3f80523c} /* (13, 6, 1) {real, imag} */,
  {32'h3f71fdbc, 32'h3fa94afa} /* (13, 6, 0) {real, imag} */,
  {32'h3d880957, 32'hbf99df1e} /* (13, 5, 15) {real, imag} */,
  {32'hbd950430, 32'hbfb96916} /* (13, 5, 14) {real, imag} */,
  {32'hbd43a00c, 32'h3f5f908b} /* (13, 5, 13) {real, imag} */,
  {32'hbee7949a, 32'hbe1a3d52} /* (13, 5, 12) {real, imag} */,
  {32'h3dc8977c, 32'hbed66ba5} /* (13, 5, 11) {real, imag} */,
  {32'hbf3b8359, 32'hbec9a849} /* (13, 5, 10) {real, imag} */,
  {32'hbe6ccacb, 32'h3db0b4ac} /* (13, 5, 9) {real, imag} */,
  {32'h3fb58e06, 32'h3eddd51f} /* (13, 5, 8) {real, imag} */,
  {32'h3f868818, 32'h3f993e50} /* (13, 5, 7) {real, imag} */,
  {32'h3d2d5420, 32'hbf548208} /* (13, 5, 6) {real, imag} */,
  {32'h3e44ced4, 32'hbf5511fa} /* (13, 5, 5) {real, imag} */,
  {32'hbede7381, 32'h3f8c8ecf} /* (13, 5, 4) {real, imag} */,
  {32'hbf0cca08, 32'h3ebf178c} /* (13, 5, 3) {real, imag} */,
  {32'h3e131094, 32'h3f18aad0} /* (13, 5, 2) {real, imag} */,
  {32'hbfd6463e, 32'h3f962a94} /* (13, 5, 1) {real, imag} */,
  {32'h3e19ea8c, 32'h3f5aa2d9} /* (13, 5, 0) {real, imag} */,
  {32'h3fada26b, 32'hbf1a5337} /* (13, 4, 15) {real, imag} */,
  {32'h3f48e533, 32'h3e800d63} /* (13, 4, 14) {real, imag} */,
  {32'hbf5a3b7a, 32'h4009941b} /* (13, 4, 13) {real, imag} */,
  {32'hbfe86c1b, 32'h3f583ce8} /* (13, 4, 12) {real, imag} */,
  {32'hbf1f3758, 32'hbe9d1d8a} /* (13, 4, 11) {real, imag} */,
  {32'h3e36bf38, 32'h3e7585b0} /* (13, 4, 10) {real, imag} */,
  {32'h3e216334, 32'h3f8ef188} /* (13, 4, 9) {real, imag} */,
  {32'hbf2ff4ef, 32'h3fac56f1} /* (13, 4, 8) {real, imag} */,
  {32'hbe40ecd6, 32'h3ffdd3b6} /* (13, 4, 7) {real, imag} */,
  {32'h3ef4fe4e, 32'h3e08ae0a} /* (13, 4, 6) {real, imag} */,
  {32'h3fabc333, 32'h3e82f84e} /* (13, 4, 5) {real, imag} */,
  {32'h3d1354f8, 32'h3f3f7a1e} /* (13, 4, 4) {real, imag} */,
  {32'hbf562822, 32'h3eb1d948} /* (13, 4, 3) {real, imag} */,
  {32'h3fe0ea4b, 32'h3e8f3890} /* (13, 4, 2) {real, imag} */,
  {32'h3f179430, 32'h3fc1c1dc} /* (13, 4, 1) {real, imag} */,
  {32'h3e577a66, 32'h3e902fa6} /* (13, 4, 0) {real, imag} */,
  {32'h3eae2783, 32'h3e6ea7d8} /* (13, 3, 15) {real, imag} */,
  {32'h3f9b861e, 32'h3fdd582e} /* (13, 3, 14) {real, imag} */,
  {32'h3e93fda6, 32'h4054652b} /* (13, 3, 13) {real, imag} */,
  {32'hc03696e4, 32'h3f918fb6} /* (13, 3, 12) {real, imag} */,
  {32'hbdae2170, 32'h3f859f22} /* (13, 3, 11) {real, imag} */,
  {32'h3f9c8fe2, 32'h3f4f259a} /* (13, 3, 10) {real, imag} */,
  {32'h3d7b4a90, 32'hbec95576} /* (13, 3, 9) {real, imag} */,
  {32'hbf46a273, 32'h3ec37596} /* (13, 3, 8) {real, imag} */,
  {32'hbe000ebe, 32'h3f9868d2} /* (13, 3, 7) {real, imag} */,
  {32'hbd816022, 32'h3e7e1674} /* (13, 3, 6) {real, imag} */,
  {32'hbedde78c, 32'h3dd2a8b0} /* (13, 3, 5) {real, imag} */,
  {32'hbf026c31, 32'h3f7ac925} /* (13, 3, 4) {real, imag} */,
  {32'hbf15fd00, 32'h3f3654e4} /* (13, 3, 3) {real, imag} */,
  {32'hbed329d2, 32'h3ea4cb99} /* (13, 3, 2) {real, imag} */,
  {32'hbf34e08f, 32'hbec60f8e} /* (13, 3, 1) {real, imag} */,
  {32'hbf436138, 32'hbf98db1d} /* (13, 3, 0) {real, imag} */,
  {32'hbfff2944, 32'h3e80c2d7} /* (13, 2, 15) {real, imag} */,
  {32'hbfdf29df, 32'h3ec8a61d} /* (13, 2, 14) {real, imag} */,
  {32'h3ef26ea2, 32'h3f6a04d2} /* (13, 2, 13) {real, imag} */,
  {32'hbfc4cd3e, 32'h3edb81c6} /* (13, 2, 12) {real, imag} */,
  {32'h3f97fbbe, 32'h3f36199b} /* (13, 2, 11) {real, imag} */,
  {32'h3ee105af, 32'hbf40d91b} /* (13, 2, 10) {real, imag} */,
  {32'h3f31fe3a, 32'hbf30e112} /* (13, 2, 9) {real, imag} */,
  {32'h3fc14da9, 32'hbf9911f2} /* (13, 2, 8) {real, imag} */,
  {32'h3fbb112a, 32'h3f8b11b6} /* (13, 2, 7) {real, imag} */,
  {32'hbef682fb, 32'h3fbe637e} /* (13, 2, 6) {real, imag} */,
  {32'h3f73aff0, 32'h3eb05294} /* (13, 2, 5) {real, imag} */,
  {32'h4000d7fb, 32'h3f73bbc3} /* (13, 2, 4) {real, imag} */,
  {32'h3f069f0e, 32'h3fac55a4} /* (13, 2, 3) {real, imag} */,
  {32'hbf96bd90, 32'hbe402898} /* (13, 2, 2) {real, imag} */,
  {32'hbf847fe1, 32'hbf8b179f} /* (13, 2, 1) {real, imag} */,
  {32'hbf3e00e1, 32'hbf68fae8} /* (13, 2, 0) {real, imag} */,
  {32'hbf531714, 32'hbe7bff2a} /* (13, 1, 15) {real, imag} */,
  {32'hbe9681a8, 32'hbf84cdb8} /* (13, 1, 14) {real, imag} */,
  {32'hbe953f79, 32'hbdc56ee2} /* (13, 1, 13) {real, imag} */,
  {32'hbfbd9459, 32'h3eab28cc} /* (13, 1, 12) {real, imag} */,
  {32'h3f0b1416, 32'hbf082cde} /* (13, 1, 11) {real, imag} */,
  {32'h3f89f7ca, 32'hbf8a403a} /* (13, 1, 10) {real, imag} */,
  {32'hbe4e9000, 32'hbf2cc8a6} /* (13, 1, 9) {real, imag} */,
  {32'h3f57cff2, 32'hbf8c20d4} /* (13, 1, 8) {real, imag} */,
  {32'h3f74a6c0, 32'h3f9ba6e4} /* (13, 1, 7) {real, imag} */,
  {32'hbd95c6b4, 32'h3ffdfef8} /* (13, 1, 6) {real, imag} */,
  {32'h3fce6f02, 32'h4018843d} /* (13, 1, 5) {real, imag} */,
  {32'h40488770, 32'h3fa35e16} /* (13, 1, 4) {real, imag} */,
  {32'h3f293737, 32'h3e5a25e8} /* (13, 1, 3) {real, imag} */,
  {32'hbf8ef69b, 32'h3cc2c780} /* (13, 1, 2) {real, imag} */,
  {32'h3f79838a, 32'h3d06464c} /* (13, 1, 1) {real, imag} */,
  {32'h3f0a4d76, 32'hbc276180} /* (13, 1, 0) {real, imag} */,
  {32'h3e96f50b, 32'hbeacbe7a} /* (13, 0, 15) {real, imag} */,
  {32'h3e2e447a, 32'hbf3d6357} /* (13, 0, 14) {real, imag} */,
  {32'hbfd75e62, 32'hbeaeb59e} /* (13, 0, 13) {real, imag} */,
  {32'hbfe48532, 32'h3f209999} /* (13, 0, 12) {real, imag} */,
  {32'hbdb507de, 32'h3e601922} /* (13, 0, 11) {real, imag} */,
  {32'h3ead8b8a, 32'hbdc1ce38} /* (13, 0, 10) {real, imag} */,
  {32'hbfa9d2b3, 32'h3f354bbe} /* (13, 0, 9) {real, imag} */,
  {32'hbf4b1776, 32'h3c144f5c} /* (13, 0, 8) {real, imag} */,
  {32'h3f0ab1fd, 32'h3f1d7a4f} /* (13, 0, 7) {real, imag} */,
  {32'hbeb50a17, 32'h3f34648a} /* (13, 0, 6) {real, imag} */,
  {32'hbee87adb, 32'h3f42c21e} /* (13, 0, 5) {real, imag} */,
  {32'h3eb0d11d, 32'h3e95dbab} /* (13, 0, 4) {real, imag} */,
  {32'h3cd8235c, 32'h3de7e9b0} /* (13, 0, 3) {real, imag} */,
  {32'hbf480586, 32'h3f4e5bdb} /* (13, 0, 2) {real, imag} */,
  {32'h3d3f59f0, 32'h3f404374} /* (13, 0, 1) {real, imag} */,
  {32'h3ee47f0c, 32'h3ebbfb0a} /* (13, 0, 0) {real, imag} */,
  {32'h3e2db84c, 32'hbefc10c2} /* (12, 15, 15) {real, imag} */,
  {32'h3c2c5490, 32'hbe1481e6} /* (12, 15, 14) {real, imag} */,
  {32'hbd9569d0, 32'h3d6a3788} /* (12, 15, 13) {real, imag} */,
  {32'h3eb1c1b4, 32'h3e8e9974} /* (12, 15, 12) {real, imag} */,
  {32'h3e97268d, 32'hbf0cda53} /* (12, 15, 11) {real, imag} */,
  {32'hbf33a30b, 32'hbf435b32} /* (12, 15, 10) {real, imag} */,
  {32'hbec2a720, 32'hbef50946} /* (12, 15, 9) {real, imag} */,
  {32'hbf2b0926, 32'h3e91f5a0} /* (12, 15, 8) {real, imag} */,
  {32'hbf8c7b14, 32'h3d59dc3c} /* (12, 15, 7) {real, imag} */,
  {32'hbdffb4e5, 32'hbefa3dc9} /* (12, 15, 6) {real, imag} */,
  {32'h3e8d8577, 32'h3b30e700} /* (12, 15, 5) {real, imag} */,
  {32'h3f83f65b, 32'h3f4d97dd} /* (12, 15, 4) {real, imag} */,
  {32'h3fd20bee, 32'h3e972cf7} /* (12, 15, 3) {real, imag} */,
  {32'h3f44c595, 32'h3edf88a8} /* (12, 15, 2) {real, imag} */,
  {32'h3f0c9136, 32'h3f15c9b4} /* (12, 15, 1) {real, imag} */,
  {32'h3e7e7fdb, 32'h3f66f0d8} /* (12, 15, 0) {real, imag} */,
  {32'hbe2b379c, 32'hbf3632ae} /* (12, 14, 15) {real, imag} */,
  {32'hbf5f24ea, 32'h3eaa1e17} /* (12, 14, 14) {real, imag} */,
  {32'hbf85c1bd, 32'h3f205c5b} /* (12, 14, 13) {real, imag} */,
  {32'hbdf5e958, 32'h3ed2900a} /* (12, 14, 12) {real, imag} */,
  {32'h3e90aef6, 32'hbf3c2666} /* (12, 14, 11) {real, imag} */,
  {32'hbff2dec1, 32'hbeaefb8a} /* (12, 14, 10) {real, imag} */,
  {32'hbf36cb64, 32'h3bf84f80} /* (12, 14, 9) {real, imag} */,
  {32'hbf4889a4, 32'hbf634fbc} /* (12, 14, 8) {real, imag} */,
  {32'hbf871877, 32'hbcb1b080} /* (12, 14, 7) {real, imag} */,
  {32'h3e49679c, 32'h3f084efe} /* (12, 14, 6) {real, imag} */,
  {32'h3e561e06, 32'h3e025bb8} /* (12, 14, 5) {real, imag} */,
  {32'h3ee518f4, 32'hbeccae62} /* (12, 14, 4) {real, imag} */,
  {32'h3fb8d18b, 32'hbfe268c4} /* (12, 14, 3) {real, imag} */,
  {32'h3fd70201, 32'hbfe43ddb} /* (12, 14, 2) {real, imag} */,
  {32'h3f893ed7, 32'h3e3a9221} /* (12, 14, 1) {real, imag} */,
  {32'h3e399382, 32'h3f60923f} /* (12, 14, 0) {real, imag} */,
  {32'hbf2be4fe, 32'hbf15cf38} /* (12, 13, 15) {real, imag} */,
  {32'hbf6ac1ca, 32'hbf0253ae} /* (12, 13, 14) {real, imag} */,
  {32'h3d645c60, 32'hbe85ca4c} /* (12, 13, 13) {real, imag} */,
  {32'h3f9c8320, 32'hbf6ea84a} /* (12, 13, 12) {real, imag} */,
  {32'hba5afe00, 32'hbf0d2bb2} /* (12, 13, 11) {real, imag} */,
  {32'hbf540a86, 32'hbcd4ca20} /* (12, 13, 10) {real, imag} */,
  {32'h3f01691a, 32'hbf08e92a} /* (12, 13, 9) {real, imag} */,
  {32'hbdabcbe2, 32'hbfb5a7cd} /* (12, 13, 8) {real, imag} */,
  {32'hbf7e18c3, 32'hbfa9a0a0} /* (12, 13, 7) {real, imag} */,
  {32'hbef736ba, 32'hbf88a3d4} /* (12, 13, 6) {real, imag} */,
  {32'h3f44881c, 32'hbf79e769} /* (12, 13, 5) {real, imag} */,
  {32'h3f550071, 32'hbfd63ef0} /* (12, 13, 4) {real, imag} */,
  {32'h3f1fb0d0, 32'hbfb9dd7e} /* (12, 13, 3) {real, imag} */,
  {32'h3f85d2dd, 32'hbf986a33} /* (12, 13, 2) {real, imag} */,
  {32'hbe267152, 32'hbfd795f6} /* (12, 13, 1) {real, imag} */,
  {32'hbedfbd90, 32'hbf17ce74} /* (12, 13, 0) {real, imag} */,
  {32'hbe99c727, 32'hbf006ad4} /* (12, 12, 15) {real, imag} */,
  {32'h3f0f994b, 32'hbdfa7c0c} /* (12, 12, 14) {real, imag} */,
  {32'h3f89d34b, 32'hbeaab8b0} /* (12, 12, 13) {real, imag} */,
  {32'h3fb4e1bd, 32'hbf82ebf8} /* (12, 12, 12) {real, imag} */,
  {32'h3f460d2c, 32'hbe222d0e} /* (12, 12, 11) {real, imag} */,
  {32'h3f1689de, 32'h3e2eca0c} /* (12, 12, 10) {real, imag} */,
  {32'h3cbe2748, 32'h3ddaabb0} /* (12, 12, 9) {real, imag} */,
  {32'hbfdb5c37, 32'hbe880129} /* (12, 12, 8) {real, imag} */,
  {32'hbfd058fa, 32'hbfb9ee4c} /* (12, 12, 7) {real, imag} */,
  {32'hbfbe932f, 32'hc0012964} /* (12, 12, 6) {real, imag} */,
  {32'hbe83991c, 32'hbf882527} /* (12, 12, 5) {real, imag} */,
  {32'hbef633f1, 32'hbed1a3f7} /* (12, 12, 4) {real, imag} */,
  {32'h3ef08cff, 32'hbe7fdabe} /* (12, 12, 3) {real, imag} */,
  {32'h3f2b2452, 32'hbf592b9e} /* (12, 12, 2) {real, imag} */,
  {32'hbd4d6df0, 32'hbf3b1521} /* (12, 12, 1) {real, imag} */,
  {32'h3cccf7d0, 32'hbf8ad4e9} /* (12, 12, 0) {real, imag} */,
  {32'hbf276ff9, 32'hbd812bbc} /* (12, 11, 15) {real, imag} */,
  {32'hbfb5dd31, 32'h3d23d5e0} /* (12, 11, 14) {real, imag} */,
  {32'hbe7b7ce0, 32'hbe95d954} /* (12, 11, 13) {real, imag} */,
  {32'hbf09a4b5, 32'hbdcb2510} /* (12, 11, 12) {real, imag} */,
  {32'h3d66df68, 32'h3c5e1fc0} /* (12, 11, 11) {real, imag} */,
  {32'h3faa73e6, 32'h3bb8b0c0} /* (12, 11, 10) {real, imag} */,
  {32'h3e9e1942, 32'h3f15ea14} /* (12, 11, 9) {real, imag} */,
  {32'hbf67276a, 32'hba6fcc40} /* (12, 11, 8) {real, imag} */,
  {32'h3f43a820, 32'hbf7da5b2} /* (12, 11, 7) {real, imag} */,
  {32'h3e5951c4, 32'hbf23e1ba} /* (12, 11, 6) {real, imag} */,
  {32'hbf641712, 32'hbf4a0153} /* (12, 11, 5) {real, imag} */,
  {32'hbffbef5e, 32'hbf03c71c} /* (12, 11, 4) {real, imag} */,
  {32'hbf7cbf5d, 32'hbf380cb3} /* (12, 11, 3) {real, imag} */,
  {32'h3e039c70, 32'hbf9cfc99} /* (12, 11, 2) {real, imag} */,
  {32'h3d0ab1d4, 32'h3e0ada10} /* (12, 11, 1) {real, imag} */,
  {32'h3e0a71b2, 32'hbf20025c} /* (12, 11, 0) {real, imag} */,
  {32'hbfa78195, 32'h3e1ae552} /* (12, 10, 15) {real, imag} */,
  {32'hbfef41fa, 32'h3f2e01c0} /* (12, 10, 14) {real, imag} */,
  {32'h3f82d79e, 32'h3d83b52c} /* (12, 10, 13) {real, imag} */,
  {32'h3e97e68d, 32'hbd8fa4b4} /* (12, 10, 12) {real, imag} */,
  {32'h3eb646ae, 32'hbea9d408} /* (12, 10, 11) {real, imag} */,
  {32'h3fa174dd, 32'hbf9ad41d} /* (12, 10, 10) {real, imag} */,
  {32'h3f74d434, 32'h3f795db3} /* (12, 10, 9) {real, imag} */,
  {32'h3eba4749, 32'h3f4b2c4d} /* (12, 10, 8) {real, imag} */,
  {32'hbdfbda50, 32'hbf391641} /* (12, 10, 7) {real, imag} */,
  {32'h3bdbd380, 32'h3ed7b3a0} /* (12, 10, 6) {real, imag} */,
  {32'hbfbecd7c, 32'hbfaa7389} /* (12, 10, 5) {real, imag} */,
  {32'hc001dbc0, 32'hbfd73b6c} /* (12, 10, 4) {real, imag} */,
  {32'hbf9ffb62, 32'hbec4bab7} /* (12, 10, 3) {real, imag} */,
  {32'hbf3d4196, 32'hbf37fdb9} /* (12, 10, 2) {real, imag} */,
  {32'hbf512517, 32'hbedc8f5f} /* (12, 10, 1) {real, imag} */,
  {32'hbf2408da, 32'hbe3de8d4} /* (12, 10, 0) {real, imag} */,
  {32'hbfbe2f69, 32'h3f75fcf2} /* (12, 9, 15) {real, imag} */,
  {32'hbfb8a0ee, 32'h3feadec5} /* (12, 9, 14) {real, imag} */,
  {32'h3e9040b6, 32'h3f1b4d21} /* (12, 9, 13) {real, imag} */,
  {32'hbea3cd44, 32'hbf123cb5} /* (12, 9, 12) {real, imag} */,
  {32'hbf613a74, 32'hbeee9847} /* (12, 9, 11) {real, imag} */,
  {32'hbeb75c20, 32'h3dcc0c20} /* (12, 9, 10) {real, imag} */,
  {32'hbf42ca87, 32'h3f2aa217} /* (12, 9, 9) {real, imag} */,
  {32'hbfe219e4, 32'h3f1cde3c} /* (12, 9, 8) {real, imag} */,
  {32'hbf8d1357, 32'h3f0807bf} /* (12, 9, 7) {real, imag} */,
  {32'h3f3de74a, 32'h3e75df64} /* (12, 9, 6) {real, imag} */,
  {32'hbf5b709e, 32'h3f08ffba} /* (12, 9, 5) {real, imag} */,
  {32'hbfb09a76, 32'h3d9c8d98} /* (12, 9, 4) {real, imag} */,
  {32'hbfcddf16, 32'h3efbfd0f} /* (12, 9, 3) {real, imag} */,
  {32'hbf291a6f, 32'h3f37bcea} /* (12, 9, 2) {real, imag} */,
  {32'h3e759948, 32'hbefda74a} /* (12, 9, 1) {real, imag} */,
  {32'hbea9d348, 32'h3ef72fb8} /* (12, 9, 0) {real, imag} */,
  {32'hbf829a10, 32'h3e42d8d8} /* (12, 8, 15) {real, imag} */,
  {32'hbf81c347, 32'h3f072f61} /* (12, 8, 14) {real, imag} */,
  {32'hbe173f5b, 32'hbd274448} /* (12, 8, 13) {real, imag} */,
  {32'h3ee37386, 32'h3e98f4c4} /* (12, 8, 12) {real, imag} */,
  {32'hbf903e8a, 32'hbe9a8aa1} /* (12, 8, 11) {real, imag} */,
  {32'hbf9d9524, 32'h3d42b0a6} /* (12, 8, 10) {real, imag} */,
  {32'hbff19486, 32'hbefce0b8} /* (12, 8, 9) {real, imag} */,
  {32'hc0061b0d, 32'h3ed690d9} /* (12, 8, 8) {real, imag} */,
  {32'hbfb32e19, 32'h3f9b9ed0} /* (12, 8, 7) {real, imag} */,
  {32'h3f4c434f, 32'hbf45c20d} /* (12, 8, 6) {real, imag} */,
  {32'hbe99d14f, 32'h3e69bd65} /* (12, 8, 5) {real, imag} */,
  {32'hc0092af7, 32'h3f0a0ca6} /* (12, 8, 4) {real, imag} */,
  {32'hc00e9740, 32'h3f01856a} /* (12, 8, 3) {real, imag} */,
  {32'hbe1c5f5a, 32'h3feb502a} /* (12, 8, 2) {real, imag} */,
  {32'h3fd67e76, 32'h3f2059ac} /* (12, 8, 1) {real, imag} */,
  {32'h3f83d8ea, 32'h3ee1a675} /* (12, 8, 0) {real, imag} */,
  {32'hbfb0a214, 32'hbe5ae239} /* (12, 7, 15) {real, imag} */,
  {32'hbf611cee, 32'h3eb8a452} /* (12, 7, 14) {real, imag} */,
  {32'hbe1740d0, 32'h3f89cf06} /* (12, 7, 13) {real, imag} */,
  {32'h3fd93d70, 32'h3fbc2860} /* (12, 7, 12) {real, imag} */,
  {32'h3dc85940, 32'hbf3fabcf} /* (12, 7, 11) {real, imag} */,
  {32'h3ea7c92a, 32'hbf81776b} /* (12, 7, 10) {real, imag} */,
  {32'h3f517032, 32'hbf43d80c} /* (12, 7, 9) {real, imag} */,
  {32'h3e9f5b82, 32'h3f185156} /* (12, 7, 8) {real, imag} */,
  {32'hbd9799d1, 32'h3f531438} /* (12, 7, 7) {real, imag} */,
  {32'h3f5a6355, 32'hbe2a56d6} /* (12, 7, 6) {real, imag} */,
  {32'h3e9b769e, 32'h3f656fe2} /* (12, 7, 5) {real, imag} */,
  {32'hbf927714, 32'h3f511f78} /* (12, 7, 4) {real, imag} */,
  {32'hbfb275a3, 32'h3ed4d2f0} /* (12, 7, 3) {real, imag} */,
  {32'hbec5da7c, 32'h3fac586e} /* (12, 7, 2) {real, imag} */,
  {32'hbdfc5644, 32'h401e8224} /* (12, 7, 1) {real, imag} */,
  {32'hbee7bcfb, 32'h3f9d8e26} /* (12, 7, 0) {real, imag} */,
  {32'hbf96189d, 32'h3f48fee3} /* (12, 6, 15) {real, imag} */,
  {32'hbf2f38e9, 32'h3fb9ab34} /* (12, 6, 14) {real, imag} */,
  {32'hbf57c8a0, 32'h3f9ac100} /* (12, 6, 13) {real, imag} */,
  {32'hbf88f430, 32'h3f6673e9} /* (12, 6, 12) {real, imag} */,
  {32'hbf329460, 32'hbe3fed50} /* (12, 6, 11) {real, imag} */,
  {32'hbf079191, 32'h3eea988c} /* (12, 6, 10) {real, imag} */,
  {32'h3df70488, 32'hbf56dbe2} /* (12, 6, 9) {real, imag} */,
  {32'h3ec0a670, 32'hbfa3525e} /* (12, 6, 8) {real, imag} */,
  {32'h3ea891d0, 32'hbe550600} /* (12, 6, 7) {real, imag} */,
  {32'h3f7d1002, 32'hbeb6a20b} /* (12, 6, 6) {real, imag} */,
  {32'h3fd2bfb7, 32'h3f5acaad} /* (12, 6, 5) {real, imag} */,
  {32'h3ef370b0, 32'h3f026f19} /* (12, 6, 4) {real, imag} */,
  {32'hbf610cb2, 32'hbf54fb79} /* (12, 6, 3) {real, imag} */,
  {32'hbf105bc6, 32'hbec324b4} /* (12, 6, 2) {real, imag} */,
  {32'hbf6aaa9f, 32'h3f6f240c} /* (12, 6, 1) {real, imag} */,
  {32'hbf960188, 32'h3fa8c918} /* (12, 6, 0) {real, imag} */,
  {32'h3dfbcf42, 32'h3eb18378} /* (12, 5, 15) {real, imag} */,
  {32'h3e914391, 32'h3f277de5} /* (12, 5, 14) {real, imag} */,
  {32'h3f0591a2, 32'h3f32153d} /* (12, 5, 13) {real, imag} */,
  {32'h3f8ec92c, 32'h3f821724} /* (12, 5, 12) {real, imag} */,
  {32'h3e1518b4, 32'h3f80a313} /* (12, 5, 11) {real, imag} */,
  {32'h3e72ff44, 32'h3f1f417f} /* (12, 5, 10) {real, imag} */,
  {32'hbd5c0fd8, 32'hbfe6dee3} /* (12, 5, 9) {real, imag} */,
  {32'hbf04c262, 32'hbfafe750} /* (12, 5, 8) {real, imag} */,
  {32'h3f30c6f6, 32'hbf74e45f} /* (12, 5, 7) {real, imag} */,
  {32'h401255d6, 32'h3ec971a0} /* (12, 5, 6) {real, imag} */,
  {32'h3fd3cb10, 32'h3f4e47c5} /* (12, 5, 5) {real, imag} */,
  {32'h3f891d7c, 32'hbe008248} /* (12, 5, 4) {real, imag} */,
  {32'h3fc54433, 32'h3e0633c6} /* (12, 5, 3) {real, imag} */,
  {32'h3f853f1f, 32'h3da11ea4} /* (12, 5, 2) {real, imag} */,
  {32'hbef8012c, 32'hbf66de34} /* (12, 5, 1) {real, imag} */,
  {32'hbedb6e83, 32'h3ea6cacf} /* (12, 5, 0) {real, imag} */,
  {32'h3e9a900a, 32'h3e5cb90c} /* (12, 4, 15) {real, imag} */,
  {32'h3f36f6bb, 32'h3ebb2ec4} /* (12, 4, 14) {real, imag} */,
  {32'h3f72be92, 32'h3fa4d4c2} /* (12, 4, 13) {real, imag} */,
  {32'h3fff3832, 32'h3f5ea6b0} /* (12, 4, 12) {real, imag} */,
  {32'h3e0fc926, 32'hbdef1566} /* (12, 4, 11) {real, imag} */,
  {32'hbcbb30b0, 32'hbe455790} /* (12, 4, 10) {real, imag} */,
  {32'h3e2f4e02, 32'hbf7affef} /* (12, 4, 9) {real, imag} */,
  {32'hbf31c845, 32'hbf6e17c1} /* (12, 4, 8) {real, imag} */,
  {32'h3f6ed550, 32'hbca8c164} /* (12, 4, 7) {real, imag} */,
  {32'h3f8fdbb5, 32'h3e53155e} /* (12, 4, 6) {real, imag} */,
  {32'h3f81e64e, 32'hbefa31d2} /* (12, 4, 5) {real, imag} */,
  {32'h3f5b4871, 32'hbf97cf97} /* (12, 4, 4) {real, imag} */,
  {32'h3f8c41f4, 32'hbef4872f} /* (12, 4, 3) {real, imag} */,
  {32'h3dd2aa13, 32'h3f1dabe9} /* (12, 4, 2) {real, imag} */,
  {32'hbf97bae2, 32'h3ec7fd2a} /* (12, 4, 1) {real, imag} */,
  {32'hbf2c6ba4, 32'h3ec35f96} /* (12, 4, 0) {real, imag} */,
  {32'h3f46c29c, 32'hbd7e01c0} /* (12, 3, 15) {real, imag} */,
  {32'h3e79f676, 32'h3eedca6c} /* (12, 3, 14) {real, imag} */,
  {32'hbf81acf2, 32'h3fab834c} /* (12, 3, 13) {real, imag} */,
  {32'h3f962c2c, 32'h3f99a216} /* (12, 3, 12) {real, imag} */,
  {32'hbdba0458, 32'h3f1105ac} /* (12, 3, 11) {real, imag} */,
  {32'hbf526218, 32'hbe7b56e7} /* (12, 3, 10) {real, imag} */,
  {32'h3f12b25c, 32'h3f77381a} /* (12, 3, 9) {real, imag} */,
  {32'h3e9afaa4, 32'h3f013ba8} /* (12, 3, 8) {real, imag} */,
  {32'h4015346e, 32'h3ee0d228} /* (12, 3, 7) {real, imag} */,
  {32'h3fb1bf54, 32'hbfc71c78} /* (12, 3, 6) {real, imag} */,
  {32'h3ea709c7, 32'hc00a5373} /* (12, 3, 5) {real, imag} */,
  {32'h3f156c82, 32'hbfc44034} /* (12, 3, 4) {real, imag} */,
  {32'hbf1782d2, 32'hbf5aa594} /* (12, 3, 3) {real, imag} */,
  {32'hbfd6e0f3, 32'h3e114f5a} /* (12, 3, 2) {real, imag} */,
  {32'hbfd8b6d2, 32'h3f7f4fa6} /* (12, 3, 1) {real, imag} */,
  {32'hbfa26b3d, 32'h3f237df2} /* (12, 3, 0) {real, imag} */,
  {32'hbdf41a28, 32'hbe7107fc} /* (12, 2, 15) {real, imag} */,
  {32'hbf584b3a, 32'h3f2f389d} /* (12, 2, 14) {real, imag} */,
  {32'hbf93ddd2, 32'h3d19f0a0} /* (12, 2, 13) {real, imag} */,
  {32'hbd5fd4f0, 32'hbe9f0614} /* (12, 2, 12) {real, imag} */,
  {32'h3e7cbfe4, 32'h3e0b27c4} /* (12, 2, 11) {real, imag} */,
  {32'hbdf98840, 32'hbf686d30} /* (12, 2, 10) {real, imag} */,
  {32'h3f622f9c, 32'h3db6ab10} /* (12, 2, 9) {real, imag} */,
  {32'h3e8b6a78, 32'h3f58a6c5} /* (12, 2, 8) {real, imag} */,
  {32'h3df5d9dc, 32'h3f8e5680} /* (12, 2, 7) {real, imag} */,
  {32'h3e880628, 32'hbed61f8a} /* (12, 2, 6) {real, imag} */,
  {32'h3fbc569e, 32'h3ea63fba} /* (12, 2, 5) {real, imag} */,
  {32'h3f46a517, 32'h3fb05afd} /* (12, 2, 4) {real, imag} */,
  {32'hbef16c5a, 32'h3f882d3e} /* (12, 2, 3) {real, imag} */,
  {32'hbdbd9c70, 32'h3f872ceb} /* (12, 2, 2) {real, imag} */,
  {32'h3f0a4ff4, 32'h3fdcd87b} /* (12, 2, 1) {real, imag} */,
  {32'hbedcd534, 32'h3ed58b90} /* (12, 2, 0) {real, imag} */,
  {32'hbefef650, 32'hbf2fbd18} /* (12, 1, 15) {real, imag} */,
  {32'hbf5c7872, 32'h3dfbc23c} /* (12, 1, 14) {real, imag} */,
  {32'hbd8a6f78, 32'h3f1ae05b} /* (12, 1, 13) {real, imag} */,
  {32'h3e9bf510, 32'h3ed08054} /* (12, 1, 12) {real, imag} */,
  {32'h3d50a1d0, 32'h3db99058} /* (12, 1, 11) {real, imag} */,
  {32'hbe2a6fe8, 32'hbeec0c1e} /* (12, 1, 10) {real, imag} */,
  {32'h3e82696e, 32'h3f2bcf6c} /* (12, 1, 9) {real, imag} */,
  {32'h3f7ec66e, 32'h3f8946ce} /* (12, 1, 8) {real, imag} */,
  {32'h3f7b8d18, 32'hbe4f3c32} /* (12, 1, 7) {real, imag} */,
  {32'h3f875444, 32'h3c00ab60} /* (12, 1, 6) {real, imag} */,
  {32'h3fddf298, 32'h3f8de5e5} /* (12, 1, 5) {real, imag} */,
  {32'hbf06871c, 32'h3e8ca3f6} /* (12, 1, 4) {real, imag} */,
  {32'hbf4fd96c, 32'hbf4c00cc} /* (12, 1, 3) {real, imag} */,
  {32'h3d5f43a0, 32'hbf6d4552} /* (12, 1, 2) {real, imag} */,
  {32'h3e082b28, 32'h3f97b0af} /* (12, 1, 1) {real, imag} */,
  {32'hbe87723b, 32'hbe199efa} /* (12, 1, 0) {real, imag} */,
  {32'hbf2e6fe8, 32'h3e3d73c5} /* (12, 0, 15) {real, imag} */,
  {32'hbe9d99ab, 32'h3cba42c0} /* (12, 0, 14) {real, imag} */,
  {32'hbe2234b6, 32'h3e0e6fb0} /* (12, 0, 13) {real, imag} */,
  {32'hbf5e080f, 32'h3eccf712} /* (12, 0, 12) {real, imag} */,
  {32'hbf8d1905, 32'hbd3082ec} /* (12, 0, 11) {real, imag} */,
  {32'hbec04b5e, 32'hbf22b0d2} /* (12, 0, 10) {real, imag} */,
  {32'h3d006c88, 32'hbe8f9d27} /* (12, 0, 9) {real, imag} */,
  {32'h3f7ef9d8, 32'h3f45767c} /* (12, 0, 8) {real, imag} */,
  {32'h3f5996e8, 32'h3ed76796} /* (12, 0, 7) {real, imag} */,
  {32'h3f5a716d, 32'h3e3a6924} /* (12, 0, 6) {real, imag} */,
  {32'h3f44096c, 32'h3e1e0815} /* (12, 0, 5) {real, imag} */,
  {32'hbd9b05a0, 32'hbf2faae8} /* (12, 0, 4) {real, imag} */,
  {32'hbd2e52a0, 32'hbe8f934e} /* (12, 0, 3) {real, imag} */,
  {32'hbe15a00b, 32'hbf389cc2} /* (12, 0, 2) {real, imag} */,
  {32'hbf1bab92, 32'hbf092017} /* (12, 0, 1) {real, imag} */,
  {32'hbf0c59de, 32'hbf162051} /* (12, 0, 0) {real, imag} */,
  {32'h3f1ad7cf, 32'h3f03733c} /* (11, 15, 15) {real, imag} */,
  {32'h3e9ca1ca, 32'h3e5add77} /* (11, 15, 14) {real, imag} */,
  {32'hbe460084, 32'h3ef8a35c} /* (11, 15, 13) {real, imag} */,
  {32'h3d92bc88, 32'hbe1acc20} /* (11, 15, 12) {real, imag} */,
  {32'h3cd89ea0, 32'h3e6ac53b} /* (11, 15, 11) {real, imag} */,
  {32'hbf6d9033, 32'hbaf57700} /* (11, 15, 10) {real, imag} */,
  {32'hbf542e51, 32'hbf65f925} /* (11, 15, 9) {real, imag} */,
  {32'h3f39f5b1, 32'hbf282775} /* (11, 15, 8) {real, imag} */,
  {32'h3f4926fe, 32'h3df15f44} /* (11, 15, 7) {real, imag} */,
  {32'h3e817e47, 32'h3f7831ce} /* (11, 15, 6) {real, imag} */,
  {32'h3eabe9fc, 32'h3f7d2f62} /* (11, 15, 5) {real, imag} */,
  {32'hbf4bd8d7, 32'hbc26e360} /* (11, 15, 4) {real, imag} */,
  {32'h3deebb64, 32'hbf347506} /* (11, 15, 3) {real, imag} */,
  {32'h3fa7614e, 32'hbf01f1fc} /* (11, 15, 2) {real, imag} */,
  {32'h3f71bd23, 32'h3e293a44} /* (11, 15, 1) {real, imag} */,
  {32'h3f3157e2, 32'h3ec21936} /* (11, 15, 0) {real, imag} */,
  {32'h3f00b2e8, 32'h3eb9620a} /* (11, 14, 15) {real, imag} */,
  {32'h3d8b70e8, 32'h3e14aff8} /* (11, 14, 14) {real, imag} */,
  {32'h3d87af4c, 32'h3e63dfd8} /* (11, 14, 13) {real, imag} */,
  {32'h3f841a36, 32'hbe70f9a8} /* (11, 14, 12) {real, imag} */,
  {32'h3ef15731, 32'h3f210817} /* (11, 14, 11) {real, imag} */,
  {32'hbf955cfe, 32'h3dad8b98} /* (11, 14, 10) {real, imag} */,
  {32'hbf991b7b, 32'hbfad62c4} /* (11, 14, 9) {real, imag} */,
  {32'h3eb023ef, 32'hbf57972a} /* (11, 14, 8) {real, imag} */,
  {32'hbcdb0190, 32'h3ebd3efe} /* (11, 14, 7) {real, imag} */,
  {32'h3d449e50, 32'h3f825386} /* (11, 14, 6) {real, imag} */,
  {32'h3f15f17a, 32'h3ed9ebaa} /* (11, 14, 5) {real, imag} */,
  {32'hbe48e7b0, 32'h3d9f8b88} /* (11, 14, 4) {real, imag} */,
  {32'hbe9d83db, 32'hbe1b8114} /* (11, 14, 3) {real, imag} */,
  {32'h3f253486, 32'hbeba4d68} /* (11, 14, 2) {real, imag} */,
  {32'h3f529e50, 32'h3eade579} /* (11, 14, 1) {real, imag} */,
  {32'h3f0306a1, 32'h3ef52f51} /* (11, 14, 0) {real, imag} */,
  {32'hbe943c78, 32'h3de34bd2} /* (11, 13, 15) {real, imag} */,
  {32'hbbc86900, 32'h3e03cdf2} /* (11, 13, 14) {real, imag} */,
  {32'h3f4190a7, 32'hbd808480} /* (11, 13, 13) {real, imag} */,
  {32'h3fe37731, 32'h3f78e5c4} /* (11, 13, 12) {real, imag} */,
  {32'h3f9a044d, 32'h3f095f74} /* (11, 13, 11) {real, imag} */,
  {32'h3d4c2c40, 32'hbddaf0ec} /* (11, 13, 10) {real, imag} */,
  {32'h3d9e926c, 32'h3ef16776} /* (11, 13, 9) {real, imag} */,
  {32'hbe9deabd, 32'h3ea48314} /* (11, 13, 8) {real, imag} */,
  {32'hbf52b14c, 32'h3f12e9be} /* (11, 13, 7) {real, imag} */,
  {32'h3eca51f2, 32'h3f91608c} /* (11, 13, 6) {real, imag} */,
  {32'h3e33efb0, 32'hbdca4f0a} /* (11, 13, 5) {real, imag} */,
  {32'hbed115ce, 32'h3ee69260} /* (11, 13, 4) {real, imag} */,
  {32'h3f12d0aa, 32'h3fa56d9a} /* (11, 13, 3) {real, imag} */,
  {32'h3f94d96a, 32'h3f03062a} /* (11, 13, 2) {real, imag} */,
  {32'h3f24da8b, 32'h3ee1691b} /* (11, 13, 1) {real, imag} */,
  {32'hbecb6caa, 32'h3ea874cc} /* (11, 13, 0) {real, imag} */,
  {32'hbe263491, 32'hbf70f61f} /* (11, 12, 15) {real, imag} */,
  {32'hbe3fc7ee, 32'hbf8035da} /* (11, 12, 14) {real, imag} */,
  {32'h3e6ecab0, 32'h3f0920ca} /* (11, 12, 13) {real, imag} */,
  {32'h3f2df548, 32'h3f0c6430} /* (11, 12, 12) {real, imag} */,
  {32'h3f4f4514, 32'hbf368910} /* (11, 12, 11) {real, imag} */,
  {32'h3df86184, 32'hbf1270e4} /* (11, 12, 10) {real, imag} */,
  {32'h3f9c32ea, 32'h3e7872e0} /* (11, 12, 9) {real, imag} */,
  {32'h3f25062a, 32'hbf20ae50} /* (11, 12, 8) {real, imag} */,
  {32'hbe81ebc8, 32'hbf155016} /* (11, 12, 7) {real, imag} */,
  {32'h3f862f13, 32'hbe6f27b8} /* (11, 12, 6) {real, imag} */,
  {32'h3f6ae5d8, 32'hbf15b311} /* (11, 12, 5) {real, imag} */,
  {32'h3bf45500, 32'hbe5241d0} /* (11, 12, 4) {real, imag} */,
  {32'h3e87621a, 32'h3f6f641e} /* (11, 12, 3) {real, imag} */,
  {32'h3d8f9f98, 32'h3f8eaa54} /* (11, 12, 2) {real, imag} */,
  {32'hbdcb0888, 32'h3f9773ff} /* (11, 12, 1) {real, imag} */,
  {32'hbe553f2d, 32'h3ec86c1b} /* (11, 12, 0) {real, imag} */,
  {32'hbee64398, 32'hbfbbb564} /* (11, 11, 15) {real, imag} */,
  {32'hbe62eaca, 32'hbecfd50e} /* (11, 11, 14) {real, imag} */,
  {32'hbe088bbc, 32'h3f979fac} /* (11, 11, 13) {real, imag} */,
  {32'hbd80b424, 32'h3eed2000} /* (11, 11, 12) {real, imag} */,
  {32'h3e4820c6, 32'hbf0486a0} /* (11, 11, 11) {real, imag} */,
  {32'h3f361a63, 32'h3c1a2b50} /* (11, 11, 10) {real, imag} */,
  {32'h3fcad500, 32'h3ef8be6b} /* (11, 11, 9) {real, imag} */,
  {32'h3f9f71fd, 32'h3e863abe} /* (11, 11, 8) {real, imag} */,
  {32'h3c68b900, 32'h3f485ab4} /* (11, 11, 7) {real, imag} */,
  {32'hbe2675d0, 32'h3ee22f14} /* (11, 11, 6) {real, imag} */,
  {32'h3f2c545a, 32'h3f6fd5ab} /* (11, 11, 5) {real, imag} */,
  {32'h3f8ed028, 32'h3f7ad5b8} /* (11, 11, 4) {real, imag} */,
  {32'h3f095af2, 32'h3d5fad54} /* (11, 11, 3) {real, imag} */,
  {32'hbf0522b0, 32'hbf51f7d4} /* (11, 11, 2) {real, imag} */,
  {32'hbf005d81, 32'hbea1a1ec} /* (11, 11, 1) {real, imag} */,
  {32'hbe0fbb80, 32'hbe526ef1} /* (11, 11, 0) {real, imag} */,
  {32'hbd61c468, 32'hbf1d53b8} /* (11, 10, 15) {real, imag} */,
  {32'hbedbdbde, 32'h3f67c6a2} /* (11, 10, 14) {real, imag} */,
  {32'hbbe3c2c0, 32'h3fee965b} /* (11, 10, 13) {real, imag} */,
  {32'h3f4fdeb9, 32'h3f8804a7} /* (11, 10, 12) {real, imag} */,
  {32'h3e031bf8, 32'hbed0fa80} /* (11, 10, 11) {real, imag} */,
  {32'h3dd2d942, 32'h3e96f5d8} /* (11, 10, 10) {real, imag} */,
  {32'h3fa1dcd6, 32'h3f0c6a31} /* (11, 10, 9) {real, imag} */,
  {32'h3ec37044, 32'h3fcaabdc} /* (11, 10, 8) {real, imag} */,
  {32'hbdf4c798, 32'h3faa1bd5} /* (11, 10, 7) {real, imag} */,
  {32'hbf6525ef, 32'h3e8a7d7c} /* (11, 10, 6) {real, imag} */,
  {32'hbf36a024, 32'h3fd24a33} /* (11, 10, 5) {real, imag} */,
  {32'h3f55da96, 32'h3f645dcc} /* (11, 10, 4) {real, imag} */,
  {32'h3f98507d, 32'h3e8e2040} /* (11, 10, 3) {real, imag} */,
  {32'hbe268b90, 32'hbf564935} /* (11, 10, 2) {real, imag} */,
  {32'hbf1046b3, 32'hbf67f88e} /* (11, 10, 1) {real, imag} */,
  {32'h3cc5b1c0, 32'hbe7305b2} /* (11, 10, 0) {real, imag} */,
  {32'h3f6866c6, 32'h3db6ad90} /* (11, 9, 15) {real, imag} */,
  {32'h3eff8b63, 32'h3e9f27cb} /* (11, 9, 14) {real, imag} */,
  {32'hbf4f5dcb, 32'h3f25a52a} /* (11, 9, 13) {real, imag} */,
  {32'h3d797bd0, 32'h3f8714a3} /* (11, 9, 12) {real, imag} */,
  {32'hbf0bcdc0, 32'hbcf8a700} /* (11, 9, 11) {real, imag} */,
  {32'hbf667e77, 32'h3f0fb0e2} /* (11, 9, 10) {real, imag} */,
  {32'h3f6128c1, 32'hbe395110} /* (11, 9, 9) {real, imag} */,
  {32'h3ec7ffa4, 32'h3ecdd8c3} /* (11, 9, 8) {real, imag} */,
  {32'hbe81203c, 32'hbe9ae352} /* (11, 9, 7) {real, imag} */,
  {32'h3f20e2a6, 32'hbf633097} /* (11, 9, 6) {real, imag} */,
  {32'hbd31fa50, 32'h3f243348} /* (11, 9, 5) {real, imag} */,
  {32'hbda151f0, 32'hbe551044} /* (11, 9, 4) {real, imag} */,
  {32'h3ed7b3d1, 32'hbe91fea6} /* (11, 9, 3) {real, imag} */,
  {32'h3f25f272, 32'hbedae5cc} /* (11, 9, 2) {real, imag} */,
  {32'h3cf7a140, 32'hbe9b7d18} /* (11, 9, 1) {real, imag} */,
  {32'h3e96fcdf, 32'h3f111f79} /* (11, 9, 0) {real, imag} */,
  {32'hbe166aa8, 32'h3e29b059} /* (11, 8, 15) {real, imag} */,
  {32'hbc6df278, 32'hbe834cad} /* (11, 8, 14) {real, imag} */,
  {32'hbe8ecfb0, 32'h3ea3ffcb} /* (11, 8, 13) {real, imag} */,
  {32'h3f3be7f3, 32'h3f0f2243} /* (11, 8, 12) {real, imag} */,
  {32'hbe2c4e2a, 32'h3ec47f52} /* (11, 8, 11) {real, imag} */,
  {32'hbf0955bc, 32'h3f6c7d60} /* (11, 8, 10) {real, imag} */,
  {32'h3f5a791f, 32'h3e7369e4} /* (11, 8, 9) {real, imag} */,
  {32'h3f13d5e4, 32'hbdecb904} /* (11, 8, 8) {real, imag} */,
  {32'hbda9ef98, 32'hbf24de18} /* (11, 8, 7) {real, imag} */,
  {32'h3f421a24, 32'hbfa8cc93} /* (11, 8, 6) {real, imag} */,
  {32'hbd9d3df0, 32'h3f1e8f99} /* (11, 8, 5) {real, imag} */,
  {32'hbf3c6399, 32'h3f359267} /* (11, 8, 4) {real, imag} */,
  {32'h3ec59350, 32'hbcadb2c0} /* (11, 8, 3) {real, imag} */,
  {32'h3f092e3f, 32'h3ee08000} /* (11, 8, 2) {real, imag} */,
  {32'hbf1a193e, 32'h3eba1d18} /* (11, 8, 1) {real, imag} */,
  {32'hbf63e7b0, 32'h3e80803f} /* (11, 8, 0) {real, imag} */,
  {32'hbf2fb868, 32'h3f0a6f6f} /* (11, 7, 15) {real, imag} */,
  {32'hbf2941cb, 32'h3e3662a0} /* (11, 7, 14) {real, imag} */,
  {32'h3eadbfe0, 32'hbee8b495} /* (11, 7, 13) {real, imag} */,
  {32'h3ecd4bdc, 32'h3dc33a6c} /* (11, 7, 12) {real, imag} */,
  {32'hbe2d95c8, 32'h3f5901e8} /* (11, 7, 11) {real, imag} */,
  {32'h3e4d2a24, 32'h3f9136da} /* (11, 7, 10) {real, imag} */,
  {32'h3ef5df42, 32'h3f1ec694} /* (11, 7, 9) {real, imag} */,
  {32'hbf166658, 32'hbdb32583} /* (11, 7, 8) {real, imag} */,
  {32'hbf35e91e, 32'hbdaa5493} /* (11, 7, 7) {real, imag} */,
  {32'hbe36a4a0, 32'hbf9f8e40} /* (11, 7, 6) {real, imag} */,
  {32'hbef9fdae, 32'hbe5193a0} /* (11, 7, 5) {real, imag} */,
  {32'hbda85818, 32'h3eaec859} /* (11, 7, 4) {real, imag} */,
  {32'h3fa55fe1, 32'h3e7a2634} /* (11, 7, 3) {real, imag} */,
  {32'h3fad9e3e, 32'h3f3a5c5a} /* (11, 7, 2) {real, imag} */,
  {32'hbe59c79c, 32'hbc40cc40} /* (11, 7, 1) {real, imag} */,
  {32'hbf94b0b1, 32'h3e22cf80} /* (11, 7, 0) {real, imag} */,
  {32'hbe89685b, 32'h3e469168} /* (11, 6, 15) {real, imag} */,
  {32'hbfa5c52a, 32'hbca74580} /* (11, 6, 14) {real, imag} */,
  {32'hbf0f3721, 32'hbef537c5} /* (11, 6, 13) {real, imag} */,
  {32'hbf1be78e, 32'hbeab6ec2} /* (11, 6, 12) {real, imag} */,
  {32'hbf30d620, 32'h3ed4a056} /* (11, 6, 11) {real, imag} */,
  {32'h3f72e098, 32'h3f06e62d} /* (11, 6, 10) {real, imag} */,
  {32'h3e7af0b4, 32'h3fa25c05} /* (11, 6, 9) {real, imag} */,
  {32'hbf93aada, 32'h3f95b607} /* (11, 6, 8) {real, imag} */,
  {32'hbf21e240, 32'h3ebf74a8} /* (11, 6, 7) {real, imag} */,
  {32'h3e81beb2, 32'hbf60909d} /* (11, 6, 6) {real, imag} */,
  {32'h3cb7b4e0, 32'hbfbd79de} /* (11, 6, 5) {real, imag} */,
  {32'hbe0152f2, 32'hbd909d68} /* (11, 6, 4) {real, imag} */,
  {32'h3e5933a6, 32'h3e9e4940} /* (11, 6, 3) {real, imag} */,
  {32'h3f5affe3, 32'h3d823c4c} /* (11, 6, 2) {real, imag} */,
  {32'h3f01eb17, 32'h3ed167d8} /* (11, 6, 1) {real, imag} */,
  {32'hbdcc2360, 32'h3f3aea15} /* (11, 6, 0) {real, imag} */,
  {32'hbe4da880, 32'hbe12d9d0} /* (11, 5, 15) {real, imag} */,
  {32'hbf9ad43d, 32'hbedbc326} /* (11, 5, 14) {real, imag} */,
  {32'hbecb28dc, 32'hbf2cd22d} /* (11, 5, 13) {real, imag} */,
  {32'hbed14e16, 32'hbeeb8dad} /* (11, 5, 12) {real, imag} */,
  {32'hbe8d2c19, 32'h3f6c80e2} /* (11, 5, 11) {real, imag} */,
  {32'h3e948b5e, 32'h3dfb1454} /* (11, 5, 10) {real, imag} */,
  {32'h3e82af4b, 32'h3f129bf2} /* (11, 5, 9) {real, imag} */,
  {32'hbe36da40, 32'h3f9fc4a6} /* (11, 5, 8) {real, imag} */,
  {32'h3c66e940, 32'h3eb51642} /* (11, 5, 7) {real, imag} */,
  {32'h3fbb4427, 32'hbd549038} /* (11, 5, 6) {real, imag} */,
  {32'h3fa8542a, 32'hbbf76f40} /* (11, 5, 5) {real, imag} */,
  {32'h3e55aeca, 32'h3f89547d} /* (11, 5, 4) {real, imag} */,
  {32'hbf041ade, 32'h3f9a579f} /* (11, 5, 3) {real, imag} */,
  {32'hbf1394bd, 32'h3ec6f89b} /* (11, 5, 2) {real, imag} */,
  {32'hbf0bad94, 32'h3f8f9f38} /* (11, 5, 1) {real, imag} */,
  {32'hbe6efa82, 32'h3f3f2165} /* (11, 5, 0) {real, imag} */,
  {32'hbea5894c, 32'hbf14c1fb} /* (11, 4, 15) {real, imag} */,
  {32'hbf364da9, 32'hbf02913e} /* (11, 4, 14) {real, imag} */,
  {32'h3f156892, 32'hbebadd58} /* (11, 4, 13) {real, imag} */,
  {32'h3f5a31aa, 32'hbee1efe3} /* (11, 4, 12) {real, imag} */,
  {32'h3e7d7b4a, 32'h3f6f74f3} /* (11, 4, 11) {real, imag} */,
  {32'hbf109600, 32'h3f023978} /* (11, 4, 10) {real, imag} */,
  {32'hbe47d120, 32'h3f7f975f} /* (11, 4, 9) {real, imag} */,
  {32'h3e878dea, 32'h3f0b520c} /* (11, 4, 8) {real, imag} */,
  {32'hbf28d12c, 32'h3bb89600} /* (11, 4, 7) {real, imag} */,
  {32'h3e1bdd63, 32'hbe8293ad} /* (11, 4, 6) {real, imag} */,
  {32'h3f29cc8a, 32'hbf473ced} /* (11, 4, 5) {real, imag} */,
  {32'hbe68f246, 32'hbdafe6e4} /* (11, 4, 4) {real, imag} */,
  {32'hbf1e1f00, 32'h3f43c100} /* (11, 4, 3) {real, imag} */,
  {32'hbf13c926, 32'h3eb4e8e6} /* (11, 4, 2) {real, imag} */,
  {32'hbf42bdd4, 32'h3f5ec0b8} /* (11, 4, 1) {real, imag} */,
  {32'hbe58a7c0, 32'h3f991e94} /* (11, 4, 0) {real, imag} */,
  {32'hbf226782, 32'hbe410d7c} /* (11, 3, 15) {real, imag} */,
  {32'hbecfcfd6, 32'h3e5fcfb4} /* (11, 3, 14) {real, imag} */,
  {32'h3f8882c8, 32'h3f21d5c4} /* (11, 3, 13) {real, imag} */,
  {32'h3ea5f240, 32'h3f33f898} /* (11, 3, 12) {real, imag} */,
  {32'hbe330120, 32'h3f44a27a} /* (11, 3, 11) {real, imag} */,
  {32'hbf498d70, 32'h3e358dc4} /* (11, 3, 10) {real, imag} */,
  {32'h3efb5760, 32'h3f0777a5} /* (11, 3, 9) {real, imag} */,
  {32'h3fbf2cba, 32'h3f03ec9c} /* (11, 3, 8) {real, imag} */,
  {32'h3f40bd62, 32'h3eda064a} /* (11, 3, 7) {real, imag} */,
  {32'hbf00e8a4, 32'hbeb6a342} /* (11, 3, 6) {real, imag} */,
  {32'h3f196104, 32'hbf817f85} /* (11, 3, 5) {real, imag} */,
  {32'h3f620785, 32'hbf4b37bd} /* (11, 3, 4) {real, imag} */,
  {32'hbf005ba4, 32'h3eb99660} /* (11, 3, 3) {real, imag} */,
  {32'hbe9b14aa, 32'hbe15647c} /* (11, 3, 2) {real, imag} */,
  {32'hbf01d385, 32'hbfbe030c} /* (11, 3, 1) {real, imag} */,
  {32'hbf59d754, 32'h3ecd3e34} /* (11, 3, 0) {real, imag} */,
  {32'hbe9d80c6, 32'h3e5e0d3e} /* (11, 2, 15) {real, imag} */,
  {32'h3e7d06d8, 32'h3db05fac} /* (11, 2, 14) {real, imag} */,
  {32'h3f9337dc, 32'h3f3526f8} /* (11, 2, 13) {real, imag} */,
  {32'h3e56d8a4, 32'h3fc9c7f0} /* (11, 2, 12) {real, imag} */,
  {32'hbeb319c1, 32'h3f065a1b} /* (11, 2, 11) {real, imag} */,
  {32'hbf05bf86, 32'h3eb007a6} /* (11, 2, 10) {real, imag} */,
  {32'hbd97c90c, 32'h3dc2f3f4} /* (11, 2, 9) {real, imag} */,
  {32'h3ed90a2c, 32'h3dab1ac8} /* (11, 2, 8) {real, imag} */,
  {32'h3f6b7b2c, 32'h3e709f54} /* (11, 2, 7) {real, imag} */,
  {32'hbe86fe79, 32'hbd429a30} /* (11, 2, 6) {real, imag} */,
  {32'h3e5a2d10, 32'h3e58a634} /* (11, 2, 5) {real, imag} */,
  {32'h3f0a5607, 32'hbee3f212} /* (11, 2, 4) {real, imag} */,
  {32'h3d895d04, 32'hbf2e88b9} /* (11, 2, 3) {real, imag} */,
  {32'h3ef69f1f, 32'hbf56f02a} /* (11, 2, 2) {real, imag} */,
  {32'h3e819200, 32'hbff22557} /* (11, 2, 1) {real, imag} */,
  {32'hbdf89560, 32'hbe2eeda8} /* (11, 2, 0) {real, imag} */,
  {32'h3e8118fb, 32'h3f693490} /* (11, 1, 15) {real, imag} */,
  {32'h3f0334b1, 32'h3e9b4368} /* (11, 1, 14) {real, imag} */,
  {32'h3f913b4c, 32'h3e7eb865} /* (11, 1, 13) {real, imag} */,
  {32'h3eb921d0, 32'h3f1c50e9} /* (11, 1, 12) {real, imag} */,
  {32'hbe88aa44, 32'hbf48e872} /* (11, 1, 11) {real, imag} */,
  {32'hbf8ecc42, 32'hbd2c7d40} /* (11, 1, 10) {real, imag} */,
  {32'hbfa17ac8, 32'hbdd6cbec} /* (11, 1, 9) {real, imag} */,
  {32'hbe846a6c, 32'hbd54e770} /* (11, 1, 8) {real, imag} */,
  {32'hbe54ad10, 32'h3e76b370} /* (11, 1, 7) {real, imag} */,
  {32'h3cc32550, 32'h3efe0836} /* (11, 1, 6) {real, imag} */,
  {32'h3f2e24e0, 32'h3f89bc7c} /* (11, 1, 5) {real, imag} */,
  {32'h3f9cd398, 32'hbeca7878} /* (11, 1, 4) {real, imag} */,
  {32'h3fa1894e, 32'hbf147a46} /* (11, 1, 3) {real, imag} */,
  {32'h3f1c7dd4, 32'hbf19df04} /* (11, 1, 2) {real, imag} */,
  {32'h3f16f7f6, 32'hbe8c3288} /* (11, 1, 1) {real, imag} */,
  {32'h3f5581ae, 32'h3f1e8adc} /* (11, 1, 0) {real, imag} */,
  {32'h3e417442, 32'h3e9f7a22} /* (11, 0, 15) {real, imag} */,
  {32'h3ec694ef, 32'h3ea9ea12} /* (11, 0, 14) {real, imag} */,
  {32'h3f82bbea, 32'h3e902260} /* (11, 0, 13) {real, imag} */,
  {32'h3f38c444, 32'hbe13ddbc} /* (11, 0, 12) {real, imag} */,
  {32'h3eb574b2, 32'hbef4ddfb} /* (11, 0, 11) {real, imag} */,
  {32'h3d45fbf4, 32'hbe964616} /* (11, 0, 10) {real, imag} */,
  {32'hbf21699a, 32'hbe3683d2} /* (11, 0, 9) {real, imag} */,
  {32'hbed57dc5, 32'h3de81a06} /* (11, 0, 8) {real, imag} */,
  {32'hbf1e01ef, 32'h3d9a4c28} /* (11, 0, 7) {real, imag} */,
  {32'hbe8369b1, 32'h3ec64a84} /* (11, 0, 6) {real, imag} */,
  {32'h3f46b45c, 32'h3f12f006} /* (11, 0, 5) {real, imag} */,
  {32'h3f351f4c, 32'hbdac9c20} /* (11, 0, 4) {real, imag} */,
  {32'h3e806b05, 32'hbee84482} /* (11, 0, 3) {real, imag} */,
  {32'h3cc80580, 32'hbf3e8f35} /* (11, 0, 2) {real, imag} */,
  {32'h3f3f4317, 32'hbd594558} /* (11, 0, 1) {real, imag} */,
  {32'h3f4b1cf4, 32'h3ef1eb4a} /* (11, 0, 0) {real, imag} */,
  {32'hbd8a394c, 32'h3eb1ca6c} /* (10, 15, 15) {real, imag} */,
  {32'hbe096ee4, 32'hbd5a8660} /* (10, 15, 14) {real, imag} */,
  {32'hbd419aea, 32'hbd9a23b4} /* (10, 15, 13) {real, imag} */,
  {32'h3cbf075c, 32'h3ebf86df} /* (10, 15, 12) {real, imag} */,
  {32'h3e164cee, 32'h3eb8f0f3} /* (10, 15, 11) {real, imag} */,
  {32'hbdca9218, 32'h3e055404} /* (10, 15, 10) {real, imag} */,
  {32'hbdb1a19a, 32'hbd134b10} /* (10, 15, 9) {real, imag} */,
  {32'hbc238f30, 32'h3d48443c} /* (10, 15, 8) {real, imag} */,
  {32'hbe9880a7, 32'hbf0c78c0} /* (10, 15, 7) {real, imag} */,
  {32'hbef90b1b, 32'hbd495238} /* (10, 15, 6) {real, imag} */,
  {32'h3e2b3a6c, 32'h3e8b982c} /* (10, 15, 5) {real, imag} */,
  {32'h3ec13388, 32'h3dedf330} /* (10, 15, 4) {real, imag} */,
  {32'h3d789b20, 32'h3f22b5aa} /* (10, 15, 3) {real, imag} */,
  {32'hbe09b7b1, 32'h3eb444b9} /* (10, 15, 2) {real, imag} */,
  {32'h3e9376ea, 32'hbf169403} /* (10, 15, 1) {real, imag} */,
  {32'h3efd7706, 32'hbed594d8} /* (10, 15, 0) {real, imag} */,
  {32'h3f155438, 32'hbe8f6552} /* (10, 14, 15) {real, imag} */,
  {32'h3ec828f6, 32'hbf0c504e} /* (10, 14, 14) {real, imag} */,
  {32'hbe7b6f7c, 32'h3e801038} /* (10, 14, 13) {real, imag} */,
  {32'h3e013644, 32'h3f2f0036} /* (10, 14, 12) {real, imag} */,
  {32'h3f83bd76, 32'h3f7f4fd8} /* (10, 14, 11) {real, imag} */,
  {32'h3f333444, 32'h3f9e15ac} /* (10, 14, 10) {real, imag} */,
  {32'h3e2be418, 32'h3f950972} /* (10, 14, 9) {real, imag} */,
  {32'h3bd4b2c0, 32'h3ead848e} /* (10, 14, 8) {real, imag} */,
  {32'hbeecedb7, 32'hbe1b2784} /* (10, 14, 7) {real, imag} */,
  {32'hbf56f19e, 32'h3e433590} /* (10, 14, 6) {real, imag} */,
  {32'hbe2b923c, 32'h3f236308} /* (10, 14, 5) {real, imag} */,
  {32'hbdbe8590, 32'h3f460408} /* (10, 14, 4) {real, imag} */,
  {32'h3d706a40, 32'h3f1eac76} /* (10, 14, 3) {real, imag} */,
  {32'hbebf7a96, 32'h3ec41b3a} /* (10, 14, 2) {real, imag} */,
  {32'hbf026bc7, 32'hbed24128} /* (10, 14, 1) {real, imag} */,
  {32'h3f10d654, 32'hbf05ca12} /* (10, 14, 0) {real, imag} */,
  {32'h3dbbf0e6, 32'hbf088342} /* (10, 13, 15) {real, imag} */,
  {32'h3d914ac2, 32'hbdf3ac70} /* (10, 13, 14) {real, imag} */,
  {32'hbc72fc30, 32'h3e831030} /* (10, 13, 13) {real, imag} */,
  {32'h3dae3468, 32'h3d857820} /* (10, 13, 12) {real, imag} */,
  {32'h3f1f1ac7, 32'h3dc3aa88} /* (10, 13, 11) {real, imag} */,
  {32'h3eff951a, 32'h3f790e61} /* (10, 13, 10) {real, imag} */,
  {32'h3e97e0c2, 32'h3f7b1e3e} /* (10, 13, 9) {real, imag} */,
  {32'hbed9eb6d, 32'h3e331708} /* (10, 13, 8) {real, imag} */,
  {32'hbea3891c, 32'hbe17a168} /* (10, 13, 7) {real, imag} */,
  {32'hbf606a08, 32'hbf06a486} /* (10, 13, 6) {real, imag} */,
  {32'hbf4555ec, 32'h3eb21a40} /* (10, 13, 5) {real, imag} */,
  {32'hbebddd1a, 32'h3f48f523} /* (10, 13, 4) {real, imag} */,
  {32'hbce9e580, 32'h3e46f5fc} /* (10, 13, 3) {real, imag} */,
  {32'h3e79b419, 32'h3e558cd2} /* (10, 13, 2) {real, imag} */,
  {32'hbea2070e, 32'h3e55cdba} /* (10, 13, 1) {real, imag} */,
  {32'hbe72e650, 32'hbb48ae00} /* (10, 13, 0) {real, imag} */,
  {32'hbe409656, 32'hbdd578bc} /* (10, 12, 15) {real, imag} */,
  {32'hbe995ac8, 32'hbea52186} /* (10, 12, 14) {real, imag} */,
  {32'h3e44834e, 32'h3e56b58a} /* (10, 12, 13) {real, imag} */,
  {32'h3e1b487e, 32'h3f4ee555} /* (10, 12, 12) {real, imag} */,
  {32'h3f223a30, 32'h3f457c21} /* (10, 12, 11) {real, imag} */,
  {32'h3d3f6c3b, 32'h3f41a21f} /* (10, 12, 10) {real, imag} */,
  {32'hbf37d116, 32'hbf29ab1a} /* (10, 12, 9) {real, imag} */,
  {32'hbf431820, 32'hbf33cc05} /* (10, 12, 8) {real, imag} */,
  {32'h3dea578c, 32'hbf6c287c} /* (10, 12, 7) {real, imag} */,
  {32'hbeff9af4, 32'hbf459bba} /* (10, 12, 6) {real, imag} */,
  {32'hbfa49f76, 32'hbebcae94} /* (10, 12, 5) {real, imag} */,
  {32'hbe3f8de1, 32'h3ed05444} /* (10, 12, 4) {real, imag} */,
  {32'h3f06a987, 32'h3f43c7a4} /* (10, 12, 3) {real, imag} */,
  {32'h3f1ee982, 32'h3ee6a2b2} /* (10, 12, 2) {real, imag} */,
  {32'h3d9cb558, 32'h3f496956} /* (10, 12, 1) {real, imag} */,
  {32'hbe604e20, 32'h3f1f1378} /* (10, 12, 0) {real, imag} */,
  {32'hbe855a9c, 32'h3f2e274f} /* (10, 11, 15) {real, imag} */,
  {32'hbf676ea6, 32'h3f2c59e7} /* (10, 11, 14) {real, imag} */,
  {32'hbf90362e, 32'h3f15cd4e} /* (10, 11, 13) {real, imag} */,
  {32'hbf4be93e, 32'h3ee2744a} /* (10, 11, 12) {real, imag} */,
  {32'h3f204c10, 32'h3e8f955e} /* (10, 11, 11) {real, imag} */,
  {32'hbe264bb0, 32'h3e8fd492} /* (10, 11, 10) {real, imag} */,
  {32'hbecdb8d4, 32'hbe9cdd30} /* (10, 11, 9) {real, imag} */,
  {32'hbeb17b32, 32'hbe8720e8} /* (10, 11, 8) {real, imag} */,
  {32'hbf2f303e, 32'hbee60bdd} /* (10, 11, 7) {real, imag} */,
  {32'hbf908a83, 32'h3d766540} /* (10, 11, 6) {real, imag} */,
  {32'hbfa2b971, 32'h3eb4b5fa} /* (10, 11, 5) {real, imag} */,
  {32'hbdbe2582, 32'h3f6b5127} /* (10, 11, 4) {real, imag} */,
  {32'h3ec1c05b, 32'h3f65a4c6} /* (10, 11, 3) {real, imag} */,
  {32'hbe937903, 32'h3f07b920} /* (10, 11, 2) {real, imag} */,
  {32'hbdb08615, 32'h3faca8cd} /* (10, 11, 1) {real, imag} */,
  {32'hbcb54a10, 32'h3f45fa5a} /* (10, 11, 0) {real, imag} */,
  {32'hbeadd685, 32'h3ec14d37} /* (10, 10, 15) {real, imag} */,
  {32'hbf870298, 32'h3e8a1662} /* (10, 10, 14) {real, imag} */,
  {32'hbf81411c, 32'hbecebdb6} /* (10, 10, 13) {real, imag} */,
  {32'hbf0a8369, 32'hbd9dfb40} /* (10, 10, 12) {real, imag} */,
  {32'hbdfcaaa0, 32'h3c2799a2} /* (10, 10, 11) {real, imag} */,
  {32'hbee26148, 32'hbdb8c42c} /* (10, 10, 10) {real, imag} */,
  {32'hbde4b1c0, 32'h3f2fb5ec} /* (10, 10, 9) {real, imag} */,
  {32'hbeda32e8, 32'h3f87de9c} /* (10, 10, 8) {real, imag} */,
  {32'hbeb6a0b8, 32'h3f014118} /* (10, 10, 7) {real, imag} */,
  {32'h3d0390d8, 32'hbf02d790} /* (10, 10, 6) {real, imag} */,
  {32'h3e89f70d, 32'hbebff4b8} /* (10, 10, 5) {real, imag} */,
  {32'h3f099682, 32'h3f430752} /* (10, 10, 4) {real, imag} */,
  {32'h3ee41e8d, 32'h3f69b389} /* (10, 10, 3) {real, imag} */,
  {32'h3cdca9c0, 32'hbe117eec} /* (10, 10, 2) {real, imag} */,
  {32'h3ee51178, 32'h3f0420ef} /* (10, 10, 1) {real, imag} */,
  {32'h3e80fb44, 32'h3e8e24de} /* (10, 10, 0) {real, imag} */,
  {32'h3eb257bd, 32'h3cce5778} /* (10, 9, 15) {real, imag} */,
  {32'h3f00c747, 32'hbf99ed0e} /* (10, 9, 14) {real, imag} */,
  {32'hbdb94bfc, 32'hbfdde7e6} /* (10, 9, 13) {real, imag} */,
  {32'hbc5f38e8, 32'h3d162ce0} /* (10, 9, 12) {real, imag} */,
  {32'h3da26b52, 32'h3f01506c} /* (10, 9, 11) {real, imag} */,
  {32'h3eda02ea, 32'hbeb242ff} /* (10, 9, 10) {real, imag} */,
  {32'h3e4dd97c, 32'hbdcc8608} /* (10, 9, 9) {real, imag} */,
  {32'hbd154650, 32'h3f5ff4c8} /* (10, 9, 8) {real, imag} */,
  {32'hbd1b9990, 32'h3f437f38} /* (10, 9, 7) {real, imag} */,
  {32'h3f2c1992, 32'h3eec002f} /* (10, 9, 6) {real, imag} */,
  {32'h3f47a1c3, 32'h3e64588e} /* (10, 9, 5) {real, imag} */,
  {32'h3f79eb66, 32'h3f05d7fe} /* (10, 9, 4) {real, imag} */,
  {32'h3e1d0a7c, 32'h3e05efc0} /* (10, 9, 3) {real, imag} */,
  {32'hbe80db6e, 32'hbf056e42} /* (10, 9, 2) {real, imag} */,
  {32'hbe88c765, 32'h3e15c2e0} /* (10, 9, 1) {real, imag} */,
  {32'hbea846ac, 32'h3ee64f11} /* (10, 9, 0) {real, imag} */,
  {32'h3e21f7f4, 32'hbe537c04} /* (10, 8, 15) {real, imag} */,
  {32'h3f058766, 32'hbfa5888d} /* (10, 8, 14) {real, imag} */,
  {32'h3c35ee20, 32'hbfce3314} /* (10, 8, 13) {real, imag} */,
  {32'h3df3d0d0, 32'hbf0ebf30} /* (10, 8, 12) {real, imag} */,
  {32'h3f0ad56f, 32'hbe4d5bf6} /* (10, 8, 11) {real, imag} */,
  {32'h3ea91636, 32'hbe895c24} /* (10, 8, 10) {real, imag} */,
  {32'hbdf8c9d0, 32'hbf1761cd} /* (10, 8, 9) {real, imag} */,
  {32'h3ef84ec8, 32'hbefaee0c} /* (10, 8, 8) {real, imag} */,
  {32'hbdd2cb80, 32'hbece19d2} /* (10, 8, 7) {real, imag} */,
  {32'hbd581f3b, 32'h3f23c0bb} /* (10, 8, 6) {real, imag} */,
  {32'h3ea4a0f0, 32'h3f47ab4a} /* (10, 8, 5) {real, imag} */,
  {32'h3eb66c1a, 32'hbd5afe92} /* (10, 8, 4) {real, imag} */,
  {32'hbf007c1a, 32'hbe8dbfce} /* (10, 8, 3) {real, imag} */,
  {32'hbed4d6e4, 32'hbedaefed} /* (10, 8, 2) {real, imag} */,
  {32'hbea62773, 32'h3e53e5ad} /* (10, 8, 1) {real, imag} */,
  {32'hbedb1e68, 32'h3f1a6756} /* (10, 8, 0) {real, imag} */,
  {32'h3f2591de, 32'hbed6b084} /* (10, 7, 15) {real, imag} */,
  {32'h3f0194f1, 32'hbf94b87b} /* (10, 7, 14) {real, imag} */,
  {32'hbed3909c, 32'hbfc7d07f} /* (10, 7, 13) {real, imag} */,
  {32'h3e83856c, 32'hbf741305} /* (10, 7, 12) {real, imag} */,
  {32'h3f3168dc, 32'hbe7faf8a} /* (10, 7, 11) {real, imag} */,
  {32'h3f769ea4, 32'hbd2462a0} /* (10, 7, 10) {real, imag} */,
  {32'h3ebc104e, 32'h3c30df80} /* (10, 7, 9) {real, imag} */,
  {32'h3edfc934, 32'hbf3925a2} /* (10, 7, 8) {real, imag} */,
  {32'hbd6d0c8a, 32'hbf0c8dba} /* (10, 7, 7) {real, imag} */,
  {32'h3e02a7dc, 32'hbd53a0e0} /* (10, 7, 6) {real, imag} */,
  {32'hbdf0cfc6, 32'hbecc8812} /* (10, 7, 5) {real, imag} */,
  {32'hbcee41d0, 32'hbf6f50e6} /* (10, 7, 4) {real, imag} */,
  {32'h3dac7f92, 32'hbe9f465c} /* (10, 7, 3) {real, imag} */,
  {32'h3d2a61fa, 32'h3d8608cc} /* (10, 7, 2) {real, imag} */,
  {32'h3f080cc2, 32'h3f438cc4} /* (10, 7, 1) {real, imag} */,
  {32'hbe31dcfc, 32'h3f3f1874} /* (10, 7, 0) {real, imag} */,
  {32'h3f333d3d, 32'hbd314420} /* (10, 6, 15) {real, imag} */,
  {32'h3ef5a4f6, 32'hbe767c23} /* (10, 6, 14) {real, imag} */,
  {32'h3dc3e5e4, 32'hbea626e8} /* (10, 6, 13) {real, imag} */,
  {32'h3f0ba7c8, 32'hbed6817c} /* (10, 6, 12) {real, imag} */,
  {32'h3ee9a0f5, 32'h3f4a8849} /* (10, 6, 11) {real, imag} */,
  {32'h3f25de52, 32'h3e47e190} /* (10, 6, 10) {real, imag} */,
  {32'hbe1c3d4c, 32'h3e206125} /* (10, 6, 9) {real, imag} */,
  {32'hbdd74e10, 32'hbe987244} /* (10, 6, 8) {real, imag} */,
  {32'hbce31180, 32'h3ea688fa} /* (10, 6, 7) {real, imag} */,
  {32'hbe836951, 32'h3df83dc4} /* (10, 6, 6) {real, imag} */,
  {32'hbee56eec, 32'hbf8c2494} /* (10, 6, 5) {real, imag} */,
  {32'hbf8f8499, 32'hbf62ccc9} /* (10, 6, 4) {real, imag} */,
  {32'hbc8378c0, 32'h3e9d9684} /* (10, 6, 3) {real, imag} */,
  {32'h3ef4f9ec, 32'h3efd3036} /* (10, 6, 2) {real, imag} */,
  {32'h3f013ec8, 32'h3f603d6f} /* (10, 6, 1) {real, imag} */,
  {32'h3c203d40, 32'h3f057077} /* (10, 6, 0) {real, imag} */,
  {32'h3e81df41, 32'h3cbd60b8} /* (10, 5, 15) {real, imag} */,
  {32'h3f0a5cb4, 32'h3d5a6470} /* (10, 5, 14) {real, imag} */,
  {32'h3e57ff02, 32'hbd3ce408} /* (10, 5, 13) {real, imag} */,
  {32'hbeb8f2e0, 32'hbe0cabcc} /* (10, 5, 12) {real, imag} */,
  {32'hbe84f456, 32'h3e596733} /* (10, 5, 11) {real, imag} */,
  {32'h3eb0a160, 32'h3eb2d20b} /* (10, 5, 10) {real, imag} */,
  {32'h3e5c2640, 32'h3e5ba563} /* (10, 5, 9) {real, imag} */,
  {32'h3edb2398, 32'h3de7fc73} /* (10, 5, 8) {real, imag} */,
  {32'h3df848f8, 32'h3f42f990} /* (10, 5, 7) {real, imag} */,
  {32'hbf2c1254, 32'h3ef2f441} /* (10, 5, 6) {real, imag} */,
  {32'hbf3ad2cb, 32'hbf4a9db6} /* (10, 5, 5) {real, imag} */,
  {32'hbee8f5ec, 32'hbea746c5} /* (10, 5, 4) {real, imag} */,
  {32'hbd287eb0, 32'h3f0568f7} /* (10, 5, 3) {real, imag} */,
  {32'hbd346d00, 32'h3f0d9b10} /* (10, 5, 2) {real, imag} */,
  {32'hbe45cc34, 32'h3f339c3d} /* (10, 5, 1) {real, imag} */,
  {32'hbd0d22e8, 32'h3f08ecef} /* (10, 5, 0) {real, imag} */,
  {32'h3f532283, 32'hbeac336a} /* (10, 4, 15) {real, imag} */,
  {32'h3f90ccfc, 32'hbe03a9cc} /* (10, 4, 14) {real, imag} */,
  {32'hbc2b4e00, 32'hbe43e7ed} /* (10, 4, 13) {real, imag} */,
  {32'hbf887206, 32'h3e9231f6} /* (10, 4, 12) {real, imag} */,
  {32'hbf58eae0, 32'hbc06f1ae} /* (10, 4, 11) {real, imag} */,
  {32'h3e5c44ea, 32'hbedf7f74} /* (10, 4, 10) {real, imag} */,
  {32'h3eb2c8bd, 32'hbf43cf90} /* (10, 4, 9) {real, imag} */,
  {32'h3f89d356, 32'hbedff993} /* (10, 4, 8) {real, imag} */,
  {32'h3f3318af, 32'h3e55f5fb} /* (10, 4, 7) {real, imag} */,
  {32'hbf347944, 32'hbf011746} /* (10, 4, 6) {real, imag} */,
  {32'hbf6a7355, 32'hbf5f1ae0} /* (10, 4, 5) {real, imag} */,
  {32'hbf3e55e2, 32'hba746bf2} /* (10, 4, 4) {real, imag} */,
  {32'h3dd30700, 32'hbe905b32} /* (10, 4, 3) {real, imag} */,
  {32'hbcd947ec, 32'hbd49c1f0} /* (10, 4, 2) {real, imag} */,
  {32'hbd6f60b6, 32'hbccf9990} /* (10, 4, 1) {real, imag} */,
  {32'hbe07d8fc, 32'h3d77bdd0} /* (10, 4, 0) {real, imag} */,
  {32'h3e705d40, 32'h3ec7c866} /* (10, 3, 15) {real, imag} */,
  {32'hbe88dd54, 32'h3e667b50} /* (10, 3, 14) {real, imag} */,
  {32'hbe94a386, 32'hbf83c306} /* (10, 3, 13) {real, imag} */,
  {32'hbf0140d3, 32'hbea00808} /* (10, 3, 12) {real, imag} */,
  {32'hbe7e6fb6, 32'h3dcbe610} /* (10, 3, 11) {real, imag} */,
  {32'hbf1fa61e, 32'hbf5d13ca} /* (10, 3, 10) {real, imag} */,
  {32'hbf182518, 32'hbec89198} /* (10, 3, 9) {real, imag} */,
  {32'h3f1a9232, 32'hbf6f21aa} /* (10, 3, 8) {real, imag} */,
  {32'h3f0c8b86, 32'hbf442eb0} /* (10, 3, 7) {real, imag} */,
  {32'hbeb0abf5, 32'hbf8608a0} /* (10, 3, 6) {real, imag} */,
  {32'h3e4f1285, 32'hbfb5e374} /* (10, 3, 5) {real, imag} */,
  {32'hbd8b3520, 32'hbf891da2} /* (10, 3, 4) {real, imag} */,
  {32'h3f5c929d, 32'hbf379da6} /* (10, 3, 3) {real, imag} */,
  {32'h3f77706c, 32'h3e3f89be} /* (10, 3, 2) {real, imag} */,
  {32'h3e14d461, 32'h3e481f9c} /* (10, 3, 1) {real, imag} */,
  {32'hbed0d515, 32'h3d764510} /* (10, 3, 0) {real, imag} */,
  {32'hbdc78f00, 32'hbb822400} /* (10, 2, 15) {real, imag} */,
  {32'hbe5226c6, 32'hbcca1700} /* (10, 2, 14) {real, imag} */,
  {32'hbea4a17c, 32'hbf4899ca} /* (10, 2, 13) {real, imag} */,
  {32'hbf21205a, 32'hbf2d59ca} /* (10, 2, 12) {real, imag} */,
  {32'hbd87c5fb, 32'h3dd75e80} /* (10, 2, 11) {real, imag} */,
  {32'hbeebdecc, 32'h3f33aef3} /* (10, 2, 10) {real, imag} */,
  {32'h3eaef8cc, 32'hbc599f30} /* (10, 2, 9) {real, imag} */,
  {32'h3e5a5b64, 32'hbf342300} /* (10, 2, 8) {real, imag} */,
  {32'hbc053e05, 32'hbf5e4c0e} /* (10, 2, 7) {real, imag} */,
  {32'h3ec7a393, 32'hbf360808} /* (10, 2, 6) {real, imag} */,
  {32'h3f61eeeb, 32'hbfe4e93c} /* (10, 2, 5) {real, imag} */,
  {32'h3f4edf1c, 32'hbf971c3b} /* (10, 2, 4) {real, imag} */,
  {32'h3f1b5ab3, 32'hbee49f2a} /* (10, 2, 3) {real, imag} */,
  {32'h3f1b7cac, 32'h3d8ab958} /* (10, 2, 2) {real, imag} */,
  {32'hbe82d947, 32'h3e0793c0} /* (10, 2, 1) {real, imag} */,
  {32'hbf0527f2, 32'h3bcf52c0} /* (10, 2, 0) {real, imag} */,
  {32'hbe175f62, 32'hbea1ca07} /* (10, 1, 15) {real, imag} */,
  {32'h3eb74810, 32'h3e1d749c} /* (10, 1, 14) {real, imag} */,
  {32'h3f191f84, 32'h3e4d9f2c} /* (10, 1, 13) {real, imag} */,
  {32'h3e5d883e, 32'hbe34ffc2} /* (10, 1, 12) {real, imag} */,
  {32'hbf63fc88, 32'hbf1c1c08} /* (10, 1, 11) {real, imag} */,
  {32'hbf03b2f0, 32'hbed6f307} /* (10, 1, 10) {real, imag} */,
  {32'h3f4dd31a, 32'hbd888180} /* (10, 1, 9) {real, imag} */,
  {32'hbe363aca, 32'h3f2a6c3f} /* (10, 1, 8) {real, imag} */,
  {32'hbf02ba92, 32'hbefcff78} /* (10, 1, 7) {real, imag} */,
  {32'h3f0e45a2, 32'hbf68fa60} /* (10, 1, 6) {real, imag} */,
  {32'h3f3b0b5e, 32'hbee958bc} /* (10, 1, 5) {real, imag} */,
  {32'hbe308598, 32'h3e741144} /* (10, 1, 4) {real, imag} */,
  {32'hbe93506c, 32'h3f01d555} /* (10, 1, 3) {real, imag} */,
  {32'h3f20eb49, 32'h3e84b156} /* (10, 1, 2) {real, imag} */,
  {32'h3e681996, 32'hbece46d4} /* (10, 1, 1) {real, imag} */,
  {32'hbe866f92, 32'hbf012db5} /* (10, 1, 0) {real, imag} */,
  {32'hbef8877a, 32'hbc8b6502} /* (10, 0, 15) {real, imag} */,
  {32'h3e20a5e2, 32'h3ebc0d3a} /* (10, 0, 14) {real, imag} */,
  {32'h3f8f7940, 32'h3e844fa8} /* (10, 0, 13) {real, imag} */,
  {32'h3f2b539c, 32'hbddf4a0c} /* (10, 0, 12) {real, imag} */,
  {32'hbeab76af, 32'hbf1e7a28} /* (10, 0, 11) {real, imag} */,
  {32'hbed55b5c, 32'hbf2aa1e0} /* (10, 0, 10) {real, imag} */,
  {32'hbdb8761e, 32'hbefb9c08} /* (10, 0, 9) {real, imag} */,
  {32'h3d94e684, 32'h3d697270} /* (10, 0, 8) {real, imag} */,
  {32'hbdecf55c, 32'hbf37d952} /* (10, 0, 7) {real, imag} */,
  {32'hbdfb8b08, 32'hbf46134b} /* (10, 0, 6) {real, imag} */,
  {32'h3ea7e885, 32'h3e0811c0} /* (10, 0, 5) {real, imag} */,
  {32'h3e54faea, 32'h3e88df10} /* (10, 0, 4) {real, imag} */,
  {32'h3e2de110, 32'hbe4a959d} /* (10, 0, 3) {real, imag} */,
  {32'h3f16816a, 32'h3e14d302} /* (10, 0, 2) {real, imag} */,
  {32'h3ea6d938, 32'hbe7f8dce} /* (10, 0, 1) {real, imag} */,
  {32'hbd2e9ed8, 32'hbee3e2a0} /* (10, 0, 0) {real, imag} */,
  {32'h3c8efd84, 32'hbea39bc0} /* (9, 15, 15) {real, imag} */,
  {32'h3d22a5b0, 32'hbeb6d5f2} /* (9, 15, 14) {real, imag} */,
  {32'hbe2add17, 32'hbe806b94} /* (9, 15, 13) {real, imag} */,
  {32'h3bead378, 32'hbe03b8ae} /* (9, 15, 12) {real, imag} */,
  {32'hbea6a608, 32'h3d8facea} /* (9, 15, 11) {real, imag} */,
  {32'hbf4669e2, 32'hbe27f44c} /* (9, 15, 10) {real, imag} */,
  {32'hbf20d265, 32'hbe39e414} /* (9, 15, 9) {real, imag} */,
  {32'hbe5cb82c, 32'h3d82c640} /* (9, 15, 8) {real, imag} */,
  {32'h3e9d2270, 32'hbdf62a70} /* (9, 15, 7) {real, imag} */,
  {32'h3f0a2c8e, 32'h3d987251} /* (9, 15, 6) {real, imag} */,
  {32'h3f384ba8, 32'h3e3cbfb2} /* (9, 15, 5) {real, imag} */,
  {32'h3ee4c29c, 32'hbdc91890} /* (9, 15, 4) {real, imag} */,
  {32'h3ec6d69a, 32'hbe5d4728} /* (9, 15, 3) {real, imag} */,
  {32'h3e9e0f36, 32'h3be0f540} /* (9, 15, 2) {real, imag} */,
  {32'hbdedf2d0, 32'hbeed1b31} /* (9, 15, 1) {real, imag} */,
  {32'hbe6567ea, 32'hbeef01a0} /* (9, 15, 0) {real, imag} */,
  {32'h3e88a803, 32'hbbed9480} /* (9, 14, 15) {real, imag} */,
  {32'h3ee98cc0, 32'h3dfc31c0} /* (9, 14, 14) {real, imag} */,
  {32'h3d8c1528, 32'hbe7d3978} /* (9, 14, 13) {real, imag} */,
  {32'hbeb8a6ca, 32'hbe308a60} /* (9, 14, 12) {real, imag} */,
  {32'hbebee42b, 32'h3ea67723} /* (9, 14, 11) {real, imag} */,
  {32'hbe9210e3, 32'hbc3e9ec0} /* (9, 14, 10) {real, imag} */,
  {32'hbe1ea812, 32'h3c66a200} /* (9, 14, 9) {real, imag} */,
  {32'hbe18ed00, 32'h3e68a018} /* (9, 14, 8) {real, imag} */,
  {32'h3e5824f8, 32'hbe0f2b2c} /* (9, 14, 7) {real, imag} */,
  {32'h3ed7ebc5, 32'h3cf39720} /* (9, 14, 6) {real, imag} */,
  {32'h3f80a3e6, 32'h3e2e2b85} /* (9, 14, 5) {real, imag} */,
  {32'h3e525ace, 32'h3d8f6398} /* (9, 14, 4) {real, imag} */,
  {32'h3e07eb19, 32'hbe9308fc} /* (9, 14, 3) {real, imag} */,
  {32'h3e6d10df, 32'hbe1488c0} /* (9, 14, 2) {real, imag} */,
  {32'h3e60a7ce, 32'hbe3ecaf0} /* (9, 14, 1) {real, imag} */,
  {32'h3e610c97, 32'hbe93d35e} /* (9, 14, 0) {real, imag} */,
  {32'hbcf95c20, 32'h3ee0180c} /* (9, 13, 15) {real, imag} */,
  {32'h3f165b90, 32'h3f26deb2} /* (9, 13, 14) {real, imag} */,
  {32'h3ef454f1, 32'h3e79ff60} /* (9, 13, 13) {real, imag} */,
  {32'hbe851e70, 32'hbd57a650} /* (9, 13, 12) {real, imag} */,
  {32'hbf033260, 32'h3ecae558} /* (9, 13, 11) {real, imag} */,
  {32'hbe8f853a, 32'h3e6d81e8} /* (9, 13, 10) {real, imag} */,
  {32'h3e2634a8, 32'h3db1b720} /* (9, 13, 9) {real, imag} */,
  {32'h3e320717, 32'hbe8a0a4b} /* (9, 13, 8) {real, imag} */,
  {32'h3e4d024e, 32'hbf601281} /* (9, 13, 7) {real, imag} */,
  {32'hbe05fff8, 32'hbd87761a} /* (9, 13, 6) {real, imag} */,
  {32'h3e3dd241, 32'hbd80aa24} /* (9, 13, 5) {real, imag} */,
  {32'h3e1532ca, 32'hbe9aa4b6} /* (9, 13, 4) {real, imag} */,
  {32'hbe389718, 32'h3e77642e} /* (9, 13, 3) {real, imag} */,
  {32'hbd9eec1f, 32'h3e3d2a3c} /* (9, 13, 2) {real, imag} */,
  {32'h3e29cccc, 32'h3d321b60} /* (9, 13, 1) {real, imag} */,
  {32'h3d98c508, 32'h3da62cac} /* (9, 13, 0) {real, imag} */,
  {32'h3d54e6b4, 32'h3ea5b470} /* (9, 12, 15) {real, imag} */,
  {32'h3e90c9bc, 32'h3f489c07} /* (9, 12, 14) {real, imag} */,
  {32'h3d99df60, 32'h3dd0f720} /* (9, 12, 13) {real, imag} */,
  {32'hbdf57378, 32'hbef32d43} /* (9, 12, 12) {real, imag} */,
  {32'hbdd186f8, 32'hbf1838e0} /* (9, 12, 11) {real, imag} */,
  {32'hbe97f8e5, 32'hbf060930} /* (9, 12, 10) {real, imag} */,
  {32'hbf042255, 32'hbee718ee} /* (9, 12, 9) {real, imag} */,
  {32'hbecbd7f2, 32'hbf1f48a3} /* (9, 12, 8) {real, imag} */,
  {32'h3e0f5ac8, 32'hbed71fab} /* (9, 12, 7) {real, imag} */,
  {32'hbeb7b0b4, 32'hbe93646a} /* (9, 12, 6) {real, imag} */,
  {32'h3dd56b80, 32'hbf37a100} /* (9, 12, 5) {real, imag} */,
  {32'h3e65cc06, 32'hbf471e47} /* (9, 12, 4) {real, imag} */,
  {32'hbe3de50c, 32'h3d4839e0} /* (9, 12, 3) {real, imag} */,
  {32'hbdc4dba8, 32'h3e9b3364} /* (9, 12, 2) {real, imag} */,
  {32'h3e9d3b2c, 32'hbede69f6} /* (9, 12, 1) {real, imag} */,
  {32'h3ec62a99, 32'hbdddc160} /* (9, 12, 0) {real, imag} */,
  {32'hbe0b1712, 32'hbead6e27} /* (9, 11, 15) {real, imag} */,
  {32'hbdf34fdf, 32'hbed3a2bf} /* (9, 11, 14) {real, imag} */,
  {32'hbe95ec84, 32'hbefb028d} /* (9, 11, 13) {real, imag} */,
  {32'hbef66258, 32'h3e4a202c} /* (9, 11, 12) {real, imag} */,
  {32'h3e21e010, 32'h3f0d776a} /* (9, 11, 11) {real, imag} */,
  {32'hbe792c9f, 32'h3ea4a42a} /* (9, 11, 10) {real, imag} */,
  {32'hbf63ad74, 32'h3f162f85} /* (9, 11, 9) {real, imag} */,
  {32'hbf22c8b1, 32'h3efbe1dc} /* (9, 11, 8) {real, imag} */,
  {32'h3d5e3e20, 32'h3dba26b0} /* (9, 11, 7) {real, imag} */,
  {32'hbe1ead48, 32'hbe7075ec} /* (9, 11, 6) {real, imag} */,
  {32'h3e965813, 32'hbf0cb390} /* (9, 11, 5) {real, imag} */,
  {32'h3ed3d11d, 32'hbdc1edf4} /* (9, 11, 4) {real, imag} */,
  {32'h3c5f8580, 32'h3e3065e7} /* (9, 11, 3) {real, imag} */,
  {32'h3ecbf215, 32'hbd97f021} /* (9, 11, 2) {real, imag} */,
  {32'h3eea0b8c, 32'hbf5e7071} /* (9, 11, 1) {real, imag} */,
  {32'h3e8c792c, 32'hbf108028} /* (9, 11, 0) {real, imag} */,
  {32'hbf05c4e6, 32'hbea0199a} /* (9, 10, 15) {real, imag} */,
  {32'hbcde8610, 32'hbf21490c} /* (9, 10, 14) {real, imag} */,
  {32'hbd8789f7, 32'hbebee9e2} /* (9, 10, 13) {real, imag} */,
  {32'hbf10e4dc, 32'h3d4d1818} /* (9, 10, 12) {real, imag} */,
  {32'h3c1e7080, 32'h3ed807a2} /* (9, 10, 11) {real, imag} */,
  {32'hbe0e1540, 32'h3f3dc871} /* (9, 10, 10) {real, imag} */,
  {32'hbeaceb4a, 32'h3f4ceda7} /* (9, 10, 9) {real, imag} */,
  {32'hbeea7ca9, 32'h3eded186} /* (9, 10, 8) {real, imag} */,
  {32'h3d870bf4, 32'hbe5e12d8} /* (9, 10, 7) {real, imag} */,
  {32'hbdfe5d04, 32'hbef1f040} /* (9, 10, 6) {real, imag} */,
  {32'h3e4e7a98, 32'hbf215adf} /* (9, 10, 5) {real, imag} */,
  {32'h3ed6dfc4, 32'hbe540b42} /* (9, 10, 4) {real, imag} */,
  {32'hbe8d55c8, 32'hbe899e46} /* (9, 10, 3) {real, imag} */,
  {32'hbe3269e8, 32'hbd602c30} /* (9, 10, 2) {real, imag} */,
  {32'hbcdbc000, 32'hbeb1217c} /* (9, 10, 1) {real, imag} */,
  {32'hbd08eb30, 32'hbebfb9e6} /* (9, 10, 0) {real, imag} */,
  {32'hbf012a1e, 32'hbe8d35f8} /* (9, 9, 15) {real, imag} */,
  {32'h3d7508fe, 32'hbea9dac1} /* (9, 9, 14) {real, imag} */,
  {32'hbdb7b9f2, 32'h3dc4f6f4} /* (9, 9, 13) {real, imag} */,
  {32'hbe9bccca, 32'h3dc85640} /* (9, 9, 12) {real, imag} */,
  {32'h3ec7a57d, 32'h3e540898} /* (9, 9, 11) {real, imag} */,
  {32'hbe0a1c20, 32'h3ef122a2} /* (9, 9, 10) {real, imag} */,
  {32'hbe7a1808, 32'h3e4d3524} /* (9, 9, 9) {real, imag} */,
  {32'hbe805c2c, 32'hbee31a88} /* (9, 9, 8) {real, imag} */,
  {32'hbe65fc32, 32'hbf2bdc2c} /* (9, 9, 7) {real, imag} */,
  {32'h3e527e34, 32'hbf13b2ce} /* (9, 9, 6) {real, imag} */,
  {32'h3f0c64e7, 32'hbf4c42c3} /* (9, 9, 5) {real, imag} */,
  {32'h3e7d93da, 32'hbefc917c} /* (9, 9, 4) {real, imag} */,
  {32'h3e750698, 32'hbf1643fd} /* (9, 9, 3) {real, imag} */,
  {32'hbcf45420, 32'hbe88e31f} /* (9, 9, 2) {real, imag} */,
  {32'h3e347bf0, 32'h3d8fdcd8} /* (9, 9, 1) {real, imag} */,
  {32'h3e394ed0, 32'h3e7eba60} /* (9, 9, 0) {real, imag} */,
  {32'hbd0ecdac, 32'hbf04f7de} /* (9, 8, 15) {real, imag} */,
  {32'h3e7a36f4, 32'hbedaa627} /* (9, 8, 14) {real, imag} */,
  {32'hbeb6ea52, 32'h3cdf7330} /* (9, 8, 13) {real, imag} */,
  {32'hbf0e005d, 32'hbeb9f7c6} /* (9, 8, 12) {real, imag} */,
  {32'h3e823e49, 32'hbd884900} /* (9, 8, 11) {real, imag} */,
  {32'h3e76134c, 32'h3f1d48d7} /* (9, 8, 10) {real, imag} */,
  {32'h3e6028a8, 32'h3f0a3b1c} /* (9, 8, 9) {real, imag} */,
  {32'h3defda3c, 32'h3f62795e} /* (9, 8, 8) {real, imag} */,
  {32'h3c1a37c0, 32'h3d7d5f10} /* (9, 8, 7) {real, imag} */,
  {32'h3ea3b3ee, 32'hbe9a72ac} /* (9, 8, 6) {real, imag} */,
  {32'h3edbb2e2, 32'hbed175dc} /* (9, 8, 5) {real, imag} */,
  {32'h3e89ea94, 32'h3e1250f8} /* (9, 8, 4) {real, imag} */,
  {32'h3f1b4f96, 32'hbdd271c0} /* (9, 8, 3) {real, imag} */,
  {32'h3eccb5ca, 32'hbea25cee} /* (9, 8, 2) {real, imag} */,
  {32'h3ea2796b, 32'h3db70630} /* (9, 8, 1) {real, imag} */,
  {32'h3ea5052d, 32'h3e097110} /* (9, 8, 0) {real, imag} */,
  {32'hbd37a648, 32'hbeeeeb6a} /* (9, 7, 15) {real, imag} */,
  {32'hbe44784e, 32'hbeb7a8fa} /* (9, 7, 14) {real, imag} */,
  {32'hbe2d3517, 32'hbd318e00} /* (9, 7, 13) {real, imag} */,
  {32'hbe79f352, 32'hbf68a99f} /* (9, 7, 12) {real, imag} */,
  {32'h3e935d4e, 32'hbebd3064} /* (9, 7, 11) {real, imag} */,
  {32'h3e8566b7, 32'h3f62bd5b} /* (9, 7, 10) {real, imag} */,
  {32'h3f458dac, 32'h3ec573d8} /* (9, 7, 9) {real, imag} */,
  {32'h3eab90e4, 32'h3f095154} /* (9, 7, 8) {real, imag} */,
  {32'hbe9e36b2, 32'hbe19dc81} /* (9, 7, 7) {real, imag} */,
  {32'h3e773ee8, 32'hbe713420} /* (9, 7, 6) {real, imag} */,
  {32'h3eadd7ae, 32'h3edbdd82} /* (9, 7, 5) {real, imag} */,
  {32'hbe41d72c, 32'h3e8d705b} /* (9, 7, 4) {real, imag} */,
  {32'hbe54527c, 32'hbf132e15} /* (9, 7, 3) {real, imag} */,
  {32'hbe50b74c, 32'hbf4e0ede} /* (9, 7, 2) {real, imag} */,
  {32'hbe82bd0e, 32'hbededd59} /* (9, 7, 1) {real, imag} */,
  {32'hbe8f13e8, 32'hbea7d038} /* (9, 7, 0) {real, imag} */,
  {32'h3d6731b4, 32'hbed6ba43} /* (9, 6, 15) {real, imag} */,
  {32'hbd47a900, 32'hbe6871a4} /* (9, 6, 14) {real, imag} */,
  {32'h3e1d8529, 32'hbe65762c} /* (9, 6, 13) {real, imag} */,
  {32'h3def22f0, 32'hbe5a2ec4} /* (9, 6, 12) {real, imag} */,
  {32'h3d20f4b8, 32'h3e8180fa} /* (9, 6, 11) {real, imag} */,
  {32'h3d656040, 32'h3ea7ea09} /* (9, 6, 10) {real, imag} */,
  {32'h3f809f4b, 32'hbea85bec} /* (9, 6, 9) {real, imag} */,
  {32'h3eb1c3c2, 32'hbe857edc} /* (9, 6, 8) {real, imag} */,
  {32'hbe95f7fc, 32'hbf4e0f86} /* (9, 6, 7) {real, imag} */,
  {32'hbdc10500, 32'hbf1edb2c} /* (9, 6, 6) {real, imag} */,
  {32'hbe5df958, 32'h3f480432} /* (9, 6, 5) {real, imag} */,
  {32'hbee17ff4, 32'h3f557004} /* (9, 6, 4) {real, imag} */,
  {32'hbef00b0e, 32'hbeb57280} /* (9, 6, 3) {real, imag} */,
  {32'hbf0a2018, 32'hbfa2437d} /* (9, 6, 2) {real, imag} */,
  {32'h3d9a7348, 32'hbf1511b8} /* (9, 6, 1) {real, imag} */,
  {32'hbdc3a688, 32'hbd6d434c} /* (9, 6, 0) {real, imag} */,
  {32'h3e56bf72, 32'hbe256c00} /* (9, 5, 15) {real, imag} */,
  {32'h3b35da00, 32'h3e7a7440} /* (9, 5, 14) {real, imag} */,
  {32'hbebdb9ca, 32'hbde2d028} /* (9, 5, 13) {real, imag} */,
  {32'hbe40ba02, 32'hbe59f560} /* (9, 5, 12) {real, imag} */,
  {32'h3e5ffa82, 32'h3d5cfd40} /* (9, 5, 11) {real, imag} */,
  {32'h3f0c07bf, 32'hbe2bc6b8} /* (9, 5, 10) {real, imag} */,
  {32'h3f8d5e2a, 32'hbf112b46} /* (9, 5, 9) {real, imag} */,
  {32'h3effd038, 32'hbf43dabe} /* (9, 5, 8) {real, imag} */,
  {32'hbcc50868, 32'hbf0b767a} /* (9, 5, 7) {real, imag} */,
  {32'h3d1ea2a0, 32'hbefadd31} /* (9, 5, 6) {real, imag} */,
  {32'hbde8c900, 32'h3dd27634} /* (9, 5, 5) {real, imag} */,
  {32'hbe0039cc, 32'hbd9d1830} /* (9, 5, 4) {real, imag} */,
  {32'hbe981762, 32'hbedc865c} /* (9, 5, 3) {real, imag} */,
  {32'hbea89648, 32'hbf5df201} /* (9, 5, 2) {real, imag} */,
  {32'h3d8fa060, 32'hbf0d52ec} /* (9, 5, 1) {real, imag} */,
  {32'hbe3e61b4, 32'h3d037696} /* (9, 5, 0) {real, imag} */,
  {32'h3ef1e344, 32'hbe30c8bc} /* (9, 4, 15) {real, imag} */,
  {32'h3deaeb00, 32'h3dae1414} /* (9, 4, 14) {real, imag} */,
  {32'hbe800cd4, 32'hbde9a610} /* (9, 4, 13) {real, imag} */,
  {32'h3dcc570e, 32'hbe23e4f4} /* (9, 4, 12) {real, imag} */,
  {32'h3eeee750, 32'h3e670f98} /* (9, 4, 11) {real, imag} */,
  {32'h3d1f1960, 32'h3e03aaf8} /* (9, 4, 10) {real, imag} */,
  {32'h3f2795a6, 32'hbef312bb} /* (9, 4, 9) {real, imag} */,
  {32'h3e24ed14, 32'hbe8c9462} /* (9, 4, 8) {real, imag} */,
  {32'hbe89623a, 32'h3e1313e8} /* (9, 4, 7) {real, imag} */,
  {32'h3e5f1c48, 32'h3d4554f8} /* (9, 4, 6) {real, imag} */,
  {32'h3ed07f50, 32'h3f205bd6} /* (9, 4, 5) {real, imag} */,
  {32'h3ae41000, 32'h3e6079ae} /* (9, 4, 4) {real, imag} */,
  {32'hbe9e1122, 32'hbeced884} /* (9, 4, 3) {real, imag} */,
  {32'hbf2bef6c, 32'hbea5efd4} /* (9, 4, 2) {real, imag} */,
  {32'hbe7d1538, 32'hbe83294e} /* (9, 4, 1) {real, imag} */,
  {32'hbe27e51f, 32'hbe5ea8a0} /* (9, 4, 0) {real, imag} */,
  {32'h3ebfaf5e, 32'h3e43f6f0} /* (9, 3, 15) {real, imag} */,
  {32'h3f2b07e7, 32'h3f15dcca} /* (9, 3, 14) {real, imag} */,
  {32'h3f03774c, 32'hbccf4418} /* (9, 3, 13) {real, imag} */,
  {32'h3dc5b088, 32'hbe9e7d71} /* (9, 3, 12) {real, imag} */,
  {32'h3e3aafb2, 32'h3e25eb40} /* (9, 3, 11) {real, imag} */,
  {32'hbe40a108, 32'h3f1fbdec} /* (9, 3, 10) {real, imag} */,
  {32'hbdb77fcc, 32'h3c919a30} /* (9, 3, 9) {real, imag} */,
  {32'hbed08b8e, 32'hbe1bd4fc} /* (9, 3, 8) {real, imag} */,
  {32'hbec6879b, 32'h3e787994} /* (9, 3, 7) {real, imag} */,
  {32'hbe7676d8, 32'h3f244b40} /* (9, 3, 6) {real, imag} */,
  {32'h3eb6d324, 32'h3f27e752} /* (9, 3, 5) {real, imag} */,
  {32'hbdb286f4, 32'h3df737e0} /* (9, 3, 4) {real, imag} */,
  {32'hbe48c0b2, 32'hbef83b24} /* (9, 3, 3) {real, imag} */,
  {32'hbed570e5, 32'hbee0871c} /* (9, 3, 2) {real, imag} */,
  {32'hbd81d83c, 32'h3e578326} /* (9, 3, 1) {real, imag} */,
  {32'hbd703440, 32'hbdd028ac} /* (9, 3, 0) {real, imag} */,
  {32'h3f156b11, 32'hbe53bb70} /* (9, 2, 15) {real, imag} */,
  {32'h3f5c4b12, 32'hbe2ea738} /* (9, 2, 14) {real, imag} */,
  {32'h3f1d5cc4, 32'hbd6de89c} /* (9, 2, 13) {real, imag} */,
  {32'h3e9e8102, 32'hbe71e741} /* (9, 2, 12) {real, imag} */,
  {32'h3e4f29ea, 32'h3d5bf4e6} /* (9, 2, 11) {real, imag} */,
  {32'h3ea97f2e, 32'h3f34e53e} /* (9, 2, 10) {real, imag} */,
  {32'hbea207ca, 32'h3f039817} /* (9, 2, 9) {real, imag} */,
  {32'hbeac40ba, 32'h3e8f2666} /* (9, 2, 8) {real, imag} */,
  {32'hbe8aba83, 32'h3d87859e} /* (9, 2, 7) {real, imag} */,
  {32'hbf127b7e, 32'h3e807172} /* (9, 2, 6) {real, imag} */,
  {32'hbdbd9a50, 32'h3f0037ac} /* (9, 2, 5) {real, imag} */,
  {32'h3d9b8df8, 32'h3e460722} /* (9, 2, 4) {real, imag} */,
  {32'hbe7850ab, 32'hbe1dd656} /* (9, 2, 3) {real, imag} */,
  {32'hbecb2519, 32'hbd9de694} /* (9, 2, 2) {real, imag} */,
  {32'h3e7ec742, 32'hbeb2a966} /* (9, 2, 1) {real, imag} */,
  {32'h3d4e1570, 32'hbe8259b3} /* (9, 2, 0) {real, imag} */,
  {32'h3e7208b3, 32'hbec5bbf8} /* (9, 1, 15) {real, imag} */,
  {32'h3edb4f13, 32'hbf17f633} /* (9, 1, 14) {real, imag} */,
  {32'h3d8096f0, 32'hbe1f9b8c} /* (9, 1, 13) {real, imag} */,
  {32'h3d714430, 32'h3f0e871f} /* (9, 1, 12) {real, imag} */,
  {32'h3ed5b19e, 32'h3f74bae9} /* (9, 1, 11) {real, imag} */,
  {32'h3edbe3cf, 32'h3eec6761} /* (9, 1, 10) {real, imag} */,
  {32'hbddbba20, 32'hbe20cc1a} /* (9, 1, 9) {real, imag} */,
  {32'hbebdc5c0, 32'h3dc00bd8} /* (9, 1, 8) {real, imag} */,
  {32'h3e78010c, 32'hbe85c2a6} /* (9, 1, 7) {real, imag} */,
  {32'hbe0c5860, 32'hbe5d0368} /* (9, 1, 6) {real, imag} */,
  {32'hbf18e598, 32'hbeb99aec} /* (9, 1, 5) {real, imag} */,
  {32'h3dd41ee0, 32'hbee584ab} /* (9, 1, 4) {real, imag} */,
  {32'hb9fb7000, 32'hbd2d13a4} /* (9, 1, 3) {real, imag} */,
  {32'hbf1f6bf0, 32'h3ebfacb8} /* (9, 1, 2) {real, imag} */,
  {32'hbecb745f, 32'h3c59b600} /* (9, 1, 1) {real, imag} */,
  {32'h3d62d74c, 32'h3c1ffe60} /* (9, 1, 0) {real, imag} */,
  {32'hbde4896e, 32'hbe0b1aac} /* (9, 0, 15) {real, imag} */,
  {32'hbec67eba, 32'h3d89f760} /* (9, 0, 14) {real, imag} */,
  {32'hbf06b304, 32'h3e94ea02} /* (9, 0, 13) {real, imag} */,
  {32'h3cbb1a40, 32'h3f0f5f0d} /* (9, 0, 12) {real, imag} */,
  {32'h3e396d7e, 32'h3f5814ca} /* (9, 0, 11) {real, imag} */,
  {32'hbdfd8f50, 32'hbba1ec20} /* (9, 0, 10) {real, imag} */,
  {32'hbe5489cc, 32'hbee679c0} /* (9, 0, 9) {real, imag} */,
  {32'hbda9cd2e, 32'hbdd5e89e} /* (9, 0, 8) {real, imag} */,
  {32'h3e0b46ca, 32'hbf14cff2} /* (9, 0, 7) {real, imag} */,
  {32'hbd2fd36a, 32'hbedbe637} /* (9, 0, 6) {real, imag} */,
  {32'hbed3ab06, 32'hbe9c015e} /* (9, 0, 5) {real, imag} */,
  {32'h3d1511a0, 32'hbe4dd2a7} /* (9, 0, 4) {real, imag} */,
  {32'h3eecd7d0, 32'hbd0315a8} /* (9, 0, 3) {real, imag} */,
  {32'h3eb77dd5, 32'h3e584dbd} /* (9, 0, 2) {real, imag} */,
  {32'hbda33cac, 32'h3e55f2b5} /* (9, 0, 1) {real, imag} */,
  {32'h3d14e870, 32'h3db974c0} /* (9, 0, 0) {real, imag} */,
  {32'h3ecfff46, 32'h00000000} /* (8, 15, 15) {real, imag} */,
  {32'h3e379b76, 32'h00000000} /* (8, 15, 14) {real, imag} */,
  {32'h3db3aa70, 32'h00000000} /* (8, 15, 13) {real, imag} */,
  {32'h3e730884, 32'h00000000} /* (8, 15, 12) {real, imag} */,
  {32'h3e53dac0, 32'h00000000} /* (8, 15, 11) {real, imag} */,
  {32'hbe2a033c, 32'h00000000} /* (8, 15, 10) {real, imag} */,
  {32'hbe652300, 32'h00000000} /* (8, 15, 9) {real, imag} */,
  {32'h3c2e0b80, 32'h00000000} /* (8, 15, 8) {real, imag} */,
  {32'hbe863630, 32'h00000000} /* (8, 15, 7) {real, imag} */,
  {32'hbdb66c40, 32'h00000000} /* (8, 15, 6) {real, imag} */,
  {32'h3d429a40, 32'h00000000} /* (8, 15, 5) {real, imag} */,
  {32'hbdb85058, 32'h00000000} /* (8, 15, 4) {real, imag} */,
  {32'h3983d000, 32'h00000000} /* (8, 15, 3) {real, imag} */,
  {32'h3e0af8b4, 32'h00000000} /* (8, 15, 2) {real, imag} */,
  {32'hbecf0087, 32'h00000000} /* (8, 15, 1) {real, imag} */,
  {32'hbedc48c4, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'h3f34e6a4, 32'h00000000} /* (8, 14, 15) {real, imag} */,
  {32'h3dcd360c, 32'h00000000} /* (8, 14, 14) {real, imag} */,
  {32'hbe328768, 32'h00000000} /* (8, 14, 13) {real, imag} */,
  {32'hbde505c8, 32'h00000000} /* (8, 14, 12) {real, imag} */,
  {32'hbb63fa00, 32'h00000000} /* (8, 14, 11) {real, imag} */,
  {32'hbf12323c, 32'h00000000} /* (8, 14, 10) {real, imag} */,
  {32'hbfb3607c, 32'h00000000} /* (8, 14, 9) {real, imag} */,
  {32'hbf366c94, 32'h00000000} /* (8, 14, 8) {real, imag} */,
  {32'hbf0168c0, 32'h00000000} /* (8, 14, 7) {real, imag} */,
  {32'hbec80654, 32'h00000000} /* (8, 14, 6) {real, imag} */,
  {32'hbf23ccde, 32'h00000000} /* (8, 14, 5) {real, imag} */,
  {32'hbe5e3ddc, 32'h00000000} /* (8, 14, 4) {real, imag} */,
  {32'h3ef3482c, 32'h00000000} /* (8, 14, 3) {real, imag} */,
  {32'h3f30ca38, 32'h00000000} /* (8, 14, 2) {real, imag} */,
  {32'h3e8b74ca, 32'h00000000} /* (8, 14, 1) {real, imag} */,
  {32'hbd77a0a0, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'h3f4bbe26, 32'h00000000} /* (8, 13, 15) {real, imag} */,
  {32'hbd6db280, 32'h00000000} /* (8, 13, 14) {real, imag} */,
  {32'hbe6e24a8, 32'h00000000} /* (8, 13, 13) {real, imag} */,
  {32'hbd022378, 32'h00000000} /* (8, 13, 12) {real, imag} */,
  {32'hbd1709ec, 32'h00000000} /* (8, 13, 11) {real, imag} */,
  {32'h3ccacce0, 32'h00000000} /* (8, 13, 10) {real, imag} */,
  {32'hbf76c0c3, 32'h00000000} /* (8, 13, 9) {real, imag} */,
  {32'hbf6fff7e, 32'h00000000} /* (8, 13, 8) {real, imag} */,
  {32'hbeabbf74, 32'h00000000} /* (8, 13, 7) {real, imag} */,
  {32'hbe0fb360, 32'h00000000} /* (8, 13, 6) {real, imag} */,
  {32'h3d31a210, 32'h00000000} /* (8, 13, 5) {real, imag} */,
  {32'h3e124c7c, 32'h00000000} /* (8, 13, 4) {real, imag} */,
  {32'h3d953b18, 32'h00000000} /* (8, 13, 3) {real, imag} */,
  {32'hbd567a00, 32'h00000000} /* (8, 13, 2) {real, imag} */,
  {32'h3e84cc60, 32'h00000000} /* (8, 13, 1) {real, imag} */,
  {32'h3eb186e0, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'h3e37d46a, 32'h00000000} /* (8, 12, 15) {real, imag} */,
  {32'h3dd521c4, 32'h00000000} /* (8, 12, 14) {real, imag} */,
  {32'hbe4550a6, 32'h00000000} /* (8, 12, 13) {real, imag} */,
  {32'hbf1a2c37, 32'h00000000} /* (8, 12, 12) {real, imag} */,
  {32'hbf331292, 32'h00000000} /* (8, 12, 11) {real, imag} */,
  {32'hbe0f28cc, 32'h00000000} /* (8, 12, 10) {real, imag} */,
  {32'h3d779040, 32'h00000000} /* (8, 12, 9) {real, imag} */,
  {32'h3d32f208, 32'h00000000} /* (8, 12, 8) {real, imag} */,
  {32'h3eb363ca, 32'h00000000} /* (8, 12, 7) {real, imag} */,
  {32'h3f640e5a, 32'h00000000} /* (8, 12, 6) {real, imag} */,
  {32'h3f27c502, 32'h00000000} /* (8, 12, 5) {real, imag} */,
  {32'hbdff4e58, 32'h00000000} /* (8, 12, 4) {real, imag} */,
  {32'h3d03e1d0, 32'h00000000} /* (8, 12, 3) {real, imag} */,
  {32'hbd54fae0, 32'h00000000} /* (8, 12, 2) {real, imag} */,
  {32'h3eceaf48, 32'h00000000} /* (8, 12, 1) {real, imag} */,
  {32'h3e92f598, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'h3d28cfd8, 32'h00000000} /* (8, 11, 15) {real, imag} */,
  {32'h3f066668, 32'h00000000} /* (8, 11, 14) {real, imag} */,
  {32'h3da1c820, 32'h00000000} /* (8, 11, 13) {real, imag} */,
  {32'hbefad9a8, 32'h00000000} /* (8, 11, 12) {real, imag} */,
  {32'hbf73a19d, 32'h00000000} /* (8, 11, 11) {real, imag} */,
  {32'hbf0c3586, 32'h00000000} /* (8, 11, 10) {real, imag} */,
  {32'h3f104818, 32'h00000000} /* (8, 11, 9) {real, imag} */,
  {32'h3f7645d2, 32'h00000000} /* (8, 11, 8) {real, imag} */,
  {32'h3f4e69a4, 32'h00000000} /* (8, 11, 7) {real, imag} */,
  {32'h3eb02e39, 32'h00000000} /* (8, 11, 6) {real, imag} */,
  {32'h3c8abec0, 32'h00000000} /* (8, 11, 5) {real, imag} */,
  {32'hbdcec300, 32'h00000000} /* (8, 11, 4) {real, imag} */,
  {32'h3e616a60, 32'h00000000} /* (8, 11, 3) {real, imag} */,
  {32'h3dcee168, 32'h00000000} /* (8, 11, 2) {real, imag} */,
  {32'h3da0e7f8, 32'h00000000} /* (8, 11, 1) {real, imag} */,
  {32'h3e0927f8, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h3ed4ca97, 32'h00000000} /* (8, 10, 15) {real, imag} */,
  {32'h3eb1c8ab, 32'h00000000} /* (8, 10, 14) {real, imag} */,
  {32'hbc4ba2c0, 32'h00000000} /* (8, 10, 13) {real, imag} */,
  {32'hbe78a010, 32'h00000000} /* (8, 10, 12) {real, imag} */,
  {32'hbee9e268, 32'h00000000} /* (8, 10, 11) {real, imag} */,
  {32'hbf069b08, 32'h00000000} /* (8, 10, 10) {real, imag} */,
  {32'hbef9af48, 32'h00000000} /* (8, 10, 9) {real, imag} */,
  {32'h3e9c60d6, 32'h00000000} /* (8, 10, 8) {real, imag} */,
  {32'hbdd41a98, 32'h00000000} /* (8, 10, 7) {real, imag} */,
  {32'h3e808ffa, 32'h00000000} /* (8, 10, 6) {real, imag} */,
  {32'hbe30afac, 32'h00000000} /* (8, 10, 5) {real, imag} */,
  {32'hbe710ee0, 32'h00000000} /* (8, 10, 4) {real, imag} */,
  {32'hbdbe1900, 32'h00000000} /* (8, 10, 3) {real, imag} */,
  {32'hbe23d132, 32'h00000000} /* (8, 10, 2) {real, imag} */,
  {32'h3e161a00, 32'h00000000} /* (8, 10, 1) {real, imag} */,
  {32'h3f146363, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'h3c6aee00, 32'h00000000} /* (8, 9, 15) {real, imag} */,
  {32'hbe58e748, 32'h00000000} /* (8, 9, 14) {real, imag} */,
  {32'h3e1bfa18, 32'h00000000} /* (8, 9, 13) {real, imag} */,
  {32'h3f1e0a33, 32'h00000000} /* (8, 9, 12) {real, imag} */,
  {32'h3f155180, 32'h00000000} /* (8, 9, 11) {real, imag} */,
  {32'h3ec93870, 32'h00000000} /* (8, 9, 10) {real, imag} */,
  {32'hbcd41580, 32'h00000000} /* (8, 9, 9) {real, imag} */,
  {32'h3e8e24f8, 32'h00000000} /* (8, 9, 8) {real, imag} */,
  {32'h3e58b3cc, 32'h00000000} /* (8, 9, 7) {real, imag} */,
  {32'h3e58ced4, 32'h00000000} /* (8, 9, 6) {real, imag} */,
  {32'hbefa739a, 32'h00000000} /* (8, 9, 5) {real, imag} */,
  {32'hbf22cc23, 32'h00000000} /* (8, 9, 4) {real, imag} */,
  {32'hbe1158c2, 32'h00000000} /* (8, 9, 3) {real, imag} */,
  {32'h3ddfe2e8, 32'h00000000} /* (8, 9, 2) {real, imag} */,
  {32'h3dbae1a0, 32'h00000000} /* (8, 9, 1) {real, imag} */,
  {32'h3eb8e450, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'h3ef76e34, 32'h00000000} /* (8, 8, 15) {real, imag} */,
  {32'h3efc6314, 32'h00000000} /* (8, 8, 14) {real, imag} */,
  {32'h3f2da0e5, 32'h00000000} /* (8, 8, 13) {real, imag} */,
  {32'h3ede2570, 32'h00000000} /* (8, 8, 12) {real, imag} */,
  {32'h3f1099e0, 32'h00000000} /* (8, 8, 11) {real, imag} */,
  {32'h3e79c7ee, 32'h00000000} /* (8, 8, 10) {real, imag} */,
  {32'hbe1125b9, 32'h00000000} /* (8, 8, 9) {real, imag} */,
  {32'h3ed17934, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'h3eaecb34, 32'h00000000} /* (8, 8, 7) {real, imag} */,
  {32'hbeef015e, 32'h00000000} /* (8, 8, 6) {real, imag} */,
  {32'hbf853786, 32'h00000000} /* (8, 8, 5) {real, imag} */,
  {32'hbf76c9d9, 32'h00000000} /* (8, 8, 4) {real, imag} */,
  {32'hbf1d9478, 32'h00000000} /* (8, 8, 3) {real, imag} */,
  {32'hbe495728, 32'h00000000} /* (8, 8, 2) {real, imag} */,
  {32'hbe112824, 32'h00000000} /* (8, 8, 1) {real, imag} */,
  {32'h3e81b249, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h3ede48ec, 32'h00000000} /* (8, 7, 15) {real, imag} */,
  {32'h3eec61e2, 32'h00000000} /* (8, 7, 14) {real, imag} */,
  {32'h3eda3f78, 32'h00000000} /* (8, 7, 13) {real, imag} */,
  {32'hbe69ebd8, 32'h00000000} /* (8, 7, 12) {real, imag} */,
  {32'h3f46f67b, 32'h00000000} /* (8, 7, 11) {real, imag} */,
  {32'h3e5527e6, 32'h00000000} /* (8, 7, 10) {real, imag} */,
  {32'h3e1b0e22, 32'h00000000} /* (8, 7, 9) {real, imag} */,
  {32'h3ecca934, 32'h00000000} /* (8, 7, 8) {real, imag} */,
  {32'h3d84d428, 32'h00000000} /* (8, 7, 7) {real, imag} */,
  {32'hbefd8e63, 32'h00000000} /* (8, 7, 6) {real, imag} */,
  {32'hbf15a27e, 32'h00000000} /* (8, 7, 5) {real, imag} */,
  {32'hbe1c1768, 32'h00000000} /* (8, 7, 4) {real, imag} */,
  {32'hbea07140, 32'h00000000} /* (8, 7, 3) {real, imag} */,
  {32'hbe480b44, 32'h00000000} /* (8, 7, 2) {real, imag} */,
  {32'hbe37d708, 32'h00000000} /* (8, 7, 1) {real, imag} */,
  {32'h3f0a883e, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h3e12e7e4, 32'h00000000} /* (8, 6, 15) {real, imag} */,
  {32'h3d3e2d80, 32'h00000000} /* (8, 6, 14) {real, imag} */,
  {32'hbe7abaf0, 32'h00000000} /* (8, 6, 13) {real, imag} */,
  {32'hbe04b060, 32'h00000000} /* (8, 6, 12) {real, imag} */,
  {32'h3f1b9f8e, 32'h00000000} /* (8, 6, 11) {real, imag} */,
  {32'hbf084167, 32'h00000000} /* (8, 6, 10) {real, imag} */,
  {32'hbf22548a, 32'h00000000} /* (8, 6, 9) {real, imag} */,
  {32'hbea98820, 32'h00000000} /* (8, 6, 8) {real, imag} */,
  {32'hbf688ef8, 32'h00000000} /* (8, 6, 7) {real, imag} */,
  {32'hbc988440, 32'h00000000} /* (8, 6, 6) {real, imag} */,
  {32'h3f23cb1f, 32'h00000000} /* (8, 6, 5) {real, imag} */,
  {32'h3f7b5743, 32'h00000000} /* (8, 6, 4) {real, imag} */,
  {32'h3ea7dd7c, 32'h00000000} /* (8, 6, 3) {real, imag} */,
  {32'h3e9a0290, 32'h00000000} /* (8, 6, 2) {real, imag} */,
  {32'hbe3a95e0, 32'h00000000} /* (8, 6, 1) {real, imag} */,
  {32'hbe365fb0, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'hbe819316, 32'h00000000} /* (8, 5, 15) {real, imag} */,
  {32'h3d221bc8, 32'h00000000} /* (8, 5, 14) {real, imag} */,
  {32'hbe8675ce, 32'h00000000} /* (8, 5, 13) {real, imag} */,
  {32'hbe345868, 32'h00000000} /* (8, 5, 12) {real, imag} */,
  {32'h3e516ec8, 32'h00000000} /* (8, 5, 11) {real, imag} */,
  {32'hbe581554, 32'h00000000} /* (8, 5, 10) {real, imag} */,
  {32'hbeec8aa0, 32'h00000000} /* (8, 5, 9) {real, imag} */,
  {32'hbefb2a1e, 32'h00000000} /* (8, 5, 8) {real, imag} */,
  {32'hbf3e05cc, 32'h00000000} /* (8, 5, 7) {real, imag} */,
  {32'hbdd61a80, 32'h00000000} /* (8, 5, 6) {real, imag} */,
  {32'h3e880450, 32'h00000000} /* (8, 5, 5) {real, imag} */,
  {32'hbd90f980, 32'h00000000} /* (8, 5, 4) {real, imag} */,
  {32'hbf06129c, 32'h00000000} /* (8, 5, 3) {real, imag} */,
  {32'hbec15170, 32'h00000000} /* (8, 5, 2) {real, imag} */,
  {32'h3e152e66, 32'h00000000} /* (8, 5, 1) {real, imag} */,
  {32'hbeef4e38, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'hbd75d160, 32'h00000000} /* (8, 4, 15) {real, imag} */,
  {32'h3e4aead4, 32'h00000000} /* (8, 4, 14) {real, imag} */,
  {32'h3e59256c, 32'h00000000} /* (8, 4, 13) {real, imag} */,
  {32'h3e955ce0, 32'h00000000} /* (8, 4, 12) {real, imag} */,
  {32'h3e588d6a, 32'h00000000} /* (8, 4, 11) {real, imag} */,
  {32'h3f0aef88, 32'h00000000} /* (8, 4, 10) {real, imag} */,
  {32'h3f171838, 32'h00000000} /* (8, 4, 9) {real, imag} */,
  {32'h3e498174, 32'h00000000} /* (8, 4, 8) {real, imag} */,
  {32'hbea80258, 32'h00000000} /* (8, 4, 7) {real, imag} */,
  {32'h3d3381e0, 32'h00000000} /* (8, 4, 6) {real, imag} */,
  {32'h3dba8abc, 32'h00000000} /* (8, 4, 5) {real, imag} */,
  {32'hbeeae9ee, 32'h00000000} /* (8, 4, 4) {real, imag} */,
  {32'hbf313ed0, 32'h00000000} /* (8, 4, 3) {real, imag} */,
  {32'hbdeaf0ac, 32'h00000000} /* (8, 4, 2) {real, imag} */,
  {32'h3f16c726, 32'h00000000} /* (8, 4, 1) {real, imag} */,
  {32'h3e28df9c, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'hbdd95ed0, 32'h00000000} /* (8, 3, 15) {real, imag} */,
  {32'hbe1fa3a2, 32'h00000000} /* (8, 3, 14) {real, imag} */,
  {32'h3e3f1a10, 32'h00000000} /* (8, 3, 13) {real, imag} */,
  {32'h3ebbcda0, 32'h00000000} /* (8, 3, 12) {real, imag} */,
  {32'hbcaf4a80, 32'h00000000} /* (8, 3, 11) {real, imag} */,
  {32'h3f42f381, 32'h00000000} /* (8, 3, 10) {real, imag} */,
  {32'h3ed12b85, 32'h00000000} /* (8, 3, 9) {real, imag} */,
  {32'hbc8910c0, 32'h00000000} /* (8, 3, 8) {real, imag} */,
  {32'h3e0c59af, 32'h00000000} /* (8, 3, 7) {real, imag} */,
  {32'h3f916782, 32'h00000000} /* (8, 3, 6) {real, imag} */,
  {32'h3f287106, 32'h00000000} /* (8, 3, 5) {real, imag} */,
  {32'h3f1b2402, 32'h00000000} /* (8, 3, 4) {real, imag} */,
  {32'hbd7ea348, 32'h00000000} /* (8, 3, 3) {real, imag} */,
  {32'h3df0c114, 32'h00000000} /* (8, 3, 2) {real, imag} */,
  {32'h3d8f4a6c, 32'h00000000} /* (8, 3, 1) {real, imag} */,
  {32'h3df03560, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'hbe11c28c, 32'h00000000} /* (8, 2, 15) {real, imag} */,
  {32'hbdcc6550, 32'h00000000} /* (8, 2, 14) {real, imag} */,
  {32'hbe87a35e, 32'h00000000} /* (8, 2, 13) {real, imag} */,
  {32'hbe361c5c, 32'h00000000} /* (8, 2, 12) {real, imag} */,
  {32'hbd2fec20, 32'h00000000} /* (8, 2, 11) {real, imag} */,
  {32'h3f718462, 32'h00000000} /* (8, 2, 10) {real, imag} */,
  {32'h3ef2c6d8, 32'h00000000} /* (8, 2, 9) {real, imag} */,
  {32'hbe646928, 32'h00000000} /* (8, 2, 8) {real, imag} */,
  {32'h3e258b54, 32'h00000000} /* (8, 2, 7) {real, imag} */,
  {32'h3ec911ff, 32'h00000000} /* (8, 2, 6) {real, imag} */,
  {32'hbe372c70, 32'h00000000} /* (8, 2, 5) {real, imag} */,
  {32'h3ed0e11a, 32'h00000000} /* (8, 2, 4) {real, imag} */,
  {32'h3ec9df02, 32'h00000000} /* (8, 2, 3) {real, imag} */,
  {32'h3e9f05b0, 32'h00000000} /* (8, 2, 2) {real, imag} */,
  {32'h3d0b8d60, 32'h00000000} /* (8, 2, 1) {real, imag} */,
  {32'hbd736c94, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'hbef289ec, 32'h00000000} /* (8, 1, 15) {real, imag} */,
  {32'hbea4d654, 32'h00000000} /* (8, 1, 14) {real, imag} */,
  {32'hbee49a80, 32'h00000000} /* (8, 1, 13) {real, imag} */,
  {32'hbefbc0b4, 32'h00000000} /* (8, 1, 12) {real, imag} */,
  {32'hbe6dda78, 32'h00000000} /* (8, 1, 11) {real, imag} */,
  {32'h3eb0ac5e, 32'h00000000} /* (8, 1, 10) {real, imag} */,
  {32'h3f859de0, 32'h00000000} /* (8, 1, 9) {real, imag} */,
  {32'hbdcc7114, 32'h00000000} /* (8, 1, 8) {real, imag} */,
  {32'hbe6bb070, 32'h00000000} /* (8, 1, 7) {real, imag} */,
  {32'hbe1489b2, 32'h00000000} /* (8, 1, 6) {real, imag} */,
  {32'hbe82883f, 32'h00000000} /* (8, 1, 5) {real, imag} */,
  {32'h3e259140, 32'h00000000} /* (8, 1, 4) {real, imag} */,
  {32'h3e8a10f4, 32'h00000000} /* (8, 1, 3) {real, imag} */,
  {32'hbdf90270, 32'h00000000} /* (8, 1, 2) {real, imag} */,
  {32'hbecb6fe0, 32'h00000000} /* (8, 1, 1) {real, imag} */,
  {32'hbe370558, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'hbe257522, 32'h00000000} /* (8, 0, 15) {real, imag} */,
  {32'hbe1fe6b0, 32'h00000000} /* (8, 0, 14) {real, imag} */,
  {32'hbb960000, 32'h00000000} /* (8, 0, 13) {real, imag} */,
  {32'h3ea6c7e2, 32'h00000000} /* (8, 0, 12) {real, imag} */,
  {32'h3e7712a4, 32'h00000000} /* (8, 0, 11) {real, imag} */,
  {32'h3e2581f4, 32'h00000000} /* (8, 0, 10) {real, imag} */,
  {32'h3edfb3fc, 32'h00000000} /* (8, 0, 9) {real, imag} */,
  {32'h3da97b80, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'hbdeb064c, 32'h00000000} /* (8, 0, 7) {real, imag} */,
  {32'hbe3d2bec, 32'h00000000} /* (8, 0, 6) {real, imag} */,
  {32'h3d034670, 32'h00000000} /* (8, 0, 5) {real, imag} */,
  {32'h3d239c20, 32'h00000000} /* (8, 0, 4) {real, imag} */,
  {32'h3e846ea4, 32'h00000000} /* (8, 0, 3) {real, imag} */,
  {32'hbe3c67b0, 32'h00000000} /* (8, 0, 2) {real, imag} */,
  {32'hbf09cf39, 32'h00000000} /* (8, 0, 1) {real, imag} */,
  {32'hbe71f092, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h3c8efd84, 32'h3ea39bc0} /* (7, 15, 15) {real, imag} */,
  {32'h3d22a5b0, 32'h3eb6d5f2} /* (7, 15, 14) {real, imag} */,
  {32'hbe2add17, 32'h3e806b94} /* (7, 15, 13) {real, imag} */,
  {32'h3bead378, 32'h3e03b8ae} /* (7, 15, 12) {real, imag} */,
  {32'hbea6a608, 32'hbd8facea} /* (7, 15, 11) {real, imag} */,
  {32'hbf4669e2, 32'h3e27f44c} /* (7, 15, 10) {real, imag} */,
  {32'hbf20d265, 32'h3e39e414} /* (7, 15, 9) {real, imag} */,
  {32'hbe5cb82c, 32'hbd82c640} /* (7, 15, 8) {real, imag} */,
  {32'h3e9d2270, 32'h3df62a70} /* (7, 15, 7) {real, imag} */,
  {32'h3f0a2c8e, 32'hbd987251} /* (7, 15, 6) {real, imag} */,
  {32'h3f384ba8, 32'hbe3cbfb2} /* (7, 15, 5) {real, imag} */,
  {32'h3ee4c29c, 32'h3dc91890} /* (7, 15, 4) {real, imag} */,
  {32'h3ec6d69a, 32'h3e5d4728} /* (7, 15, 3) {real, imag} */,
  {32'h3e9e0f36, 32'hbbe0f540} /* (7, 15, 2) {real, imag} */,
  {32'hbdedf2d0, 32'h3eed1b31} /* (7, 15, 1) {real, imag} */,
  {32'hbe6567ea, 32'h3eef01a0} /* (7, 15, 0) {real, imag} */,
  {32'h3e88a803, 32'h3bed9480} /* (7, 14, 15) {real, imag} */,
  {32'h3ee98cc0, 32'hbdfc31c0} /* (7, 14, 14) {real, imag} */,
  {32'h3d8c1528, 32'h3e7d3978} /* (7, 14, 13) {real, imag} */,
  {32'hbeb8a6ca, 32'h3e308a60} /* (7, 14, 12) {real, imag} */,
  {32'hbebee42b, 32'hbea67723} /* (7, 14, 11) {real, imag} */,
  {32'hbe9210e3, 32'h3c3e9ec0} /* (7, 14, 10) {real, imag} */,
  {32'hbe1ea812, 32'hbc66a200} /* (7, 14, 9) {real, imag} */,
  {32'hbe18ed00, 32'hbe68a018} /* (7, 14, 8) {real, imag} */,
  {32'h3e5824f8, 32'h3e0f2b2c} /* (7, 14, 7) {real, imag} */,
  {32'h3ed7ebc5, 32'hbcf39720} /* (7, 14, 6) {real, imag} */,
  {32'h3f80a3e6, 32'hbe2e2b85} /* (7, 14, 5) {real, imag} */,
  {32'h3e525ace, 32'hbd8f6398} /* (7, 14, 4) {real, imag} */,
  {32'h3e07eb19, 32'h3e9308fc} /* (7, 14, 3) {real, imag} */,
  {32'h3e6d10df, 32'h3e1488c0} /* (7, 14, 2) {real, imag} */,
  {32'h3e60a7ce, 32'h3e3ecaf0} /* (7, 14, 1) {real, imag} */,
  {32'h3e610c97, 32'h3e93d35e} /* (7, 14, 0) {real, imag} */,
  {32'hbcf95c20, 32'hbee0180c} /* (7, 13, 15) {real, imag} */,
  {32'h3f165b90, 32'hbf26deb2} /* (7, 13, 14) {real, imag} */,
  {32'h3ef454f1, 32'hbe79ff60} /* (7, 13, 13) {real, imag} */,
  {32'hbe851e70, 32'h3d57a650} /* (7, 13, 12) {real, imag} */,
  {32'hbf033260, 32'hbecae558} /* (7, 13, 11) {real, imag} */,
  {32'hbe8f853a, 32'hbe6d81e8} /* (7, 13, 10) {real, imag} */,
  {32'h3e2634a8, 32'hbdb1b720} /* (7, 13, 9) {real, imag} */,
  {32'h3e320717, 32'h3e8a0a4b} /* (7, 13, 8) {real, imag} */,
  {32'h3e4d024e, 32'h3f601281} /* (7, 13, 7) {real, imag} */,
  {32'hbe05fff8, 32'h3d87761a} /* (7, 13, 6) {real, imag} */,
  {32'h3e3dd241, 32'h3d80aa24} /* (7, 13, 5) {real, imag} */,
  {32'h3e1532ca, 32'h3e9aa4b6} /* (7, 13, 4) {real, imag} */,
  {32'hbe389718, 32'hbe77642e} /* (7, 13, 3) {real, imag} */,
  {32'hbd9eec1f, 32'hbe3d2a3c} /* (7, 13, 2) {real, imag} */,
  {32'h3e29cccc, 32'hbd321b60} /* (7, 13, 1) {real, imag} */,
  {32'h3d98c508, 32'hbda62cac} /* (7, 13, 0) {real, imag} */,
  {32'h3d54e6b4, 32'hbea5b470} /* (7, 12, 15) {real, imag} */,
  {32'h3e90c9bc, 32'hbf489c07} /* (7, 12, 14) {real, imag} */,
  {32'h3d99df60, 32'hbdd0f720} /* (7, 12, 13) {real, imag} */,
  {32'hbdf57378, 32'h3ef32d43} /* (7, 12, 12) {real, imag} */,
  {32'hbdd186f8, 32'h3f1838e0} /* (7, 12, 11) {real, imag} */,
  {32'hbe97f8e5, 32'h3f060930} /* (7, 12, 10) {real, imag} */,
  {32'hbf042255, 32'h3ee718ee} /* (7, 12, 9) {real, imag} */,
  {32'hbecbd7f2, 32'h3f1f48a3} /* (7, 12, 8) {real, imag} */,
  {32'h3e0f5ac8, 32'h3ed71fab} /* (7, 12, 7) {real, imag} */,
  {32'hbeb7b0b4, 32'h3e93646a} /* (7, 12, 6) {real, imag} */,
  {32'h3dd56b80, 32'h3f37a100} /* (7, 12, 5) {real, imag} */,
  {32'h3e65cc06, 32'h3f471e47} /* (7, 12, 4) {real, imag} */,
  {32'hbe3de50c, 32'hbd4839e0} /* (7, 12, 3) {real, imag} */,
  {32'hbdc4dba8, 32'hbe9b3364} /* (7, 12, 2) {real, imag} */,
  {32'h3e9d3b2c, 32'h3ede69f6} /* (7, 12, 1) {real, imag} */,
  {32'h3ec62a99, 32'h3dddc160} /* (7, 12, 0) {real, imag} */,
  {32'hbe0b1712, 32'h3ead6e27} /* (7, 11, 15) {real, imag} */,
  {32'hbdf34fdf, 32'h3ed3a2bf} /* (7, 11, 14) {real, imag} */,
  {32'hbe95ec84, 32'h3efb028d} /* (7, 11, 13) {real, imag} */,
  {32'hbef66258, 32'hbe4a202c} /* (7, 11, 12) {real, imag} */,
  {32'h3e21e010, 32'hbf0d776a} /* (7, 11, 11) {real, imag} */,
  {32'hbe792c9f, 32'hbea4a42a} /* (7, 11, 10) {real, imag} */,
  {32'hbf63ad74, 32'hbf162f85} /* (7, 11, 9) {real, imag} */,
  {32'hbf22c8b1, 32'hbefbe1dc} /* (7, 11, 8) {real, imag} */,
  {32'h3d5e3e20, 32'hbdba26b0} /* (7, 11, 7) {real, imag} */,
  {32'hbe1ead48, 32'h3e7075ec} /* (7, 11, 6) {real, imag} */,
  {32'h3e965813, 32'h3f0cb390} /* (7, 11, 5) {real, imag} */,
  {32'h3ed3d11d, 32'h3dc1edf4} /* (7, 11, 4) {real, imag} */,
  {32'h3c5f8580, 32'hbe3065e7} /* (7, 11, 3) {real, imag} */,
  {32'h3ecbf215, 32'h3d97f021} /* (7, 11, 2) {real, imag} */,
  {32'h3eea0b8c, 32'h3f5e7071} /* (7, 11, 1) {real, imag} */,
  {32'h3e8c792c, 32'h3f108028} /* (7, 11, 0) {real, imag} */,
  {32'hbf05c4e6, 32'h3ea0199a} /* (7, 10, 15) {real, imag} */,
  {32'hbcde8610, 32'h3f21490c} /* (7, 10, 14) {real, imag} */,
  {32'hbd8789f7, 32'h3ebee9e2} /* (7, 10, 13) {real, imag} */,
  {32'hbf10e4dc, 32'hbd4d1818} /* (7, 10, 12) {real, imag} */,
  {32'h3c1e7080, 32'hbed807a2} /* (7, 10, 11) {real, imag} */,
  {32'hbe0e1540, 32'hbf3dc871} /* (7, 10, 10) {real, imag} */,
  {32'hbeaceb4a, 32'hbf4ceda7} /* (7, 10, 9) {real, imag} */,
  {32'hbeea7ca9, 32'hbeded186} /* (7, 10, 8) {real, imag} */,
  {32'h3d870bf4, 32'h3e5e12d8} /* (7, 10, 7) {real, imag} */,
  {32'hbdfe5d04, 32'h3ef1f040} /* (7, 10, 6) {real, imag} */,
  {32'h3e4e7a98, 32'h3f215adf} /* (7, 10, 5) {real, imag} */,
  {32'h3ed6dfc4, 32'h3e540b42} /* (7, 10, 4) {real, imag} */,
  {32'hbe8d55c8, 32'h3e899e46} /* (7, 10, 3) {real, imag} */,
  {32'hbe3269e8, 32'h3d602c30} /* (7, 10, 2) {real, imag} */,
  {32'hbcdbc000, 32'h3eb1217c} /* (7, 10, 1) {real, imag} */,
  {32'hbd08eb30, 32'h3ebfb9e6} /* (7, 10, 0) {real, imag} */,
  {32'hbf012a1e, 32'h3e8d35f8} /* (7, 9, 15) {real, imag} */,
  {32'h3d7508fe, 32'h3ea9dac1} /* (7, 9, 14) {real, imag} */,
  {32'hbdb7b9f2, 32'hbdc4f6f4} /* (7, 9, 13) {real, imag} */,
  {32'hbe9bccca, 32'hbdc85640} /* (7, 9, 12) {real, imag} */,
  {32'h3ec7a57d, 32'hbe540898} /* (7, 9, 11) {real, imag} */,
  {32'hbe0a1c20, 32'hbef122a2} /* (7, 9, 10) {real, imag} */,
  {32'hbe7a1808, 32'hbe4d3524} /* (7, 9, 9) {real, imag} */,
  {32'hbe805c2c, 32'h3ee31a88} /* (7, 9, 8) {real, imag} */,
  {32'hbe65fc32, 32'h3f2bdc2c} /* (7, 9, 7) {real, imag} */,
  {32'h3e527e34, 32'h3f13b2ce} /* (7, 9, 6) {real, imag} */,
  {32'h3f0c64e7, 32'h3f4c42c3} /* (7, 9, 5) {real, imag} */,
  {32'h3e7d93da, 32'h3efc917c} /* (7, 9, 4) {real, imag} */,
  {32'h3e750698, 32'h3f1643fd} /* (7, 9, 3) {real, imag} */,
  {32'hbcf45420, 32'h3e88e31f} /* (7, 9, 2) {real, imag} */,
  {32'h3e347bf0, 32'hbd8fdcd8} /* (7, 9, 1) {real, imag} */,
  {32'h3e394ed0, 32'hbe7eba60} /* (7, 9, 0) {real, imag} */,
  {32'hbd0ecdac, 32'h3f04f7de} /* (7, 8, 15) {real, imag} */,
  {32'h3e7a36f4, 32'h3edaa627} /* (7, 8, 14) {real, imag} */,
  {32'hbeb6ea52, 32'hbcdf7330} /* (7, 8, 13) {real, imag} */,
  {32'hbf0e005d, 32'h3eb9f7c6} /* (7, 8, 12) {real, imag} */,
  {32'h3e823e49, 32'h3d884900} /* (7, 8, 11) {real, imag} */,
  {32'h3e76134c, 32'hbf1d48d7} /* (7, 8, 10) {real, imag} */,
  {32'h3e6028a8, 32'hbf0a3b1c} /* (7, 8, 9) {real, imag} */,
  {32'h3defda3c, 32'hbf62795e} /* (7, 8, 8) {real, imag} */,
  {32'h3c1a37c0, 32'hbd7d5f10} /* (7, 8, 7) {real, imag} */,
  {32'h3ea3b3ee, 32'h3e9a72ac} /* (7, 8, 6) {real, imag} */,
  {32'h3edbb2e2, 32'h3ed175dc} /* (7, 8, 5) {real, imag} */,
  {32'h3e89ea94, 32'hbe1250f8} /* (7, 8, 4) {real, imag} */,
  {32'h3f1b4f96, 32'h3dd271c0} /* (7, 8, 3) {real, imag} */,
  {32'h3eccb5ca, 32'h3ea25cee} /* (7, 8, 2) {real, imag} */,
  {32'h3ea2796b, 32'hbdb70630} /* (7, 8, 1) {real, imag} */,
  {32'h3ea5052d, 32'hbe097110} /* (7, 8, 0) {real, imag} */,
  {32'hbd37a648, 32'h3eeeeb6a} /* (7, 7, 15) {real, imag} */,
  {32'hbe44784e, 32'h3eb7a8fa} /* (7, 7, 14) {real, imag} */,
  {32'hbe2d3517, 32'h3d318e00} /* (7, 7, 13) {real, imag} */,
  {32'hbe79f352, 32'h3f68a99f} /* (7, 7, 12) {real, imag} */,
  {32'h3e935d4e, 32'h3ebd3064} /* (7, 7, 11) {real, imag} */,
  {32'h3e8566b7, 32'hbf62bd5b} /* (7, 7, 10) {real, imag} */,
  {32'h3f458dac, 32'hbec573d8} /* (7, 7, 9) {real, imag} */,
  {32'h3eab90e4, 32'hbf095154} /* (7, 7, 8) {real, imag} */,
  {32'hbe9e36b2, 32'h3e19dc81} /* (7, 7, 7) {real, imag} */,
  {32'h3e773ee8, 32'h3e713420} /* (7, 7, 6) {real, imag} */,
  {32'h3eadd7ae, 32'hbedbdd82} /* (7, 7, 5) {real, imag} */,
  {32'hbe41d72c, 32'hbe8d705b} /* (7, 7, 4) {real, imag} */,
  {32'hbe54527c, 32'h3f132e15} /* (7, 7, 3) {real, imag} */,
  {32'hbe50b74c, 32'h3f4e0ede} /* (7, 7, 2) {real, imag} */,
  {32'hbe82bd0e, 32'h3ededd59} /* (7, 7, 1) {real, imag} */,
  {32'hbe8f13e8, 32'h3ea7d038} /* (7, 7, 0) {real, imag} */,
  {32'h3d6731b4, 32'h3ed6ba43} /* (7, 6, 15) {real, imag} */,
  {32'hbd47a900, 32'h3e6871a4} /* (7, 6, 14) {real, imag} */,
  {32'h3e1d8529, 32'h3e65762c} /* (7, 6, 13) {real, imag} */,
  {32'h3def22f0, 32'h3e5a2ec4} /* (7, 6, 12) {real, imag} */,
  {32'h3d20f4b8, 32'hbe8180fa} /* (7, 6, 11) {real, imag} */,
  {32'h3d656040, 32'hbea7ea09} /* (7, 6, 10) {real, imag} */,
  {32'h3f809f4b, 32'h3ea85bec} /* (7, 6, 9) {real, imag} */,
  {32'h3eb1c3c2, 32'h3e857edc} /* (7, 6, 8) {real, imag} */,
  {32'hbe95f7fc, 32'h3f4e0f86} /* (7, 6, 7) {real, imag} */,
  {32'hbdc10500, 32'h3f1edb2c} /* (7, 6, 6) {real, imag} */,
  {32'hbe5df958, 32'hbf480432} /* (7, 6, 5) {real, imag} */,
  {32'hbee17ff4, 32'hbf557004} /* (7, 6, 4) {real, imag} */,
  {32'hbef00b0e, 32'h3eb57280} /* (7, 6, 3) {real, imag} */,
  {32'hbf0a2018, 32'h3fa2437d} /* (7, 6, 2) {real, imag} */,
  {32'h3d9a7348, 32'h3f1511b8} /* (7, 6, 1) {real, imag} */,
  {32'hbdc3a688, 32'h3d6d434c} /* (7, 6, 0) {real, imag} */,
  {32'h3e56bf72, 32'h3e256c00} /* (7, 5, 15) {real, imag} */,
  {32'h3b35da00, 32'hbe7a7440} /* (7, 5, 14) {real, imag} */,
  {32'hbebdb9ca, 32'h3de2d028} /* (7, 5, 13) {real, imag} */,
  {32'hbe40ba02, 32'h3e59f560} /* (7, 5, 12) {real, imag} */,
  {32'h3e5ffa82, 32'hbd5cfd40} /* (7, 5, 11) {real, imag} */,
  {32'h3f0c07bf, 32'h3e2bc6b8} /* (7, 5, 10) {real, imag} */,
  {32'h3f8d5e2a, 32'h3f112b46} /* (7, 5, 9) {real, imag} */,
  {32'h3effd038, 32'h3f43dabe} /* (7, 5, 8) {real, imag} */,
  {32'hbcc50868, 32'h3f0b767a} /* (7, 5, 7) {real, imag} */,
  {32'h3d1ea2a0, 32'h3efadd31} /* (7, 5, 6) {real, imag} */,
  {32'hbde8c900, 32'hbdd27634} /* (7, 5, 5) {real, imag} */,
  {32'hbe0039cc, 32'h3d9d1830} /* (7, 5, 4) {real, imag} */,
  {32'hbe981762, 32'h3edc865c} /* (7, 5, 3) {real, imag} */,
  {32'hbea89648, 32'h3f5df201} /* (7, 5, 2) {real, imag} */,
  {32'h3d8fa060, 32'h3f0d52ec} /* (7, 5, 1) {real, imag} */,
  {32'hbe3e61b4, 32'hbd037696} /* (7, 5, 0) {real, imag} */,
  {32'h3ef1e344, 32'h3e30c8bc} /* (7, 4, 15) {real, imag} */,
  {32'h3deaeb00, 32'hbdae1414} /* (7, 4, 14) {real, imag} */,
  {32'hbe800cd4, 32'h3de9a610} /* (7, 4, 13) {real, imag} */,
  {32'h3dcc570e, 32'h3e23e4f4} /* (7, 4, 12) {real, imag} */,
  {32'h3eeee750, 32'hbe670f98} /* (7, 4, 11) {real, imag} */,
  {32'h3d1f1960, 32'hbe03aaf8} /* (7, 4, 10) {real, imag} */,
  {32'h3f2795a6, 32'h3ef312bb} /* (7, 4, 9) {real, imag} */,
  {32'h3e24ed14, 32'h3e8c9462} /* (7, 4, 8) {real, imag} */,
  {32'hbe89623a, 32'hbe1313e8} /* (7, 4, 7) {real, imag} */,
  {32'h3e5f1c48, 32'hbd4554f8} /* (7, 4, 6) {real, imag} */,
  {32'h3ed07f50, 32'hbf205bd6} /* (7, 4, 5) {real, imag} */,
  {32'h3ae41000, 32'hbe6079ae} /* (7, 4, 4) {real, imag} */,
  {32'hbe9e1122, 32'h3eced884} /* (7, 4, 3) {real, imag} */,
  {32'hbf2bef6c, 32'h3ea5efd4} /* (7, 4, 2) {real, imag} */,
  {32'hbe7d1538, 32'h3e83294e} /* (7, 4, 1) {real, imag} */,
  {32'hbe27e51f, 32'h3e5ea8a0} /* (7, 4, 0) {real, imag} */,
  {32'h3ebfaf5e, 32'hbe43f6f0} /* (7, 3, 15) {real, imag} */,
  {32'h3f2b07e7, 32'hbf15dcca} /* (7, 3, 14) {real, imag} */,
  {32'h3f03774c, 32'h3ccf4418} /* (7, 3, 13) {real, imag} */,
  {32'h3dc5b088, 32'h3e9e7d71} /* (7, 3, 12) {real, imag} */,
  {32'h3e3aafb2, 32'hbe25eb40} /* (7, 3, 11) {real, imag} */,
  {32'hbe40a108, 32'hbf1fbdec} /* (7, 3, 10) {real, imag} */,
  {32'hbdb77fcc, 32'hbc919a30} /* (7, 3, 9) {real, imag} */,
  {32'hbed08b8e, 32'h3e1bd4fc} /* (7, 3, 8) {real, imag} */,
  {32'hbec6879b, 32'hbe787994} /* (7, 3, 7) {real, imag} */,
  {32'hbe7676d8, 32'hbf244b40} /* (7, 3, 6) {real, imag} */,
  {32'h3eb6d324, 32'hbf27e752} /* (7, 3, 5) {real, imag} */,
  {32'hbdb286f4, 32'hbdf737e0} /* (7, 3, 4) {real, imag} */,
  {32'hbe48c0b2, 32'h3ef83b24} /* (7, 3, 3) {real, imag} */,
  {32'hbed570e5, 32'h3ee0871c} /* (7, 3, 2) {real, imag} */,
  {32'hbd81d83c, 32'hbe578326} /* (7, 3, 1) {real, imag} */,
  {32'hbd703440, 32'h3dd028ac} /* (7, 3, 0) {real, imag} */,
  {32'h3f156b11, 32'h3e53bb70} /* (7, 2, 15) {real, imag} */,
  {32'h3f5c4b12, 32'h3e2ea738} /* (7, 2, 14) {real, imag} */,
  {32'h3f1d5cc4, 32'h3d6de89c} /* (7, 2, 13) {real, imag} */,
  {32'h3e9e8102, 32'h3e71e741} /* (7, 2, 12) {real, imag} */,
  {32'h3e4f29ea, 32'hbd5bf4e6} /* (7, 2, 11) {real, imag} */,
  {32'h3ea97f2e, 32'hbf34e53e} /* (7, 2, 10) {real, imag} */,
  {32'hbea207ca, 32'hbf039817} /* (7, 2, 9) {real, imag} */,
  {32'hbeac40ba, 32'hbe8f2666} /* (7, 2, 8) {real, imag} */,
  {32'hbe8aba83, 32'hbd87859e} /* (7, 2, 7) {real, imag} */,
  {32'hbf127b7e, 32'hbe807172} /* (7, 2, 6) {real, imag} */,
  {32'hbdbd9a50, 32'hbf0037ac} /* (7, 2, 5) {real, imag} */,
  {32'h3d9b8df8, 32'hbe460722} /* (7, 2, 4) {real, imag} */,
  {32'hbe7850ab, 32'h3e1dd656} /* (7, 2, 3) {real, imag} */,
  {32'hbecb2519, 32'h3d9de694} /* (7, 2, 2) {real, imag} */,
  {32'h3e7ec742, 32'h3eb2a966} /* (7, 2, 1) {real, imag} */,
  {32'h3d4e1570, 32'h3e8259b3} /* (7, 2, 0) {real, imag} */,
  {32'h3e7208b3, 32'h3ec5bbf8} /* (7, 1, 15) {real, imag} */,
  {32'h3edb4f13, 32'h3f17f633} /* (7, 1, 14) {real, imag} */,
  {32'h3d8096f0, 32'h3e1f9b8c} /* (7, 1, 13) {real, imag} */,
  {32'h3d714430, 32'hbf0e871f} /* (7, 1, 12) {real, imag} */,
  {32'h3ed5b19e, 32'hbf74bae9} /* (7, 1, 11) {real, imag} */,
  {32'h3edbe3cf, 32'hbeec6761} /* (7, 1, 10) {real, imag} */,
  {32'hbddbba20, 32'h3e20cc1a} /* (7, 1, 9) {real, imag} */,
  {32'hbebdc5c0, 32'hbdc00bd8} /* (7, 1, 8) {real, imag} */,
  {32'h3e78010c, 32'h3e85c2a6} /* (7, 1, 7) {real, imag} */,
  {32'hbe0c5860, 32'h3e5d0368} /* (7, 1, 6) {real, imag} */,
  {32'hbf18e598, 32'h3eb99aec} /* (7, 1, 5) {real, imag} */,
  {32'h3dd41ee0, 32'h3ee584ab} /* (7, 1, 4) {real, imag} */,
  {32'hb9fb7000, 32'h3d2d13a4} /* (7, 1, 3) {real, imag} */,
  {32'hbf1f6bf0, 32'hbebfacb8} /* (7, 1, 2) {real, imag} */,
  {32'hbecb745f, 32'hbc59b600} /* (7, 1, 1) {real, imag} */,
  {32'h3d62d74c, 32'hbc1ffe60} /* (7, 1, 0) {real, imag} */,
  {32'hbde4896e, 32'h3e0b1aac} /* (7, 0, 15) {real, imag} */,
  {32'hbec67eba, 32'hbd89f760} /* (7, 0, 14) {real, imag} */,
  {32'hbf06b304, 32'hbe94ea02} /* (7, 0, 13) {real, imag} */,
  {32'h3cbb1a40, 32'hbf0f5f0d} /* (7, 0, 12) {real, imag} */,
  {32'h3e396d7e, 32'hbf5814ca} /* (7, 0, 11) {real, imag} */,
  {32'hbdfd8f50, 32'h3ba1ec20} /* (7, 0, 10) {real, imag} */,
  {32'hbe5489cc, 32'h3ee679c0} /* (7, 0, 9) {real, imag} */,
  {32'hbda9cd2e, 32'h3dd5e89e} /* (7, 0, 8) {real, imag} */,
  {32'h3e0b46ca, 32'h3f14cff2} /* (7, 0, 7) {real, imag} */,
  {32'hbd2fd36a, 32'h3edbe637} /* (7, 0, 6) {real, imag} */,
  {32'hbed3ab06, 32'h3e9c015e} /* (7, 0, 5) {real, imag} */,
  {32'h3d1511a0, 32'h3e4dd2a7} /* (7, 0, 4) {real, imag} */,
  {32'h3eecd7d0, 32'h3d0315a8} /* (7, 0, 3) {real, imag} */,
  {32'h3eb77dd5, 32'hbe584dbd} /* (7, 0, 2) {real, imag} */,
  {32'hbda33cac, 32'hbe55f2b5} /* (7, 0, 1) {real, imag} */,
  {32'h3d14e870, 32'hbdb974c0} /* (7, 0, 0) {real, imag} */,
  {32'hbd8a394c, 32'hbeb1ca6c} /* (6, 15, 15) {real, imag} */,
  {32'hbe096ee4, 32'h3d5a8660} /* (6, 15, 14) {real, imag} */,
  {32'hbd419aea, 32'h3d9a23b4} /* (6, 15, 13) {real, imag} */,
  {32'h3cbf075c, 32'hbebf86df} /* (6, 15, 12) {real, imag} */,
  {32'h3e164cee, 32'hbeb8f0f3} /* (6, 15, 11) {real, imag} */,
  {32'hbdca9218, 32'hbe055404} /* (6, 15, 10) {real, imag} */,
  {32'hbdb1a19a, 32'h3d134b10} /* (6, 15, 9) {real, imag} */,
  {32'hbc238f30, 32'hbd48443c} /* (6, 15, 8) {real, imag} */,
  {32'hbe9880a7, 32'h3f0c78c0} /* (6, 15, 7) {real, imag} */,
  {32'hbef90b1b, 32'h3d495238} /* (6, 15, 6) {real, imag} */,
  {32'h3e2b3a6c, 32'hbe8b982c} /* (6, 15, 5) {real, imag} */,
  {32'h3ec13388, 32'hbdedf330} /* (6, 15, 4) {real, imag} */,
  {32'h3d789b20, 32'hbf22b5aa} /* (6, 15, 3) {real, imag} */,
  {32'hbe09b7b1, 32'hbeb444b9} /* (6, 15, 2) {real, imag} */,
  {32'h3e9376ea, 32'h3f169403} /* (6, 15, 1) {real, imag} */,
  {32'h3efd7706, 32'h3ed594d8} /* (6, 15, 0) {real, imag} */,
  {32'h3f155438, 32'h3e8f6552} /* (6, 14, 15) {real, imag} */,
  {32'h3ec828f6, 32'h3f0c504e} /* (6, 14, 14) {real, imag} */,
  {32'hbe7b6f7c, 32'hbe801038} /* (6, 14, 13) {real, imag} */,
  {32'h3e013644, 32'hbf2f0036} /* (6, 14, 12) {real, imag} */,
  {32'h3f83bd76, 32'hbf7f4fd8} /* (6, 14, 11) {real, imag} */,
  {32'h3f333444, 32'hbf9e15ac} /* (6, 14, 10) {real, imag} */,
  {32'h3e2be418, 32'hbf950972} /* (6, 14, 9) {real, imag} */,
  {32'h3bd4b2c0, 32'hbead848e} /* (6, 14, 8) {real, imag} */,
  {32'hbeecedb7, 32'h3e1b2784} /* (6, 14, 7) {real, imag} */,
  {32'hbf56f19e, 32'hbe433590} /* (6, 14, 6) {real, imag} */,
  {32'hbe2b923c, 32'hbf236308} /* (6, 14, 5) {real, imag} */,
  {32'hbdbe8590, 32'hbf460408} /* (6, 14, 4) {real, imag} */,
  {32'h3d706a40, 32'hbf1eac76} /* (6, 14, 3) {real, imag} */,
  {32'hbebf7a96, 32'hbec41b3a} /* (6, 14, 2) {real, imag} */,
  {32'hbf026bc7, 32'h3ed24128} /* (6, 14, 1) {real, imag} */,
  {32'h3f10d654, 32'h3f05ca12} /* (6, 14, 0) {real, imag} */,
  {32'h3dbbf0e6, 32'h3f088342} /* (6, 13, 15) {real, imag} */,
  {32'h3d914ac2, 32'h3df3ac70} /* (6, 13, 14) {real, imag} */,
  {32'hbc72fc30, 32'hbe831030} /* (6, 13, 13) {real, imag} */,
  {32'h3dae3468, 32'hbd857820} /* (6, 13, 12) {real, imag} */,
  {32'h3f1f1ac7, 32'hbdc3aa88} /* (6, 13, 11) {real, imag} */,
  {32'h3eff951a, 32'hbf790e61} /* (6, 13, 10) {real, imag} */,
  {32'h3e97e0c2, 32'hbf7b1e3e} /* (6, 13, 9) {real, imag} */,
  {32'hbed9eb6d, 32'hbe331708} /* (6, 13, 8) {real, imag} */,
  {32'hbea3891c, 32'h3e17a168} /* (6, 13, 7) {real, imag} */,
  {32'hbf606a08, 32'h3f06a486} /* (6, 13, 6) {real, imag} */,
  {32'hbf4555ec, 32'hbeb21a40} /* (6, 13, 5) {real, imag} */,
  {32'hbebddd1a, 32'hbf48f523} /* (6, 13, 4) {real, imag} */,
  {32'hbce9e580, 32'hbe46f5fc} /* (6, 13, 3) {real, imag} */,
  {32'h3e79b419, 32'hbe558cd2} /* (6, 13, 2) {real, imag} */,
  {32'hbea2070e, 32'hbe55cdba} /* (6, 13, 1) {real, imag} */,
  {32'hbe72e650, 32'h3b48ae00} /* (6, 13, 0) {real, imag} */,
  {32'hbe409656, 32'h3dd578bc} /* (6, 12, 15) {real, imag} */,
  {32'hbe995ac8, 32'h3ea52186} /* (6, 12, 14) {real, imag} */,
  {32'h3e44834e, 32'hbe56b58a} /* (6, 12, 13) {real, imag} */,
  {32'h3e1b487e, 32'hbf4ee555} /* (6, 12, 12) {real, imag} */,
  {32'h3f223a30, 32'hbf457c21} /* (6, 12, 11) {real, imag} */,
  {32'h3d3f6c3b, 32'hbf41a21f} /* (6, 12, 10) {real, imag} */,
  {32'hbf37d116, 32'h3f29ab1a} /* (6, 12, 9) {real, imag} */,
  {32'hbf431820, 32'h3f33cc05} /* (6, 12, 8) {real, imag} */,
  {32'h3dea578c, 32'h3f6c287c} /* (6, 12, 7) {real, imag} */,
  {32'hbeff9af4, 32'h3f459bba} /* (6, 12, 6) {real, imag} */,
  {32'hbfa49f76, 32'h3ebcae94} /* (6, 12, 5) {real, imag} */,
  {32'hbe3f8de1, 32'hbed05444} /* (6, 12, 4) {real, imag} */,
  {32'h3f06a987, 32'hbf43c7a4} /* (6, 12, 3) {real, imag} */,
  {32'h3f1ee982, 32'hbee6a2b2} /* (6, 12, 2) {real, imag} */,
  {32'h3d9cb558, 32'hbf496956} /* (6, 12, 1) {real, imag} */,
  {32'hbe604e20, 32'hbf1f1378} /* (6, 12, 0) {real, imag} */,
  {32'hbe855a9c, 32'hbf2e274f} /* (6, 11, 15) {real, imag} */,
  {32'hbf676ea6, 32'hbf2c59e7} /* (6, 11, 14) {real, imag} */,
  {32'hbf90362e, 32'hbf15cd4e} /* (6, 11, 13) {real, imag} */,
  {32'hbf4be93e, 32'hbee2744a} /* (6, 11, 12) {real, imag} */,
  {32'h3f204c10, 32'hbe8f955e} /* (6, 11, 11) {real, imag} */,
  {32'hbe264bb0, 32'hbe8fd492} /* (6, 11, 10) {real, imag} */,
  {32'hbecdb8d4, 32'h3e9cdd30} /* (6, 11, 9) {real, imag} */,
  {32'hbeb17b32, 32'h3e8720e8} /* (6, 11, 8) {real, imag} */,
  {32'hbf2f303e, 32'h3ee60bdd} /* (6, 11, 7) {real, imag} */,
  {32'hbf908a83, 32'hbd766540} /* (6, 11, 6) {real, imag} */,
  {32'hbfa2b971, 32'hbeb4b5fa} /* (6, 11, 5) {real, imag} */,
  {32'hbdbe2582, 32'hbf6b5127} /* (6, 11, 4) {real, imag} */,
  {32'h3ec1c05b, 32'hbf65a4c6} /* (6, 11, 3) {real, imag} */,
  {32'hbe937903, 32'hbf07b920} /* (6, 11, 2) {real, imag} */,
  {32'hbdb08615, 32'hbfaca8cd} /* (6, 11, 1) {real, imag} */,
  {32'hbcb54a10, 32'hbf45fa5a} /* (6, 11, 0) {real, imag} */,
  {32'hbeadd685, 32'hbec14d37} /* (6, 10, 15) {real, imag} */,
  {32'hbf870298, 32'hbe8a1662} /* (6, 10, 14) {real, imag} */,
  {32'hbf81411c, 32'h3ecebdb6} /* (6, 10, 13) {real, imag} */,
  {32'hbf0a8369, 32'h3d9dfb40} /* (6, 10, 12) {real, imag} */,
  {32'hbdfcaaa0, 32'hbc2799a2} /* (6, 10, 11) {real, imag} */,
  {32'hbee26148, 32'h3db8c42c} /* (6, 10, 10) {real, imag} */,
  {32'hbde4b1c0, 32'hbf2fb5ec} /* (6, 10, 9) {real, imag} */,
  {32'hbeda32e8, 32'hbf87de9c} /* (6, 10, 8) {real, imag} */,
  {32'hbeb6a0b8, 32'hbf014118} /* (6, 10, 7) {real, imag} */,
  {32'h3d0390d8, 32'h3f02d790} /* (6, 10, 6) {real, imag} */,
  {32'h3e89f70d, 32'h3ebff4b8} /* (6, 10, 5) {real, imag} */,
  {32'h3f099682, 32'hbf430752} /* (6, 10, 4) {real, imag} */,
  {32'h3ee41e8d, 32'hbf69b389} /* (6, 10, 3) {real, imag} */,
  {32'h3cdca9c0, 32'h3e117eec} /* (6, 10, 2) {real, imag} */,
  {32'h3ee51178, 32'hbf0420ef} /* (6, 10, 1) {real, imag} */,
  {32'h3e80fb44, 32'hbe8e24de} /* (6, 10, 0) {real, imag} */,
  {32'h3eb257bd, 32'hbcce5778} /* (6, 9, 15) {real, imag} */,
  {32'h3f00c747, 32'h3f99ed0e} /* (6, 9, 14) {real, imag} */,
  {32'hbdb94bfc, 32'h3fdde7e6} /* (6, 9, 13) {real, imag} */,
  {32'hbc5f38e8, 32'hbd162ce0} /* (6, 9, 12) {real, imag} */,
  {32'h3da26b52, 32'hbf01506c} /* (6, 9, 11) {real, imag} */,
  {32'h3eda02ea, 32'h3eb242ff} /* (6, 9, 10) {real, imag} */,
  {32'h3e4dd97c, 32'h3dcc8608} /* (6, 9, 9) {real, imag} */,
  {32'hbd154650, 32'hbf5ff4c8} /* (6, 9, 8) {real, imag} */,
  {32'hbd1b9990, 32'hbf437f38} /* (6, 9, 7) {real, imag} */,
  {32'h3f2c1992, 32'hbeec002f} /* (6, 9, 6) {real, imag} */,
  {32'h3f47a1c3, 32'hbe64588e} /* (6, 9, 5) {real, imag} */,
  {32'h3f79eb66, 32'hbf05d7fe} /* (6, 9, 4) {real, imag} */,
  {32'h3e1d0a7c, 32'hbe05efc0} /* (6, 9, 3) {real, imag} */,
  {32'hbe80db6e, 32'h3f056e42} /* (6, 9, 2) {real, imag} */,
  {32'hbe88c765, 32'hbe15c2e0} /* (6, 9, 1) {real, imag} */,
  {32'hbea846ac, 32'hbee64f11} /* (6, 9, 0) {real, imag} */,
  {32'h3e21f7f4, 32'h3e537c04} /* (6, 8, 15) {real, imag} */,
  {32'h3f058766, 32'h3fa5888d} /* (6, 8, 14) {real, imag} */,
  {32'h3c35ee20, 32'h3fce3314} /* (6, 8, 13) {real, imag} */,
  {32'h3df3d0d0, 32'h3f0ebf30} /* (6, 8, 12) {real, imag} */,
  {32'h3f0ad56f, 32'h3e4d5bf6} /* (6, 8, 11) {real, imag} */,
  {32'h3ea91636, 32'h3e895c24} /* (6, 8, 10) {real, imag} */,
  {32'hbdf8c9d0, 32'h3f1761cd} /* (6, 8, 9) {real, imag} */,
  {32'h3ef84ec8, 32'h3efaee0c} /* (6, 8, 8) {real, imag} */,
  {32'hbdd2cb80, 32'h3ece19d2} /* (6, 8, 7) {real, imag} */,
  {32'hbd581f3b, 32'hbf23c0bb} /* (6, 8, 6) {real, imag} */,
  {32'h3ea4a0f0, 32'hbf47ab4a} /* (6, 8, 5) {real, imag} */,
  {32'h3eb66c1a, 32'h3d5afe92} /* (6, 8, 4) {real, imag} */,
  {32'hbf007c1a, 32'h3e8dbfce} /* (6, 8, 3) {real, imag} */,
  {32'hbed4d6e4, 32'h3edaefed} /* (6, 8, 2) {real, imag} */,
  {32'hbea62773, 32'hbe53e5ad} /* (6, 8, 1) {real, imag} */,
  {32'hbedb1e68, 32'hbf1a6756} /* (6, 8, 0) {real, imag} */,
  {32'h3f2591de, 32'h3ed6b084} /* (6, 7, 15) {real, imag} */,
  {32'h3f0194f1, 32'h3f94b87b} /* (6, 7, 14) {real, imag} */,
  {32'hbed3909c, 32'h3fc7d07f} /* (6, 7, 13) {real, imag} */,
  {32'h3e83856c, 32'h3f741305} /* (6, 7, 12) {real, imag} */,
  {32'h3f3168dc, 32'h3e7faf8a} /* (6, 7, 11) {real, imag} */,
  {32'h3f769ea4, 32'h3d2462a0} /* (6, 7, 10) {real, imag} */,
  {32'h3ebc104e, 32'hbc30df80} /* (6, 7, 9) {real, imag} */,
  {32'h3edfc934, 32'h3f3925a2} /* (6, 7, 8) {real, imag} */,
  {32'hbd6d0c8a, 32'h3f0c8dba} /* (6, 7, 7) {real, imag} */,
  {32'h3e02a7dc, 32'h3d53a0e0} /* (6, 7, 6) {real, imag} */,
  {32'hbdf0cfc6, 32'h3ecc8812} /* (6, 7, 5) {real, imag} */,
  {32'hbcee41d0, 32'h3f6f50e6} /* (6, 7, 4) {real, imag} */,
  {32'h3dac7f92, 32'h3e9f465c} /* (6, 7, 3) {real, imag} */,
  {32'h3d2a61fa, 32'hbd8608cc} /* (6, 7, 2) {real, imag} */,
  {32'h3f080cc2, 32'hbf438cc4} /* (6, 7, 1) {real, imag} */,
  {32'hbe31dcfc, 32'hbf3f1874} /* (6, 7, 0) {real, imag} */,
  {32'h3f333d3d, 32'h3d314420} /* (6, 6, 15) {real, imag} */,
  {32'h3ef5a4f6, 32'h3e767c23} /* (6, 6, 14) {real, imag} */,
  {32'h3dc3e5e4, 32'h3ea626e8} /* (6, 6, 13) {real, imag} */,
  {32'h3f0ba7c8, 32'h3ed6817c} /* (6, 6, 12) {real, imag} */,
  {32'h3ee9a0f5, 32'hbf4a8849} /* (6, 6, 11) {real, imag} */,
  {32'h3f25de52, 32'hbe47e190} /* (6, 6, 10) {real, imag} */,
  {32'hbe1c3d4c, 32'hbe206125} /* (6, 6, 9) {real, imag} */,
  {32'hbdd74e10, 32'h3e987244} /* (6, 6, 8) {real, imag} */,
  {32'hbce31180, 32'hbea688fa} /* (6, 6, 7) {real, imag} */,
  {32'hbe836951, 32'hbdf83dc4} /* (6, 6, 6) {real, imag} */,
  {32'hbee56eec, 32'h3f8c2494} /* (6, 6, 5) {real, imag} */,
  {32'hbf8f8499, 32'h3f62ccc9} /* (6, 6, 4) {real, imag} */,
  {32'hbc8378c0, 32'hbe9d9684} /* (6, 6, 3) {real, imag} */,
  {32'h3ef4f9ec, 32'hbefd3036} /* (6, 6, 2) {real, imag} */,
  {32'h3f013ec8, 32'hbf603d6f} /* (6, 6, 1) {real, imag} */,
  {32'h3c203d40, 32'hbf057077} /* (6, 6, 0) {real, imag} */,
  {32'h3e81df41, 32'hbcbd60b8} /* (6, 5, 15) {real, imag} */,
  {32'h3f0a5cb4, 32'hbd5a6470} /* (6, 5, 14) {real, imag} */,
  {32'h3e57ff02, 32'h3d3ce408} /* (6, 5, 13) {real, imag} */,
  {32'hbeb8f2e0, 32'h3e0cabcc} /* (6, 5, 12) {real, imag} */,
  {32'hbe84f456, 32'hbe596733} /* (6, 5, 11) {real, imag} */,
  {32'h3eb0a160, 32'hbeb2d20b} /* (6, 5, 10) {real, imag} */,
  {32'h3e5c2640, 32'hbe5ba563} /* (6, 5, 9) {real, imag} */,
  {32'h3edb2398, 32'hbde7fc73} /* (6, 5, 8) {real, imag} */,
  {32'h3df848f8, 32'hbf42f990} /* (6, 5, 7) {real, imag} */,
  {32'hbf2c1254, 32'hbef2f441} /* (6, 5, 6) {real, imag} */,
  {32'hbf3ad2cb, 32'h3f4a9db6} /* (6, 5, 5) {real, imag} */,
  {32'hbee8f5ec, 32'h3ea746c5} /* (6, 5, 4) {real, imag} */,
  {32'hbd287eb0, 32'hbf0568f7} /* (6, 5, 3) {real, imag} */,
  {32'hbd346d00, 32'hbf0d9b10} /* (6, 5, 2) {real, imag} */,
  {32'hbe45cc34, 32'hbf339c3d} /* (6, 5, 1) {real, imag} */,
  {32'hbd0d22e8, 32'hbf08ecef} /* (6, 5, 0) {real, imag} */,
  {32'h3f532283, 32'h3eac336a} /* (6, 4, 15) {real, imag} */,
  {32'h3f90ccfc, 32'h3e03a9cc} /* (6, 4, 14) {real, imag} */,
  {32'hbc2b4e00, 32'h3e43e7ed} /* (6, 4, 13) {real, imag} */,
  {32'hbf887206, 32'hbe9231f6} /* (6, 4, 12) {real, imag} */,
  {32'hbf58eae0, 32'h3c06f1ae} /* (6, 4, 11) {real, imag} */,
  {32'h3e5c44ea, 32'h3edf7f74} /* (6, 4, 10) {real, imag} */,
  {32'h3eb2c8bd, 32'h3f43cf90} /* (6, 4, 9) {real, imag} */,
  {32'h3f89d356, 32'h3edff993} /* (6, 4, 8) {real, imag} */,
  {32'h3f3318af, 32'hbe55f5fb} /* (6, 4, 7) {real, imag} */,
  {32'hbf347944, 32'h3f011746} /* (6, 4, 6) {real, imag} */,
  {32'hbf6a7355, 32'h3f5f1ae0} /* (6, 4, 5) {real, imag} */,
  {32'hbf3e55e2, 32'h3a746bf2} /* (6, 4, 4) {real, imag} */,
  {32'h3dd30700, 32'h3e905b32} /* (6, 4, 3) {real, imag} */,
  {32'hbcd947ec, 32'h3d49c1f0} /* (6, 4, 2) {real, imag} */,
  {32'hbd6f60b6, 32'h3ccf9990} /* (6, 4, 1) {real, imag} */,
  {32'hbe07d8fc, 32'hbd77bdd0} /* (6, 4, 0) {real, imag} */,
  {32'h3e705d40, 32'hbec7c866} /* (6, 3, 15) {real, imag} */,
  {32'hbe88dd54, 32'hbe667b50} /* (6, 3, 14) {real, imag} */,
  {32'hbe94a386, 32'h3f83c306} /* (6, 3, 13) {real, imag} */,
  {32'hbf0140d3, 32'h3ea00808} /* (6, 3, 12) {real, imag} */,
  {32'hbe7e6fb6, 32'hbdcbe610} /* (6, 3, 11) {real, imag} */,
  {32'hbf1fa61e, 32'h3f5d13ca} /* (6, 3, 10) {real, imag} */,
  {32'hbf182518, 32'h3ec89198} /* (6, 3, 9) {real, imag} */,
  {32'h3f1a9232, 32'h3f6f21aa} /* (6, 3, 8) {real, imag} */,
  {32'h3f0c8b86, 32'h3f442eb0} /* (6, 3, 7) {real, imag} */,
  {32'hbeb0abf5, 32'h3f8608a0} /* (6, 3, 6) {real, imag} */,
  {32'h3e4f1285, 32'h3fb5e374} /* (6, 3, 5) {real, imag} */,
  {32'hbd8b3520, 32'h3f891da2} /* (6, 3, 4) {real, imag} */,
  {32'h3f5c929d, 32'h3f379da6} /* (6, 3, 3) {real, imag} */,
  {32'h3f77706c, 32'hbe3f89be} /* (6, 3, 2) {real, imag} */,
  {32'h3e14d461, 32'hbe481f9c} /* (6, 3, 1) {real, imag} */,
  {32'hbed0d515, 32'hbd764510} /* (6, 3, 0) {real, imag} */,
  {32'hbdc78f00, 32'h3b822400} /* (6, 2, 15) {real, imag} */,
  {32'hbe5226c6, 32'h3cca1700} /* (6, 2, 14) {real, imag} */,
  {32'hbea4a17c, 32'h3f4899ca} /* (6, 2, 13) {real, imag} */,
  {32'hbf21205a, 32'h3f2d59ca} /* (6, 2, 12) {real, imag} */,
  {32'hbd87c5fb, 32'hbdd75e80} /* (6, 2, 11) {real, imag} */,
  {32'hbeebdecc, 32'hbf33aef3} /* (6, 2, 10) {real, imag} */,
  {32'h3eaef8cc, 32'h3c599f30} /* (6, 2, 9) {real, imag} */,
  {32'h3e5a5b64, 32'h3f342300} /* (6, 2, 8) {real, imag} */,
  {32'hbc053e05, 32'h3f5e4c0e} /* (6, 2, 7) {real, imag} */,
  {32'h3ec7a393, 32'h3f360808} /* (6, 2, 6) {real, imag} */,
  {32'h3f61eeeb, 32'h3fe4e93c} /* (6, 2, 5) {real, imag} */,
  {32'h3f4edf1c, 32'h3f971c3b} /* (6, 2, 4) {real, imag} */,
  {32'h3f1b5ab3, 32'h3ee49f2a} /* (6, 2, 3) {real, imag} */,
  {32'h3f1b7cac, 32'hbd8ab958} /* (6, 2, 2) {real, imag} */,
  {32'hbe82d947, 32'hbe0793c0} /* (6, 2, 1) {real, imag} */,
  {32'hbf0527f2, 32'hbbcf52c0} /* (6, 2, 0) {real, imag} */,
  {32'hbe175f62, 32'h3ea1ca07} /* (6, 1, 15) {real, imag} */,
  {32'h3eb74810, 32'hbe1d749c} /* (6, 1, 14) {real, imag} */,
  {32'h3f191f84, 32'hbe4d9f2c} /* (6, 1, 13) {real, imag} */,
  {32'h3e5d883e, 32'h3e34ffc2} /* (6, 1, 12) {real, imag} */,
  {32'hbf63fc88, 32'h3f1c1c08} /* (6, 1, 11) {real, imag} */,
  {32'hbf03b2f0, 32'h3ed6f307} /* (6, 1, 10) {real, imag} */,
  {32'h3f4dd31a, 32'h3d888180} /* (6, 1, 9) {real, imag} */,
  {32'hbe363aca, 32'hbf2a6c3f} /* (6, 1, 8) {real, imag} */,
  {32'hbf02ba92, 32'h3efcff78} /* (6, 1, 7) {real, imag} */,
  {32'h3f0e45a2, 32'h3f68fa60} /* (6, 1, 6) {real, imag} */,
  {32'h3f3b0b5e, 32'h3ee958bc} /* (6, 1, 5) {real, imag} */,
  {32'hbe308598, 32'hbe741144} /* (6, 1, 4) {real, imag} */,
  {32'hbe93506c, 32'hbf01d555} /* (6, 1, 3) {real, imag} */,
  {32'h3f20eb49, 32'hbe84b156} /* (6, 1, 2) {real, imag} */,
  {32'h3e681996, 32'h3ece46d4} /* (6, 1, 1) {real, imag} */,
  {32'hbe866f92, 32'h3f012db5} /* (6, 1, 0) {real, imag} */,
  {32'hbef8877a, 32'h3c8b6502} /* (6, 0, 15) {real, imag} */,
  {32'h3e20a5e2, 32'hbebc0d3a} /* (6, 0, 14) {real, imag} */,
  {32'h3f8f7940, 32'hbe844fa8} /* (6, 0, 13) {real, imag} */,
  {32'h3f2b539c, 32'h3ddf4a0c} /* (6, 0, 12) {real, imag} */,
  {32'hbeab76af, 32'h3f1e7a28} /* (6, 0, 11) {real, imag} */,
  {32'hbed55b5c, 32'h3f2aa1e0} /* (6, 0, 10) {real, imag} */,
  {32'hbdb8761e, 32'h3efb9c08} /* (6, 0, 9) {real, imag} */,
  {32'h3d94e684, 32'hbd697270} /* (6, 0, 8) {real, imag} */,
  {32'hbdecf55c, 32'h3f37d952} /* (6, 0, 7) {real, imag} */,
  {32'hbdfb8b08, 32'h3f46134b} /* (6, 0, 6) {real, imag} */,
  {32'h3ea7e885, 32'hbe0811c0} /* (6, 0, 5) {real, imag} */,
  {32'h3e54faea, 32'hbe88df10} /* (6, 0, 4) {real, imag} */,
  {32'h3e2de110, 32'h3e4a959d} /* (6, 0, 3) {real, imag} */,
  {32'h3f16816a, 32'hbe14d302} /* (6, 0, 2) {real, imag} */,
  {32'h3ea6d938, 32'h3e7f8dce} /* (6, 0, 1) {real, imag} */,
  {32'hbd2e9ed8, 32'h3ee3e2a0} /* (6, 0, 0) {real, imag} */,
  {32'h3f1ad7cf, 32'hbf03733c} /* (5, 15, 15) {real, imag} */,
  {32'h3e9ca1ca, 32'hbe5add77} /* (5, 15, 14) {real, imag} */,
  {32'hbe460084, 32'hbef8a35c} /* (5, 15, 13) {real, imag} */,
  {32'h3d92bc88, 32'h3e1acc20} /* (5, 15, 12) {real, imag} */,
  {32'h3cd89ea0, 32'hbe6ac53b} /* (5, 15, 11) {real, imag} */,
  {32'hbf6d9033, 32'h3af57700} /* (5, 15, 10) {real, imag} */,
  {32'hbf542e51, 32'h3f65f925} /* (5, 15, 9) {real, imag} */,
  {32'h3f39f5b1, 32'h3f282775} /* (5, 15, 8) {real, imag} */,
  {32'h3f4926fe, 32'hbdf15f44} /* (5, 15, 7) {real, imag} */,
  {32'h3e817e47, 32'hbf7831ce} /* (5, 15, 6) {real, imag} */,
  {32'h3eabe9fc, 32'hbf7d2f62} /* (5, 15, 5) {real, imag} */,
  {32'hbf4bd8d7, 32'h3c26e360} /* (5, 15, 4) {real, imag} */,
  {32'h3deebb64, 32'h3f347506} /* (5, 15, 3) {real, imag} */,
  {32'h3fa7614e, 32'h3f01f1fc} /* (5, 15, 2) {real, imag} */,
  {32'h3f71bd23, 32'hbe293a44} /* (5, 15, 1) {real, imag} */,
  {32'h3f3157e2, 32'hbec21936} /* (5, 15, 0) {real, imag} */,
  {32'h3f00b2e8, 32'hbeb9620a} /* (5, 14, 15) {real, imag} */,
  {32'h3d8b70e8, 32'hbe14aff8} /* (5, 14, 14) {real, imag} */,
  {32'h3d87af4c, 32'hbe63dfd8} /* (5, 14, 13) {real, imag} */,
  {32'h3f841a36, 32'h3e70f9a8} /* (5, 14, 12) {real, imag} */,
  {32'h3ef15731, 32'hbf210817} /* (5, 14, 11) {real, imag} */,
  {32'hbf955cfe, 32'hbdad8b98} /* (5, 14, 10) {real, imag} */,
  {32'hbf991b7b, 32'h3fad62c4} /* (5, 14, 9) {real, imag} */,
  {32'h3eb023ef, 32'h3f57972a} /* (5, 14, 8) {real, imag} */,
  {32'hbcdb0190, 32'hbebd3efe} /* (5, 14, 7) {real, imag} */,
  {32'h3d449e50, 32'hbf825386} /* (5, 14, 6) {real, imag} */,
  {32'h3f15f17a, 32'hbed9ebaa} /* (5, 14, 5) {real, imag} */,
  {32'hbe48e7b0, 32'hbd9f8b88} /* (5, 14, 4) {real, imag} */,
  {32'hbe9d83db, 32'h3e1b8114} /* (5, 14, 3) {real, imag} */,
  {32'h3f253486, 32'h3eba4d68} /* (5, 14, 2) {real, imag} */,
  {32'h3f529e50, 32'hbeade579} /* (5, 14, 1) {real, imag} */,
  {32'h3f0306a1, 32'hbef52f51} /* (5, 14, 0) {real, imag} */,
  {32'hbe943c78, 32'hbde34bd2} /* (5, 13, 15) {real, imag} */,
  {32'hbbc86900, 32'hbe03cdf2} /* (5, 13, 14) {real, imag} */,
  {32'h3f4190a7, 32'h3d808480} /* (5, 13, 13) {real, imag} */,
  {32'h3fe37731, 32'hbf78e5c4} /* (5, 13, 12) {real, imag} */,
  {32'h3f9a044d, 32'hbf095f74} /* (5, 13, 11) {real, imag} */,
  {32'h3d4c2c40, 32'h3ddaf0ec} /* (5, 13, 10) {real, imag} */,
  {32'h3d9e926c, 32'hbef16776} /* (5, 13, 9) {real, imag} */,
  {32'hbe9deabd, 32'hbea48314} /* (5, 13, 8) {real, imag} */,
  {32'hbf52b14c, 32'hbf12e9be} /* (5, 13, 7) {real, imag} */,
  {32'h3eca51f2, 32'hbf91608c} /* (5, 13, 6) {real, imag} */,
  {32'h3e33efb0, 32'h3dca4f0a} /* (5, 13, 5) {real, imag} */,
  {32'hbed115ce, 32'hbee69260} /* (5, 13, 4) {real, imag} */,
  {32'h3f12d0aa, 32'hbfa56d9a} /* (5, 13, 3) {real, imag} */,
  {32'h3f94d96a, 32'hbf03062a} /* (5, 13, 2) {real, imag} */,
  {32'h3f24da8b, 32'hbee1691b} /* (5, 13, 1) {real, imag} */,
  {32'hbecb6caa, 32'hbea874cc} /* (5, 13, 0) {real, imag} */,
  {32'hbe263491, 32'h3f70f61f} /* (5, 12, 15) {real, imag} */,
  {32'hbe3fc7ee, 32'h3f8035da} /* (5, 12, 14) {real, imag} */,
  {32'h3e6ecab0, 32'hbf0920ca} /* (5, 12, 13) {real, imag} */,
  {32'h3f2df548, 32'hbf0c6430} /* (5, 12, 12) {real, imag} */,
  {32'h3f4f4514, 32'h3f368910} /* (5, 12, 11) {real, imag} */,
  {32'h3df86184, 32'h3f1270e4} /* (5, 12, 10) {real, imag} */,
  {32'h3f9c32ea, 32'hbe7872e0} /* (5, 12, 9) {real, imag} */,
  {32'h3f25062a, 32'h3f20ae50} /* (5, 12, 8) {real, imag} */,
  {32'hbe81ebc8, 32'h3f155016} /* (5, 12, 7) {real, imag} */,
  {32'h3f862f13, 32'h3e6f27b8} /* (5, 12, 6) {real, imag} */,
  {32'h3f6ae5d8, 32'h3f15b311} /* (5, 12, 5) {real, imag} */,
  {32'h3bf45500, 32'h3e5241d0} /* (5, 12, 4) {real, imag} */,
  {32'h3e87621a, 32'hbf6f641e} /* (5, 12, 3) {real, imag} */,
  {32'h3d8f9f98, 32'hbf8eaa54} /* (5, 12, 2) {real, imag} */,
  {32'hbdcb0888, 32'hbf9773ff} /* (5, 12, 1) {real, imag} */,
  {32'hbe553f2d, 32'hbec86c1b} /* (5, 12, 0) {real, imag} */,
  {32'hbee64398, 32'h3fbbb564} /* (5, 11, 15) {real, imag} */,
  {32'hbe62eaca, 32'h3ecfd50e} /* (5, 11, 14) {real, imag} */,
  {32'hbe088bbc, 32'hbf979fac} /* (5, 11, 13) {real, imag} */,
  {32'hbd80b424, 32'hbeed2000} /* (5, 11, 12) {real, imag} */,
  {32'h3e4820c6, 32'h3f0486a0} /* (5, 11, 11) {real, imag} */,
  {32'h3f361a63, 32'hbc1a2b50} /* (5, 11, 10) {real, imag} */,
  {32'h3fcad500, 32'hbef8be6b} /* (5, 11, 9) {real, imag} */,
  {32'h3f9f71fd, 32'hbe863abe} /* (5, 11, 8) {real, imag} */,
  {32'h3c68b900, 32'hbf485ab4} /* (5, 11, 7) {real, imag} */,
  {32'hbe2675d0, 32'hbee22f14} /* (5, 11, 6) {real, imag} */,
  {32'h3f2c545a, 32'hbf6fd5ab} /* (5, 11, 5) {real, imag} */,
  {32'h3f8ed028, 32'hbf7ad5b8} /* (5, 11, 4) {real, imag} */,
  {32'h3f095af2, 32'hbd5fad54} /* (5, 11, 3) {real, imag} */,
  {32'hbf0522b0, 32'h3f51f7d4} /* (5, 11, 2) {real, imag} */,
  {32'hbf005d81, 32'h3ea1a1ec} /* (5, 11, 1) {real, imag} */,
  {32'hbe0fbb80, 32'h3e526ef1} /* (5, 11, 0) {real, imag} */,
  {32'hbd61c468, 32'h3f1d53b8} /* (5, 10, 15) {real, imag} */,
  {32'hbedbdbde, 32'hbf67c6a2} /* (5, 10, 14) {real, imag} */,
  {32'hbbe3c2c0, 32'hbfee965b} /* (5, 10, 13) {real, imag} */,
  {32'h3f4fdeb9, 32'hbf8804a7} /* (5, 10, 12) {real, imag} */,
  {32'h3e031bf8, 32'h3ed0fa80} /* (5, 10, 11) {real, imag} */,
  {32'h3dd2d942, 32'hbe96f5d8} /* (5, 10, 10) {real, imag} */,
  {32'h3fa1dcd6, 32'hbf0c6a31} /* (5, 10, 9) {real, imag} */,
  {32'h3ec37044, 32'hbfcaabdc} /* (5, 10, 8) {real, imag} */,
  {32'hbdf4c798, 32'hbfaa1bd5} /* (5, 10, 7) {real, imag} */,
  {32'hbf6525ef, 32'hbe8a7d7c} /* (5, 10, 6) {real, imag} */,
  {32'hbf36a024, 32'hbfd24a33} /* (5, 10, 5) {real, imag} */,
  {32'h3f55da96, 32'hbf645dcc} /* (5, 10, 4) {real, imag} */,
  {32'h3f98507d, 32'hbe8e2040} /* (5, 10, 3) {real, imag} */,
  {32'hbe268b90, 32'h3f564935} /* (5, 10, 2) {real, imag} */,
  {32'hbf1046b3, 32'h3f67f88e} /* (5, 10, 1) {real, imag} */,
  {32'h3cc5b1c0, 32'h3e7305b2} /* (5, 10, 0) {real, imag} */,
  {32'h3f6866c6, 32'hbdb6ad90} /* (5, 9, 15) {real, imag} */,
  {32'h3eff8b63, 32'hbe9f27cb} /* (5, 9, 14) {real, imag} */,
  {32'hbf4f5dcb, 32'hbf25a52a} /* (5, 9, 13) {real, imag} */,
  {32'h3d797bd0, 32'hbf8714a3} /* (5, 9, 12) {real, imag} */,
  {32'hbf0bcdc0, 32'h3cf8a700} /* (5, 9, 11) {real, imag} */,
  {32'hbf667e77, 32'hbf0fb0e2} /* (5, 9, 10) {real, imag} */,
  {32'h3f6128c1, 32'h3e395110} /* (5, 9, 9) {real, imag} */,
  {32'h3ec7ffa4, 32'hbecdd8c3} /* (5, 9, 8) {real, imag} */,
  {32'hbe81203c, 32'h3e9ae352} /* (5, 9, 7) {real, imag} */,
  {32'h3f20e2a6, 32'h3f633097} /* (5, 9, 6) {real, imag} */,
  {32'hbd31fa50, 32'hbf243348} /* (5, 9, 5) {real, imag} */,
  {32'hbda151f0, 32'h3e551044} /* (5, 9, 4) {real, imag} */,
  {32'h3ed7b3d1, 32'h3e91fea6} /* (5, 9, 3) {real, imag} */,
  {32'h3f25f272, 32'h3edae5cc} /* (5, 9, 2) {real, imag} */,
  {32'h3cf7a140, 32'h3e9b7d18} /* (5, 9, 1) {real, imag} */,
  {32'h3e96fcdf, 32'hbf111f79} /* (5, 9, 0) {real, imag} */,
  {32'hbe166aa8, 32'hbe29b059} /* (5, 8, 15) {real, imag} */,
  {32'hbc6df278, 32'h3e834cad} /* (5, 8, 14) {real, imag} */,
  {32'hbe8ecfb0, 32'hbea3ffcb} /* (5, 8, 13) {real, imag} */,
  {32'h3f3be7f3, 32'hbf0f2243} /* (5, 8, 12) {real, imag} */,
  {32'hbe2c4e2a, 32'hbec47f52} /* (5, 8, 11) {real, imag} */,
  {32'hbf0955bc, 32'hbf6c7d60} /* (5, 8, 10) {real, imag} */,
  {32'h3f5a791f, 32'hbe7369e4} /* (5, 8, 9) {real, imag} */,
  {32'h3f13d5e4, 32'h3decb904} /* (5, 8, 8) {real, imag} */,
  {32'hbda9ef98, 32'h3f24de18} /* (5, 8, 7) {real, imag} */,
  {32'h3f421a24, 32'h3fa8cc93} /* (5, 8, 6) {real, imag} */,
  {32'hbd9d3df0, 32'hbf1e8f99} /* (5, 8, 5) {real, imag} */,
  {32'hbf3c6399, 32'hbf359267} /* (5, 8, 4) {real, imag} */,
  {32'h3ec59350, 32'h3cadb2c0} /* (5, 8, 3) {real, imag} */,
  {32'h3f092e3f, 32'hbee08000} /* (5, 8, 2) {real, imag} */,
  {32'hbf1a193e, 32'hbeba1d18} /* (5, 8, 1) {real, imag} */,
  {32'hbf63e7b0, 32'hbe80803f} /* (5, 8, 0) {real, imag} */,
  {32'hbf2fb868, 32'hbf0a6f6f} /* (5, 7, 15) {real, imag} */,
  {32'hbf2941cb, 32'hbe3662a0} /* (5, 7, 14) {real, imag} */,
  {32'h3eadbfe0, 32'h3ee8b495} /* (5, 7, 13) {real, imag} */,
  {32'h3ecd4bdc, 32'hbdc33a6c} /* (5, 7, 12) {real, imag} */,
  {32'hbe2d95c8, 32'hbf5901e8} /* (5, 7, 11) {real, imag} */,
  {32'h3e4d2a24, 32'hbf9136da} /* (5, 7, 10) {real, imag} */,
  {32'h3ef5df42, 32'hbf1ec694} /* (5, 7, 9) {real, imag} */,
  {32'hbf166658, 32'h3db32583} /* (5, 7, 8) {real, imag} */,
  {32'hbf35e91e, 32'h3daa5493} /* (5, 7, 7) {real, imag} */,
  {32'hbe36a4a0, 32'h3f9f8e40} /* (5, 7, 6) {real, imag} */,
  {32'hbef9fdae, 32'h3e5193a0} /* (5, 7, 5) {real, imag} */,
  {32'hbda85818, 32'hbeaec859} /* (5, 7, 4) {real, imag} */,
  {32'h3fa55fe1, 32'hbe7a2634} /* (5, 7, 3) {real, imag} */,
  {32'h3fad9e3e, 32'hbf3a5c5a} /* (5, 7, 2) {real, imag} */,
  {32'hbe59c79c, 32'h3c40cc40} /* (5, 7, 1) {real, imag} */,
  {32'hbf94b0b1, 32'hbe22cf80} /* (5, 7, 0) {real, imag} */,
  {32'hbe89685b, 32'hbe469168} /* (5, 6, 15) {real, imag} */,
  {32'hbfa5c52a, 32'h3ca74580} /* (5, 6, 14) {real, imag} */,
  {32'hbf0f3721, 32'h3ef537c5} /* (5, 6, 13) {real, imag} */,
  {32'hbf1be78e, 32'h3eab6ec2} /* (5, 6, 12) {real, imag} */,
  {32'hbf30d620, 32'hbed4a056} /* (5, 6, 11) {real, imag} */,
  {32'h3f72e098, 32'hbf06e62d} /* (5, 6, 10) {real, imag} */,
  {32'h3e7af0b4, 32'hbfa25c05} /* (5, 6, 9) {real, imag} */,
  {32'hbf93aada, 32'hbf95b607} /* (5, 6, 8) {real, imag} */,
  {32'hbf21e240, 32'hbebf74a8} /* (5, 6, 7) {real, imag} */,
  {32'h3e81beb2, 32'h3f60909d} /* (5, 6, 6) {real, imag} */,
  {32'h3cb7b4e0, 32'h3fbd79de} /* (5, 6, 5) {real, imag} */,
  {32'hbe0152f2, 32'h3d909d68} /* (5, 6, 4) {real, imag} */,
  {32'h3e5933a6, 32'hbe9e4940} /* (5, 6, 3) {real, imag} */,
  {32'h3f5affe3, 32'hbd823c4c} /* (5, 6, 2) {real, imag} */,
  {32'h3f01eb17, 32'hbed167d8} /* (5, 6, 1) {real, imag} */,
  {32'hbdcc2360, 32'hbf3aea15} /* (5, 6, 0) {real, imag} */,
  {32'hbe4da880, 32'h3e12d9d0} /* (5, 5, 15) {real, imag} */,
  {32'hbf9ad43d, 32'h3edbc326} /* (5, 5, 14) {real, imag} */,
  {32'hbecb28dc, 32'h3f2cd22d} /* (5, 5, 13) {real, imag} */,
  {32'hbed14e16, 32'h3eeb8dad} /* (5, 5, 12) {real, imag} */,
  {32'hbe8d2c19, 32'hbf6c80e2} /* (5, 5, 11) {real, imag} */,
  {32'h3e948b5e, 32'hbdfb1454} /* (5, 5, 10) {real, imag} */,
  {32'h3e82af4b, 32'hbf129bf2} /* (5, 5, 9) {real, imag} */,
  {32'hbe36da40, 32'hbf9fc4a6} /* (5, 5, 8) {real, imag} */,
  {32'h3c66e940, 32'hbeb51642} /* (5, 5, 7) {real, imag} */,
  {32'h3fbb4427, 32'h3d549038} /* (5, 5, 6) {real, imag} */,
  {32'h3fa8542a, 32'h3bf76f40} /* (5, 5, 5) {real, imag} */,
  {32'h3e55aeca, 32'hbf89547d} /* (5, 5, 4) {real, imag} */,
  {32'hbf041ade, 32'hbf9a579f} /* (5, 5, 3) {real, imag} */,
  {32'hbf1394bd, 32'hbec6f89b} /* (5, 5, 2) {real, imag} */,
  {32'hbf0bad94, 32'hbf8f9f38} /* (5, 5, 1) {real, imag} */,
  {32'hbe6efa82, 32'hbf3f2165} /* (5, 5, 0) {real, imag} */,
  {32'hbea5894c, 32'h3f14c1fb} /* (5, 4, 15) {real, imag} */,
  {32'hbf364da9, 32'h3f02913e} /* (5, 4, 14) {real, imag} */,
  {32'h3f156892, 32'h3ebadd58} /* (5, 4, 13) {real, imag} */,
  {32'h3f5a31aa, 32'h3ee1efe3} /* (5, 4, 12) {real, imag} */,
  {32'h3e7d7b4a, 32'hbf6f74f3} /* (5, 4, 11) {real, imag} */,
  {32'hbf109600, 32'hbf023978} /* (5, 4, 10) {real, imag} */,
  {32'hbe47d120, 32'hbf7f975f} /* (5, 4, 9) {real, imag} */,
  {32'h3e878dea, 32'hbf0b520c} /* (5, 4, 8) {real, imag} */,
  {32'hbf28d12c, 32'hbbb89600} /* (5, 4, 7) {real, imag} */,
  {32'h3e1bdd63, 32'h3e8293ad} /* (5, 4, 6) {real, imag} */,
  {32'h3f29cc8a, 32'h3f473ced} /* (5, 4, 5) {real, imag} */,
  {32'hbe68f246, 32'h3dafe6e4} /* (5, 4, 4) {real, imag} */,
  {32'hbf1e1f00, 32'hbf43c100} /* (5, 4, 3) {real, imag} */,
  {32'hbf13c926, 32'hbeb4e8e6} /* (5, 4, 2) {real, imag} */,
  {32'hbf42bdd4, 32'hbf5ec0b8} /* (5, 4, 1) {real, imag} */,
  {32'hbe58a7c0, 32'hbf991e94} /* (5, 4, 0) {real, imag} */,
  {32'hbf226782, 32'h3e410d7c} /* (5, 3, 15) {real, imag} */,
  {32'hbecfcfd6, 32'hbe5fcfb4} /* (5, 3, 14) {real, imag} */,
  {32'h3f8882c8, 32'hbf21d5c4} /* (5, 3, 13) {real, imag} */,
  {32'h3ea5f240, 32'hbf33f898} /* (5, 3, 12) {real, imag} */,
  {32'hbe330120, 32'hbf44a27a} /* (5, 3, 11) {real, imag} */,
  {32'hbf498d70, 32'hbe358dc4} /* (5, 3, 10) {real, imag} */,
  {32'h3efb5760, 32'hbf0777a5} /* (5, 3, 9) {real, imag} */,
  {32'h3fbf2cba, 32'hbf03ec9c} /* (5, 3, 8) {real, imag} */,
  {32'h3f40bd62, 32'hbeda064a} /* (5, 3, 7) {real, imag} */,
  {32'hbf00e8a4, 32'h3eb6a342} /* (5, 3, 6) {real, imag} */,
  {32'h3f196104, 32'h3f817f85} /* (5, 3, 5) {real, imag} */,
  {32'h3f620785, 32'h3f4b37bd} /* (5, 3, 4) {real, imag} */,
  {32'hbf005ba4, 32'hbeb99660} /* (5, 3, 3) {real, imag} */,
  {32'hbe9b14aa, 32'h3e15647c} /* (5, 3, 2) {real, imag} */,
  {32'hbf01d385, 32'h3fbe030c} /* (5, 3, 1) {real, imag} */,
  {32'hbf59d754, 32'hbecd3e34} /* (5, 3, 0) {real, imag} */,
  {32'hbe9d80c6, 32'hbe5e0d3e} /* (5, 2, 15) {real, imag} */,
  {32'h3e7d06d8, 32'hbdb05fac} /* (5, 2, 14) {real, imag} */,
  {32'h3f9337dc, 32'hbf3526f8} /* (5, 2, 13) {real, imag} */,
  {32'h3e56d8a4, 32'hbfc9c7f0} /* (5, 2, 12) {real, imag} */,
  {32'hbeb319c1, 32'hbf065a1b} /* (5, 2, 11) {real, imag} */,
  {32'hbf05bf86, 32'hbeb007a6} /* (5, 2, 10) {real, imag} */,
  {32'hbd97c90c, 32'hbdc2f3f4} /* (5, 2, 9) {real, imag} */,
  {32'h3ed90a2c, 32'hbdab1ac8} /* (5, 2, 8) {real, imag} */,
  {32'h3f6b7b2c, 32'hbe709f54} /* (5, 2, 7) {real, imag} */,
  {32'hbe86fe79, 32'h3d429a30} /* (5, 2, 6) {real, imag} */,
  {32'h3e5a2d10, 32'hbe58a634} /* (5, 2, 5) {real, imag} */,
  {32'h3f0a5607, 32'h3ee3f212} /* (5, 2, 4) {real, imag} */,
  {32'h3d895d04, 32'h3f2e88b9} /* (5, 2, 3) {real, imag} */,
  {32'h3ef69f1f, 32'h3f56f02a} /* (5, 2, 2) {real, imag} */,
  {32'h3e819200, 32'h3ff22557} /* (5, 2, 1) {real, imag} */,
  {32'hbdf89560, 32'h3e2eeda8} /* (5, 2, 0) {real, imag} */,
  {32'h3e8118fb, 32'hbf693490} /* (5, 1, 15) {real, imag} */,
  {32'h3f0334b1, 32'hbe9b4368} /* (5, 1, 14) {real, imag} */,
  {32'h3f913b4c, 32'hbe7eb865} /* (5, 1, 13) {real, imag} */,
  {32'h3eb921d0, 32'hbf1c50e9} /* (5, 1, 12) {real, imag} */,
  {32'hbe88aa44, 32'h3f48e872} /* (5, 1, 11) {real, imag} */,
  {32'hbf8ecc42, 32'h3d2c7d40} /* (5, 1, 10) {real, imag} */,
  {32'hbfa17ac8, 32'h3dd6cbec} /* (5, 1, 9) {real, imag} */,
  {32'hbe846a6c, 32'h3d54e770} /* (5, 1, 8) {real, imag} */,
  {32'hbe54ad10, 32'hbe76b370} /* (5, 1, 7) {real, imag} */,
  {32'h3cc32550, 32'hbefe0836} /* (5, 1, 6) {real, imag} */,
  {32'h3f2e24e0, 32'hbf89bc7c} /* (5, 1, 5) {real, imag} */,
  {32'h3f9cd398, 32'h3eca7878} /* (5, 1, 4) {real, imag} */,
  {32'h3fa1894e, 32'h3f147a46} /* (5, 1, 3) {real, imag} */,
  {32'h3f1c7dd4, 32'h3f19df04} /* (5, 1, 2) {real, imag} */,
  {32'h3f16f7f6, 32'h3e8c3288} /* (5, 1, 1) {real, imag} */,
  {32'h3f5581ae, 32'hbf1e8adc} /* (5, 1, 0) {real, imag} */,
  {32'h3e417442, 32'hbe9f7a22} /* (5, 0, 15) {real, imag} */,
  {32'h3ec694ef, 32'hbea9ea12} /* (5, 0, 14) {real, imag} */,
  {32'h3f82bbea, 32'hbe902260} /* (5, 0, 13) {real, imag} */,
  {32'h3f38c444, 32'h3e13ddbc} /* (5, 0, 12) {real, imag} */,
  {32'h3eb574b2, 32'h3ef4ddfb} /* (5, 0, 11) {real, imag} */,
  {32'h3d45fbf4, 32'h3e964616} /* (5, 0, 10) {real, imag} */,
  {32'hbf21699a, 32'h3e3683d2} /* (5, 0, 9) {real, imag} */,
  {32'hbed57dc5, 32'hbde81a06} /* (5, 0, 8) {real, imag} */,
  {32'hbf1e01ef, 32'hbd9a4c28} /* (5, 0, 7) {real, imag} */,
  {32'hbe8369b1, 32'hbec64a84} /* (5, 0, 6) {real, imag} */,
  {32'h3f46b45c, 32'hbf12f006} /* (5, 0, 5) {real, imag} */,
  {32'h3f351f4c, 32'h3dac9c20} /* (5, 0, 4) {real, imag} */,
  {32'h3e806b05, 32'h3ee84482} /* (5, 0, 3) {real, imag} */,
  {32'h3cc80580, 32'h3f3e8f35} /* (5, 0, 2) {real, imag} */,
  {32'h3f3f4317, 32'h3d594558} /* (5, 0, 1) {real, imag} */,
  {32'h3f4b1cf4, 32'hbef1eb4a} /* (5, 0, 0) {real, imag} */,
  {32'h3e2db84c, 32'h3efc10c2} /* (4, 15, 15) {real, imag} */,
  {32'h3c2c5490, 32'h3e1481e6} /* (4, 15, 14) {real, imag} */,
  {32'hbd9569d0, 32'hbd6a3788} /* (4, 15, 13) {real, imag} */,
  {32'h3eb1c1b4, 32'hbe8e9974} /* (4, 15, 12) {real, imag} */,
  {32'h3e97268d, 32'h3f0cda53} /* (4, 15, 11) {real, imag} */,
  {32'hbf33a30b, 32'h3f435b32} /* (4, 15, 10) {real, imag} */,
  {32'hbec2a720, 32'h3ef50946} /* (4, 15, 9) {real, imag} */,
  {32'hbf2b0926, 32'hbe91f5a0} /* (4, 15, 8) {real, imag} */,
  {32'hbf8c7b14, 32'hbd59dc3c} /* (4, 15, 7) {real, imag} */,
  {32'hbdffb4e5, 32'h3efa3dc9} /* (4, 15, 6) {real, imag} */,
  {32'h3e8d8577, 32'hbb30e700} /* (4, 15, 5) {real, imag} */,
  {32'h3f83f65b, 32'hbf4d97dd} /* (4, 15, 4) {real, imag} */,
  {32'h3fd20bee, 32'hbe972cf7} /* (4, 15, 3) {real, imag} */,
  {32'h3f44c595, 32'hbedf88a8} /* (4, 15, 2) {real, imag} */,
  {32'h3f0c9136, 32'hbf15c9b4} /* (4, 15, 1) {real, imag} */,
  {32'h3e7e7fdb, 32'hbf66f0d8} /* (4, 15, 0) {real, imag} */,
  {32'hbe2b379c, 32'h3f3632ae} /* (4, 14, 15) {real, imag} */,
  {32'hbf5f24ea, 32'hbeaa1e17} /* (4, 14, 14) {real, imag} */,
  {32'hbf85c1bd, 32'hbf205c5b} /* (4, 14, 13) {real, imag} */,
  {32'hbdf5e958, 32'hbed2900a} /* (4, 14, 12) {real, imag} */,
  {32'h3e90aef6, 32'h3f3c2666} /* (4, 14, 11) {real, imag} */,
  {32'hbff2dec1, 32'h3eaefb8a} /* (4, 14, 10) {real, imag} */,
  {32'hbf36cb64, 32'hbbf84f80} /* (4, 14, 9) {real, imag} */,
  {32'hbf4889a4, 32'h3f634fbc} /* (4, 14, 8) {real, imag} */,
  {32'hbf871877, 32'h3cb1b080} /* (4, 14, 7) {real, imag} */,
  {32'h3e49679c, 32'hbf084efe} /* (4, 14, 6) {real, imag} */,
  {32'h3e561e06, 32'hbe025bb8} /* (4, 14, 5) {real, imag} */,
  {32'h3ee518f4, 32'h3eccae62} /* (4, 14, 4) {real, imag} */,
  {32'h3fb8d18b, 32'h3fe268c4} /* (4, 14, 3) {real, imag} */,
  {32'h3fd70201, 32'h3fe43ddb} /* (4, 14, 2) {real, imag} */,
  {32'h3f893ed7, 32'hbe3a9221} /* (4, 14, 1) {real, imag} */,
  {32'h3e399382, 32'hbf60923f} /* (4, 14, 0) {real, imag} */,
  {32'hbf2be4fe, 32'h3f15cf38} /* (4, 13, 15) {real, imag} */,
  {32'hbf6ac1ca, 32'h3f0253ae} /* (4, 13, 14) {real, imag} */,
  {32'h3d645c60, 32'h3e85ca4c} /* (4, 13, 13) {real, imag} */,
  {32'h3f9c8320, 32'h3f6ea84a} /* (4, 13, 12) {real, imag} */,
  {32'hba5afe00, 32'h3f0d2bb2} /* (4, 13, 11) {real, imag} */,
  {32'hbf540a86, 32'h3cd4ca20} /* (4, 13, 10) {real, imag} */,
  {32'h3f01691a, 32'h3f08e92a} /* (4, 13, 9) {real, imag} */,
  {32'hbdabcbe2, 32'h3fb5a7cd} /* (4, 13, 8) {real, imag} */,
  {32'hbf7e18c3, 32'h3fa9a0a0} /* (4, 13, 7) {real, imag} */,
  {32'hbef736ba, 32'h3f88a3d4} /* (4, 13, 6) {real, imag} */,
  {32'h3f44881c, 32'h3f79e769} /* (4, 13, 5) {real, imag} */,
  {32'h3f550071, 32'h3fd63ef0} /* (4, 13, 4) {real, imag} */,
  {32'h3f1fb0d0, 32'h3fb9dd7e} /* (4, 13, 3) {real, imag} */,
  {32'h3f85d2dd, 32'h3f986a33} /* (4, 13, 2) {real, imag} */,
  {32'hbe267152, 32'h3fd795f6} /* (4, 13, 1) {real, imag} */,
  {32'hbedfbd90, 32'h3f17ce74} /* (4, 13, 0) {real, imag} */,
  {32'hbe99c727, 32'h3f006ad4} /* (4, 12, 15) {real, imag} */,
  {32'h3f0f994b, 32'h3dfa7c0c} /* (4, 12, 14) {real, imag} */,
  {32'h3f89d34b, 32'h3eaab8b0} /* (4, 12, 13) {real, imag} */,
  {32'h3fb4e1bd, 32'h3f82ebf8} /* (4, 12, 12) {real, imag} */,
  {32'h3f460d2c, 32'h3e222d0e} /* (4, 12, 11) {real, imag} */,
  {32'h3f1689de, 32'hbe2eca0c} /* (4, 12, 10) {real, imag} */,
  {32'h3cbe2748, 32'hbddaabb0} /* (4, 12, 9) {real, imag} */,
  {32'hbfdb5c37, 32'h3e880129} /* (4, 12, 8) {real, imag} */,
  {32'hbfd058fa, 32'h3fb9ee4c} /* (4, 12, 7) {real, imag} */,
  {32'hbfbe932f, 32'h40012964} /* (4, 12, 6) {real, imag} */,
  {32'hbe83991c, 32'h3f882527} /* (4, 12, 5) {real, imag} */,
  {32'hbef633f1, 32'h3ed1a3f7} /* (4, 12, 4) {real, imag} */,
  {32'h3ef08cff, 32'h3e7fdabe} /* (4, 12, 3) {real, imag} */,
  {32'h3f2b2452, 32'h3f592b9e} /* (4, 12, 2) {real, imag} */,
  {32'hbd4d6df0, 32'h3f3b1521} /* (4, 12, 1) {real, imag} */,
  {32'h3cccf7d0, 32'h3f8ad4e9} /* (4, 12, 0) {real, imag} */,
  {32'hbf276ff9, 32'h3d812bbc} /* (4, 11, 15) {real, imag} */,
  {32'hbfb5dd31, 32'hbd23d5e0} /* (4, 11, 14) {real, imag} */,
  {32'hbe7b7ce0, 32'h3e95d954} /* (4, 11, 13) {real, imag} */,
  {32'hbf09a4b5, 32'h3dcb2510} /* (4, 11, 12) {real, imag} */,
  {32'h3d66df68, 32'hbc5e1fc0} /* (4, 11, 11) {real, imag} */,
  {32'h3faa73e6, 32'hbbb8b0c0} /* (4, 11, 10) {real, imag} */,
  {32'h3e9e1942, 32'hbf15ea14} /* (4, 11, 9) {real, imag} */,
  {32'hbf67276a, 32'h3a6fcc40} /* (4, 11, 8) {real, imag} */,
  {32'h3f43a820, 32'h3f7da5b2} /* (4, 11, 7) {real, imag} */,
  {32'h3e5951c4, 32'h3f23e1ba} /* (4, 11, 6) {real, imag} */,
  {32'hbf641712, 32'h3f4a0153} /* (4, 11, 5) {real, imag} */,
  {32'hbffbef5e, 32'h3f03c71c} /* (4, 11, 4) {real, imag} */,
  {32'hbf7cbf5d, 32'h3f380cb3} /* (4, 11, 3) {real, imag} */,
  {32'h3e039c70, 32'h3f9cfc99} /* (4, 11, 2) {real, imag} */,
  {32'h3d0ab1d4, 32'hbe0ada10} /* (4, 11, 1) {real, imag} */,
  {32'h3e0a71b2, 32'h3f20025c} /* (4, 11, 0) {real, imag} */,
  {32'hbfa78195, 32'hbe1ae552} /* (4, 10, 15) {real, imag} */,
  {32'hbfef41fa, 32'hbf2e01c0} /* (4, 10, 14) {real, imag} */,
  {32'h3f82d79e, 32'hbd83b52c} /* (4, 10, 13) {real, imag} */,
  {32'h3e97e68d, 32'h3d8fa4b4} /* (4, 10, 12) {real, imag} */,
  {32'h3eb646ae, 32'h3ea9d408} /* (4, 10, 11) {real, imag} */,
  {32'h3fa174dd, 32'h3f9ad41d} /* (4, 10, 10) {real, imag} */,
  {32'h3f74d434, 32'hbf795db3} /* (4, 10, 9) {real, imag} */,
  {32'h3eba4749, 32'hbf4b2c4d} /* (4, 10, 8) {real, imag} */,
  {32'hbdfbda50, 32'h3f391641} /* (4, 10, 7) {real, imag} */,
  {32'h3bdbd380, 32'hbed7b3a0} /* (4, 10, 6) {real, imag} */,
  {32'hbfbecd7c, 32'h3faa7389} /* (4, 10, 5) {real, imag} */,
  {32'hc001dbc0, 32'h3fd73b6c} /* (4, 10, 4) {real, imag} */,
  {32'hbf9ffb62, 32'h3ec4bab7} /* (4, 10, 3) {real, imag} */,
  {32'hbf3d4196, 32'h3f37fdb9} /* (4, 10, 2) {real, imag} */,
  {32'hbf512517, 32'h3edc8f5f} /* (4, 10, 1) {real, imag} */,
  {32'hbf2408da, 32'h3e3de8d4} /* (4, 10, 0) {real, imag} */,
  {32'hbfbe2f69, 32'hbf75fcf2} /* (4, 9, 15) {real, imag} */,
  {32'hbfb8a0ee, 32'hbfeadec5} /* (4, 9, 14) {real, imag} */,
  {32'h3e9040b6, 32'hbf1b4d21} /* (4, 9, 13) {real, imag} */,
  {32'hbea3cd44, 32'h3f123cb5} /* (4, 9, 12) {real, imag} */,
  {32'hbf613a74, 32'h3eee9847} /* (4, 9, 11) {real, imag} */,
  {32'hbeb75c20, 32'hbdcc0c20} /* (4, 9, 10) {real, imag} */,
  {32'hbf42ca87, 32'hbf2aa217} /* (4, 9, 9) {real, imag} */,
  {32'hbfe219e4, 32'hbf1cde3c} /* (4, 9, 8) {real, imag} */,
  {32'hbf8d1357, 32'hbf0807bf} /* (4, 9, 7) {real, imag} */,
  {32'h3f3de74a, 32'hbe75df64} /* (4, 9, 6) {real, imag} */,
  {32'hbf5b709e, 32'hbf08ffba} /* (4, 9, 5) {real, imag} */,
  {32'hbfb09a76, 32'hbd9c8d98} /* (4, 9, 4) {real, imag} */,
  {32'hbfcddf16, 32'hbefbfd0f} /* (4, 9, 3) {real, imag} */,
  {32'hbf291a6f, 32'hbf37bcea} /* (4, 9, 2) {real, imag} */,
  {32'h3e759948, 32'h3efda74a} /* (4, 9, 1) {real, imag} */,
  {32'hbea9d348, 32'hbef72fb8} /* (4, 9, 0) {real, imag} */,
  {32'hbf829a10, 32'hbe42d8d8} /* (4, 8, 15) {real, imag} */,
  {32'hbf81c347, 32'hbf072f61} /* (4, 8, 14) {real, imag} */,
  {32'hbe173f5b, 32'h3d274448} /* (4, 8, 13) {real, imag} */,
  {32'h3ee37386, 32'hbe98f4c4} /* (4, 8, 12) {real, imag} */,
  {32'hbf903e8a, 32'h3e9a8aa1} /* (4, 8, 11) {real, imag} */,
  {32'hbf9d9524, 32'hbd42b0a6} /* (4, 8, 10) {real, imag} */,
  {32'hbff19486, 32'h3efce0b8} /* (4, 8, 9) {real, imag} */,
  {32'hc0061b0d, 32'hbed690d9} /* (4, 8, 8) {real, imag} */,
  {32'hbfb32e19, 32'hbf9b9ed0} /* (4, 8, 7) {real, imag} */,
  {32'h3f4c434f, 32'h3f45c20d} /* (4, 8, 6) {real, imag} */,
  {32'hbe99d14f, 32'hbe69bd65} /* (4, 8, 5) {real, imag} */,
  {32'hc0092af7, 32'hbf0a0ca6} /* (4, 8, 4) {real, imag} */,
  {32'hc00e9740, 32'hbf01856a} /* (4, 8, 3) {real, imag} */,
  {32'hbe1c5f5a, 32'hbfeb502a} /* (4, 8, 2) {real, imag} */,
  {32'h3fd67e76, 32'hbf2059ac} /* (4, 8, 1) {real, imag} */,
  {32'h3f83d8ea, 32'hbee1a675} /* (4, 8, 0) {real, imag} */,
  {32'hbfb0a214, 32'h3e5ae239} /* (4, 7, 15) {real, imag} */,
  {32'hbf611cee, 32'hbeb8a452} /* (4, 7, 14) {real, imag} */,
  {32'hbe1740d0, 32'hbf89cf06} /* (4, 7, 13) {real, imag} */,
  {32'h3fd93d70, 32'hbfbc2860} /* (4, 7, 12) {real, imag} */,
  {32'h3dc85940, 32'h3f3fabcf} /* (4, 7, 11) {real, imag} */,
  {32'h3ea7c92a, 32'h3f81776b} /* (4, 7, 10) {real, imag} */,
  {32'h3f517032, 32'h3f43d80c} /* (4, 7, 9) {real, imag} */,
  {32'h3e9f5b82, 32'hbf185156} /* (4, 7, 8) {real, imag} */,
  {32'hbd9799d1, 32'hbf531438} /* (4, 7, 7) {real, imag} */,
  {32'h3f5a6355, 32'h3e2a56d6} /* (4, 7, 6) {real, imag} */,
  {32'h3e9b769e, 32'hbf656fe2} /* (4, 7, 5) {real, imag} */,
  {32'hbf927714, 32'hbf511f78} /* (4, 7, 4) {real, imag} */,
  {32'hbfb275a3, 32'hbed4d2f0} /* (4, 7, 3) {real, imag} */,
  {32'hbec5da7c, 32'hbfac586e} /* (4, 7, 2) {real, imag} */,
  {32'hbdfc5644, 32'hc01e8224} /* (4, 7, 1) {real, imag} */,
  {32'hbee7bcfb, 32'hbf9d8e26} /* (4, 7, 0) {real, imag} */,
  {32'hbf96189d, 32'hbf48fee3} /* (4, 6, 15) {real, imag} */,
  {32'hbf2f38e9, 32'hbfb9ab34} /* (4, 6, 14) {real, imag} */,
  {32'hbf57c8a0, 32'hbf9ac100} /* (4, 6, 13) {real, imag} */,
  {32'hbf88f430, 32'hbf6673e9} /* (4, 6, 12) {real, imag} */,
  {32'hbf329460, 32'h3e3fed50} /* (4, 6, 11) {real, imag} */,
  {32'hbf079191, 32'hbeea988c} /* (4, 6, 10) {real, imag} */,
  {32'h3df70488, 32'h3f56dbe2} /* (4, 6, 9) {real, imag} */,
  {32'h3ec0a670, 32'h3fa3525e} /* (4, 6, 8) {real, imag} */,
  {32'h3ea891d0, 32'h3e550600} /* (4, 6, 7) {real, imag} */,
  {32'h3f7d1002, 32'h3eb6a20b} /* (4, 6, 6) {real, imag} */,
  {32'h3fd2bfb7, 32'hbf5acaad} /* (4, 6, 5) {real, imag} */,
  {32'h3ef370b0, 32'hbf026f19} /* (4, 6, 4) {real, imag} */,
  {32'hbf610cb2, 32'h3f54fb79} /* (4, 6, 3) {real, imag} */,
  {32'hbf105bc6, 32'h3ec324b4} /* (4, 6, 2) {real, imag} */,
  {32'hbf6aaa9f, 32'hbf6f240c} /* (4, 6, 1) {real, imag} */,
  {32'hbf960188, 32'hbfa8c918} /* (4, 6, 0) {real, imag} */,
  {32'h3dfbcf42, 32'hbeb18378} /* (4, 5, 15) {real, imag} */,
  {32'h3e914391, 32'hbf277de5} /* (4, 5, 14) {real, imag} */,
  {32'h3f0591a2, 32'hbf32153d} /* (4, 5, 13) {real, imag} */,
  {32'h3f8ec92c, 32'hbf821724} /* (4, 5, 12) {real, imag} */,
  {32'h3e1518b4, 32'hbf80a313} /* (4, 5, 11) {real, imag} */,
  {32'h3e72ff44, 32'hbf1f417f} /* (4, 5, 10) {real, imag} */,
  {32'hbd5c0fd8, 32'h3fe6dee3} /* (4, 5, 9) {real, imag} */,
  {32'hbf04c262, 32'h3fafe750} /* (4, 5, 8) {real, imag} */,
  {32'h3f30c6f6, 32'h3f74e45f} /* (4, 5, 7) {real, imag} */,
  {32'h401255d6, 32'hbec971a0} /* (4, 5, 6) {real, imag} */,
  {32'h3fd3cb10, 32'hbf4e47c5} /* (4, 5, 5) {real, imag} */,
  {32'h3f891d7c, 32'h3e008248} /* (4, 5, 4) {real, imag} */,
  {32'h3fc54433, 32'hbe0633c6} /* (4, 5, 3) {real, imag} */,
  {32'h3f853f1f, 32'hbda11ea4} /* (4, 5, 2) {real, imag} */,
  {32'hbef8012c, 32'h3f66de34} /* (4, 5, 1) {real, imag} */,
  {32'hbedb6e83, 32'hbea6cacf} /* (4, 5, 0) {real, imag} */,
  {32'h3e9a900a, 32'hbe5cb90c} /* (4, 4, 15) {real, imag} */,
  {32'h3f36f6bb, 32'hbebb2ec4} /* (4, 4, 14) {real, imag} */,
  {32'h3f72be92, 32'hbfa4d4c2} /* (4, 4, 13) {real, imag} */,
  {32'h3fff3832, 32'hbf5ea6b0} /* (4, 4, 12) {real, imag} */,
  {32'h3e0fc926, 32'h3def1566} /* (4, 4, 11) {real, imag} */,
  {32'hbcbb30b0, 32'h3e455790} /* (4, 4, 10) {real, imag} */,
  {32'h3e2f4e02, 32'h3f7affef} /* (4, 4, 9) {real, imag} */,
  {32'hbf31c845, 32'h3f6e17c1} /* (4, 4, 8) {real, imag} */,
  {32'h3f6ed550, 32'h3ca8c164} /* (4, 4, 7) {real, imag} */,
  {32'h3f8fdbb5, 32'hbe53155e} /* (4, 4, 6) {real, imag} */,
  {32'h3f81e64e, 32'h3efa31d2} /* (4, 4, 5) {real, imag} */,
  {32'h3f5b4871, 32'h3f97cf97} /* (4, 4, 4) {real, imag} */,
  {32'h3f8c41f4, 32'h3ef4872f} /* (4, 4, 3) {real, imag} */,
  {32'h3dd2aa13, 32'hbf1dabe9} /* (4, 4, 2) {real, imag} */,
  {32'hbf97bae2, 32'hbec7fd2a} /* (4, 4, 1) {real, imag} */,
  {32'hbf2c6ba4, 32'hbec35f96} /* (4, 4, 0) {real, imag} */,
  {32'h3f46c29c, 32'h3d7e01c0} /* (4, 3, 15) {real, imag} */,
  {32'h3e79f676, 32'hbeedca6c} /* (4, 3, 14) {real, imag} */,
  {32'hbf81acf2, 32'hbfab834c} /* (4, 3, 13) {real, imag} */,
  {32'h3f962c2c, 32'hbf99a216} /* (4, 3, 12) {real, imag} */,
  {32'hbdba0458, 32'hbf1105ac} /* (4, 3, 11) {real, imag} */,
  {32'hbf526218, 32'h3e7b56e7} /* (4, 3, 10) {real, imag} */,
  {32'h3f12b25c, 32'hbf77381a} /* (4, 3, 9) {real, imag} */,
  {32'h3e9afaa4, 32'hbf013ba8} /* (4, 3, 8) {real, imag} */,
  {32'h4015346e, 32'hbee0d228} /* (4, 3, 7) {real, imag} */,
  {32'h3fb1bf54, 32'h3fc71c78} /* (4, 3, 6) {real, imag} */,
  {32'h3ea709c7, 32'h400a5373} /* (4, 3, 5) {real, imag} */,
  {32'h3f156c82, 32'h3fc44034} /* (4, 3, 4) {real, imag} */,
  {32'hbf1782d2, 32'h3f5aa594} /* (4, 3, 3) {real, imag} */,
  {32'hbfd6e0f3, 32'hbe114f5a} /* (4, 3, 2) {real, imag} */,
  {32'hbfd8b6d2, 32'hbf7f4fa6} /* (4, 3, 1) {real, imag} */,
  {32'hbfa26b3d, 32'hbf237df2} /* (4, 3, 0) {real, imag} */,
  {32'hbdf41a28, 32'h3e7107fc} /* (4, 2, 15) {real, imag} */,
  {32'hbf584b3a, 32'hbf2f389d} /* (4, 2, 14) {real, imag} */,
  {32'hbf93ddd2, 32'hbd19f0a0} /* (4, 2, 13) {real, imag} */,
  {32'hbd5fd4f0, 32'h3e9f0614} /* (4, 2, 12) {real, imag} */,
  {32'h3e7cbfe4, 32'hbe0b27c4} /* (4, 2, 11) {real, imag} */,
  {32'hbdf98840, 32'h3f686d30} /* (4, 2, 10) {real, imag} */,
  {32'h3f622f9c, 32'hbdb6ab10} /* (4, 2, 9) {real, imag} */,
  {32'h3e8b6a78, 32'hbf58a6c5} /* (4, 2, 8) {real, imag} */,
  {32'h3df5d9dc, 32'hbf8e5680} /* (4, 2, 7) {real, imag} */,
  {32'h3e880628, 32'h3ed61f8a} /* (4, 2, 6) {real, imag} */,
  {32'h3fbc569e, 32'hbea63fba} /* (4, 2, 5) {real, imag} */,
  {32'h3f46a517, 32'hbfb05afd} /* (4, 2, 4) {real, imag} */,
  {32'hbef16c5a, 32'hbf882d3e} /* (4, 2, 3) {real, imag} */,
  {32'hbdbd9c70, 32'hbf872ceb} /* (4, 2, 2) {real, imag} */,
  {32'h3f0a4ff4, 32'hbfdcd87b} /* (4, 2, 1) {real, imag} */,
  {32'hbedcd534, 32'hbed58b90} /* (4, 2, 0) {real, imag} */,
  {32'hbefef650, 32'h3f2fbd18} /* (4, 1, 15) {real, imag} */,
  {32'hbf5c7872, 32'hbdfbc23c} /* (4, 1, 14) {real, imag} */,
  {32'hbd8a6f78, 32'hbf1ae05b} /* (4, 1, 13) {real, imag} */,
  {32'h3e9bf510, 32'hbed08054} /* (4, 1, 12) {real, imag} */,
  {32'h3d50a1d0, 32'hbdb99058} /* (4, 1, 11) {real, imag} */,
  {32'hbe2a6fe8, 32'h3eec0c1e} /* (4, 1, 10) {real, imag} */,
  {32'h3e82696e, 32'hbf2bcf6c} /* (4, 1, 9) {real, imag} */,
  {32'h3f7ec66e, 32'hbf8946ce} /* (4, 1, 8) {real, imag} */,
  {32'h3f7b8d18, 32'h3e4f3c32} /* (4, 1, 7) {real, imag} */,
  {32'h3f875444, 32'hbc00ab60} /* (4, 1, 6) {real, imag} */,
  {32'h3fddf298, 32'hbf8de5e5} /* (4, 1, 5) {real, imag} */,
  {32'hbf06871c, 32'hbe8ca3f6} /* (4, 1, 4) {real, imag} */,
  {32'hbf4fd96c, 32'h3f4c00cc} /* (4, 1, 3) {real, imag} */,
  {32'h3d5f43a0, 32'h3f6d4552} /* (4, 1, 2) {real, imag} */,
  {32'h3e082b28, 32'hbf97b0af} /* (4, 1, 1) {real, imag} */,
  {32'hbe87723b, 32'h3e199efa} /* (4, 1, 0) {real, imag} */,
  {32'hbf2e6fe8, 32'hbe3d73c5} /* (4, 0, 15) {real, imag} */,
  {32'hbe9d99ab, 32'hbcba42c0} /* (4, 0, 14) {real, imag} */,
  {32'hbe2234b6, 32'hbe0e6fb0} /* (4, 0, 13) {real, imag} */,
  {32'hbf5e080f, 32'hbeccf712} /* (4, 0, 12) {real, imag} */,
  {32'hbf8d1905, 32'h3d3082ec} /* (4, 0, 11) {real, imag} */,
  {32'hbec04b5e, 32'h3f22b0d2} /* (4, 0, 10) {real, imag} */,
  {32'h3d006c88, 32'h3e8f9d27} /* (4, 0, 9) {real, imag} */,
  {32'h3f7ef9d8, 32'hbf45767c} /* (4, 0, 8) {real, imag} */,
  {32'h3f5996e8, 32'hbed76796} /* (4, 0, 7) {real, imag} */,
  {32'h3f5a716d, 32'hbe3a6924} /* (4, 0, 6) {real, imag} */,
  {32'h3f44096c, 32'hbe1e0815} /* (4, 0, 5) {real, imag} */,
  {32'hbd9b05a0, 32'h3f2faae8} /* (4, 0, 4) {real, imag} */,
  {32'hbd2e52a0, 32'h3e8f934e} /* (4, 0, 3) {real, imag} */,
  {32'hbe15a00b, 32'h3f389cc2} /* (4, 0, 2) {real, imag} */,
  {32'hbf1bab92, 32'h3f092017} /* (4, 0, 1) {real, imag} */,
  {32'hbf0c59de, 32'h3f162051} /* (4, 0, 0) {real, imag} */,
  {32'hbe8ab3fa, 32'hbf33eb10} /* (3, 15, 15) {real, imag} */,
  {32'h3eaf2c72, 32'hbf08622a} /* (3, 15, 14) {real, imag} */,
  {32'hbe28b414, 32'h3fa5a8c9} /* (3, 15, 13) {real, imag} */,
  {32'hbe42ee9a, 32'h3fb44e04} /* (3, 15, 12) {real, imag} */,
  {32'hbf3ecc43, 32'h3dc8f06a} /* (3, 15, 11) {real, imag} */,
  {32'h3ddb94c8, 32'h3f30bf62} /* (3, 15, 10) {real, imag} */,
  {32'hbe76f8fc, 32'hbe18c184} /* (3, 15, 9) {real, imag} */,
  {32'hbf29d2d5, 32'hbf2bc001} /* (3, 15, 8) {real, imag} */,
  {32'hbe5046a6, 32'hbf4a2994} /* (3, 15, 7) {real, imag} */,
  {32'h3ea1b065, 32'hbe138a16} /* (3, 15, 6) {real, imag} */,
  {32'hbe3bca3c, 32'h3f9a121b} /* (3, 15, 5) {real, imag} */,
  {32'h3f9fba21, 32'h3f1cd670} /* (3, 15, 4) {real, imag} */,
  {32'h3ec76719, 32'hbe92de88} /* (3, 15, 3) {real, imag} */,
  {32'hbf6bc195, 32'h3e26862a} /* (3, 15, 2) {real, imag} */,
  {32'h3e9e7976, 32'hbece91c2} /* (3, 15, 1) {real, imag} */,
  {32'h3dd2daac, 32'hbdd6d910} /* (3, 15, 0) {real, imag} */,
  {32'hbe6ee96a, 32'hbf9d9972} /* (3, 14, 15) {real, imag} */,
  {32'h3f693a0b, 32'hbe745450} /* (3, 14, 14) {real, imag} */,
  {32'h3f463444, 32'h401480dc} /* (3, 14, 13) {real, imag} */,
  {32'hbefa795c, 32'h402308d6} /* (3, 14, 12) {real, imag} */,
  {32'h3e29ceca, 32'h3f1bffd5} /* (3, 14, 11) {real, imag} */,
  {32'h3fb7ee7a, 32'h3faacbe2} /* (3, 14, 10) {real, imag} */,
  {32'h3f6b1dc2, 32'hbe103184} /* (3, 14, 9) {real, imag} */,
  {32'hbf4575a6, 32'hbf3db862} /* (3, 14, 8) {real, imag} */,
  {32'h3f332d1a, 32'hbf328fe9} /* (3, 14, 7) {real, imag} */,
  {32'h3f89f4ee, 32'hbf3f1460} /* (3, 14, 6) {real, imag} */,
  {32'h3da30ae4, 32'h3f632043} /* (3, 14, 5) {real, imag} */,
  {32'h3fa54301, 32'h3e9b018c} /* (3, 14, 4) {real, imag} */,
  {32'h3eaa4eb5, 32'hbf84a748} /* (3, 14, 3) {real, imag} */,
  {32'hbeb8432b, 32'hbf176d9c} /* (3, 14, 2) {real, imag} */,
  {32'h3fde22ba, 32'hbcb5e870} /* (3, 14, 1) {real, imag} */,
  {32'h3eac49a6, 32'h3e86cdef} /* (3, 14, 0) {real, imag} */,
  {32'hbe88df6c, 32'hbf1ac332} /* (3, 13, 15) {real, imag} */,
  {32'h40248dba, 32'h3ecfd29f} /* (3, 13, 14) {real, imag} */,
  {32'h3f4d79d9, 32'h3f85c04e} /* (3, 13, 13) {real, imag} */,
  {32'hbf9c24b9, 32'h3f0a40ca} /* (3, 13, 12) {real, imag} */,
  {32'h3f6d72b2, 32'hbf58b756} /* (3, 13, 11) {real, imag} */,
  {32'h3fb604e0, 32'hbf2b9e4c} /* (3, 13, 10) {real, imag} */,
  {32'hbf0f685a, 32'hbfa8673e} /* (3, 13, 9) {real, imag} */,
  {32'hbeb2540f, 32'h3da7e1f6} /* (3, 13, 8) {real, imag} */,
  {32'h400696f5, 32'h3f3208fe} /* (3, 13, 7) {real, imag} */,
  {32'hbf1a521a, 32'h3e6d4d90} /* (3, 13, 6) {real, imag} */,
  {32'hbfc71aa6, 32'h3e75dbe1} /* (3, 13, 5) {real, imag} */,
  {32'hbf085865, 32'hbee62132} /* (3, 13, 4) {real, imag} */,
  {32'h3f44fdaa, 32'hbd10f910} /* (3, 13, 3) {real, imag} */,
  {32'h3f0f92fc, 32'h3e099704} /* (3, 13, 2) {real, imag} */,
  {32'h3f5feb97, 32'h3f404bb8} /* (3, 13, 1) {real, imag} */,
  {32'hbf0f5639, 32'h3eaef546} /* (3, 13, 0) {real, imag} */,
  {32'hbeb2d7dc, 32'hbf0a0869} /* (3, 12, 15) {real, imag} */,
  {32'h3eba97a7, 32'h3e2def36} /* (3, 12, 14) {real, imag} */,
  {32'hbf57ca84, 32'hbea97e67} /* (3, 12, 13) {real, imag} */,
  {32'hbf627d58, 32'hbf8a4c2d} /* (3, 12, 12) {real, imag} */,
  {32'h3faaa4c6, 32'hbf93f3dc} /* (3, 12, 11) {real, imag} */,
  {32'hbf31f822, 32'hbf1bf634} /* (3, 12, 10) {real, imag} */,
  {32'hc025dcd2, 32'hbef4ff7c} /* (3, 12, 9) {real, imag} */,
  {32'hbf885a9b, 32'h3f37a20a} /* (3, 12, 8) {real, imag} */,
  {32'h3f898306, 32'h3fd575e5} /* (3, 12, 7) {real, imag} */,
  {32'h3e6b88f8, 32'h400796d0} /* (3, 12, 6) {real, imag} */,
  {32'hbf7206e8, 32'h3fadf80a} /* (3, 12, 5) {real, imag} */,
  {32'h3e9e3926, 32'hbf0c766e} /* (3, 12, 4) {real, imag} */,
  {32'h3fc6b56a, 32'hbf9b5b71} /* (3, 12, 3) {real, imag} */,
  {32'h3fd9d638, 32'hbd8ea3a8} /* (3, 12, 2) {real, imag} */,
  {32'h3f81d7a0, 32'h3f524b23} /* (3, 12, 1) {real, imag} */,
  {32'h3f18590f, 32'hbe89f79f} /* (3, 12, 0) {real, imag} */,
  {32'h3e5f3fb4, 32'hbee6c7f6} /* (3, 11, 15) {real, imag} */,
  {32'hbdd84353, 32'hbf101f09} /* (3, 11, 14) {real, imag} */,
  {32'hbfc6d120, 32'hbfd61516} /* (3, 11, 13) {real, imag} */,
  {32'h3f3805c2, 32'hbff8c328} /* (3, 11, 12) {real, imag} */,
  {32'h3e9b33eb, 32'hbfa30f52} /* (3, 11, 11) {real, imag} */,
  {32'hbf09fc4f, 32'hbea3e6f8} /* (3, 11, 10) {real, imag} */,
  {32'hbfb8c620, 32'h3e4d61ca} /* (3, 11, 9) {real, imag} */,
  {32'hbf99774b, 32'hbf4b5ab9} /* (3, 11, 8) {real, imag} */,
  {32'h3fc3737a, 32'h3f16b924} /* (3, 11, 7) {real, imag} */,
  {32'h404890c1, 32'h40192b50} /* (3, 11, 6) {real, imag} */,
  {32'h3fa7488d, 32'h4003bc2a} /* (3, 11, 5) {real, imag} */,
  {32'hbe48f41e, 32'h3fb26456} /* (3, 11, 4) {real, imag} */,
  {32'h3de31b9c, 32'h3e020175} /* (3, 11, 3) {real, imag} */,
  {32'h3f663014, 32'h3f4217f8} /* (3, 11, 2) {real, imag} */,
  {32'h3f93d43c, 32'h3e891de8} /* (3, 11, 1) {real, imag} */,
  {32'h3efb30de, 32'hbea5890a} /* (3, 11, 0) {real, imag} */,
  {32'h3ef52c31, 32'hbf3da638} /* (3, 10, 15) {real, imag} */,
  {32'h3f76cb93, 32'hbdb0b498} /* (3, 10, 14) {real, imag} */,
  {32'hbf3af132, 32'hbf43ace2} /* (3, 10, 13) {real, imag} */,
  {32'h3e106aa8, 32'hbfe86621} /* (3, 10, 12) {real, imag} */,
  {32'hbdaf5fcf, 32'hbfd18d78} /* (3, 10, 11) {real, imag} */,
  {32'h3e86a026, 32'hbfd472e6} /* (3, 10, 10) {real, imag} */,
  {32'h3ec97cda, 32'hbfa13028} /* (3, 10, 9) {real, imag} */,
  {32'h3f3cd786, 32'hbe835b6a} /* (3, 10, 8) {real, imag} */,
  {32'h3fda06b8, 32'h3ec9e9e5} /* (3, 10, 7) {real, imag} */,
  {32'h3f6fe303, 32'hbe5b90a3} /* (3, 10, 6) {real, imag} */,
  {32'h3f8f8136, 32'h3eb98274} /* (3, 10, 5) {real, imag} */,
  {32'h3f708ece, 32'h3f2b358c} /* (3, 10, 4) {real, imag} */,
  {32'h3f1d5f10, 32'hbefb579e} /* (3, 10, 3) {real, imag} */,
  {32'h3f8f02a8, 32'h3e21b98c} /* (3, 10, 2) {real, imag} */,
  {32'h3f5f7551, 32'h3edd083c} /* (3, 10, 1) {real, imag} */,
  {32'hbe9594de, 32'h3ef770bf} /* (3, 10, 0) {real, imag} */,
  {32'h3ed035cc, 32'hbfbac715} /* (3, 9, 15) {real, imag} */,
  {32'hbf5d5292, 32'hbf3728f6} /* (3, 9, 14) {real, imag} */,
  {32'hbf6c6445, 32'h3c28d420} /* (3, 9, 13) {real, imag} */,
  {32'hbf134b6b, 32'hc01bf926} /* (3, 9, 12) {real, imag} */,
  {32'h3f027c18, 32'hc00b64b9} /* (3, 9, 11) {real, imag} */,
  {32'h3fd042f8, 32'hbfe4d605} /* (3, 9, 10) {real, imag} */,
  {32'h40052cf4, 32'hc00df8cf} /* (3, 9, 9) {real, imag} */,
  {32'h3f73eb8a, 32'h3ec430f7} /* (3, 9, 8) {real, imag} */,
  {32'h3fac0153, 32'h3ed4bd3a} /* (3, 9, 7) {real, imag} */,
  {32'hbf383f96, 32'hbfba9a10} /* (3, 9, 6) {real, imag} */,
  {32'hbfd17e04, 32'hbfd2395e} /* (3, 9, 5) {real, imag} */,
  {32'hbf02fcca, 32'hbf892e6c} /* (3, 9, 4) {real, imag} */,
  {32'hbdf84e6c, 32'hbeabf526} /* (3, 9, 3) {real, imag} */,
  {32'h3fb7de8d, 32'hbebf957e} /* (3, 9, 2) {real, imag} */,
  {32'h3f96a043, 32'hbf06e0df} /* (3, 9, 1) {real, imag} */,
  {32'h3d8f95eb, 32'h3f56c565} /* (3, 9, 0) {real, imag} */,
  {32'h3fd51aaf, 32'hbdff28e2} /* (3, 8, 15) {real, imag} */,
  {32'hbdd0749f, 32'hbf45090e} /* (3, 8, 14) {real, imag} */,
  {32'hc0086eca, 32'hbdf0b494} /* (3, 8, 13) {real, imag} */,
  {32'hc000ed25, 32'hbf9bc008} /* (3, 8, 12) {real, imag} */,
  {32'hbf31b9e4, 32'hbf671a49} /* (3, 8, 11) {real, imag} */,
  {32'h3f7e6ac4, 32'hbe8f54cc} /* (3, 8, 10) {real, imag} */,
  {32'h3f8858b8, 32'hbf55987d} /* (3, 8, 9) {real, imag} */,
  {32'hbf4e905c, 32'hbf3705ce} /* (3, 8, 8) {real, imag} */,
  {32'h3d871ce8, 32'hbe9e52fd} /* (3, 8, 7) {real, imag} */,
  {32'hbfd66200, 32'h3ec0c640} /* (3, 8, 6) {real, imag} */,
  {32'hbf6f0bcc, 32'h3f2f8feb} /* (3, 8, 5) {real, imag} */,
  {32'h3ebe4f7e, 32'hbe8d69f4} /* (3, 8, 4) {real, imag} */,
  {32'h3f2b17f4, 32'hbf8ccb3d} /* (3, 8, 3) {real, imag} */,
  {32'h3fd7bdce, 32'hbececd90} /* (3, 8, 2) {real, imag} */,
  {32'h3f88d2ac, 32'h3ed8f95c} /* (3, 8, 1) {real, imag} */,
  {32'h3f68b058, 32'h3e97b013} /* (3, 8, 0) {real, imag} */,
  {32'h3fa870ea, 32'h3ffcde20} /* (3, 7, 15) {real, imag} */,
  {32'h3f9522f4, 32'h4020f5a4} /* (3, 7, 14) {real, imag} */,
  {32'hc0008905, 32'h3f477280} /* (3, 7, 13) {real, imag} */,
  {32'hc04e711e, 32'hbf40247a} /* (3, 7, 12) {real, imag} */,
  {32'hc00ad2c0, 32'hc01f2ee8} /* (3, 7, 11) {real, imag} */,
  {32'hbea66ac6, 32'hbf4594f9} /* (3, 7, 10) {real, imag} */,
  {32'hbfa82638, 32'h3fa7813a} /* (3, 7, 9) {real, imag} */,
  {32'hbfaee6a9, 32'hbe500d72} /* (3, 7, 8) {real, imag} */,
  {32'h3dd1b060, 32'hbe9d15f0} /* (3, 7, 7) {real, imag} */,
  {32'hbf95d224, 32'h3f99a5da} /* (3, 7, 6) {real, imag} */,
  {32'hbd6eef2c, 32'h4000ab89} /* (3, 7, 5) {real, imag} */,
  {32'h3fa16720, 32'h3f0ad65c} /* (3, 7, 4) {real, imag} */,
  {32'h3fd6320b, 32'hbf71cbab} /* (3, 7, 3) {real, imag} */,
  {32'h3fdc104e, 32'hbf65edc4} /* (3, 7, 2) {real, imag} */,
  {32'h3fdb1d92, 32'hbf8318ea} /* (3, 7, 1) {real, imag} */,
  {32'h3fdaa221, 32'hbf9a446c} /* (3, 7, 0) {real, imag} */,
  {32'h3e93aa27, 32'h3fec3b6b} /* (3, 6, 15) {real, imag} */,
  {32'h3f73a43c, 32'h3fe29afa} /* (3, 6, 14) {real, imag} */,
  {32'hbbae8f80, 32'hbe99916f} /* (3, 6, 13) {real, imag} */,
  {32'hbfba2bef, 32'hbe0e5454} /* (3, 6, 12) {real, imag} */,
  {32'hbf4099f4, 32'hbfbd3074} /* (3, 6, 11) {real, imag} */,
  {32'hbd2d0f88, 32'hbf363cbb} /* (3, 6, 10) {real, imag} */,
  {32'hbf19a4f7, 32'h3f06f904} /* (3, 6, 9) {real, imag} */,
  {32'h3f0b8b91, 32'hbf66abe7} /* (3, 6, 8) {real, imag} */,
  {32'h3f63ccf2, 32'hbfa87c34} /* (3, 6, 7) {real, imag} */,
  {32'hbf0c54eb, 32'h3f3ff70d} /* (3, 6, 6) {real, imag} */,
  {32'hbf14fdc1, 32'h3f1768a0} /* (3, 6, 5) {real, imag} */,
  {32'h3ebd6aef, 32'hbe433508} /* (3, 6, 4) {real, imag} */,
  {32'h3ea21a5d, 32'hbda658a6} /* (3, 6, 3) {real, imag} */,
  {32'hbea6803e, 32'hbf48ad38} /* (3, 6, 2) {real, imag} */,
  {32'hbf7c5ddd, 32'hbf80523c} /* (3, 6, 1) {real, imag} */,
  {32'h3f71fdbc, 32'hbfa94afa} /* (3, 6, 0) {real, imag} */,
  {32'h3d880957, 32'h3f99df1e} /* (3, 5, 15) {real, imag} */,
  {32'hbd950430, 32'h3fb96916} /* (3, 5, 14) {real, imag} */,
  {32'hbd43a00c, 32'hbf5f908b} /* (3, 5, 13) {real, imag} */,
  {32'hbee7949a, 32'h3e1a3d52} /* (3, 5, 12) {real, imag} */,
  {32'h3dc8977c, 32'h3ed66ba5} /* (3, 5, 11) {real, imag} */,
  {32'hbf3b8359, 32'h3ec9a849} /* (3, 5, 10) {real, imag} */,
  {32'hbe6ccacb, 32'hbdb0b4ac} /* (3, 5, 9) {real, imag} */,
  {32'h3fb58e06, 32'hbeddd51f} /* (3, 5, 8) {real, imag} */,
  {32'h3f868818, 32'hbf993e50} /* (3, 5, 7) {real, imag} */,
  {32'h3d2d5420, 32'h3f548208} /* (3, 5, 6) {real, imag} */,
  {32'h3e44ced4, 32'h3f5511fa} /* (3, 5, 5) {real, imag} */,
  {32'hbede7381, 32'hbf8c8ecf} /* (3, 5, 4) {real, imag} */,
  {32'hbf0cca08, 32'hbebf178c} /* (3, 5, 3) {real, imag} */,
  {32'h3e131094, 32'hbf18aad0} /* (3, 5, 2) {real, imag} */,
  {32'hbfd6463e, 32'hbf962a94} /* (3, 5, 1) {real, imag} */,
  {32'h3e19ea8c, 32'hbf5aa2d9} /* (3, 5, 0) {real, imag} */,
  {32'h3fada26b, 32'h3f1a5337} /* (3, 4, 15) {real, imag} */,
  {32'h3f48e533, 32'hbe800d63} /* (3, 4, 14) {real, imag} */,
  {32'hbf5a3b7a, 32'hc009941b} /* (3, 4, 13) {real, imag} */,
  {32'hbfe86c1b, 32'hbf583ce8} /* (3, 4, 12) {real, imag} */,
  {32'hbf1f3758, 32'h3e9d1d8a} /* (3, 4, 11) {real, imag} */,
  {32'h3e36bf38, 32'hbe7585b0} /* (3, 4, 10) {real, imag} */,
  {32'h3e216334, 32'hbf8ef188} /* (3, 4, 9) {real, imag} */,
  {32'hbf2ff4ef, 32'hbfac56f1} /* (3, 4, 8) {real, imag} */,
  {32'hbe40ecd6, 32'hbffdd3b6} /* (3, 4, 7) {real, imag} */,
  {32'h3ef4fe4e, 32'hbe08ae0a} /* (3, 4, 6) {real, imag} */,
  {32'h3fabc333, 32'hbe82f84e} /* (3, 4, 5) {real, imag} */,
  {32'h3d1354f8, 32'hbf3f7a1e} /* (3, 4, 4) {real, imag} */,
  {32'hbf562822, 32'hbeb1d948} /* (3, 4, 3) {real, imag} */,
  {32'h3fe0ea4b, 32'hbe8f3890} /* (3, 4, 2) {real, imag} */,
  {32'h3f179430, 32'hbfc1c1dc} /* (3, 4, 1) {real, imag} */,
  {32'h3e577a66, 32'hbe902fa6} /* (3, 4, 0) {real, imag} */,
  {32'h3eae2783, 32'hbe6ea7d8} /* (3, 3, 15) {real, imag} */,
  {32'h3f9b861e, 32'hbfdd582e} /* (3, 3, 14) {real, imag} */,
  {32'h3e93fda6, 32'hc054652b} /* (3, 3, 13) {real, imag} */,
  {32'hc03696e4, 32'hbf918fb6} /* (3, 3, 12) {real, imag} */,
  {32'hbdae2170, 32'hbf859f22} /* (3, 3, 11) {real, imag} */,
  {32'h3f9c8fe2, 32'hbf4f259a} /* (3, 3, 10) {real, imag} */,
  {32'h3d7b4a90, 32'h3ec95576} /* (3, 3, 9) {real, imag} */,
  {32'hbf46a273, 32'hbec37596} /* (3, 3, 8) {real, imag} */,
  {32'hbe000ebe, 32'hbf9868d2} /* (3, 3, 7) {real, imag} */,
  {32'hbd816022, 32'hbe7e1674} /* (3, 3, 6) {real, imag} */,
  {32'hbedde78c, 32'hbdd2a8b0} /* (3, 3, 5) {real, imag} */,
  {32'hbf026c31, 32'hbf7ac925} /* (3, 3, 4) {real, imag} */,
  {32'hbf15fd00, 32'hbf3654e4} /* (3, 3, 3) {real, imag} */,
  {32'hbed329d2, 32'hbea4cb99} /* (3, 3, 2) {real, imag} */,
  {32'hbf34e08f, 32'h3ec60f8e} /* (3, 3, 1) {real, imag} */,
  {32'hbf436138, 32'h3f98db1d} /* (3, 3, 0) {real, imag} */,
  {32'hbfff2944, 32'hbe80c2d7} /* (3, 2, 15) {real, imag} */,
  {32'hbfdf29df, 32'hbec8a61d} /* (3, 2, 14) {real, imag} */,
  {32'h3ef26ea2, 32'hbf6a04d2} /* (3, 2, 13) {real, imag} */,
  {32'hbfc4cd3e, 32'hbedb81c6} /* (3, 2, 12) {real, imag} */,
  {32'h3f97fbbe, 32'hbf36199b} /* (3, 2, 11) {real, imag} */,
  {32'h3ee105af, 32'h3f40d91b} /* (3, 2, 10) {real, imag} */,
  {32'h3f31fe3a, 32'h3f30e112} /* (3, 2, 9) {real, imag} */,
  {32'h3fc14da9, 32'h3f9911f2} /* (3, 2, 8) {real, imag} */,
  {32'h3fbb112a, 32'hbf8b11b6} /* (3, 2, 7) {real, imag} */,
  {32'hbef682fb, 32'hbfbe637e} /* (3, 2, 6) {real, imag} */,
  {32'h3f73aff0, 32'hbeb05294} /* (3, 2, 5) {real, imag} */,
  {32'h4000d7fb, 32'hbf73bbc3} /* (3, 2, 4) {real, imag} */,
  {32'h3f069f0e, 32'hbfac55a4} /* (3, 2, 3) {real, imag} */,
  {32'hbf96bd90, 32'h3e402898} /* (3, 2, 2) {real, imag} */,
  {32'hbf847fe1, 32'h3f8b179f} /* (3, 2, 1) {real, imag} */,
  {32'hbf3e00e1, 32'h3f68fae8} /* (3, 2, 0) {real, imag} */,
  {32'hbf531714, 32'h3e7bff2a} /* (3, 1, 15) {real, imag} */,
  {32'hbe9681a8, 32'h3f84cdb8} /* (3, 1, 14) {real, imag} */,
  {32'hbe953f79, 32'h3dc56ee2} /* (3, 1, 13) {real, imag} */,
  {32'hbfbd9459, 32'hbeab28cc} /* (3, 1, 12) {real, imag} */,
  {32'h3f0b1416, 32'h3f082cde} /* (3, 1, 11) {real, imag} */,
  {32'h3f89f7ca, 32'h3f8a403a} /* (3, 1, 10) {real, imag} */,
  {32'hbe4e9000, 32'h3f2cc8a6} /* (3, 1, 9) {real, imag} */,
  {32'h3f57cff2, 32'h3f8c20d4} /* (3, 1, 8) {real, imag} */,
  {32'h3f74a6c0, 32'hbf9ba6e4} /* (3, 1, 7) {real, imag} */,
  {32'hbd95c6b4, 32'hbffdfef8} /* (3, 1, 6) {real, imag} */,
  {32'h3fce6f02, 32'hc018843d} /* (3, 1, 5) {real, imag} */,
  {32'h40488770, 32'hbfa35e16} /* (3, 1, 4) {real, imag} */,
  {32'h3f293737, 32'hbe5a25e8} /* (3, 1, 3) {real, imag} */,
  {32'hbf8ef69b, 32'hbcc2c780} /* (3, 1, 2) {real, imag} */,
  {32'h3f79838a, 32'hbd06464c} /* (3, 1, 1) {real, imag} */,
  {32'h3f0a4d76, 32'h3c276180} /* (3, 1, 0) {real, imag} */,
  {32'h3e96f50b, 32'h3eacbe7a} /* (3, 0, 15) {real, imag} */,
  {32'h3e2e447a, 32'h3f3d6357} /* (3, 0, 14) {real, imag} */,
  {32'hbfd75e62, 32'h3eaeb59e} /* (3, 0, 13) {real, imag} */,
  {32'hbfe48532, 32'hbf209999} /* (3, 0, 12) {real, imag} */,
  {32'hbdb507de, 32'hbe601922} /* (3, 0, 11) {real, imag} */,
  {32'h3ead8b8a, 32'h3dc1ce38} /* (3, 0, 10) {real, imag} */,
  {32'hbfa9d2b3, 32'hbf354bbe} /* (3, 0, 9) {real, imag} */,
  {32'hbf4b1776, 32'hbc144f5c} /* (3, 0, 8) {real, imag} */,
  {32'h3f0ab1fd, 32'hbf1d7a4f} /* (3, 0, 7) {real, imag} */,
  {32'hbeb50a17, 32'hbf34648a} /* (3, 0, 6) {real, imag} */,
  {32'hbee87adb, 32'hbf42c21e} /* (3, 0, 5) {real, imag} */,
  {32'h3eb0d11d, 32'hbe95dbab} /* (3, 0, 4) {real, imag} */,
  {32'h3cd8235c, 32'hbde7e9b0} /* (3, 0, 3) {real, imag} */,
  {32'hbf480586, 32'hbf4e5bdb} /* (3, 0, 2) {real, imag} */,
  {32'h3d3f59f0, 32'hbf404374} /* (3, 0, 1) {real, imag} */,
  {32'h3ee47f0c, 32'hbebbfb0a} /* (3, 0, 0) {real, imag} */,
  {32'h3f3d3f60, 32'hbe8a8b26} /* (2, 15, 15) {real, imag} */,
  {32'h3f6ef991, 32'hbf145b34} /* (2, 15, 14) {real, imag} */,
  {32'h3dc94b89, 32'hbf1f0ebc} /* (2, 15, 13) {real, imag} */,
  {32'hbdf470ff, 32'hbf628f20} /* (2, 15, 12) {real, imag} */,
  {32'h3f2590b0, 32'hbf8f7e46} /* (2, 15, 11) {real, imag} */,
  {32'h3faa1e0e, 32'hbfde5ae0} /* (2, 15, 10) {real, imag} */,
  {32'h3e7d3989, 32'hbee177a4} /* (2, 15, 9) {real, imag} */,
  {32'h3ea92fee, 32'h3ebab11a} /* (2, 15, 8) {real, imag} */,
  {32'h3e78e48e, 32'hbf5bff3a} /* (2, 15, 7) {real, imag} */,
  {32'h3e7f0ffa, 32'hbebafdaf} /* (2, 15, 6) {real, imag} */,
  {32'hbf7f840b, 32'hbcef8758} /* (2, 15, 5) {real, imag} */,
  {32'hc025ba54, 32'hbec73604} /* (2, 15, 4) {real, imag} */,
  {32'hc0112e82, 32'h3ec73788} /* (2, 15, 3) {real, imag} */,
  {32'hbedc6fe4, 32'hbf129bde} /* (2, 15, 2) {real, imag} */,
  {32'h3c2e4990, 32'hbec59b69} /* (2, 15, 1) {real, imag} */,
  {32'hbf37a027, 32'h3fa0d8aa} /* (2, 15, 0) {real, imag} */,
  {32'h3f0d505c, 32'hbf8f6d78} /* (2, 14, 15) {real, imag} */,
  {32'h40048b71, 32'hc02db0d8} /* (2, 14, 14) {real, imag} */,
  {32'h3fbc6230, 32'hc0227609} /* (2, 14, 13) {real, imag} */,
  {32'h3fc34ba6, 32'hc0098e1a} /* (2, 14, 12) {real, imag} */,
  {32'h3f93f600, 32'hbf984dba} /* (2, 14, 11) {real, imag} */,
  {32'h40078a26, 32'hbf81e78c} /* (2, 14, 10) {real, imag} */,
  {32'h3fc29478, 32'hbe064484} /* (2, 14, 9) {real, imag} */,
  {32'h3f6429b0, 32'hbe2f6e50} /* (2, 14, 8) {real, imag} */,
  {32'hbf8bf688, 32'hbf381db6} /* (2, 14, 7) {real, imag} */,
  {32'h3f091530, 32'hbf54c23e} /* (2, 14, 6) {real, imag} */,
  {32'h3f35e1bc, 32'hc02aba28} /* (2, 14, 5) {real, imag} */,
  {32'hc00d4802, 32'hbfa89d2a} /* (2, 14, 4) {real, imag} */,
  {32'hc000ddc4, 32'h3ea7fea1} /* (2, 14, 3) {real, imag} */,
  {32'h3e729850, 32'h3e97c36e} /* (2, 14, 2) {real, imag} */,
  {32'h3e233c81, 32'h3e1c3930} /* (2, 14, 1) {real, imag} */,
  {32'hbf7e4662, 32'h3f50b3c4} /* (2, 14, 0) {real, imag} */,
  {32'hbef6b7e4, 32'hbe8a1b22} /* (2, 13, 15) {real, imag} */,
  {32'h3ee14698, 32'hbf56c201} /* (2, 13, 14) {real, imag} */,
  {32'h3ed56290, 32'hbfa8b14a} /* (2, 13, 13) {real, imag} */,
  {32'h3fcf76b8, 32'hc028eef5} /* (2, 13, 12) {real, imag} */,
  {32'h3f875d68, 32'hbf9ea0dc} /* (2, 13, 11) {real, imag} */,
  {32'h3eb371be, 32'h3f5ff8b3} /* (2, 13, 10) {real, imag} */,
  {32'h3fd99c98, 32'h3f8b886b} /* (2, 13, 9) {real, imag} */,
  {32'h3f29283c, 32'hbf5ab86c} /* (2, 13, 8) {real, imag} */,
  {32'hbfc801f3, 32'hbfefb1af} /* (2, 13, 7) {real, imag} */,
  {32'h3f536e92, 32'h3dcb5b80} /* (2, 13, 6) {real, imag} */,
  {32'h3fa95842, 32'hbfe576e8} /* (2, 13, 5) {real, imag} */,
  {32'hbf23c9dd, 32'hbfdcd4ee} /* (2, 13, 4) {real, imag} */,
  {32'hbfddcb14, 32'hbf0222cb} /* (2, 13, 3) {real, imag} */,
  {32'h3f2c5611, 32'h3f3a5486} /* (2, 13, 2) {real, imag} */,
  {32'h3fbbe7c4, 32'hbf99bb2b} /* (2, 13, 1) {real, imag} */,
  {32'h3f69e73c, 32'hbfaf0255} /* (2, 13, 0) {real, imag} */,
  {32'hbe0e9a2e, 32'h3f2f9bc4} /* (2, 12, 15) {real, imag} */,
  {32'h3e0728bc, 32'h3fe52eb8} /* (2, 12, 14) {real, imag} */,
  {32'hbec8f80b, 32'h3ef4cec5} /* (2, 12, 13) {real, imag} */,
  {32'hbf42e1ec, 32'hbfecf978} /* (2, 12, 12) {real, imag} */,
  {32'hbe79631a, 32'hbfb73436} /* (2, 12, 11) {real, imag} */,
  {32'h3e095c25, 32'hbec63502} /* (2, 12, 10) {real, imag} */,
  {32'h3f4aa780, 32'hbf03fe1c} /* (2, 12, 9) {real, imag} */,
  {32'hbe980317, 32'hbf473203} /* (2, 12, 8) {real, imag} */,
  {32'hbf1d424a, 32'hbfea0e9e} /* (2, 12, 7) {real, imag} */,
  {32'hbf462cb2, 32'hbfcc4615} /* (2, 12, 6) {real, imag} */,
  {32'hbff4d480, 32'hbff7dfdb} /* (2, 12, 5) {real, imag} */,
  {32'hbe4e183f, 32'hbfb6dff7} /* (2, 12, 4) {real, imag} */,
  {32'h3f834706, 32'hbcb46ef0} /* (2, 12, 3) {real, imag} */,
  {32'h4010b3d2, 32'hbe04970c} /* (2, 12, 2) {real, imag} */,
  {32'h3fa1ed3a, 32'hbfd49f45} /* (2, 12, 1) {real, imag} */,
  {32'h3f5060d0, 32'hbfc10a5e} /* (2, 12, 0) {real, imag} */,
  {32'h3f6ae236, 32'h3fb58516} /* (2, 11, 15) {real, imag} */,
  {32'h40286cf4, 32'h3f7a4dd9} /* (2, 11, 14) {real, imag} */,
  {32'h3f8a763c, 32'hbff775ff} /* (2, 11, 13) {real, imag} */,
  {32'hbfecc81f, 32'hbf89432a} /* (2, 11, 12) {real, imag} */,
  {32'hbfeea524, 32'hbf732857} /* (2, 11, 11) {real, imag} */,
  {32'h3fa6155d, 32'hc0040c58} /* (2, 11, 10) {real, imag} */,
  {32'h3fcf8b4f, 32'hc0288662} /* (2, 11, 9) {real, imag} */,
  {32'hbbd18320, 32'hbf4b8170} /* (2, 11, 8) {real, imag} */,
  {32'hbf85e5c1, 32'hbe8757d3} /* (2, 11, 7) {real, imag} */,
  {32'hbf714c1a, 32'hbfa0fbf2} /* (2, 11, 6) {real, imag} */,
  {32'hbfb586cd, 32'hc00be4a1} /* (2, 11, 5) {real, imag} */,
  {32'h3e553541, 32'hbf88468c} /* (2, 11, 4) {real, imag} */,
  {32'h3e8877b9, 32'h3f5fb92e} /* (2, 11, 3) {real, imag} */,
  {32'h3dd56074, 32'hbf353296} /* (2, 11, 2) {real, imag} */,
  {32'h3e9e09de, 32'hbf77e47f} /* (2, 11, 1) {real, imag} */,
  {32'hbebe7297, 32'hbf8dd525} /* (2, 11, 0) {real, imag} */,
  {32'h3eaccbbf, 32'hbed91ff7} /* (2, 10, 15) {real, imag} */,
  {32'h401a7c18, 32'hbf85ad02} /* (2, 10, 14) {real, imag} */,
  {32'h3f812054, 32'hbf01648d} /* (2, 10, 13) {real, imag} */,
  {32'hbfc6ec4c, 32'hbf588a7d} /* (2, 10, 12) {real, imag} */,
  {32'hbf7dd158, 32'h3d6be6ac} /* (2, 10, 11) {real, imag} */,
  {32'h3e96b178, 32'hbec99397} /* (2, 10, 10) {real, imag} */,
  {32'h40133a16, 32'hbfb60bf4} /* (2, 10, 9) {real, imag} */,
  {32'h3fbcb976, 32'hbf2ac954} /* (2, 10, 8) {real, imag} */,
  {32'hbf4fd2b6, 32'hbf39288c} /* (2, 10, 7) {real, imag} */,
  {32'h3e993e79, 32'hbe5fc5e4} /* (2, 10, 6) {real, imag} */,
  {32'hbf10f41e, 32'h3e858718} /* (2, 10, 5) {real, imag} */,
  {32'hbe912ae7, 32'h3f4cd5f6} /* (2, 10, 4) {real, imag} */,
  {32'h3f409e34, 32'h4007ce2e} /* (2, 10, 3) {real, imag} */,
  {32'h3f5f8a4f, 32'hbeef4d36} /* (2, 10, 2) {real, imag} */,
  {32'hbea63d6c, 32'hbf2a2b19} /* (2, 10, 1) {real, imag} */,
  {32'hbf917a51, 32'hbd761fec} /* (2, 10, 0) {real, imag} */,
  {32'hbf46059e, 32'hbea74cf4} /* (2, 9, 15) {real, imag} */,
  {32'hbf6900bf, 32'hbff2d218} /* (2, 9, 14) {real, imag} */,
  {32'hbf289c12, 32'hbf1cf427} /* (2, 9, 13) {real, imag} */,
  {32'h3df7d729, 32'h3f450d27} /* (2, 9, 12) {real, imag} */,
  {32'h3ec5a4de, 32'h3f957fd2} /* (2, 9, 11) {real, imag} */,
  {32'hbe9ab212, 32'h3ec05bc5} /* (2, 9, 10) {real, imag} */,
  {32'h3e9598de, 32'hbfb70dd0} /* (2, 9, 9) {real, imag} */,
  {32'h3eff1f64, 32'hbf265eda} /* (2, 9, 8) {real, imag} */,
  {32'hbef37d1a, 32'hc008eb2a} /* (2, 9, 7) {real, imag} */,
  {32'h4018cb4a, 32'hbea2d115} /* (2, 9, 6) {real, imag} */,
  {32'h4011ff64, 32'h3f8cb800} /* (2, 9, 5) {real, imag} */,
  {32'h3fde547b, 32'hbeffbbe3} /* (2, 9, 4) {real, imag} */,
  {32'h3ffec19e, 32'hbf4d79a7} /* (2, 9, 3) {real, imag} */,
  {32'h3f885b3c, 32'hbeb69803} /* (2, 9, 2) {real, imag} */,
  {32'h3f09c4bc, 32'hbffd1862} /* (2, 9, 1) {real, imag} */,
  {32'h3e2585fc, 32'hbf95d05a} /* (2, 9, 0) {real, imag} */,
  {32'hbfb1f350, 32'hbfb2d16e} /* (2, 8, 15) {real, imag} */,
  {32'hbfac85ca, 32'hc0870c9d} /* (2, 8, 14) {real, imag} */,
  {32'h3f413e62, 32'hc0182bdb} /* (2, 8, 13) {real, imag} */,
  {32'h4021128c, 32'hbea86ec4} /* (2, 8, 12) {real, imag} */,
  {32'h3ed6b492, 32'hbe409882} /* (2, 8, 11) {real, imag} */,
  {32'hbeba6832, 32'h3f4e3da2} /* (2, 8, 10) {real, imag} */,
  {32'hbfe2d90e, 32'hbf3720f5} /* (2, 8, 9) {real, imag} */,
  {32'hbf46e04c, 32'hbed68e1e} /* (2, 8, 8) {real, imag} */,
  {32'h3e809c6b, 32'hbf9b42ca} /* (2, 8, 7) {real, imag} */,
  {32'h3d15a0bb, 32'h3dc31738} /* (2, 8, 6) {real, imag} */,
  {32'h3f78eb60, 32'h3f23274a} /* (2, 8, 5) {real, imag} */,
  {32'h3f392ac9, 32'h3d3c83b2} /* (2, 8, 4) {real, imag} */,
  {32'h401e75e8, 32'h3ee30210} /* (2, 8, 3) {real, imag} */,
  {32'h3ff3e60b, 32'h3fb26bdc} /* (2, 8, 2) {real, imag} */,
  {32'h3f26ec78, 32'h3e9d6058} /* (2, 8, 1) {real, imag} */,
  {32'h3ef8bc20, 32'hbf1b7d36} /* (2, 8, 0) {real, imag} */,
  {32'h3f1f692a, 32'hbfbb9f74} /* (2, 7, 15) {real, imag} */,
  {32'h3f0d925f, 32'hc059a264} /* (2, 7, 14) {real, imag} */,
  {32'h40069c06, 32'hc058a4b0} /* (2, 7, 13) {real, imag} */,
  {32'h402d99bc, 32'hc0306e87} /* (2, 7, 12) {real, imag} */,
  {32'h3eb0cc24, 32'hbf770c30} /* (2, 7, 11) {real, imag} */,
  {32'hbef48374, 32'h4006fa80} /* (2, 7, 10) {real, imag} */,
  {32'hc005b92b, 32'h3f425a5d} /* (2, 7, 9) {real, imag} */,
  {32'hbf82e0b3, 32'hbf3362e6} /* (2, 7, 8) {real, imag} */,
  {32'h3e6c2620, 32'hbf23d7b2} /* (2, 7, 7) {real, imag} */,
  {32'hbf1a3437, 32'h4024c82e} /* (2, 7, 6) {real, imag} */,
  {32'hbee19b92, 32'h3fbf8aec} /* (2, 7, 5) {real, imag} */,
  {32'h3ef52a89, 32'hbec5b72f} /* (2, 7, 4) {real, imag} */,
  {32'hbde93da2, 32'hbddd4f61} /* (2, 7, 3) {real, imag} */,
  {32'hbd99d33d, 32'h3f5f8432} /* (2, 7, 2) {real, imag} */,
  {32'h3ea9e26d, 32'h3f8c21da} /* (2, 7, 1) {real, imag} */,
  {32'h3fcdc39c, 32'hbfab2b62} /* (2, 7, 0) {real, imag} */,
  {32'h3f44c8a1, 32'hbf8e2ee0} /* (2, 6, 15) {real, imag} */,
  {32'h3f28578d, 32'hbe5da825} /* (2, 6, 14) {real, imag} */,
  {32'h3f8bbdc4, 32'hc02541fd} /* (2, 6, 13) {real, imag} */,
  {32'h4000d2be, 32'hc06361d2} /* (2, 6, 12) {real, imag} */,
  {32'h3f9af807, 32'h3f1c287f} /* (2, 6, 11) {real, imag} */,
  {32'hbec2d341, 32'h4017d23f} /* (2, 6, 10) {real, imag} */,
  {32'hbfa9e33e, 32'h3f236b35} /* (2, 6, 9) {real, imag} */,
  {32'hbf440dac, 32'h3f223124} /* (2, 6, 8) {real, imag} */,
  {32'hc028ed73, 32'h3eae78b2} /* (2, 6, 7) {real, imag} */,
  {32'hbf9dbccf, 32'h3ed2f949} /* (2, 6, 6) {real, imag} */,
  {32'hbe93d0b8, 32'h3e9cec2e} /* (2, 6, 5) {real, imag} */,
  {32'h3f2f6d9a, 32'hbf12a707} /* (2, 6, 4) {real, imag} */,
  {32'hbff1759d, 32'h3d63dd04} /* (2, 6, 3) {real, imag} */,
  {32'hbe9d5050, 32'h3faaf2a0} /* (2, 6, 2) {real, imag} */,
  {32'h403f1a3d, 32'h3ec50a56} /* (2, 6, 1) {real, imag} */,
  {32'h3fcc95dc, 32'hbf3b00c9} /* (2, 6, 0) {real, imag} */,
  {32'h3df14941, 32'hbe91418e} /* (2, 5, 15) {real, imag} */,
  {32'hbcdf6df0, 32'h3f96d0ee} /* (2, 5, 14) {real, imag} */,
  {32'h3f725218, 32'hbf383c20} /* (2, 5, 13) {real, imag} */,
  {32'h3fc3ad85, 32'hbfd70cfc} /* (2, 5, 12) {real, imag} */,
  {32'h3fdc424e, 32'h3cf508a8} /* (2, 5, 11) {real, imag} */,
  {32'h3e0810d2, 32'h3ef23159} /* (2, 5, 10) {real, imag} */,
  {32'hbf9d4798, 32'h3e8f3f60} /* (2, 5, 9) {real, imag} */,
  {32'hbf0f971d, 32'hbeb76ee0} /* (2, 5, 8) {real, imag} */,
  {32'hbffb019a, 32'hbf0115a2} /* (2, 5, 7) {real, imag} */,
  {32'hbf0a8384, 32'hbdeadf84} /* (2, 5, 6) {real, imag} */,
  {32'h3f5e098f, 32'hbe9fab19} /* (2, 5, 5) {real, imag} */,
  {32'h3e45b1c8, 32'hbe384f5a} /* (2, 5, 4) {real, imag} */,
  {32'hbfb153e6, 32'h3e6e4c4f} /* (2, 5, 3) {real, imag} */,
  {32'h3e38bab2, 32'h3e6ce9df} /* (2, 5, 2) {real, imag} */,
  {32'h3fa77666, 32'hbfac91e4} /* (2, 5, 1) {real, imag} */,
  {32'h3f296bfe, 32'hbf85f914} /* (2, 5, 0) {real, imag} */,
  {32'hbfa9faa2, 32'h3f56bb23} /* (2, 4, 15) {real, imag} */,
  {32'h3f11c595, 32'h3fbf3b90} /* (2, 4, 14) {real, imag} */,
  {32'h3ff5cf3a, 32'hbe7815b9} /* (2, 4, 13) {real, imag} */,
  {32'hbe11da34, 32'h3f985e42} /* (2, 4, 12) {real, imag} */,
  {32'hbead7831, 32'hbd8499e2} /* (2, 4, 11) {real, imag} */,
  {32'hbf749106, 32'h3f1cb7ec} /* (2, 4, 10) {real, imag} */,
  {32'hbecbc41f, 32'h401c2963} /* (2, 4, 9) {real, imag} */,
  {32'hbf4b81ea, 32'h3f230090} /* (2, 4, 8) {real, imag} */,
  {32'h3e878916, 32'hbd2d91c4} /* (2, 4, 7) {real, imag} */,
  {32'h3f63f21e, 32'h3f7830da} /* (2, 4, 6) {real, imag} */,
  {32'hbed9b872, 32'h3f3cc040} /* (2, 4, 5) {real, imag} */,
  {32'h3f851c6b, 32'h3adab3f9} /* (2, 4, 4) {real, imag} */,
  {32'h3eda8ba0, 32'hc009c653} /* (2, 4, 3) {real, imag} */,
  {32'h3e85a62f, 32'hbff059ca} /* (2, 4, 2) {real, imag} */,
  {32'hbe903222, 32'hbf804332} /* (2, 4, 1) {real, imag} */,
  {32'hbeb9a2bd, 32'hbf29b50e} /* (2, 4, 0) {real, imag} */,
  {32'hbe03fac0, 32'h3f428171} /* (2, 3, 15) {real, imag} */,
  {32'h3ff3efbb, 32'h401ebee9} /* (2, 3, 14) {real, imag} */,
  {32'h3ed10b3a, 32'h4052e44b} /* (2, 3, 13) {real, imag} */,
  {32'hbfba5476, 32'h40343ae1} /* (2, 3, 12) {real, imag} */,
  {32'hbf510ee0, 32'h3fb8c11e} /* (2, 3, 11) {real, imag} */,
  {32'hbeb2ca7e, 32'h3f236644} /* (2, 3, 10) {real, imag} */,
  {32'h3f264b74, 32'h3e192775} /* (2, 3, 9) {real, imag} */,
  {32'h3dca34a8, 32'hbec5c395} /* (2, 3, 8) {real, imag} */,
  {32'h3ebbd6d7, 32'hbe5f40e0} /* (2, 3, 7) {real, imag} */,
  {32'h3f46a5ec, 32'h3f80071e} /* (2, 3, 6) {real, imag} */,
  {32'h3e93a8a4, 32'h3faa38c8} /* (2, 3, 5) {real, imag} */,
  {32'h3fb343fe, 32'hbfb97e9e} /* (2, 3, 4) {real, imag} */,
  {32'hbeaacdfa, 32'hbf9f895e} /* (2, 3, 3) {real, imag} */,
  {32'h3eb8ed89, 32'hbf73c216} /* (2, 3, 2) {real, imag} */,
  {32'hbe9aee6a, 32'hbf5665eb} /* (2, 3, 1) {real, imag} */,
  {32'hbec5ecc9, 32'h3ec3248e} /* (2, 3, 0) {real, imag} */,
  {32'h3f3c76c5, 32'h3f876e09} /* (2, 2, 15) {real, imag} */,
  {32'h3f4b402a, 32'h4007078a} /* (2, 2, 14) {real, imag} */,
  {32'hbff22585, 32'h4042dabe} /* (2, 2, 13) {real, imag} */,
  {32'hbfd737cf, 32'h3fc2adb5} /* (2, 2, 12) {real, imag} */,
  {32'hbe8c1f38, 32'hc00c0ea4} /* (2, 2, 11) {real, imag} */,
  {32'h3f9bc1d2, 32'hbfe12394} /* (2, 2, 10) {real, imag} */,
  {32'h3f5a7c9e, 32'h3ef0b2ee} /* (2, 2, 9) {real, imag} */,
  {32'h3eca07f6, 32'hbfa21018} /* (2, 2, 8) {real, imag} */,
  {32'hbd1629bf, 32'hbff28989} /* (2, 2, 7) {real, imag} */,
  {32'h3f3e5946, 32'hbf87ad3c} /* (2, 2, 6) {real, imag} */,
  {32'h400b5d49, 32'hbe119d78} /* (2, 2, 5) {real, imag} */,
  {32'h4027d2f3, 32'h3dc053b0} /* (2, 2, 4) {real, imag} */,
  {32'h3f1bfe87, 32'h3f4eb04d} /* (2, 2, 3) {real, imag} */,
  {32'hbd1e4ea0, 32'h3f422a73} /* (2, 2, 2) {real, imag} */,
  {32'hbf73c6d8, 32'hbf8c1656} /* (2, 2, 1) {real, imag} */,
  {32'h3e00abe8, 32'hbf576d2c} /* (2, 2, 0) {real, imag} */,
  {32'hbdd1f7cc, 32'h3f1f91fa} /* (2, 1, 15) {real, imag} */,
  {32'hbfcb949e, 32'h3fe20bc6} /* (2, 1, 14) {real, imag} */,
  {32'hc04617fd, 32'h3f831d86} /* (2, 1, 13) {real, imag} */,
  {32'h3ea3b0f7, 32'hbd5c40a8} /* (2, 1, 12) {real, imag} */,
  {32'hbcff2f90, 32'hc07d11e2} /* (2, 1, 11) {real, imag} */,
  {32'hbf90ac0e, 32'hbfa9e774} /* (2, 1, 10) {real, imag} */,
  {32'h3e88e8a8, 32'h4017ba9e} /* (2, 1, 9) {real, imag} */,
  {32'hbd953b05, 32'h3de5af88} /* (2, 1, 8) {real, imag} */,
  {32'h3f7bc2c2, 32'hc0568383} /* (2, 1, 7) {real, imag} */,
  {32'h3f8a3fc2, 32'hc0414c94} /* (2, 1, 6) {real, imag} */,
  {32'h3ed018e8, 32'hbf1dd222} /* (2, 1, 5) {real, imag} */,
  {32'h3fc48ba7, 32'hbf5199ed} /* (2, 1, 4) {real, imag} */,
  {32'h3f5f87fa, 32'hbf3f418f} /* (2, 1, 3) {real, imag} */,
  {32'hbf6642b3, 32'h3d23cdae} /* (2, 1, 2) {real, imag} */,
  {32'h3db04f13, 32'hc01c7438} /* (2, 1, 1) {real, imag} */,
  {32'h3e40d054, 32'hc009df71} /* (2, 1, 0) {real, imag} */,
  {32'hbdba27ea, 32'hbde48640} /* (2, 0, 15) {real, imag} */,
  {32'hbf3ad4d4, 32'h3ebeed98} /* (2, 0, 14) {real, imag} */,
  {32'hbfaa3c5c, 32'hbe51540d} /* (2, 0, 13) {real, imag} */,
  {32'h3fab45ce, 32'hbf4c18ca} /* (2, 0, 12) {real, imag} */,
  {32'h3fa752e8, 32'hbfce99c8} /* (2, 0, 11) {real, imag} */,
  {32'hbe834a94, 32'hbfa70f20} /* (2, 0, 10) {real, imag} */,
  {32'hbed9a0ba, 32'h3fa3f402} /* (2, 0, 9) {real, imag} */,
  {32'hbf5fdc2a, 32'h3ff2771c} /* (2, 0, 8) {real, imag} */,
  {32'h3f47fd20, 32'hbfa66fcf} /* (2, 0, 7) {real, imag} */,
  {32'h3f74ed57, 32'hbf570731} /* (2, 0, 6) {real, imag} */,
  {32'hbf10af66, 32'h3faaa620} /* (2, 0, 5) {real, imag} */,
  {32'hbf95dc2f, 32'hbe47519d} /* (2, 0, 4) {real, imag} */,
  {32'hbf3ef01a, 32'hbd13c91c} /* (2, 0, 3) {real, imag} */,
  {32'hbf091c06, 32'hbed15047} /* (2, 0, 2) {real, imag} */,
  {32'hbeb1d168, 32'hbf90b1e0} /* (2, 0, 1) {real, imag} */,
  {32'hbf1aca4c, 32'hbe7eb2b3} /* (2, 0, 0) {real, imag} */,
  {32'hbddce957, 32'h3fd03ae4} /* (1, 15, 15) {real, imag} */,
  {32'hbf42cbd1, 32'h3f144999} /* (1, 15, 14) {real, imag} */,
  {32'hbe5b6e19, 32'hbf02a37a} /* (1, 15, 13) {real, imag} */,
  {32'hbd860cf0, 32'h3ee06bd9} /* (1, 15, 12) {real, imag} */,
  {32'h3d31f09c, 32'h3e413c9f} /* (1, 15, 11) {real, imag} */,
  {32'hbdcb8f34, 32'hbfd6470c} /* (1, 15, 10) {real, imag} */,
  {32'hbe5fd664, 32'hbfea310e} /* (1, 15, 9) {real, imag} */,
  {32'h3fc865f2, 32'hc02e56dc} /* (1, 15, 8) {real, imag} */,
  {32'h3f85fb02, 32'hbf06d42b} /* (1, 15, 7) {real, imag} */,
  {32'hbe8c1c14, 32'hbe0e0b54} /* (1, 15, 6) {real, imag} */,
  {32'hbf64c87c, 32'hbdb61c14} /* (1, 15, 5) {real, imag} */,
  {32'h3de3c068, 32'h3fa165aa} /* (1, 15, 4) {real, imag} */,
  {32'hbdddb576, 32'h3f9e336e} /* (1, 15, 3) {real, imag} */,
  {32'hbe893456, 32'h3f4f3cec} /* (1, 15, 2) {real, imag} */,
  {32'hbf8afe46, 32'h3dd4a2dc} /* (1, 15, 1) {real, imag} */,
  {32'hbf5d92f6, 32'h3eeb98ec} /* (1, 15, 0) {real, imag} */,
  {32'hbe413a1a, 32'h3f975b16} /* (1, 14, 15) {real, imag} */,
  {32'hc009584c, 32'h3fe3bf25} /* (1, 14, 14) {real, imag} */,
  {32'hbfde3372, 32'h3fe39f05} /* (1, 14, 13) {real, imag} */,
  {32'hbf45b899, 32'h3e2c5798} /* (1, 14, 12) {real, imag} */,
  {32'h3f724c80, 32'hbe4476e6} /* (1, 14, 11) {real, imag} */,
  {32'h3f9a23d8, 32'hbf4494f5} /* (1, 14, 10) {real, imag} */,
  {32'hbe4266f2, 32'hbd4efc00} /* (1, 14, 9) {real, imag} */,
  {32'h3fd34c82, 32'hc010338a} /* (1, 14, 8) {real, imag} */,
  {32'h3f7564ca, 32'h3f6b1f93} /* (1, 14, 7) {real, imag} */,
  {32'hbf69e52e, 32'h3f86a9e4} /* (1, 14, 6) {real, imag} */,
  {32'hc0183169, 32'h3f0e3f5a} /* (1, 14, 5) {real, imag} */,
  {32'h3f89f6f7, 32'h3f721139} /* (1, 14, 4) {real, imag} */,
  {32'h3f059cb4, 32'h3ecb36dc} /* (1, 14, 3) {real, imag} */,
  {32'hbda9c35a, 32'h3d2108f8} /* (1, 14, 2) {real, imag} */,
  {32'hbeb38c7f, 32'hbfa24976} /* (1, 14, 1) {real, imag} */,
  {32'hbe0f180d, 32'hbfdf6edc} /* (1, 14, 0) {real, imag} */,
  {32'h3fbcd73e, 32'h3f48610e} /* (1, 13, 15) {real, imag} */,
  {32'hbf673ff8, 32'h403da6f0} /* (1, 13, 14) {real, imag} */,
  {32'hbf944b2a, 32'h3f81d694} /* (1, 13, 13) {real, imag} */,
  {32'hbeee4a5a, 32'hbfe96f10} /* (1, 13, 12) {real, imag} */,
  {32'h3e1be196, 32'h3ddd8f3a} /* (1, 13, 11) {real, imag} */,
  {32'hbed04fa6, 32'h3f50ec2c} /* (1, 13, 10) {real, imag} */,
  {32'hbfffae79, 32'h4009005b} /* (1, 13, 9) {real, imag} */,
  {32'h3e8d7b95, 32'hbf351512} /* (1, 13, 8) {real, imag} */,
  {32'hbea223e5, 32'hbd989158} /* (1, 13, 7) {real, imag} */,
  {32'hbfa7b48b, 32'h3ef0f244} /* (1, 13, 6) {real, imag} */,
  {32'hbf1ea63c, 32'h3ee19af9} /* (1, 13, 5) {real, imag} */,
  {32'h3f07de0a, 32'h3fd333a6} /* (1, 13, 4) {real, imag} */,
  {32'h3fa1fc63, 32'hbf93e868} /* (1, 13, 3) {real, imag} */,
  {32'hbdd46489, 32'hbf247e6e} /* (1, 13, 2) {real, imag} */,
  {32'h3e9fbdae, 32'h3f22a5fc} /* (1, 13, 1) {real, imag} */,
  {32'h3fc57d38, 32'hbeb18521} /* (1, 13, 0) {real, imag} */,
  {32'h3ea33948, 32'h3f88287c} /* (1, 12, 15) {real, imag} */,
  {32'h3e55eb90, 32'h3dc5c570} /* (1, 12, 14) {real, imag} */,
  {32'h3facad40, 32'hc03f3e93} /* (1, 12, 13) {real, imag} */,
  {32'h3fb24a14, 32'hbf1113ce} /* (1, 12, 12) {real, imag} */,
  {32'hbf632b24, 32'h3f983af8} /* (1, 12, 11) {real, imag} */,
  {32'hbf7bcb4e, 32'h3fcb01c0} /* (1, 12, 10) {real, imag} */,
  {32'hc00c5c1d, 32'h401c9bdd} /* (1, 12, 9) {real, imag} */,
  {32'hbfd9ee9e, 32'h3ea9e262} /* (1, 12, 8) {real, imag} */,
  {32'hbfdaaaaf, 32'hbea987bd} /* (1, 12, 7) {real, imag} */,
  {32'hbef3a57c, 32'hbf69c163} /* (1, 12, 6) {real, imag} */,
  {32'h3fa75c05, 32'hbfa0d6ee} /* (1, 12, 5) {real, imag} */,
  {32'hbf2a2c50, 32'h3f8d57b0} /* (1, 12, 4) {real, imag} */,
  {32'h3d4934d0, 32'hbf1e695c} /* (1, 12, 3) {real, imag} */,
  {32'h3f057ba2, 32'hbfb98222} /* (1, 12, 2) {real, imag} */,
  {32'h3f9c89ff, 32'h3f8acefe} /* (1, 12, 1) {real, imag} */,
  {32'h3ea02d2b, 32'h3f80fc2e} /* (1, 12, 0) {real, imag} */,
  {32'hbf28f806, 32'hbf2b9774} /* (1, 11, 15) {real, imag} */,
  {32'hbcef92ac, 32'hbedca1e1} /* (1, 11, 14) {real, imag} */,
  {32'h4021334c, 32'hbf56f80e} /* (1, 11, 13) {real, imag} */,
  {32'h40445e15, 32'h3e36d53c} /* (1, 11, 12) {real, imag} */,
  {32'h3fb7bedc, 32'h3fad558d} /* (1, 11, 11) {real, imag} */,
  {32'hbec4ce80, 32'h3f8f9a9a} /* (1, 11, 10) {real, imag} */,
  {32'hbf678232, 32'h4023a585} /* (1, 11, 9) {real, imag} */,
  {32'h3f920e18, 32'h3ff3a9f5} /* (1, 11, 8) {real, imag} */,
  {32'hbefc6f68, 32'h3fc325e1} /* (1, 11, 7) {real, imag} */,
  {32'hbf60988e, 32'hbf0b4873} /* (1, 11, 6) {real, imag} */,
  {32'hbf01274e, 32'hbfc29ebe} /* (1, 11, 5) {real, imag} */,
  {32'hbf8d43c9, 32'hbe54f306} /* (1, 11, 4) {real, imag} */,
  {32'hbfe6e698, 32'hbf0afcb5} /* (1, 11, 3) {real, imag} */,
  {32'hbf9ccab5, 32'h3e6296e8} /* (1, 11, 2) {real, imag} */,
  {32'hbdcae7a0, 32'h3f90697c} /* (1, 11, 1) {real, imag} */,
  {32'h3d887886, 32'hbd57f890} /* (1, 11, 0) {real, imag} */,
  {32'h3efdb21c, 32'hbebfe6ec} /* (1, 10, 15) {real, imag} */,
  {32'h3f160f74, 32'h3fb1aa8a} /* (1, 10, 14) {real, imag} */,
  {32'h3ea1c956, 32'h3f38f50d} /* (1, 10, 13) {real, imag} */,
  {32'h3feeabf2, 32'h3f171a3a} /* (1, 10, 12) {real, imag} */,
  {32'h4011acb6, 32'h3e7b563c} /* (1, 10, 11) {real, imag} */,
  {32'h3f926d24, 32'hbf8e3fe7} /* (1, 10, 10) {real, imag} */,
  {32'hbfe7e2c0, 32'h3ea324e6} /* (1, 10, 9) {real, imag} */,
  {32'hbfb08e42, 32'h3fad3dec} /* (1, 10, 8) {real, imag} */,
  {32'hbf41c3f2, 32'h404bb998} /* (1, 10, 7) {real, imag} */,
  {32'hbecd34bb, 32'h3f6132b2} /* (1, 10, 6) {real, imag} */,
  {32'hbff47b57, 32'hbf9501bc} /* (1, 10, 5) {real, imag} */,
  {32'hc02550fc, 32'hbf356682} /* (1, 10, 4) {real, imag} */,
  {32'hc0292071, 32'h3e0c7555} /* (1, 10, 3) {real, imag} */,
  {32'hc059132c, 32'h3f6fefbd} /* (1, 10, 2) {real, imag} */,
  {32'hc001f86e, 32'h3f980441} /* (1, 10, 1) {real, imag} */,
  {32'h3ef0e84e, 32'h3e8e62aa} /* (1, 10, 0) {real, imag} */,
  {32'h3f0986c6, 32'hbe3553a3} /* (1, 9, 15) {real, imag} */,
  {32'hbdf71211, 32'h3eee68df} /* (1, 9, 14) {real, imag} */,
  {32'h3e130b15, 32'hbeb82619} /* (1, 9, 13) {real, imag} */,
  {32'h3fd90d1e, 32'h3fb3a6f6} /* (1, 9, 12) {real, imag} */,
  {32'h3e75f1a6, 32'h3fd489ab} /* (1, 9, 11) {real, imag} */,
  {32'h3fe993f5, 32'hbf4423af} /* (1, 9, 10) {real, imag} */,
  {32'hbfc23180, 32'hc00062c8} /* (1, 9, 9) {real, imag} */,
  {32'hc013fada, 32'hbfaeb4b2} /* (1, 9, 8) {real, imag} */,
  {32'hbe643e80, 32'hbf0e7f22} /* (1, 9, 7) {real, imag} */,
  {32'h3f564217, 32'hbf983905} /* (1, 9, 6) {real, imag} */,
  {32'h3e3a3768, 32'hc01bb2e6} /* (1, 9, 5) {real, imag} */,
  {32'h3d878de8, 32'hbfc198d9} /* (1, 9, 4) {real, imag} */,
  {32'h3eb3be7e, 32'hbe43688d} /* (1, 9, 3) {real, imag} */,
  {32'hbf7900fb, 32'h3f91dd0c} /* (1, 9, 2) {real, imag} */,
  {32'hbfda3832, 32'h3f0459ee} /* (1, 9, 1) {real, imag} */,
  {32'h3f780130, 32'h3f0033da} /* (1, 9, 0) {real, imag} */,
  {32'hbf00f561, 32'hc005a3cc} /* (1, 8, 15) {real, imag} */,
  {32'hbee9ee98, 32'hbf90ecf0} /* (1, 8, 14) {real, imag} */,
  {32'hbf232305, 32'h3ecaad65} /* (1, 8, 13) {real, imag} */,
  {32'hbe18a1f4, 32'h3ec48946} /* (1, 8, 12) {real, imag} */,
  {32'hbb1c6980, 32'h3faed098} /* (1, 8, 11) {real, imag} */,
  {32'h3fce115a, 32'hbf14bf69} /* (1, 8, 10) {real, imag} */,
  {32'h3ebfd930, 32'hbf49e5ee} /* (1, 8, 9) {real, imag} */,
  {32'hbf741c0a, 32'h3e077018} /* (1, 8, 8) {real, imag} */,
  {32'hbfa6229a, 32'hbfe779c6} /* (1, 8, 7) {real, imag} */,
  {32'hbf4c3313, 32'hc04e4f34} /* (1, 8, 6) {real, imag} */,
  {32'h3e41dda8, 32'hc0524e34} /* (1, 8, 5) {real, imag} */,
  {32'h402f61ae, 32'hbfd7767d} /* (1, 8, 4) {real, imag} */,
  {32'h401040dc, 32'hbfaf4004} /* (1, 8, 3) {real, imag} */,
  {32'h3f7493df, 32'h3f4378d3} /* (1, 8, 2) {real, imag} */,
  {32'hbf5d1100, 32'h3eedafa0} /* (1, 8, 1) {real, imag} */,
  {32'h3e953955, 32'hbfd3b40c} /* (1, 8, 0) {real, imag} */,
  {32'hbf5a8342, 32'hbfcd61ba} /* (1, 7, 15) {real, imag} */,
  {32'hbf9726e0, 32'hbf7d712d} /* (1, 7, 14) {real, imag} */,
  {32'hbefa222c, 32'hbf9111ca} /* (1, 7, 13) {real, imag} */,
  {32'hbf9d9d2e, 32'h3fbbbbe6} /* (1, 7, 12) {real, imag} */,
  {32'hbe7bc3c4, 32'h403a34b8} /* (1, 7, 11) {real, imag} */,
  {32'h3f407460, 32'hbd91f768} /* (1, 7, 10) {real, imag} */,
  {32'h3f78b51e, 32'hbf033e1c} /* (1, 7, 9) {real, imag} */,
  {32'h3f480d34, 32'h3e9a843a} /* (1, 7, 8) {real, imag} */,
  {32'hbeadd4ee, 32'h3f056ec6} /* (1, 7, 7) {real, imag} */,
  {32'hbfc6ffc1, 32'h3ee97d58} /* (1, 7, 6) {real, imag} */,
  {32'hbe774fb4, 32'hbddadee8} /* (1, 7, 5) {real, imag} */,
  {32'h3fa7a2a0, 32'h3f009a3e} /* (1, 7, 4) {real, imag} */,
  {32'hbc2232c0, 32'h3f3a411f} /* (1, 7, 3) {real, imag} */,
  {32'hbf0520bd, 32'h3fa25111} /* (1, 7, 2) {real, imag} */,
  {32'h3f9a9836, 32'hbee835b3} /* (1, 7, 1) {real, imag} */,
  {32'h3fce3dee, 32'hbfda9158} /* (1, 7, 0) {real, imag} */,
  {32'hbea186a0, 32'hbf37d958} /* (1, 6, 15) {real, imag} */,
  {32'hbf8d372a, 32'h3f8ef550} /* (1, 6, 14) {real, imag} */,
  {32'hbe9b78da, 32'h3fb28eda} /* (1, 6, 13) {real, imag} */,
  {32'h3f807bd7, 32'h40001b78} /* (1, 6, 12) {real, imag} */,
  {32'h3df818dc, 32'h3fdacce6} /* (1, 6, 11) {real, imag} */,
  {32'h3fca218c, 32'h3f173a58} /* (1, 6, 10) {real, imag} */,
  {32'h3e984551, 32'h40245570} /* (1, 6, 9) {real, imag} */,
  {32'h3ed972ea, 32'h3f012477} /* (1, 6, 8) {real, imag} */,
  {32'h3ff149b7, 32'h40187c10} /* (1, 6, 7) {real, imag} */,
  {32'hbf9832c5, 32'h3f947108} /* (1, 6, 6) {real, imag} */,
  {32'hc015bb08, 32'h3fc0a27f} /* (1, 6, 5) {real, imag} */,
  {32'hbf2c0256, 32'h3f87b2b8} /* (1, 6, 4) {real, imag} */,
  {32'h3ed012a6, 32'h3fdde004} /* (1, 6, 3) {real, imag} */,
  {32'hbf86cdec, 32'h3fc31053} /* (1, 6, 2) {real, imag} */,
  {32'h3ee5d73a, 32'hbfc7646c} /* (1, 6, 1) {real, imag} */,
  {32'h3f9d8e4e, 32'hbee7885e} /* (1, 6, 0) {real, imag} */,
  {32'hbebd6383, 32'h3fc82aca} /* (1, 5, 15) {real, imag} */,
  {32'hbfb1667b, 32'h40166ccc} /* (1, 5, 14) {real, imag} */,
  {32'hbee2d63a, 32'h3e8ee6ca} /* (1, 5, 13) {real, imag} */,
  {32'h3f346c24, 32'hbde16b68} /* (1, 5, 12) {real, imag} */,
  {32'h3f4dc4a0, 32'hbf194376} /* (1, 5, 11) {real, imag} */,
  {32'h3ff97554, 32'hbf35ddf3} /* (1, 5, 10) {real, imag} */,
  {32'hbf81171e, 32'h3f7ea2ca} /* (1, 5, 9) {real, imag} */,
  {32'h3f630c40, 32'hbfa3e505} /* (1, 5, 8) {real, imag} */,
  {32'h3e57178f, 32'h3ed6344c} /* (1, 5, 7) {real, imag} */,
  {32'hc0189f20, 32'hbc81ccf0} /* (1, 5, 6) {real, imag} */,
  {32'hc0778c04, 32'h3f3b23da} /* (1, 5, 5) {real, imag} */,
  {32'hbfda30be, 32'h3fc649f7} /* (1, 5, 4) {real, imag} */,
  {32'h3fad6898, 32'h401504a8} /* (1, 5, 3) {real, imag} */,
  {32'h4006c8a8, 32'h4007990e} /* (1, 5, 2) {real, imag} */,
  {32'h4064966f, 32'hbeaa8a0b} /* (1, 5, 1) {real, imag} */,
  {32'h3f84cfe6, 32'hbe65fafc} /* (1, 5, 0) {real, imag} */,
  {32'hbf47728c, 32'h3fb9d202} /* (1, 4, 15) {real, imag} */,
  {32'hc0247742, 32'h3f62b116} /* (1, 4, 14) {real, imag} */,
  {32'hbfaaea25, 32'hbeb32e60} /* (1, 4, 13) {real, imag} */,
  {32'h3d900a16, 32'h3eb86dd2} /* (1, 4, 12) {real, imag} */,
  {32'h3e29486b, 32'hc0031728} /* (1, 4, 11) {real, imag} */,
  {32'h401f367e, 32'hc03ae798} /* (1, 4, 10) {real, imag} */,
  {32'hbfa5d034, 32'hbfbaac40} /* (1, 4, 9) {real, imag} */,
  {32'h3fa91b54, 32'h3f1dfd8b} /* (1, 4, 8) {real, imag} */,
  {32'h3f4a4a37, 32'h3fe1efb7} /* (1, 4, 7) {real, imag} */,
  {32'hc03a096c, 32'h3f430522} /* (1, 4, 6) {real, imag} */,
  {32'hc0706b1a, 32'hbff08703} /* (1, 4, 5) {real, imag} */,
  {32'hc01ea482, 32'h3f6a4456} /* (1, 4, 4) {real, imag} */,
  {32'h3e982c5e, 32'h4069e406} /* (1, 4, 3) {real, imag} */,
  {32'h3fd1edfa, 32'h3fe8379d} /* (1, 4, 2) {real, imag} */,
  {32'h3fd0d09d, 32'h3f3de33e} /* (1, 4, 1) {real, imag} */,
  {32'hbd61b45c, 32'h3f1b1cb8} /* (1, 4, 0) {real, imag} */,
  {32'h3de90ae0, 32'h3f05f7a9} /* (1, 3, 15) {real, imag} */,
  {32'hbeba578e, 32'hbf49f18c} /* (1, 3, 14) {real, imag} */,
  {32'h3fae5c3a, 32'hbc39f850} /* (1, 3, 13) {real, imag} */,
  {32'h3fd82592, 32'h3f99ad40} /* (1, 3, 12) {real, imag} */,
  {32'h3e50e37a, 32'hbfd98e87} /* (1, 3, 11) {real, imag} */,
  {32'h3fe03dfd, 32'hbf83d670} /* (1, 3, 10) {real, imag} */,
  {32'h3f4055d2, 32'hbf35c02a} /* (1, 3, 9) {real, imag} */,
  {32'h3f2f355d, 32'h3fb5d758} /* (1, 3, 8) {real, imag} */,
  {32'h3eb5d4bf, 32'h3fb424e2} /* (1, 3, 7) {real, imag} */,
  {32'hc01022d8, 32'h3f9c29c1} /* (1, 3, 6) {real, imag} */,
  {32'hc04e5738, 32'hbf6aeb24} /* (1, 3, 5) {real, imag} */,
  {32'h3d08533c, 32'h3fb2841b} /* (1, 3, 4) {real, imag} */,
  {32'h3f8d607c, 32'h405a6f42} /* (1, 3, 3) {real, imag} */,
  {32'h3d2e2468, 32'h3ed456b4} /* (1, 3, 2) {real, imag} */,
  {32'hbf4401e8, 32'h3e9aa051} /* (1, 3, 1) {real, imag} */,
  {32'h3f33a094, 32'h3ee9fe71} /* (1, 3, 0) {real, imag} */,
  {32'h3f110423, 32'h3fe7ae2e} /* (1, 2, 15) {real, imag} */,
  {32'h3fdf0243, 32'h3eb6c472} /* (1, 2, 14) {real, imag} */,
  {32'h4036c0f5, 32'hbe5f7911} /* (1, 2, 13) {real, imag} */,
  {32'h400d7868, 32'hbe4d36d9} /* (1, 2, 12) {real, imag} */,
  {32'h3f7995ae, 32'hbe36e6c6} /* (1, 2, 11) {real, imag} */,
  {32'h3fcf91e6, 32'h3ff6da95} /* (1, 2, 10) {real, imag} */,
  {32'h3fc5c834, 32'hbe445d59} /* (1, 2, 9) {real, imag} */,
  {32'h3f872a9a, 32'h3dae501e} /* (1, 2, 8) {real, imag} */,
  {32'h3ecc2a27, 32'h3d517e6c} /* (1, 2, 7) {real, imag} */,
  {32'hc01745b6, 32'hbf9dab3c} /* (1, 2, 6) {real, imag} */,
  {32'hbfdaf8fb, 32'hc01ddeba} /* (1, 2, 5) {real, imag} */,
  {32'hbf95475a, 32'hbe43aebe} /* (1, 2, 4) {real, imag} */,
  {32'hbed527d8, 32'h3f39d1ae} /* (1, 2, 3) {real, imag} */,
  {32'hbf0d90be, 32'h3e5c9612} /* (1, 2, 2) {real, imag} */,
  {32'hbee66807, 32'h3f8d5e84} /* (1, 2, 1) {real, imag} */,
  {32'h3f986950, 32'h3f1f3f7e} /* (1, 2, 0) {real, imag} */,
  {32'hbf38f11a, 32'h3fc6b26b} /* (1, 1, 15) {real, imag} */,
  {32'hbf7cf252, 32'h3ecfadd8} /* (1, 1, 14) {real, imag} */,
  {32'h3f6c896d, 32'hbedec9c8} /* (1, 1, 13) {real, imag} */,
  {32'h3fa3a264, 32'hbf23b86b} /* (1, 1, 12) {real, imag} */,
  {32'h3f1c720b, 32'h3f3d991f} /* (1, 1, 11) {real, imag} */,
  {32'hbe6f99fe, 32'h3f98758c} /* (1, 1, 10) {real, imag} */,
  {32'h3d42d0d0, 32'h3f801163} /* (1, 1, 9) {real, imag} */,
  {32'h3e547750, 32'h3fb80e2a} /* (1, 1, 8) {real, imag} */,
  {32'hbf76c161, 32'h3f2260a9} /* (1, 1, 7) {real, imag} */,
  {32'hbfa8e45e, 32'hbff96ef7} /* (1, 1, 6) {real, imag} */,
  {32'hbf6145fc, 32'hc0330d92} /* (1, 1, 5) {real, imag} */,
  {32'hc084ce48, 32'hbe0d8c36} /* (1, 1, 4) {real, imag} */,
  {32'hbfec5327, 32'hbef0697c} /* (1, 1, 3) {real, imag} */,
  {32'h3f795920, 32'hbeb53774} /* (1, 1, 2) {real, imag} */,
  {32'h3f4bc28c, 32'h3f61eccc} /* (1, 1, 1) {real, imag} */,
  {32'h3e13638d, 32'h3f625a7a} /* (1, 1, 0) {real, imag} */,
  {32'hbeedf410, 32'h3f842654} /* (1, 0, 15) {real, imag} */,
  {32'hbdd92efc, 32'hbd7a9a00} /* (1, 0, 14) {real, imag} */,
  {32'h3f187760, 32'hbf0a8f11} /* (1, 0, 13) {real, imag} */,
  {32'h3f9d39df, 32'h3eaa4ace} /* (1, 0, 12) {real, imag} */,
  {32'h3e0e545a, 32'h3f2a52ac} /* (1, 0, 11) {real, imag} */,
  {32'hbfad071a, 32'h3e6ae869} /* (1, 0, 10) {real, imag} */,
  {32'hbf8cb960, 32'h3e99a2a2} /* (1, 0, 9) {real, imag} */,
  {32'hbeccabf4, 32'h3dd05aea} /* (1, 0, 8) {real, imag} */,
  {32'hbf73290e, 32'h3ebf1209} /* (1, 0, 7) {real, imag} */,
  {32'hbe137076, 32'hbfada07c} /* (1, 0, 6) {real, imag} */,
  {32'hbece395c, 32'hbffb62ea} /* (1, 0, 5) {real, imag} */,
  {32'hbf7a0334, 32'h3e8742fe} /* (1, 0, 4) {real, imag} */,
  {32'hbdf7fe7e, 32'h3f16ce5a} /* (1, 0, 3) {real, imag} */,
  {32'h3f46f216, 32'h3de21ece} /* (1, 0, 2) {real, imag} */,
  {32'h3eeb609f, 32'h3e281bb3} /* (1, 0, 1) {real, imag} */,
  {32'hbf0a98bd, 32'h3f30228c} /* (1, 0, 0) {real, imag} */,
  {32'h3ebc6776, 32'h00000000} /* (0, 15, 15) {real, imag} */,
  {32'hbf39f7a8, 32'h00000000} /* (0, 15, 14) {real, imag} */,
  {32'hbf06d77d, 32'h00000000} /* (0, 15, 13) {real, imag} */,
  {32'h3f4c7fd9, 32'h00000000} /* (0, 15, 12) {real, imag} */,
  {32'h400df503, 32'h00000000} /* (0, 15, 11) {real, imag} */,
  {32'hbfa0ee86, 32'h00000000} /* (0, 15, 10) {real, imag} */,
  {32'hc0316ac2, 32'h00000000} /* (0, 15, 9) {real, imag} */,
  {32'hc025d500, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'h3eb4a3ec, 32'h00000000} /* (0, 15, 7) {real, imag} */,
  {32'h3f4d52bf, 32'h00000000} /* (0, 15, 6) {real, imag} */,
  {32'hba94b000, 32'h00000000} /* (0, 15, 5) {real, imag} */,
  {32'hbf87dbf4, 32'h00000000} /* (0, 15, 4) {real, imag} */,
  {32'hbfb24759, 32'h00000000} /* (0, 15, 3) {real, imag} */,
  {32'hbfc81756, 32'h00000000} /* (0, 15, 2) {real, imag} */,
  {32'hbe3f5286, 32'h00000000} /* (0, 15, 1) {real, imag} */,
  {32'h3ecb35fc, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h400657d1, 32'h00000000} /* (0, 14, 15) {real, imag} */,
  {32'hbf11789e, 32'h00000000} /* (0, 14, 14) {real, imag} */,
  {32'hc018f254, 32'h00000000} /* (0, 14, 13) {real, imag} */,
  {32'hbeccf96e, 32'h00000000} /* (0, 14, 12) {real, imag} */,
  {32'h403668fa, 32'h00000000} /* (0, 14, 11) {real, imag} */,
  {32'hc06a118d, 32'h00000000} /* (0, 14, 10) {real, imag} */,
  {32'hc081d23c, 32'h00000000} /* (0, 14, 9) {real, imag} */,
  {32'hbff27d2e, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'h3fbac10a, 32'h00000000} /* (0, 14, 7) {real, imag} */,
  {32'h4058fd26, 32'h00000000} /* (0, 14, 6) {real, imag} */,
  {32'h3fc4d543, 32'h00000000} /* (0, 14, 5) {real, imag} */,
  {32'hbfaf6e38, 32'h00000000} /* (0, 14, 4) {real, imag} */,
  {32'hc03ac852, 32'h00000000} /* (0, 14, 3) {real, imag} */,
  {32'hc09ae35f, 32'h00000000} /* (0, 14, 2) {real, imag} */,
  {32'hbf51b765, 32'h00000000} /* (0, 14, 1) {real, imag} */,
  {32'h400af674, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h3e4076fa, 32'h00000000} /* (0, 13, 15) {real, imag} */,
  {32'hbf957e96, 32'h00000000} /* (0, 13, 14) {real, imag} */,
  {32'hc00c65b6, 32'h00000000} /* (0, 13, 13) {real, imag} */,
  {32'hbf278de6, 32'h00000000} /* (0, 13, 12) {real, imag} */,
  {32'h3db4a63e, 32'h00000000} /* (0, 13, 11) {real, imag} */,
  {32'hbf9a4b9a, 32'h00000000} /* (0, 13, 10) {real, imag} */,
  {32'hbeb6af92, 32'h00000000} /* (0, 13, 9) {real, imag} */,
  {32'h3f28b63e, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'h3fb4e620, 32'h00000000} /* (0, 13, 7) {real, imag} */,
  {32'h40846c46, 32'h00000000} /* (0, 13, 6) {real, imag} */,
  {32'h3fd38f7c, 32'h00000000} /* (0, 13, 5) {real, imag} */,
  {32'hbef65242, 32'h00000000} /* (0, 13, 4) {real, imag} */,
  {32'hbfc68592, 32'h00000000} /* (0, 13, 3) {real, imag} */,
  {32'hc028a9fb, 32'h00000000} /* (0, 13, 2) {real, imag} */,
  {32'h3f9b674c, 32'h00000000} /* (0, 13, 1) {real, imag} */,
  {32'h40193cc4, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'hbf03aeea, 32'h00000000} /* (0, 12, 15) {real, imag} */,
  {32'hbf672fc8, 32'h00000000} /* (0, 12, 14) {real, imag} */,
  {32'h3f87d399, 32'h00000000} /* (0, 12, 13) {real, imag} */,
  {32'h3e7ef83c, 32'h00000000} /* (0, 12, 12) {real, imag} */,
  {32'hc01d41ae, 32'h00000000} /* (0, 12, 11) {real, imag} */,
  {32'hbfee6c02, 32'h00000000} /* (0, 12, 10) {real, imag} */,
  {32'h3f4221e4, 32'h00000000} /* (0, 12, 9) {real, imag} */,
  {32'hbf6dceec, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'hc0027587, 32'h00000000} /* (0, 12, 7) {real, imag} */,
  {32'hbf78a59e, 32'h00000000} /* (0, 12, 6) {real, imag} */,
  {32'h3f7e7f92, 32'h00000000} /* (0, 12, 5) {real, imag} */,
  {32'h3d84f960, 32'h00000000} /* (0, 12, 4) {real, imag} */,
  {32'hbf44fd56, 32'h00000000} /* (0, 12, 3) {real, imag} */,
  {32'hc01c2918, 32'h00000000} /* (0, 12, 2) {real, imag} */,
  {32'h3fcaf24b, 32'h00000000} /* (0, 12, 1) {real, imag} */,
  {32'h3f9909be, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h3f5de0b0, 32'h00000000} /* (0, 11, 15) {real, imag} */,
  {32'h3f9cce2a, 32'h00000000} /* (0, 11, 14) {real, imag} */,
  {32'h3fc55606, 32'h00000000} /* (0, 11, 13) {real, imag} */,
  {32'h3e0bc181, 32'h00000000} /* (0, 11, 12) {real, imag} */,
  {32'hbf72c8b7, 32'h00000000} /* (0, 11, 11) {real, imag} */,
  {32'hc00ee6d6, 32'h00000000} /* (0, 11, 10) {real, imag} */,
  {32'h4000acd0, 32'h00000000} /* (0, 11, 9) {real, imag} */,
  {32'h3f3f8062, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'hbf1de964, 32'h00000000} /* (0, 11, 7) {real, imag} */,
  {32'hbea0efa1, 32'h00000000} /* (0, 11, 6) {real, imag} */,
  {32'h40308e30, 32'h00000000} /* (0, 11, 5) {real, imag} */,
  {32'h405536a2, 32'h00000000} /* (0, 11, 4) {real, imag} */,
  {32'h3f56633e, 32'h00000000} /* (0, 11, 3) {real, imag} */,
  {32'hbfc973d4, 32'h00000000} /* (0, 11, 2) {real, imag} */,
  {32'h3f4cc57b, 32'h00000000} /* (0, 11, 1) {real, imag} */,
  {32'h3ea52a96, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h3f93cf20, 32'h00000000} /* (0, 10, 15) {real, imag} */,
  {32'h3ed24639, 32'h00000000} /* (0, 10, 14) {real, imag} */,
  {32'hbfa6b468, 32'h00000000} /* (0, 10, 13) {real, imag} */,
  {32'h3f083c2b, 32'h00000000} /* (0, 10, 12) {real, imag} */,
  {32'h3fa27508, 32'h00000000} /* (0, 10, 11) {real, imag} */,
  {32'h3de06f5c, 32'h00000000} /* (0, 10, 10) {real, imag} */,
  {32'h3fdcb29e, 32'h00000000} /* (0, 10, 9) {real, imag} */,
  {32'h3f4097e1, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'h3fc59bb6, 32'h00000000} /* (0, 10, 7) {real, imag} */,
  {32'h3f849e86, 32'h00000000} /* (0, 10, 6) {real, imag} */,
  {32'h3f0ad591, 32'h00000000} /* (0, 10, 5) {real, imag} */,
  {32'h40723012, 32'h00000000} /* (0, 10, 4) {real, imag} */,
  {32'h401ca25e, 32'h00000000} /* (0, 10, 3) {real, imag} */,
  {32'h3f71b312, 32'h00000000} /* (0, 10, 2) {real, imag} */,
  {32'h4010a30c, 32'h00000000} /* (0, 10, 1) {real, imag} */,
  {32'h3f6a8871, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'h40084a19, 32'h00000000} /* (0, 9, 15) {real, imag} */,
  {32'h3f123862, 32'h00000000} /* (0, 9, 14) {real, imag} */,
  {32'hbf9e56a4, 32'h00000000} /* (0, 9, 13) {real, imag} */,
  {32'hbe6787c3, 32'h00000000} /* (0, 9, 12) {real, imag} */,
  {32'h404c8e3e, 32'h00000000} /* (0, 9, 11) {real, imag} */,
  {32'h401955e2, 32'h00000000} /* (0, 9, 10) {real, imag} */,
  {32'hbf1d12c2, 32'h00000000} /* (0, 9, 9) {real, imag} */,
  {32'hbfb4aabe, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'h3ffb7578, 32'h00000000} /* (0, 9, 7) {real, imag} */,
  {32'hbfb72bd0, 32'h00000000} /* (0, 9, 6) {real, imag} */,
  {32'hbedceddc, 32'h00000000} /* (0, 9, 5) {real, imag} */,
  {32'h3f7c0ed3, 32'h00000000} /* (0, 9, 4) {real, imag} */,
  {32'h3f3c00d0, 32'h00000000} /* (0, 9, 3) {real, imag} */,
  {32'h3f3a26dd, 32'h00000000} /* (0, 9, 2) {real, imag} */,
  {32'h4091d35c, 32'h00000000} /* (0, 9, 1) {real, imag} */,
  {32'h402cd9dc, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'h4053c87c, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'h402e2e56, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'hbf3ddeab, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'hc0242894, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'h3e9ab60d, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'h3f5464ce, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hbd71e3dc, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'hbfd0ce5d, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'h3f8f3621, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hbfda7c40, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'hbe9f5c66, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'hbf4eb1e1, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'hc0062da7, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'hbff5b195, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'h3f2735f3, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'h3f4a7dc8, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h3f329ebc, 32'h00000000} /* (0, 7, 15) {real, imag} */,
  {32'h3e481c3c, 32'h00000000} /* (0, 7, 14) {real, imag} */,
  {32'hbfe7bf7e, 32'h00000000} /* (0, 7, 13) {real, imag} */,
  {32'hbfd01cd4, 32'h00000000} /* (0, 7, 12) {real, imag} */,
  {32'hbf4ddf2f, 32'h00000000} /* (0, 7, 11) {real, imag} */,
  {32'hbeee76b7, 32'h00000000} /* (0, 7, 10) {real, imag} */,
  {32'h3f80c624, 32'h00000000} /* (0, 7, 9) {real, imag} */,
  {32'hbf2c62f2, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'h3efc9b0a, 32'h00000000} /* (0, 7, 7) {real, imag} */,
  {32'hbf8b811a, 32'h00000000} /* (0, 7, 6) {real, imag} */,
  {32'hc02abeec, 32'h00000000} /* (0, 7, 5) {real, imag} */,
  {32'hbff153eb, 32'h00000000} /* (0, 7, 4) {real, imag} */,
  {32'h3f214b18, 32'h00000000} /* (0, 7, 3) {real, imag} */,
  {32'hbf62431f, 32'h00000000} /* (0, 7, 2) {real, imag} */,
  {32'hbfe068c7, 32'h00000000} /* (0, 7, 1) {real, imag} */,
  {32'h3ee0fa61, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'hbec73f82, 32'h00000000} /* (0, 6, 15) {real, imag} */,
  {32'hc00b573e, 32'h00000000} /* (0, 6, 14) {real, imag} */,
  {32'hc01982b3, 32'h00000000} /* (0, 6, 13) {real, imag} */,
  {32'hbdb8c1f0, 32'h00000000} /* (0, 6, 12) {real, imag} */,
  {32'h3da10c1c, 32'h00000000} /* (0, 6, 11) {real, imag} */,
  {32'hbed71c4e, 32'h00000000} /* (0, 6, 10) {real, imag} */,
  {32'h40396c60, 32'h00000000} /* (0, 6, 9) {real, imag} */,
  {32'hbf6ed934, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'h3fbbb97a, 32'h00000000} /* (0, 6, 7) {real, imag} */,
  {32'h401f8b5c, 32'h00000000} /* (0, 6, 6) {real, imag} */,
  {32'hbeba9c8e, 32'h00000000} /* (0, 6, 5) {real, imag} */,
  {32'hbed88fb6, 32'h00000000} /* (0, 6, 4) {real, imag} */,
  {32'hc0196404, 32'h00000000} /* (0, 6, 3) {real, imag} */,
  {32'hc0dbbe93, 32'h00000000} /* (0, 6, 2) {real, imag} */,
  {32'hc031bbd4, 32'h00000000} /* (0, 6, 1) {real, imag} */,
  {32'h4002e993, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hbf0c1bc9, 32'h00000000} /* (0, 5, 15) {real, imag} */,
  {32'hbe7b0ff6, 32'h00000000} /* (0, 5, 14) {real, imag} */,
  {32'hbfe2e816, 32'h00000000} /* (0, 5, 13) {real, imag} */,
  {32'hbf7011e4, 32'h00000000} /* (0, 5, 12) {real, imag} */,
  {32'hbfa66eed, 32'h00000000} /* (0, 5, 11) {real, imag} */,
  {32'hbffc7aae, 32'h00000000} /* (0, 5, 10) {real, imag} */,
  {32'h3fce8c42, 32'h00000000} /* (0, 5, 9) {real, imag} */,
  {32'hbf03e381, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'h402c3149, 32'h00000000} /* (0, 5, 7) {real, imag} */,
  {32'h4096308a, 32'h00000000} /* (0, 5, 6) {real, imag} */,
  {32'h3fa85c7f, 32'h00000000} /* (0, 5, 5) {real, imag} */,
  {32'h4041cebc, 32'h00000000} /* (0, 5, 4) {real, imag} */,
  {32'hbdf04e04, 32'h00000000} /* (0, 5, 3) {real, imag} */,
  {32'hbfd1e576, 32'h00000000} /* (0, 5, 2) {real, imag} */,
  {32'h3f5a8142, 32'h00000000} /* (0, 5, 1) {real, imag} */,
  {32'h3fc135b2, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hbf8ab1ec, 32'h00000000} /* (0, 4, 15) {real, imag} */,
  {32'h3fa55efc, 32'h00000000} /* (0, 4, 14) {real, imag} */,
  {32'h3f217471, 32'h00000000} /* (0, 4, 13) {real, imag} */,
  {32'h3ecf0ccc, 32'h00000000} /* (0, 4, 12) {real, imag} */,
  {32'hbed7c72f, 32'h00000000} /* (0, 4, 11) {real, imag} */,
  {32'hbfa44dd4, 32'h00000000} /* (0, 4, 10) {real, imag} */,
  {32'h3dc5ad74, 32'h00000000} /* (0, 4, 9) {real, imag} */,
  {32'h3d710d30, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'hbe0745f0, 32'h00000000} /* (0, 4, 7) {real, imag} */,
  {32'h3f8a6eb3, 32'h00000000} /* (0, 4, 6) {real, imag} */,
  {32'h3e761356, 32'h00000000} /* (0, 4, 5) {real, imag} */,
  {32'h3fc515a2, 32'h00000000} /* (0, 4, 4) {real, imag} */,
  {32'h3f8457e8, 32'h00000000} /* (0, 4, 3) {real, imag} */,
  {32'hbef8c8e7, 32'h00000000} /* (0, 4, 2) {real, imag} */,
  {32'h3f7b65cc, 32'h00000000} /* (0, 4, 1) {real, imag} */,
  {32'h3f9379e4, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hc010c3c0, 32'h00000000} /* (0, 3, 15) {real, imag} */,
  {32'hbd400488, 32'h00000000} /* (0, 3, 14) {real, imag} */,
  {32'h40174b65, 32'h00000000} /* (0, 3, 13) {real, imag} */,
  {32'h400ee01a, 32'h00000000} /* (0, 3, 12) {real, imag} */,
  {32'h4080cc3e, 32'h00000000} /* (0, 3, 11) {real, imag} */,
  {32'hbf2eaa27, 32'h00000000} /* (0, 3, 10) {real, imag} */,
  {32'hbf3ebe7a, 32'h00000000} /* (0, 3, 9) {real, imag} */,
  {32'h3f1a1354, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h3ee12168, 32'h00000000} /* (0, 3, 7) {real, imag} */,
  {32'hbfafbe3a, 32'h00000000} /* (0, 3, 6) {real, imag} */,
  {32'hc0418f3e, 32'h00000000} /* (0, 3, 5) {real, imag} */,
  {32'hc0744814, 32'h00000000} /* (0, 3, 4) {real, imag} */,
  {32'h3db2f5a4, 32'h00000000} /* (0, 3, 3) {real, imag} */,
  {32'hbeb5605d, 32'h00000000} /* (0, 3, 2) {real, imag} */,
  {32'hbe7d9256, 32'h00000000} /* (0, 3, 1) {real, imag} */,
  {32'h3fe834a0, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hc002f2e3, 32'h00000000} /* (0, 2, 15) {real, imag} */,
  {32'hc0299642, 32'h00000000} /* (0, 2, 14) {real, imag} */,
  {32'h3f647005, 32'h00000000} /* (0, 2, 13) {real, imag} */,
  {32'h3fd1683c, 32'h00000000} /* (0, 2, 12) {real, imag} */,
  {32'h3fcb9eec, 32'h00000000} /* (0, 2, 11) {real, imag} */,
  {32'hbfdec863, 32'h00000000} /* (0, 2, 10) {real, imag} */,
  {32'hc01dcbf4, 32'h00000000} /* (0, 2, 9) {real, imag} */,
  {32'hbf6a86b0, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'h40048761, 32'h00000000} /* (0, 2, 7) {real, imag} */,
  {32'hbd9dc2b8, 32'h00000000} /* (0, 2, 6) {real, imag} */,
  {32'hc037fc0f, 32'h00000000} /* (0, 2, 5) {real, imag} */,
  {32'hbfbb2004, 32'h00000000} /* (0, 2, 4) {real, imag} */,
  {32'hbf839b42, 32'h00000000} /* (0, 2, 3) {real, imag} */,
  {32'hc081392b, 32'h00000000} /* (0, 2, 2) {real, imag} */,
  {32'hc06fab58, 32'h00000000} /* (0, 2, 1) {real, imag} */,
  {32'h3e51ad05, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hbff1f5eb, 32'h00000000} /* (0, 1, 15) {real, imag} */,
  {32'hc00a7710, 32'h00000000} /* (0, 1, 14) {real, imag} */,
  {32'h4025f44e, 32'h00000000} /* (0, 1, 13) {real, imag} */,
  {32'h40474282, 32'h00000000} /* (0, 1, 12) {real, imag} */,
  {32'hbf1ee148, 32'h00000000} /* (0, 1, 11) {real, imag} */,
  {32'hbc06cc40, 32'h00000000} /* (0, 1, 10) {real, imag} */,
  {32'h402828b0, 32'h00000000} /* (0, 1, 9) {real, imag} */,
  {32'h3f17698e, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'hbed3dfc6, 32'h00000000} /* (0, 1, 7) {real, imag} */,
  {32'h3ddc1cf4, 32'h00000000} /* (0, 1, 6) {real, imag} */,
  {32'h3e630b76, 32'h00000000} /* (0, 1, 5) {real, imag} */,
  {32'h40144eb4, 32'h00000000} /* (0, 1, 4) {real, imag} */,
  {32'hbf0a2832, 32'h00000000} /* (0, 1, 3) {real, imag} */,
  {32'hc04d3a3c, 32'h00000000} /* (0, 1, 2) {real, imag} */,
  {32'hc02c839f, 32'h00000000} /* (0, 1, 1) {real, imag} */,
  {32'hbe1d9ea4, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hbf3a77be, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'hbeb61d92, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'h40081651, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h3fff2d0c, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'hbf05754d, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'hbf7e35b3, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'h3f042403, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'h3f8b2f3e, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'hbf294e9c, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'hbf05d3eb, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'h3f8aac9c, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'h4016fb4c, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'h3f6a4e6a, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'h3f578ab0, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'h3f28f1ad, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'h3f944dff, 32'h00000000} /* (0, 0, 0) {real, imag} */};
