-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
l4uSVVE4wIVxeFRVCxZv8SJAH8TpPxTgd8A1S+fdXqDfPIeBW0f2nAzSyPs5XTAr
EDrT2T6qRtSJK7ruM6ngEISVtUWDJP3hYc0cdQ7S6/mwR+8OP0c9sV10HFB3MvAI
3PqosdqYwWx9KUn2S98mSbco443yfmJqC+S45QRiAARXUbcftITcqg==
--pragma protect end_key_block
--pragma protect digest_block
PfBFNFzVn3FFh/p4Wmsn8VZuGhA=
--pragma protect end_digest_block
--pragma protect data_block
c1P1xfixNL+uPylx5neiQY3zgSeNlXCzwS6SjbA99BPb9QttEn/cA6xmSi3RZFRp
Nr1pTuhwJ25Ve7v8G8ajV07P34NPBu9WECsF7t5hmP7j/f+bGFWnUnbAJJ4rXQcO
/i5aBwVb25i5So1wBBLRor6xRhPKI/ujMNxu5Ra7ebdC8rO2plKOTeJk0ED/BIYP
dKtI28HYRWsDERExBbS6sfvTrAR0JdqsopiJsNOjXWgGCgV6GfKXONzRz88e26yO
HDApk9VqdBJce53Os+jnoRi1fh0R0dxrw247P4gJZP7VfGJv9GwzCRyVA9hdRisA
gtw7CMozi1Vap+7jWWoFptdFNh17pZiULzx0iKe/5YBd9fBB4vngvE+aGaXQa5VO
ZHa3hM0TmoPM0DrCVPaZRMXkjC3njjti9PFdsrv9Smy8Lbp+mdGuAxMLQ+d78SOe
b+rqow3taBC0gVJH4uy0Ebdodw8cWjxpEQZ70YNcKM1iAhB8CmeTqSOYZ6aQ1ANg
PLcV5t2mOSa2SZ0uI/9KIllH2KoZmwI/woZUcqMDQpNtPh2M4o2sVa+1CS0DCcnT
LDi5YqbEuDwzB/qf4diJNGiuyHlOVl3v42BosTX4tg9vhyyyxKUksiWKnRnfrkJH
ELq1BeaA9CZdGHr+V95AXtzfmeVzj0W1WmZ27Z5ZZucUMH4J63iyhEc1C7PQuhXz
MWYGoisjq2x6J0UQ4s76u/SoiSvVcPcVTQtNb1zivCSmuqf8JsHnddhchDPclgyl
Ypv93TQVpi/rXL+ySfnmYhE38u9IICqyx35MTWHCkYWor5yyVzmASzGOMvG44Kg5
a037JeriKc62+8AYR/+7uvJ9QIoqWQrYmRW4rCGWVb5gkUoFG61XtnD6wF2gyH25
U5Epr9omiphBA/j9gfKApJUqH8ZEWV5JmKvBAREQoxHIy9LvBXeoBReuTgipsjU/
nmFRbMhDyCoXzfrhx1DSLWIjscO9AiS12d+yvLr4KXVgHl9bCCLDAwh7r1tabOOU
hsKUkzzN7nyhW6XF1MFWJNrjziSl/8C6NyYC1Z8QH4MuNAeLBc3OeMa+tnzfrbEo
41Ii7eaNqNMwTRnYRDzj0vOxd9RULP1759zT5tmv3AzeL7VWBye1vz1lAWZ1AYy7
nNTc5325gByFN1Oh6X21NT5T3u0HMjSYIBjZxofZhuckVTFk/pMpsqQVrNxGil4f
xznY0IbnbvdzIqL2JlX3FvE9fL1cDcK9MDEOWwMVqRGL4B7ucv2LwhT3+l9/ps+m
DfEXO+snxX9FQ/4JzQWzk9q4W6UDOwyO0EWjoUEzLQACMfRlw6OC/NSqRWYVQAcO
EwksIEIAo0a8vVf7jbqhDWo7FTbrrFykOSXx4seI45zOsCkBZdSgWp5u/8MLnLND
H5PqIEFSt9E3+HWNsYq54kntUkSrWsUxq3TcUJaRsZhnesctacjygdySAIek/GeX
MdNgksWDjc4t4GvSEO3f3w/sZ+QqF9ipA3gUwwASfFaa2ZMT5Ugpbm9GOA4+WC+3
W/sYr2BwLN2yPqoFEWrSoIHPbA9H+MycWtBM+R+vQKDdvbY22oudix2+7NPPi2XZ
JFpo2KeYm6yGNQ9NCbsnS5BjGOV5rlVh2AGsdImMPqR1HzkZ2qVdMGjpFtZNEQly
K0isqiThqJBn89Y8v0A1L90w78b6krv2bAXDlucaVNRrJDhzK/0KVxomInRPwvd4
k6wGA6Qz4YBF5MDp6cuCrC2c8qiXHYegU8I9JA/uhiLmHt17QeTw4tOPq6gOgIMm
DjsuMWwuBCxNAUTZn9VcLUsF+CfagJ/zNi8/FJob4BlzUglvu81ITT42eHPuVDcv
bvjmkkNpsBHGM6A4zvGkxQdn2jPcmN9C1xaBIzEo7/KlrtDkSwP3hEWA4Cbhkk8o
pJx4IaEjAr6Tukr78H9n+JJwSyab5wHFVHtTLFbXDu1J52QyeEkQ7m7qo0IT2pC4
CSeOXwP6a/H2AF5DONHcfQ8py+mHQWdjp4v034k30rYkGMBLPmfGS6/uGZCxiId7
EFIKV4S1d2OdrHFdWPDMF0bQDvF1R1pJa3NS6ZAgzioKM/cV0IirE/bU23PUM7qM
+Cm7YLyu2Xvi1k2Z540KFXF1tLp5nm1AwrQ+KCXdF5sAhyTxgHGP/zXWAgDvmXXz
I7g93RAwFBdViV/DAgEZMoN2OSyciAlVIC3tOF4p3/LhGb/FUlf9klqVJ6o+2iy5
18Tf+zaAIVLgURIYW0dW8xw+CeC7T5EPAAgL8loMQPLKUTI2zWC10nV4nZ1y5/B7
DAkG0vAmRCxzTt/tzfxk33OpAO2Vqh/G/qfkbtZkPAYlXZP8V1sUsHbnhn1jj7l9
GhOp0q5yJsZChBVVVdf9CaeV45+k499YT6kiR3Sdh+tzbu4BWzlMNAYPa3eP+SDf
Vz2Cl+0ZlRlUJ629oQz97KeYE6NZv4c24sKWbpkMqg+ME57hBThZbUs0tQDCUX2r

--pragma protect end_data_block
--pragma protect digest_block
M5+KkvrGgeyeFNNCxnSzZI6u22M=
--pragma protect end_digest_block
--pragma protect end_protected
