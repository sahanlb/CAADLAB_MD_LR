// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7tt/qlBVWloKZpl9vgA1tsiLIZv98UH2w/4QZ8GQ/ScoeGClPQfs7q+t8bnP4mfI
SQfsks7uPams3732+cUnMkutPPpD8L3m77/VxSOkzioEL2EyuFZl6dAZ6bgGV3R1
x0sT9RJCmyXBxFaqgm218c5hxA/v4jLvv3jseWCpGWHRnYc5kQBMTg==
//pragma protect end_key_block
//pragma protect digest_block
bfg1Vsr8gEhRh4InTaosbzWYbh8=
//pragma protect end_digest_block
//pragma protect data_block
KH+kU8joB+qRy5HKpuGvb8AxqIS181m0QXTHsUwZzOslFnLEWTb7vLk+XXSNOw+R
70ygcl2T5ziuxghvMJVuw+T5aIKeRjIF4dbpL/HGBzO84+la647d1p7xuNX+HYKO
B15t5Q4eq+7qs2tvl6NlTxLgqSC4TH8x7TezJoyTwQiHc9y4MWMGZs8TppFyG20X
mOuiDDvVhAFUJ+8wePfHVAraZ0G8ycuMGgia2poTW9afLlVrC7HdZ+GZBtpHZ+S3
fKEe9zxmeaiyi/1TeDXjuIysh8Tu8AodNWI8o9Djl2+z7DCKYBqSb39y0OaLIcKi
+xwWY6EuhKT9A82xwXi1JVyRjBzz8UR6kJWI80wn+QigQb8eGDee1QaqI32WHoGy
uqGZWFdPAqTQTgpp/Fq8sfSNgp2KQpr9IZROvVgaZN5FjaPfI7TGycm7HcWfrEkT
rNfNMlvOLtLaM17IOp40AhKL+xs2GTP7pFVVtdp0bLuIBzQjLxl8Qyf8bCVu1vqP
NKB3bAsnt8Tr8m2EQUtU0G8yl8MqhcO8bj5k1cJshhf/3ilekZlgXRVFKtWmso/k
PlQTLP7ZCUL4Jk67JWFfi+UQXegGfpYxGhfqpGUP0AS7vUNWeLSbG7BqZ4BsivMF
UgOVrW/JbnDGTKDsEHLJRHfiY3zj1VjnI8ITamN32OB9YfkQ19G+KNf4BSFuwOxh
oONNoM9ZKNSFSNNA+rICl7zJGtZPgsZaPl8mgMZT0b8Qs7gUfuHkH0xJHayMzA7E
mhCq14RigT26zjxwFOki6LtaeahnqBiZVCB/5K93N8ilPOM0v6iO1sPB/7/aQlsP
h+MgaoClQy6sxzk38mcgveVs4niTtB6tqC7bd4qk5Ff8gUEbQByvRMWk/zdx072S
Hjn2qN4Et2fWoLx5F93ppZlpMl9y+9aD5oG3mJZ3K+UzqUTex/uPwby0ixFPMAeS
6W89dVePjMmOGXvMpZYndEaaa8pRzclEd+PgCROLWhKK5KuD1Lq6wPoX407W/ffG
EZsLsl4h81zlrc0x+n3R51dtLxMo1QkYZeGTyiyoRgqtkDUKtw2cl623TZara5Pg
tVWxWRs2slvR9UZOgDLPYraXuScTzfovxRsn2MDAuQFcBygWZOICHfS1lhKH0brQ
37eCsYM0PoL31YLgyfqeuoN/UbGhSpyond+0J1JvfKCUM/qt5ma4W8rqiUKiEW3f
/C2rMRzB77XfS6yRFBRZnlrr8hk7593fkejPFmx1Kjy5OIxRlNydJYmFtQkGP/zT
1Tg+KcKIn0exxJz5Ov4PxmqZ8kDLNj0OB/o0aBU8gkB0zQV3W4mVz8VCIRyFp/T+
FLp8DjYh8i7HRIPc4VBPwaIB0jiP2+EnBeCjcaxLTuVd+sh8R+vlyzwe48gD+g+W
KqmGGadYAyRle8+HllmupyoFh4T0ENZUudaJtyYgvx6EyarZdXTLWXNxtPe+GjIC
aky+bLrnWgdjVTtiKDGRABs0jus6hETzmBELon3pace/gPafgOaWIiqdn9trWtk0
rhTS9iBPUHrjvjFmSxRBSVxFt5rWZeU5bJMQ4ktmLQXrc1M5gr4BITW+8WpC0wBk
ZCDbitOCKGGJXhzw3QnICltmpkO0jWZel+p35gbYcNuWXp8wcMYMArdr4e/qK6Yw
PoscUKI1qVEwXglvh0mXVnWgQRHzzADgfxA51X7+yZxlisl2U2JsLi80jsV0gxA0
ukx+RyObhWjPpDZmjXm1QKRX0V5sG+DboGcpbXJG6SklgJbHdFgKeGGC0+EuGQ0o
SFSrROpW5TqePQg5tsWK6ovsyAcl2gfCM3WcknclW+PFOnMXLIhtpZgFT3/1/pA5
VelGadn6XpGv5ScaMu1jBPfqezqfAXk7r++q0tHgwKQ1uyHo/9ZSnIvmG8tQWaJF
CD3UKIZYRO2o/WR+xNY/Ff0PW5rj/iqgsv5ZVoLVV84OfGweVwNPSuC52yN9ZQvJ
DF1PrePNnpSvDTqTLbyq98KlLOOxWuPYQsBBimNT6N/i+FFTEhEB1puHqjXk3Le9
THwOyvA8RMqqkcwQ3tMD0t4OcX7hM6qAyYYJV+pnA3ux0QVQ/UsIrtrB5UiskvND
dpD6JctM5F3XkngzSjs3HDBLxdt6Jhw5Svw6CiPAgW0gOnfZccK2Azu4fuj31Af/
4h7ZFsqwJmhNgnIm2fogglQl0msA5B12IhOkvTd6C/CHsFJ32Bbs2jHyeOqM/OCW
KhlddcPy3dWNZDggAo8dxYXO49cUiUc7kzScgPL2dzoDYK9VfakjF63n4VrDCh0R
lnZUAiJIQKslBYr8e7KX6GOI8kXCTtAZdWnSDNX2D9+36cwwoXfBhaARnEAMqXxs
pE2CCm8RLZ2wlt4ivbkSvYOvTAXPeouzPWjUsSLWgmBo4WDn71bN4PLKjmnm4IoO
husZRrxmMqUxg1IqHNLuucbzYu0n8YlnmAvEhoesEulB1ABORktGLlPpjIbC01pV
ep08ZI/sHk37Z3sLxWj6cZdyvuXavg/bQe9/IbARiMj52agoWhvwSUrTLvW/r8Fn
4NBlh+ydzW77aC+xyW37e3Q3SaCv+0XLML2nfnjVxpg/VoKvB82e5KLvqFkhYPcp
XdZdbZntDnGpDcd90N07lMNY7dqO+g6Wy61I0yzXsmTNeB+i4WLhpAMfFzWk8Bn0
qgPS+406/7t/3RJ+U8L0nfKSvvMGfFRxumZYnjtp+Eafl1vvv+9WAIWohxQJBKc9
9WHUzbsodhktOudNBq/aVUIB3g7iUgBboaCs2XwHI1OINuNqzNg9y14nIRocaivW
DjyOP2uGP7KAGE2EjvrrvuAyBtzIgEJ7Il+300K0bw58VWyWfXhvBgPoijVY41LJ
q/aCoNSuF+szwQLIby0gRj2t3xI74XygU5RULdVyBIliM6w+o6+ToR1/yp4ykvbJ
4qZ8qYvN850gUgqy0yyHVOuVJMI2S1SfRsLADNfboGK4WjujLp4/fFvGi6h0GPG7
+/px8KICQkgdM5PSO9l4c5218B4Ee/hsXzI3YCvf9anolAgYF/JF3ECDKXyHbQww
NqevCuL+EZytoOYcd9ASYXdaRG/zV2mcUM9u7mcamkXNEKiZYsUYjYseTfGeCo0Z
Rqlrh5CAM5M/yvDiAjyMlR4lIHwGP5trvl8CsJmOXAqTmLApaCX5jJzp1rsgbLTC
P6dUWoE2prkfWg5q9eLLA2tihDe5LFVKqP1f52NgyG7nVvyfpHgLXtgQrkgTSBz3
pdk5veVoLtjXuHoXsJwkGlLRaxGLEv9sPJ9Wb+KJuhBYRV0rmuHDwE2g+p3EF/oT
dkc2qTbZxegN4p8IGtdEkwuPfHMiEFeck09xb7qdspU67h8W+JNYvL4XBC8KtwVM
H9b8YrZOlm46fcR1ejURAQx8mR4pI4/YlrX7OEYav3PYnxAHDCco9OH8JiPc7gaM
14+FJmzAxdg+gZI3XWk8aOaMzcCXcX4Oym+hLLAHVynGWCFy0RqGBxP5QN8Adwid
QKk5cTZrldETEBgMgsxV9+3Wkc9wt2uNASjHtNaJjy7Kouh8C4b2dDj3CZGLm5kn
yX1ZFWWE136umi2ltTUSnkhjEB7L5BWteUfjok0FVKSIMYehhZxWOBervKlzztLT
q4HlA6/dDtk5LgUG0837x6iATsUF2gp1JqPscnNmmOqFdoZO1DNiq9NM8urGvU7T
cKx0bki3I4hvwETec82/W/Fh1GVCwu/HKsSx2F5vF6dm8xLaz6hqSFBmhBrf1jFF
FeDRvV2Rfe/+uNGghITagA07c76rOX4NGH6ObJQRiLBfKqRHwJ7TaqhF9z1nhCBI
YSkpOsakeskb5HkyM6xFineGpPTpP7EZIEjOXfuMgPzO4PVazPjtlyfGcPpR0/Jq
RZyt6pyrzOWPiCYBYXjNZzp9k0EMZftX7AyuDVVbSVI1qqEVnp8QGBLq5l8A9DPL
TaKfRqWn1Dy376oHT8N79J72UVXI+Mk0O0DzwqVvXTeRplzyypZWf3+H+Mnm69yW
5FFAF5z4M9ZVb9ypBQb8yMPaKSwNJOyDraPCuMHqxk4JywX2o6J20VPoBsWHKdIJ
usID8I8zhkG9iGpz3FtthRpeENTaGm244ciN8TO5A6YJF/QpDRKThUluFlOG3l/s
fuoe6WxZ1qOH9S8PcZ+71M7SF9sYvgGRYjZhBim/AGji6YmXrqxDc2ZPvSOLpPkM
c8kdHqD8PUmTM+nhWcsRBMH+KkZ7umXd1FjtYzc+CizEqkuo4uDWkcBobYB2zzvu
Na5jeDJXXPWMxqfSd/2JZdttF1PhGNagx0Bu/q/CmyCFmZDiuso3tq5o4yxhoKMS
/GTzZrUI6YSPXe8LN4O6h7OZsUMa3/jSH9+Lhfz5kATni8EXr6m5Inmit4rnab/2
PFNoyocS3Uha+PPQx9k0BsW3cWXIywfommEiSh1fD2Zw4OYHw8xd4+sJJf6YTG/D
MqzFxOBi/3d0HCb06ECbH0KkpETMqowUeQfm/tQR5W3SmOXkCi+dsDuIyByYyj41
cICCjNp6zYvIHdYzkS8NYgtKFhf+ofKJH8LSah2FoFnamLK1XDYHIq2gsStk3OMT
N6n9omSxD9hekxPbz/LsVasw1Tv8/ZXyVLQwC25p6tYSLpq4fStCyeX/p2NNFovw
0ctZrgwEv7a4JskHvMn3MCO91Dzq23DpjOx1oWDfexUcdhoYTUX1UuGQP4RhqgUo
4WnAdfmXhG5vob/6lasqUH6H4hqKg1oTM/EkhJQ7Kakpcs68zoSEWzsi40Ymc/o/
Ng+hPegy3UDDY8YASfzTBsdoT85Zd75TMrCx0EByGBw7mIso8S5CFV//n2yw8VK9
ZbdJ9Fbrj7VjFtY3ZYcPgI3XL1HZIx5SdwoglSCV6h6U+DCV4veg74Fox68FGT4A
e4epStL8YWOaVt2BHNkBCuhLe++SbUO6rO8dN8c/MJSHMafEn+b9RmDYmBB38doQ
Y6e74KfHKNVwJ47ek+pNbtORGYZqEWrI5l4+ytFPdStSLc3ncOlvT0hmhKcg8hBl
WB/wuN0rlTcpVL8GJO9kH0n7Iec7inS+NdKYtP0FvHt7Q4egckCZto2L54neGz5Q
Jqhc5pnD6tsGFjaTUbDDFCR1veG6mSkOFjkMg4N4fSHDMNiVSSDFtjQHCJnhTBXC
LAwO0S5cfOZLyNYnvjXPMuUZaozxf0bN7jzfWe/IXO+3QRnUPSucmhqM04GMiJk+
ySOOuCCdR3WbrCcBLghhYBSoDwu+5BB9jvZaxs/9ucdKRVWj9aRMV4aPsWQFBJIC
4/IgFziIc9XjeIz7RDwvuNVXD07oR+l9lGc0VHQP3KID8OwOoES0B6Hd/r+nxFsu
Ji57Wlm3O1MStn3wbAZbasCLjfuRQP6XwfQ7GYSpHfbtoBakPSKQk9W82TYn+UNO
8SEqNk65xJGkzdJ1EoOB3+cNVNgsUdhLCi3fq+oLPBrTTHnmT//Zwt2CTkAJrTRj
feiAuSVFREQ6P0VXP8zNEXdO4uDXz42xXfogy4N6wHGs2ei1zu79Dq4l+Zb2oyAA
qfKgtjpAO87DySTBnUPM+j6j+o9P9Jb/PMDZ49eG46ROOzND23YhAl4UyQD1hfpV
uA/i/7ocZyI+6tPQk4ugPVSpNNLv0VWiXb+67+fcpRJPEEA7nrmU2Kli+bKzXWSf
S+2hTzxI2Ps5Fvzn3inB/4SoGgkKeT/KEWGkkzyY9XIKWNvnbT7Gd/20KAmWZ5VM
O9SM9fbYhpGn63rQnKdX75XmjqhOEY+uKT5XBvS7ccoMvJsd+HiHuCpvQ/oO7KE7
oyIID7JmTETjxjbImdswxI02n/aqhK4O9I1zwjtzksn1uJJ4dZa11P+WI5OxDT6b
uPlV6PFbCddbpeC6/RjNB8oHb5jGxqFzPEiXVPcv6tQF8cnUotGVZ98y+yZoKeu5
/FM/lxp9wjygcf6FymNACz4O/JMVABUDskFs6e4oUiN1RxDQ0JkW2MXTOZJsj3Js
H4L7HFwBm5Ae71RkJ9pH5m99AFcZV9acd29t08vkg7nEyT8l5SKrxTKxEGm2yfmp
tzRtonik83t0GHOPJktOo40zfXsKkrUrjI2tNO/rDvsc/d0EzCqrBKGMCFd3ve8o
DOo38A4HAZx/VfyK/jenczfYAHGeJPHOHfrxryA/m3LnEw8lcZRFR+4iR9U3KaRJ
ulQeq6g8B39TldfAU00AovtNIO68h8d3n0nUHffHGuVV+BN+ScptPhAen9je/pzR
nW2LWhAfeGk9YtMJNe5dAbtmvCKUfZV6DYBTooZ6Q4xk1P7xeizcRqjArU/mrLOX
Uz/bkjXPCRyUchJvZxyyz6DxAzDEsrRuAr42AIWcF3IbB5BORVr1j/HRLZAwnr13
OqErJ7hk9rRfzAf0x46U4f69Qm5FmNxHEkXOc844S1wDn+nlDGk/yj8qj/VABHzS
DOagN1tMz5a9w+hWolp11D10v2cuV8K0l32BIB4AHb3cGSgqez0L6ZaV2pCe9xnH
PSeFq56GN1RfFrRlP4SY2sGdIjfNdJOFtWKR70Fxmdhyf1jcov6eA+WIjyYjm6SI
WnxX3Rnpnp8IUDzE6iwKgk09GSskSzoX/Z31i8C0vQk/c/ZHE89zqIL2R8zgsyPd
GOFPSYDhogiIkh4Zs9sqjzceC1mi3eXEDCujaJzqdSoMKVjT66jtylGI/AUveJg1
N3v8fiBpx6NXXAzy5Rai3+4DU3WhTrKdFAUVFDH871FQDdCsXqOuDBbHtPFR79rp
kLypLxe0UkG3Wrm85Eel+NP7Yy+8dMbLp76Exq/4crXKp9dfbQHXTM2P5X2jZVUf
WBXZdzGfu/dDfveoVEqqt8GuPhiohfT45B8spe8skcIWNjNg418ccQpkB4Ws0cSF
B5jNHyZ+3ppcf3+hyA13bwy2ZE5+U2TMMdmbxaFYKbc7+O8k7jo7wv2eIGSVkMbc
/BeL104QPdT5MagtIQD6RyeC+1fKcFenW/eM1PwEPSLW3DoA4LIqELH4evfA+uBT
DpWx/EYpI1kgZOVkDSe7zz+pvCrdHqcexhyT/KT8lTtNY5ope3Avutwu5hosjUqE
RPu/aoAYiksC96I0CBEqJVUd3t4tkGTrRtG2zTp71qa7yWGJBo8UGb/hID3XDpQf
WI46gB643DB9n0YCJMjguHsRjXcqT2tCDKKeb8CnxwKU8YCm+7dxJQTHg7UCBqv5
Omqin0U0bCAzviE8aOccjL9qMxyI9G7+vBSvca0tIxZuw2wf6xsysxzHgahXKp0F
WhWBhVu/8pUglkhAmOvGxlNRjFfECEhO2464jjOaRgjeoZVl1itX7aJqVSGG3PU/
hOqx9gLehK+iQAOLRXCDkHnsbHYLeD2V3UDq241nuxStpanOWQ92Pjn3yHNsv+C9
k7F5WOlTj67PlP9bdFO2PlxcTKX8RKX/cT0Lc78yeAPmfdz+WMhm14ogpbKQs+OZ
X6G3Gq8HvayaLg2QTks5SpcWUNhzRqYX9c+LqEEFrHIZTtu6O3fal4wJATmPR8HI
Uw4YvhzulPj4/iyQmGbIvjqueB/bJjdOdjfYHFvT7vQJCyxK+Ok5ZFGPTn9CV8BV
+FS47x3f+w/vk2+WPUymJTsM8c7s/PQ6K0JzrGdxxSyX8DY8C/4PS5ID20OtL22w
H2RjlJ4uhCoS8Dq3eaeVoRM5CGSkCNTowyZTBaTiTfVKCY9o5eZB3n/yHSOhSriB
65U56DKmVmLOpkJcB/gFXzc1s0w0KtkQCj8HqFzlPe0SelBbQBajMuBL3toI5Czi
VcJV0a419MyC6TebHfqRFr+millmckp6umXUe2YSO08/YjcIEaRqjZCRq+UpOftl
XySHMGIPJU/cSclzWGbGRpPUg4ndJ/wGaM728KV1UdRAdkfqlljTIBNPUE8TblPe
rXzjPHljcj6vuJUJ3o5WFITp8wD8/UfdnPCkh5ppK0VhqDgxvYtZPugQfmsAfeUr
srnnP+TghkP+DtdwPewmGkFRm7IM0zmJ40ImtM+IVA//sEbE1WEfVyASPderVGY4
/x6eeYWMQQZux4v6aN68IlIog4ANSrG8emnk0JsqSRW19d3FqA+SOhSDUEPe2CaM
eHmLIY+oieNNx+sh70QOwgH1JTSg1zz47q/nvXSL6ggRPw/3ShFNBr/bTpeu/cm/
DkpWmOfhvJgWOSkKn8xnyEZOnQ/m5i4wkpiHBY3EKx4JzHRj/K0AsXdFTJEFIMHU
tMrIYxG6CY0/fMK4fZbxSBc6l5s1gqo8nFf+sSO/3ctUfof9uU8eBA9StwXoKC4u
nN3OGZvKmHJPiOxp7MYnX8zwUlDGv4hJzqxIACRzp19QF4mnclU5BKPTw/TEH9Hx
9SvSZbStobN+msaNlPR+oY4LIh+46iHY95juJhP6lm9hw5UCaLcm+ezRULGZBOi2
8SbgJHrEon5Pgqw9Fbc340r5dThr43MfHKAYN0TaOn0YswP8i8osCy2U2YYJ6aVK
Hj8e1wUQYkjMi2m5+x60cDEfm9IgaACnPeutDjgzEo1bmsbTQuIivciLOtgPUchd
31yT4/vOfHjhesqL9Atitwdn3bd8OnSsSyJazV4ubLJ/Bo3TzT5y9PuQi/SZCWAk
+dEfjlkk6KT4TNP9AJX5MmPhFJIkB+q4gUa1vdfYJ0L0o+OKxSFd93rs6bGOEeAN
BYpyeWOWoZccDvkcdZZIm6C2ryy8gifgFJZ6WPDDpBn5bxPCQQbAjCE76xqDtrj3
hC9ZOq/dZ91X5jsjmPSEO9YuQLZwkl2lZbxlhrMD05XEpDIpYN0AQgDlqsh94IJ1
agArnDOv+2TbCGYLz6jcMoujXzYF2hv6/PUl3QRAUGnEIxmKcebYEZ+kjGykGXTP
LgdBP6sm6vb8BhZBSOdLZ7eOQ4UcwsBCIXDU8Gl/JohPHbKOv+VNecqU6tj20xyZ
Pk+eVAwyJoooAWYzEFI3aeW+k55MxGGMU8QfrarNzqcDojaVNSuP75kKsaVVmKNI
4yWJ+HoO+CixhmvqC1PiDM4NmBb15bymPoK3ygYw3FYHNE3nik1oGkYcBk3jhUz6
B4Nibb52ZYriYPI1AKID/2vnwAsYW0AG4mWvIjtMrGHningOudu81Y9Xen08lmmR
ausZx2NxEX4lvhUrBRiLfkM/CzFVvh9fuWSwq4pjqG5tnu0wINwRNyvAjf1mxB3y
dks8p8gECtKpP6G5T/y/X/Sl7nsEhC3tBt1GocpU1Nc6ThYriMguD9OBYy1BcJvM
/gItCG2y5xHG/ZNIQMnkwOb3BrrecOwwz+nCVdCmnJNTHblmM+i+Qb6pFwUVHtDX
/QL0uij/3g8sCrn6SlQDRiZ/ELgLrbrHO19psQnhLy7FD0auwVYa5iTzu+WNg1rp
r74cT7Vcn67ylILVpB9gTO21PpHAniSpmMgszBuNFqP8gU190YonaKXLYW0ar+z6
ddF5tmiOzwrZwvmnQVEHn8CEXyYXzcvpzW9BtCAEsiGvsnvJUGEbi0fWLmxsIIyp
2c+33es9kjNqXmLewXyGMPjLvN+ik7tj70abEq+U0kNaJze0wIzcf5t3oE4xvBTh
TTFs7TvWIOqjHNfZLzkzpIHqYLqKXbHz3VoiYBtmYNmqq67voFYF5cqqODFf/2it
cGrpB3bMJ+5pOclc31/Md4MJtwON/UWx8Uda8BE24cX2pEuWKVDE42m0QU55FcAr
p0u1AItwp1QRFP9J4xqn923QGnMHcJ6TSnlFqIFhOveaeY3o6c1bkjdUogTGkkPo
hPWLkssM+GD/jUYvi9SqisUi+FdenFIP16JmIHp2eWybtBNiO+CfjW1goBhtFoY2
cIj7L/d1azxAPW1uJpBQVv+vzShYB8nieGiOMqMJnj8NtIA67iFfj3xHl+7sXyHL
l6JmgfFxufCbBUFdc+iJOIqov35VaGRj3z5ikVlVx0Xpkct0lsp7qdf4hL2GEIOf
cwlfEj3r3wYtNIOznLgd3/ED5pnFmte/+zUx6wN3n3/gNUdvfOE4ZGBR7QUqexbm
WRo04Nkc+dcKgbxisC84ZXGgB5nsvd256Uw8MwoGMwBKRiW6hVVgImfnKT9LFZJD
hYVaRJ3M+n7TM6Huey5rEo6gsxnC6EqwRBCSzRHlrftv8ZQ02IVV1YT+JwxVKf4q
GPPkz9eoSRc+HXPV1Z6c504J04OmvHo+W/C9c6s+cfcmc88QfaPeYPDxy2gr10/G
1SCEoM2it8PetPBffmWk9f09sNV/MTH12KkNxRMm6xqECUIzYKICBMplPg+TfrQD
MYh6BXNWw8yROU8L69QwDIHU/jjhngb4MsJG7SDAGeRzqkuU2ebLgN548eTee5fF
NsSoq9bLLVMZHzlnFzd9yVCeliK5avJ6VlYGSkwp4O8Qbx6tWJo5hcSNN3JFI2I5
VbNrrlgK92Xn63L4QTqshTYGwRfJCAXtJ/wYDOZ2DT81OHF1DhL/WPzxtMQ+Kd5f
8wV9x+RVza12DE/V7GqMqHvFI3gH7KjbYfNC8rXv78aKKTlHmWozlNIa8nRLgXNf
x/zvECq/GJ0Gve7Gfp/6Jk9FscJ7TQf/KOLnWES7k573+n5d3zBEWQ4XgG3yv2Aa
P+t/+cRZaBnsnwQVUSIMwy8vXyiUsO5UozJeyD1/YQqLg4i01RiniZtCzNWgQwY+
9vp+6WnKxRhsSMx4aJxh9POcMQlnjxaB3nTadik6pKwXICm5cZWvjeHNow8rfONa
ju+NObDbTIGEPu176hoMuCEK7eX0fOasDA9J9u+K+/GhEXYN/DiEP2E19fjbLBUA
vvxxcDE4gCWnxs4Rw/D1FpbFTmEXPaXsd+yz/gJbqezqE5FDqKYxznM2eQTQxXVm
USerXTA55O26+yiJSOb/jhlx9BcVbO9tu1rOlRa/GIdm3JzFajfsT1u+3ZIvJw0A
H5ePG5f8WDKgpe3e6M71unZOzXR8LaaKV5HkSX5+TVpMenUNyblNOzhlHxGP6smR
YWhdP+6p/MicbqpdkvQJBQMMj/DSXVtzXyeGWePurriw1ZGWV6xcBXolnysJJJqx
0/DVMTvcpxqwdGYru2ST3KzBJ/8v6yuYNOm2zMNSAvoQr4yXG/rriOqeN1AdcyG3
QNrCK3skvXkYws8NWGPtzlPVf+MTAZKQ93pTIbi2TNRwKtWPMMougYfo7cZHBeIm
zj7L+CLbvd69MvC7jO/LmlZMUbfTHIiEXCxTN2OD4EJv+AZiZZinOFsA0TEY6Pmd
P6weSagju11Gw+HkwtA5DGim/m3LPd4rcVt7rOJrEZRH39zHj+nu3/JwqgHwwD7r
pkZdw4yHwa3P0BLvmX0WWyyocnAyyhhP2FPjZJkwabkauVvJwHUfRUkCRTQuzfJW
qwlFFlAY7pkiB7QnM1WIE0U7q4B6cciSZtvh35HMwB+FGfUWUEPD0onPLxoDxJLv
+Rhu8fXn5nT43y7oXQdtH/sxAoJRZW6yKnv1fT+N1WhhrbGReqwQGo3CtytPswov
TM47Iu3oUc5CkomJE+z+/gd3I1jDdOvkbQUSyTWtRgDfGuGsC/WMJ5nQmlbCg8s1
jEXdLEF3FCIdkegZB3Rc0/bCcs/6Z+6j2c6/BAB4BxG738XjAi4ict5tn1f1luRe
qt6qJu1p+Hj1+0aKqx1AZpUnKPN6mmsyyp7UIe/0D//LqB0JbIH6sAqnv0pFf3xl
1puUTYXSOuh/VyvGbk3Wuwb9qCtj9H3jfCmga0Z9TBvsdSDHRPS8gPZocdwh7n6c
+8wdhWprWeT66CMj2wE5awV7wtBQIaWsaA3IApt8/EtN6wB6HS+Si93qywzFVZyM
01yAOt/JwXe7RaZ5u9nnxZ0q4U70R8oohCOVA2ixDmNvmrQAirqXQ9BHKT7deIeQ
DsKGXhlIGDgEqpLN/lvmREcW3QYykmwCYJypNGGdYOJ0J1FMhG4F3pktG+CsGg7k
6U9iYbKxMsp4r1cejPVCSOfvbFZl483Xacfcfny4fTrq/TpqrA6zjUpbikiriSbG
bMnp/6XEeXH2v58Zr8fOp3dmPEvaKp6Yd26FZiYAR14nFQFlNmA8QUCoo+DIBMWM
tRHHjHdOA6UEs3/W/dqlnL3wiVjbzutpq4ZANR3gXKZ5vMMAZv085CTP8uPNWgkn
YQlpHhhMevO73ePiKDTDmi5u8qC6ZcguXqhBTpyZcfBSFLyVG+yZYQIGRHqTU8MI
SxT3TCoMBQsW1FGuIHVsVCYJY+7tDgHv72LpREX5HLb6V3nBNtcSIGu7xiwCaoLM
j03h6WBeQi1I6Y/dVJCpLlUv05vyCv8djReDQVefIkn60dWYYraOTNhunAO+R3DS
79iGlplkTdTgl679DqgYX3nBkjVXB0ZTwSb29QbClffvy8Cq19i0TeHfILwq+O/8
w5+FDW1EJO8yOVVX6Awfaln4l0AOdvZvGsSgDND9RLwIvqVHXd8UlrsIfS27HAzm
Pwkyp9DIFNTx4wnBQbM+PYgNJI5i1oD533hQ+H4iA+0FCLmcBzecvx9GugBBvhgI
jD2B5MKunN6pQGQJRhOLXkCynjTKYWEX/rZWEH+saQ2eKmOkmcQlTk9x9lUj5Z9R
TpktZEdE8gtLVDgg6YNLBUnJOF01QJqmMo/krDE2smmRmnOBzzKfNV9ZVErQFdyD
eU6bm7YwixKA1MMSHCL81GwuBWhQSQbG7u9AxhazlGNxnZk7cwyxlWqZZq8nznyE
/eOqej/JohigrCHjcswisUiqyoCsm5NTLmgc21D3AZklWBWJBK9N35sjrzBEMFOl
VN9Fb3IvsdbzBBZmPVdqx8EIMmuXnx/+BkNrD6VtrvkuWeYm6ORicSFhXw0B5ytG
//UsskUGpbcv6B7O0X34JuxwJFBKcn5bWy57C2AOm8IqgsgKPsMeZ1u1gXAt58T+
gB+iGlPDu39g6BrJGIp8TDE4uJ+AZ/bJ7RWgTifKJr6egMYz5nu6DmwSs9BxR/vp
ziFAMQ0GM+qLM3B2sY0biz+WuUYwpnORyWrgAWp4kY7wpyvi4cHOf9adsRGWTJjh
4n1wi0hBlfRx3N2PeDuOGeiCnGj7SWXvYKgRSbpary+1G4+TZ6ShBs22R83eM7DT
AEX1mhLXxJF2D3s/kEjTEG2/jI/oLExovdriYccaIRBWa9wTXXF8Nv8H70Amxxn6
mzZahjxXqECJFo3j6WG77BmIXqFjC4L6YP0U2gkihhQPSPvWZ5ukzMNtBRGcjBYU
oWYyVC2md9BcwzPfgmszmbYAs2KtbUAGMzGSyaRtNWlLDV1F1KqXdOWgv1O+hrn8
FNv5yfVYDLhtBsnAWPP92eMMPWVlr7TsiGxUx+4fC85pgeFNAxgDKHljPu3Z6SwI
j7OEni15ezdANWFDmLe2WDWWlj6qMLseNP9du5ipuNVOGi/CUCy/2C9NvpyQ3h21
5TszS5cD/TcHuS4tPGYtwGhBzPxc/SKGxfqJLNSDWgGg21AaBYN9T819wqL9OelX
7roG81Lv/dfF4aJ23AFKeLTwN2GdH5nteQCocXy4VFcft8IzHgCmGyOYDwXkRYmv
GKN1gPuXAWBQXvxKALmu+f9oEQ9OGeuHgMLiarBCukKy9lah+G2nLxcfVYoJeWr+
4qVzUn+WqmQWj/lXqT35zNDZUmTrl6vcSzrnqx5bfcD076Efum0GibAwUikDOgka
nhVabrhfnGFQFpSnWBf471baOqZl8SB2//PXWWExGN6dA0HB0tJKeqpXt2+0JqYZ
v/r/icidkSgBAEPCVNsfreiUY3W3Ply1c0/s6kErOgZ8SUl0fiO2cPazisSXjxjA
PpClEsdKF+70G+8rCr8KN2XlHf1BSkilUYggBBAlNdMOr9I/Y5wNROrOiODbSMXb
TiKOaC4Z3U1wfFCldx4qW9OldNb4abgHGwQZ8NHtzqMRgg23aUzKM6ny2fUUXnnC
ULLVuTvdZCb5PVm2NwlNwdZ0E3PUdfR2+tJpxlf/HMHvaGwxCxY+lq6ukZiNx9/y
jyMsT3j/gTL6L1Gy7F9X7Uj7tXCPkV4hm90OK2Ic+gLeQVp6Kq1hby+qV+bELd4V
SU6Ht0IfoTvsT9r1wDaVxfvwthAh4k04XbvDY+fCKQR2Syow4LqJFSFMjrQNf/WY
r3U7OMVhlTrjVrZfbdjJ2a9cz3T0qFp5L5AoMOaUJgljK0hTOrqWu9RC62HdI2Lg
YdTeKWsr8bwl35uuQDtm69Us0B/gtd6lPo9gcB2z65DLf5fvC4y5HGJTWXN2mmIk
Gs3UEsPU/LSayqs20uK+pFPNfBq1l/nuGLSmWfjEM4z3W0ZwOpjPOer+YO5qAKB+
swLljL2BHf/Qvxi3ct+d81cVDWGpVzh0v9edIbjn4tEYS7yDnWgX1fkDmX2ppNCO
wDGMJeXOS69BZ4N9xpBOXvA+h2I+T63eY40mKc+sM54Gakh77q6kywdBJaGYxrKw
ksSjneBEt8/kFiZd5To2BOkO31kbvQ66Wy7id8F+ufWLcrNJ/51HUBGYSlk52KZT
rlcfR5X0NLJvbByAKlYModnR1NpLfSujxu7N40wansWYOQnKhNk2sYiHFjNBx/yU
nqpwOhKeeheIEmkCGxe/yEYgy8bC0x3DJArcRrgYRK/HMKa85s95pUPT7enH1+Ws
DuVI5zeLDRT2TaHAAt00qwZtBB7iTNdVKG4OWLsdwmrX9lta9yczyysVufU9wUbG
mE12ySBboRrml4f4nY0O8CytNe21zO9mr94WSbWxdTSqWnDIw6eAR4JryIfEKmIS
rE8ov+mkeew4PPq3kHoW0RnBjVF+5cco8+bYyds+emR9CIspTyFoCqGxT70hzdTL
pFiseQlUrr10LgLso2XW3OUoAqho7cknFeTsByv9J6w6J04xqZ7vm2NuIFqTlUNq
cY//I9usqaqiiuDnx54XkFnPmLxYn8VkApEySFZANF9w+tT4FTdexyp1hb9+ewJo

//pragma protect end_data_block
//pragma protect digest_block
tbuZMWDFqhvhEeyB4rwX2lzGp18=
//pragma protect end_digest_block
//pragma protect end_protected
