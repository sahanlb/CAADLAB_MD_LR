-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
4sBqnaGzPQaLzOE25lAG/Dhq7i+7BAzM/1+PmGWNS9sNtrOYHoXil5XvqQhKuPJ9
26Q+Hp4qE0cAXr1USYKtDkW770uE4Zu9cflrrAip5z456MClyOAGba+vEZkXVBDX
bi0qEjq7/ki/dOpR0Yvra8YAglGTukYhtBxbDEGuUQg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5168)
`protect data_block
tplAy4FRdVSEcDWQqyoIemGbFlwJUQYucYp+ny5vt624rQPuIQDwpO0hGK3Fkx2b
W3ajFs5BoG45rmr2aE5y2wVh3tjm8CZw+kyzjCYFK8I3wyzAem8EEj//qz+mRjm/
JQeEVYxn4mtsfFv0paC/rP16775k1GoAcix0+qN8g8P3tl/+sfrJ8fe7wj4DctML
q0kCg5igoufmp/7Rz/NRwdlq9gXGlfZ4+BjgDAsIfCVt6KIVCfbVVglcAsalqvZo
GeYck0BZ08bh4fM78JrZ1Ijf+eYNvFBTJxStWJwI/fLf1Ew3/oMyXbItG/gHFII3
5HH0gTJ0TDG0TZlhma8EHNkGu+r8WLDWXZRIGklcyRIQw3vpaN2M900/rb1yRmSk
3ph/aAJXJ+3XfeFJXlsI/aVUugxsFXv9jgOhGbXpwbUEY5Ej5oY0xZwAzZpvMEWH
ryqKU1fAEoJBEXN4KD/fE5PU0WDzp+X+9RBT0FFPAUG3iFzWBSEDlmGBWGMG6O7u
63Rk+13GjeQ0svCfaml4zBObOz5XhSu8SyAaaXVaVDKE3oBa3EVssxkYqfn+ncm1
EHELHaVUX5ZH1V4OTYQ/a8roeYRpOMZ/zvSX0hjD63hvvWjw35lt6M4EEFu/XfGq
+BNZbklQiM9VFwo/hy6JzeBe0ahoM6sdKFLbL2u3YedU4UG7m8Z9N+1K8x3ynTYl
t33W74rSedvOnQuNKmvsP94j7FRlohq3jzOOElwNN3vdiavzOfAhyMW4ZJ9kYyFc
MV6QTLGhIeaksAM7bkelhFAZUip5oFv27IWVy28x+yDtpp5KDXEx0M2xMVWJm0vW
NhAq92w0EyCf7awrZ+NHsyr5XhSBS5nQmdiR3vMc9o3lCV3a9ycZLLBlD4QZVHA/
t9NQ2LX5VsnOyU86HGJ2b0p1AreZXoX3dErUL++g/RsusfvZBt7qqfRitKIoLrKK
qrlmohtyuzfn+2Dl0Svw8t/JrZXMwN+EuRWRNMJlMnT+rkYVStnHEWplyBK12s8V
La1g5aWKK1S/vwBXbZeE8hTEOgAymuzKEhvFl6zss+L3eC47K3kOZ2OTPWjICtJb
aAyR7+Hnwq0Mhfnz6QIhFNm8KYanFODr+Iz1rNkhKkZMORfHuvcb8FEp3MRISLyN
HdJR2W8UlJFxYd0nyZLZAF4vnxq4EVDBXMdGfsemm0TZwmoh1EZOISl45O/HpNDR
bIB8xLlOB+2f9omZzZRyXKkQHbR42nzhMwkUiTBVqDSN9G3/OKDScS/tVUiEel8c
dI4IlxR0en64890zozhsm+TuEavbxazGmjLAlwOFoEHm5o2i9URSoWJiovTdH119
ibSROzEK6F/ghsRxD4gmr58OQZmBss2fXadHH/5VFCfy5lUDoizY5PujcWo4PgIi
mQfdT52g9NhXQgTq6to4oecGBYdSoQVY+glvp6bFKJ9+P1+v+DWzl1rRWEu3Cj8o
tjoh+J4NwVpYvwe4Ow81ywGU2+XXgHbrzcewazeCdXrQBNyFh4B8VHEN/KXU8B8N
Tvc2n+Tz5HePReNSzRFdApWlMClo7VLR/Hsr4A8VoUP75dtC0VxvzGSyrHRuW72l
7kufVp9vEpnbGigG8PIndip4SosQki5SNQo2AIWYRV+NMnhHbS1xYnSPGikJQeMU
rwfbh6lUBqtPbZpLz+PMF0fjuib0WwbhUBFl+fAUMIbKIWQaPXzTdrBhR4OUOoNj
k868Mr8KpMUmeopNRzmLQWvfKiffVIDnCPtVs8yo8BOhCCJuALtJ52HzpoI8R7/M
+UBeZqc0rCOUTwyvpdQLkXoSslTcFfiZ/HOFiS+JDPGOiELx1Du2EM6Y5TE+0reh
y3fce76FTVF6FYvKXrgcRwco7LtEPh8q1w8RqBkAl/D0e7/zk4mgcLNe3VA23E9o
+TKCFjlJSN3U1QsbkGO+u82n7dcUmeDrlNtpHg1seo+tcU77YhBs3hVU2GT7gH8V
xQqbSG7euruxMA5C5mpkWPEanEsOyiY4qDf1Txn9ifmQc4dh7jLigjwQbDp+5kLg
Z7lW8EsP/jN7M/QmP6HENIn0Kt0YpUZQr+Jkf22uBB4mwz67WIxCCZ1drQH9pxJH
BOnFFowK5KG8iXvr/Lyv3JyqOMRdYhjFMjBv06DfkDSj3iZ4KMzzUsOYT8LnKUgs
JqcebfgMKws8k9oOI3IAA+3DBRNKCGRq0hRJqNFKuY3jBm3TpX89d16Vwud0wjGz
gUEbvAi4gW15Pdr9eV0Jb2jZ39pwUWiMOb+5cBmryZj+89wBBQCjTZjb4qla0wVg
pm+o8TTNBcqQtNXK3MmDBFIgpp9UlEAbFxjpckkK75B9yY7q1Yx3v5iqjRezGXyQ
y8D+SgtjQ7HS3wiLxH2MXfpo4X9yGPc78n2l1pTTvwLpCtcHQ2JGjeUngKw6Fk1n
iycYIMIKyj4XWkvPQDPnzklLppaIjlT2qoCqR9Sor1HKGvwd7J8KvvszmkY/mbbN
lUUYo5NH6j0//1BJjm5hittspCzoJNOFGssJmVNBwP0aQA7J8qi3nIZ0EkppYPnB
Iar7xoe0d7VNLUPhXjcifzzeNVwhEiJD8BASsAcs/asEglHS/EZHBojhR7Op185V
vnGU5ZZQrYaZjHni29mrFRSyPsGziTIPUDeeFoizgxE6Jl+CjKuLraHWw1ealigQ
0bvl/Op7yodg2DMe25uG4S3ZcL55AhkXibXod70EiXH5BZOT//85PHG6IC7Bx5ls
rEqCNB00a2tSY+AEONQYDGRn2SIJBUqXmj/I72bUd36D/kmgjq8QfWY8Saq1wSla
VHfNb87GQkFWNWvoo1aVfAon0VxzVGlHQ8wngE+KQXsdzv3+JE25pNVYtsqS2AV6
xIZ6E4PYYXqctx/fy7XfWSsZrpDy3+12pBaRXVcAX1DSedHkX0s+NtJYwsXVziqO
VUHnj5xHbYTKmydsL5BAMoc2lCZGUfy665tHo/rSIQ7/XCecCS+faT3av+c4muHB
ViZcgQM6sYVIUtC/rjEhukMGX+dvTtKp4398bzQBk9R2VsmVe0A5k0G9YqxOMMfK
uAFI9HFXyESx/2ZtNN40+isFuvN27oWrHtW7SLZWLM/4nH6ZXdMl78+kPl1wpc5N
c+/hSh5CUfgeT4VUsXziLDJQAxPzc8f9MabDzei75Lj8VDspg3/FNDOvdk3rFIkf
50S7jIMYVAtxKO0xurpiOCIDgAktEnpQacdo54sVTyPb8Co4ngjWmLqjcw92+jkB
//rlimw/fW0L578eJyMn/vlj9HkyqMj5vFnNupK8AZK5aBL8X14/mcxWkm89GHBO
no03ubRTZz8Xjghto3kBi2ZbR5QFfODXiXXlucmoBPZzkq6lD/M8eIiHiuuoXaCo
xV4Twp24ttRImk7mTFOKEB4C13A85Mk3CDGAKGSTFX+Ew1nv8+zc4CiOXpn/z+sG
Mbb3/8QkJyrsXbY8hjHJhugmKQw/Gxu+uMC6UmMo+7p1McnhaCWmceyTHksq4tGp
Zjm1HsfINsTZOPP6kBUnhtTiU8kZAiubtkXjMqDVI65OQg1CSgT6E7545jsR45CM
gfIO3lmUQKUR69tHZMbqSvNh/yVlOfhL6oCZ4hP15hpAlGu9LXAPiKdwYx1CzZLy
5/s4TMTkmpoz10xOGJ352s0REGpTcBxA9R0KD4I8AJ39QOrNX3ki/8wGVW8H6Ihq
lA4b1g14xXW1jPIof9mnym49yeA7MUTGCYLkW2SGYTVohypgzBP9ttJl87IwpNik
D/0zwD3siUa1E+5tzpoI24Q+0oomSTua/kcQsAh6vfP/zO+13fUNe0QhmAzNOWu+
69W56T+8UKm/Z041KR6URfSOfmFbmMabN/Xb1wkyCu9Vugzo5yFvhKTFQe+D0M/V
wuUg7a9tpR7XxkGsjHbqfDnKQDKj1W1jL2MBnJOvVD7Tv72rxBCV9lXJIEuQzB+3
35sV2S7SV4Nh/Lcemg02q1UNUDRTt1SnYOoSCpPPPh5jZk73gfgJCzwxCixHYU0O
aAZmhFHiiJzNHusUQuXb9JXj5cfBQAK4uUr98D0bHYuhSZgGuK/YtQ5weR8lCZ8C
WJfkaPhsvW/AuJb6SRcxjY27LS2z+Ktgpq/iQjhGM2LgjCNCrx6xxK3gEBK3PDIv
pXmnvxATABE7MukrkqOjZm2LVPaPwnkLMWFXFETq9GvQpVmK4FsC3VdkhZITpGPG
MGnezT9N5KcUhT7+aRQvpCHsK/xBLVVt5uWKOSvgjuX5rRxIr+onWsJNvaJC5VLg
PZvdHqMvp4rh4dDv74NHMeuXdn/Z2l1+0E/uYs3k3lTYGjmSE0gH+qL/QAWfZNNC
RR84aLnF1ECMD9Z3llDpL2ccLCkiEmR+w7HZI7bJ1BwcyGkIqzgQQ0r4FvlNtfu1
Uh7I4vebcqO3iTMAwzZe0tRdGX6ggdY4QQJ2sB7IWUWvMudmFEa/R2j9NnXIZEfH
uGPu5aAlbYtyVq8Vbuzn1sMaPa2hsGIa1xYuc8mvWLW4KnSHcxWJIbrYSAKEIjlZ
OZ6xY8v348QiQ37VliuhJqxGawVomyZpMAfXoW8LocdAUAhptBxWrasAvBmWYw4e
dou7D4wIBTWUUyJrSoaQEJKZoA5IT4d+dLnZlkvbuIzBaARvNRDoB/PHrLtumvdT
BmNJGuGJZu8we9ldN73iBMN91nsLuwCcMUVI6RVgk1NiSygaMxApDoigMEZCUZUJ
kecxeCxvDBqEWwLXAzsM2AFXL/pvJ3yk4FropWiRlr0/cxiSS8Li6TfwRRYZ2nzk
8BLmiOTpv91pmnQXZa+tBPgcfbyVcHp+HXrzAEZfzzyOIzr2rWIecQMhv1yus9f4
0O2kYLupfIgZpnfyNvBn3KXrP3v4Hs49yYj83QXHWYp3lYrnHGEr8ui17qpO7s00
R/psaSTR5Y8tFKNlK17BdqP+qnq2TwzHb3VVsJPoNQcvLgZXbau8ifkv3AQ0/N7Y
CO3UPAgarSZAwdeUcPtpLkktSB2wKuuvPZ1xcZb+FwefDPkc4xGeXvmvX0PLaBWA
F1CraBDJx7O5asAfM/HrUUeEbyhmXmZ2IV91LiCO9oeYuq6qUTFenLLziEJS4eML
SoviKzIGkc2MZ+fUFj5N1e+fZAeFZiOHhAOavVlr2P71PYB72yFxd8cX2ePbyDnD
eU5bMgulw5k3hdDQeHhBwHxbKkcebAafb00GspEbQJw3GiF3lkA26ZbZc0bUIu/K
D0qUIH55gMtOBD5R7V5eDtHP7ys/nsAYTB1EXB/gRpE/niTVRZqqzL57nScSeQu6
JhZtmX81DoRLDcG78HgfgcmJFqCvFHzYXtK73ApvBycPBkJlG0Pk/lAI7ejLpjX3
KwXzTSal3HyTaHYBMiK+NSFlAcywwfFaIyxEJOuMOLZqtFTsRuOrswG2LG7f21F1
9btawZVOWv+V3iS3kDecffYOhHV8q7+Xff1Fem7fTgvgx6UjM6nvCYHb/iXG0nwA
KAZ4bD0sR/EVJmK5rpqFIcH+Uf8L3PeYMfMTAJdyXXnuXNxPHCQSiC95sRwMNkbJ
HgS1HvU38FTmivnLSPyWKiVK0lNC2KnRXu7zRKGd9Ud5q0+ktLGYb+1NoJI8LXUM
oMTD3ly8NcSVzC2w9FjAS25rgNJmZgSBARKzhGhPKMIrq8RCQYGZ/fJ7AN0mIWet
fpgzOZjQefT0SKW/L0iEOrHgYr7ryPsgjJ7DuZc/Q2LHhvUHQfUEgI0gQ2/tpIFr
DA31tf37DeSjf1dlq5d/7TwOURLQvx2N46FA5Z6g4gq2DllJJmPLqWrjZN6MQXHS
uACW7c7k7IwA0pMAHPFjIs2VrhVGP4KlHZVhHbWJLperLUAM1Jep+xmmsCW0V48f
4KoQlaAWI6I8QkYkqLThb76YisILSIsciHZBP32Pj+TsS1pW+E1tLCW+NZ4tj0ly
3zccXo4xiqAs1DW0zhiFFpjdxh4jG6dTNjWHvuvuSkVO07ycufTpOuZAly5fVobs
IZnC+r+PoEigKYkwq04r1oeP+e3qx4M40HInSLbv8P3UP+RSyZ/VsofeRRQb/mn/
Nm/XzgIqb1Jyu8UGQIKMHJtSfDfIPngQpIbHQuM8K+acQOcwwTBaXQ9voQw4fS0m
Dc2Fh+cFTtGXvPWmeb4kASmHwLqRhelx9kf15zR2TcmvMUcLwXa8FW6krf6Q9zmG
PgfXAeYBR6hSwfcpXLr6jilzLuX3dEGUpOjXk42Zs/l87YZPxTVdRSxZpwD8E8eH
uH7BT4OsTrjFLYl8OHFVcLmLoVK7Yc8zcdwWR+46Rcrj1pCc5R3J6Uay5NYu3J/2
RH4ZVi6llLMp7lKd1Cfx1jHdjEn2sa97rAQ0trKm4/w1bh7MS6YBuSeE4bRL8vvg
oagKiytcM9WC8XJVOvhrLW6XNfGQR0OxRgk1x8EFfC8LntbOBS+7b/B6NhW0kUIA
m/LDo32BINBkmrayp5m99GHvM7L2lhR+By1KS8TqIgZ+cxBk0e/KhOWP0HQ2/Hrr
DfXhuCT4IO87Vr03rcDoqcC4kIX1+17fKYTHM1Ki8x2aoWfJEbje2orNBk0JY3tm
YgkVcZEhsSX8MaIGRExkzBJqKokIJM29GCya2SxSa/r6CeVyxmkaIj0jXhYgcj5D
hQVeaNoeOr63NOwVUcNWOaPvHgun7UKMdfJUxywUhaXclnBKwobVEUaWHupBPiMC
zdIjc9Nmsi7JKTMjtW49/1RRhrgxQznl/s7dObq2XTa20+M3QA+N85XTZgrBfDJG
Gmc7LFQJmiZhTVQevNZMr8Mn1asaeGOJVl1PYnZSOCVRlYkJJ3S4n81mFGtLqPX0
APPac3dVwoWQ3psR/nG64Dz9jlZ+sdUD/ZPjs24g6rw=
`protect end_protected
