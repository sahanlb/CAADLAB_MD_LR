-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
PFtz95flJDDLfoqbm3Ay6wbd7w7U12sjT0Z/wxBX0OWmeU40uO/Hy7NHYZUCluvo
DYdv6xLQXdHj/1XFvDYCsLnec6kXdtcs9syuLfMJxds4flOXwDFYCyydau3y9M0S
FKIS23+cW0cGxINQl8wDT/6iSLjDztk+VS5mmi0Q0ilepx4u0yT+Ag==
--pragma protect end_key_block
--pragma protect digest_block
nJlwgkiZhJvXEMdTDoeQFQIiBTY=
--pragma protect end_digest_block
--pragma protect data_block
D9f8JdWpoJxiyPstQTlji215iMrzttcPPj1mEEJMhr2CH0jA1IvPeHRRDpqGja9t
cf04B0SwaMYQ642D58pIW39jB0edD7iAuWCAq3pB85LD3OVNGxUDdSY7vXVkqg5b
cY/TjVBGswHN0MfDnjJT8ik9yFezRgSNb2twUyQe1e//xiSUm/F3a5EUlVkH1qsR
PE1G45izpcjBbY5dtuKeefpFr4TxeH5rQ3/9Fh/CepOIDxJaexn48Zs+TbRyGZZB
jRSNYOFTwhS4SNuwqV8TBJWoiPBRvRqMbu289pvSj6UfR79f1kzy0H1Aw/1VOOrS
u/0Zs0022mCm3Gx/ZEp1JvUz+cSvGBUZWDpNu64FteFp1ayUyx08bKYdpqOwm2Jr
DAmuThFrxVf1ONBvuz/A62I2qQTZQ1uox3nrujJ5ZIBINJ6bBlFjenN0mawCoglx
Uh1WbGIjgzhAMI6MVc2MREPm6OIm2s+puHQdbKMApAF+ULai0RbFu4z6NdXibZcf
U+/oSjuIjzZeZCgulWZQIMzEwG1Y8SLYLPAAzMmeADjzT6E2jvynCLJiAzK/pAzY
xWvfr7eTZm+dinysi4CBpiXmcLkB13bc8oiJGsKVc1NEW0easOI5VsIq/u+/dOBN
xlCH1SJouN5MjjveVjcEYaCSqPUT78D/uUEGKYv4824rQfJ0RpsFF/yYfyKtyOMm
vrPXv5yhhEn3u+tsvAUMhQ/Ly/2kv6zqn7p/rEbfd1z6mrbdBur4s8k+zFt4HKoF
sDOIY0JAazwQl/dOVV7jI5+A/LGCoZlb5F8HIRHgBRWGFf5Uj7ZBL7sX8+Aj0IMp
Xn6x/zlvAjcwa9H4AgPyKD6JRKH+Ues/nuvJNxt3IECx/WVatMltUR4Z5z96Tfeo
t7IP+zHbvPYZlEoj7N77WkkpB08i50F0G1Nr0Jt8dfUlJ545pC1Ze/eg4cERWpJ/
DlvJTy7Sw98gIdF2tqRJ8G+i4c49okQSyG4cJo/vbS6T0cTZ5LmJ0Z13miPOGpkD
pxaDsRzKgNOh4WdP1rLfxWcLBGA6lJ1US7b3gB1Ifk9TxHWYV2ptbPbPdooGAkm9
eRwAdGVC6zUl1KJrOtQHOfkPhiGSEH7dMvnnZyL8UWuT1y/5hOQ7/yiFEUeQU3Tl
6OscEFAP9drMrzCIXf0UzjRxmNkExtBwLAh5HZlHGTAVNv2yayL6TP7XvYSpCjm0
MotvQlJJjFnRA+SLbL40oahLcxFQD3N1ja5s0xKNe0bfAvJVEPr230OXdbV7LbCB
8ZC7c0PA0EwopGn5kIXQg0K9bcnBzSkEuRJ97/7T2UzAxlqulwcMOSXb2hQrMwBj
Cibw+DWtdfEmJER0hLDJuvtEO7W51m+aNmpHYHwauXoWGB7OTSEsH/R9Y7Nl523a
5TcuYQv80Hbkg09bmuEU+7CEmnYaGIavTrgOkyGOFTzKshMjbCZCdFhW6tpKGDwP
1yZZ3/Iuh7x3GGi+3Dw11oYPZ6hQuShyJSVvE4NsDr0geynVkdFbd0EBzwHYNtQl
9aOQRfSsx72/hrE7fDak0P2lcg6BSgma+/VzNCt6sCvfAOcuDSL3Ef8JedhUTTh3
+PCoPFxFIP2baS6W6tvAxZWL4Om8P4XTdD0ZyqO5CPRhUk2NJ2+/5wuuKPS4RlE9
vMbF3SFPEKHBCWxv31L7Osj8OPlC6nUnxnmTaUBHrUs7JBvecFFNPpth4rAYnFI3
HJTJjA7tShcfsGqMvVIll62KIlOriq9F9IHHKuagV7BEGHljkvTItvpUV/XmmZVd
pdjjMY4+Jb6jaIJkMWssxc/YdG+5NrByNqBj746Fll6+tN84fzv9q/y2JWlRwflM
Ywcnzq44+fc9aZBQI0u9muSmw5HO7PG7G9zefecuphd9k8e71moac577+qm6g8Ho
to7SvzEKAStCe2gQSDi0nhx8YgQT3cS1dzriW7HyDb3BHFmejfNSBLqDzNlCQhZ7
HYuoCSsUrpTlkRnQ4gWW1RDVwRwnQr385SVuBAia4wsVZujHYl0pKUiqhvw1sWw9
phqvf6/beDJ3h4Ltu8Ntb3Y7qN3K8Xe4lRbqL7fZd9BngD/UZZJ3nZ5cQYJEa9hM
DpHW9uJ+aFcgU6u5h4P7fhkhZKRqB97lBV5aHNxeUiPbKr2xU0NfAQ//hern64Rb
pv6IJllZoFNT6lyBPI/68DNPL5Q5lrxL/Y5d6pJcZ5uWSVpN1Nugbsty3FA+rK+T
IpnfhfvdWafvHG0zAS8+Cl87Usksr5j07ABjbMrR1GH/+RjD8qgG3j2xlbAT+g9w
D1mx6DqwxYU+V/E7hknkNNM3josgUpSlwi5ex9JnDTuonc46gvmfLtaFdoAkSnph
4jfM++uLUtYddeM+dnZ9ZrHI9L1R/dgMrMr+QPcp3qT0qRBhAg8XoplnTlK4dixT
uTTYgSMbqYdVp4ukW05XRsLioBCUPJm5iStZ5tDYhnQ0oKpfQaVTUVnKNOJRdDmT
Z6NbcsRCsIJmBXxvIcVQVPmccNv5obL3GntWpSM0UfmehrHqogRQYdAm8bbWJz/o
6iN3lmfKMYFQi1hOlx1/SEazf9jk0Teh+bGhoRBYEayKKfwmxgM/odRZcTzp1e9f
ZphwcskWnnz7gaJ8krOt34Er/qt5GO/BNJZ0+N/eOAzmlpLijeQSWZ3oujM4/gVU
CQOd419altAVx4RG7aMVyVoXPqgT1/h4dqOlAkZZcsud20/BdiaKBNY1aQIApJ2z
KYs4yCF0dKhN9QnNedzYb++hWts51Tycw66OyJtpTnAt19e2VE4sFCDHGbyHPTrP
kFTc/6hJPUix4RBZuANa3c6VCIIyxRd5tEuTWfeAs5LYNbjd/07BsFoduls8jl+a
cUe0VQcvcphDqvZ93EuCMlQpOHr95iJ7Roz1l12M1ehwJ9OSD6SsaH7QzutNDlzt
OlsEWRuDshdym4a75Bnx4n/otXmGg/a9r1eI+gvc0aAH1xtp/m8H+l8PWATmkMqJ
VIYVMNhIGBHk8caeJymVjAkWkgM+UK7lrHCshDawsk0UDTZLecS5XGJcx+Rx+Low
uELPWA+N/6srpz7N57B2jAQQuIZGiEhoZmQv7kIYTllzUWJxoj4dKTckNnfDZ+Qp
WBqNPcwGVWEWqFSI7oEA3YgPqUJq/3kTl4856fj38xTYaiDGWAatFVnZ0Cmbj+U/
BdCHKLD+02qiiU6XdSSKtjD4gdq/XBij0t+eqNaoMAiVRLWxN+CN6xrrTH35Yzs3
xOEtmJZ//8RGDb1xSBQguSftKoXrMJ/PJWCGubzkbyn7uyZo+9hbwpH4WqII4dVc
FiiGNqmPk58M/ePdY6eC5ACvfv9W5Bx/2L9Qj3eURcoX/cmARKLsmRKA4O/HjjvT
JfvtTlgNNUzPs2lhjOxDXk2M4I8xvIpasFBhcYFNM69WYqm6++pCagF2YCKtHw9L
ZwF6UGJ+rEGMp5Lgo7XoxmGoViCLnqfJMZY92TpYWvupVbjsKuCmDruqNIzPQm+8
5R5FVchpGQ/HWTf06KvAvhJptzQszhs58Z2LIu+9KIgH8SG+wriDsHPJ4c2v/MHH
oNQ6kHIj8Kxgmn0b+6ad1eyTPuYEDm30U84P5Kfp0wjNeZ7hR9i7ul2ZyHB4zq7F
oHJY03sWNPKDSGlGCtAQRkMCSnm93Myg1nSjeQl1U9fUHsI1bYkOlqXrDq4dyOF+
dlIDWBL/U80viB/PfRM/pzcjSMEPeMNENnq7t4Lp1Z2V5Zdbh293ZyCoGfFI1X8e
Hw7qmAwGSH6LBJ447+EJTVSeStiej9579p1CUfih/19ySPXg3CQirTI9LF2yTnlk
Y0B7a336v0NKSURjwPU8xwNeDp5Tqgcv+ltOEzSxhMuTPGM2fvLbD2K0X4iMdJO4
OINhsxhefE4HRkpygU/i0RHJCSofFyWo2aB38n+8mdIFD7DoCB3SlKV1kfhilnVI
c3JD6k5JcgIiS7mVchOJO8itW/7+vDEFzkiEkdAUqwrS+XBuGnYc6E4EfHgy6B6B
Udj0FntzaucYaDf0C4KS6GA7xpsmHlcmgJxGfcr1AiXCVdX0ps//RVg/kOPovfT6
dNLPVKmF7oskbR/daPc/BHIvsB6+M8o6JlULQo8DDKB8Xd5GTQbqFXzR51UK4qEP
ukTFQz+0NtboJTlLUz8Sc3xH8HL1Hr9Ut7hSvZyhRZ9aomunFYQpLAixB4/dKN9p
y62xRAWLIRZZ1Kakmu2kKQn55kaoHsqWAsqdqt383bjUIHgIKddgZi1opK/iHyVi
1WGQr5k0RPCD4fTIlavIfZ3ycE6b1FtaantsQ2H6yhbsiLXS652ZIeBNNximcIz5
50ae1lpBMWeyCC+epJOx5/HuUZoDO5hkUH2Z4goqcs/PkkuKG3YT+q0zXCZdKLpV
cvtre0zTU9i33y8cfsmDuZqJsaBiUyxwwjbSEUlk5JF7Q00a1lqTaWQuSHxxrFJA
OeWQ6COohcwaAPm1zJ2DL2NcM7HS9jjGkyfQQ2XkIKs/NeDogmvaEl0wgAcIw0qj
7Jt+ude1zwV2BGjTB/zc4KiJh4MVTpkJua4F7+k8e/L0D/wkISz6+AkF6UUjTOdC
TGN5RDwXER/7xOTYZey+gInvpwIuW6ORWiU40pPAIQceHedLDl071f0uh6Y4L/tY
W6l3OXNnanJgm1jz+bn2GYRsg5F5xopYy0ZXkDG4xXb+iR80UmtRFM5yETDG1wv/
6P4WdWC21QF9nG97f6XpJ04dv2Q0PYYLP2Xi+4Z4JwJ+LGPIjnJyUQqyVepz6eRl
N5FqASrO4tVjAeb0Kz40gaGPnB8al2AtmnzhjjW3Nz04vpH8smNXMBPnKKQkHeO7
GVc4wciA+jpETChhm8YxVQCCJzh+CTOIgiJOQOFNkTeV03jVuFdD/NbiMPM51TbW
Tqr5Qo4uEMBFfWaQerb21Fel4/voY4gar+cWn0bt9rJduoO6WsBVRF4VyqwZjAsN
lYdeU69fg8whoUWNsO1GtMNTIUbhQ5z1at2xiqbDybo9sj3PpGOOD3Udd841HQzu
YtwtySgH/Rh6QErwlKQaCIbqO2m5AouzQWx9tqkJALaZ/FdjxrwRfNQ2V3Sj9lCs
m9aD3t3NyEOplLF5KFRWEGLsm+Jt5Gitm0OWdQquWTyaMzI4Ascx2cjQiYhKw/3r
oaPE6I/Eux/CZtKcIjfuTpmb4PLK7H8jGPtBTHAVmUdsxhgqNNEW/oXJBHBpNCTA
5VsnRHdUiOv5DbUGQQCHzvYzR1lmbifKmGaLw+FtOOjamqkOJ2Yaeoc6M4rzCfLA
ihtKtqPxefrdKQRqZxF3oSUBkX3k9V+8nQwwbH/77uMA0W1cYgYZArJTakXX0cag
y8WhIb/TMw5U16hTvuj+MeTTd+TlPhk1z396xtijfo1BWNpzqfHuhmkzV5k08vAU
F34HcnmdFpo235yzMTtjbr8ayN9/DpLBmVsDV2cMAeewJ0xOfQam2dmzM11p3bfv
5NeGaVafq5CZx1WWuvWrLrNiGwY2NEpJo8GtWIvSixHp+bOVTLjRoVKjl3BTSLZO
fhAHQjGjsQmiGceYT/kbNRBSs1xtf5W0qGl1wxzRisxr9BqVtAuzCHXY2QgUy5Ux
iMZqUjXhKEyhRumZDT6OCxqmMZrSEeq9m1yoBWeUe4mnTtGCt/v/kTaxWYUMOa9c
XfSIJOGXqYvp4PvVWLEvJdnWPY7z7cUHBDYmkuNOIYn4HJKTteGacpX2YEkDjveW
j6+oy3/9FTdUKdvnVrQhCdv+6xRJ7hoCtqRbbAVjV4mTUzs1CLddsYTfdse0J9A0
TLidx5Wyu+Xs8i7eQhnF/UJRMSY7H1cDdfe4DZFdfNkPoNWMlZKbPRAECA0rY3su
02HnhheP6mLXWC39vmIqsKq1gMbnj4Sa5k08YJaJaz6z5WKMX3cmn/N/C6yZ9apH
m+MY0GIDd0Uzz+qEh8skRPRzYCzX75WfUSI0SjuGt7MJKXWIBpmbeet2zCxX14l2
78whhwZ/qtph2xYSiu+dY6/0qTHQkjoNfIZIE+ZrUI0t+zp0qC/QGPVmnpigz3Hn
Hpagzb16ruCn8TrNMDbkjYihOR8FFimAgPdLf2OcBKsghkl3lF+dFmwYHn4k5gty
QCjyuFpk1jyMliu1CG0i6AY569ptYZpaM3rDkLXfhrTP0qgrg02Azs8wyUmkY90y
Bh2CDqhGvqII6ca9PoZ+oeMUaul+yfxe2svDoTdQ6qrCij8P27y63B/s6bWEp3YC
vEKVXtilx2DRIyfBIMEeHAHhk0a3oRCjZoghNOdxSQibtDnEqhZWCRt/2cTLJjyd
ocU4qDxWFR4ufllhg7niUIcoHpdbwPtX7u92zKAtqApN+QCSxGzf3vzhzeTlrxkh
zD7c2GKtxEsDYDv7tsAGgSRy6GLZV4HpOdD046rVCeGsTS8VUSXv7JyBHH/y1J2/
sq/hW8f2E9+n+t08K6nDJQmDsgXYuLb6RMI39z8fDLMznyVkN8qL+16mByOP/+l0
UBubkknKw95zaSDbrlrgmZa43awOm4MVk1J9Hp4Wd5Apneh6i7w7FBWaFValgagL
5VkczFEmWcsfuul5I42X+DrIs7yFwlNznjv+QGTDYfTsA7DMBxGoMXXMzx2w/go5
/rMIvDOcipqQ0CUsosgaZ6+3Vs9AhmVsIx9Bdh1QuOqTmNW6rMVIItt32PPbzui7
OxSBrAkSuR3JgJPHF9kSiNlDLCdAnLoVBRGIZ9wT1uLgMB+1rzk3SWSDDaHt7x40
IIA+QaRPiyCkPbV/Dp6APQgT2U9vY4Jrq18FI+7fXyhCsJIXoqPa9k0ksrl3wLsI
VOsGFyP3f5C+iNbIzM+Mvd2etYs/U+WDeKFFyTkBejpzJUSHVcgTDUWOqa7FYgqt
UTLS2KUyMOVw2dSDfr+TZW8Q1ZwVBJbQB4SlfaHEFhAzCO4zU71wlVV7XM+9kf9a
rgRNrRFmc91MYJoHDsc+k5DWahEjJl99Nm1FokyLR5aiDNWb0LnCAo3geQ87W4u7
uqVyl4k7jfMBAOhA2MxbdliLMv48TxbELXXhxeBUVYLXj0HEUP0s4eYSs2lhsu5S
uacFk20bYWxoHYIsyyS3B8Sw7P01jgaF0KOVFNYeLsZVNvWtEcHm2a6aP3IpG7lR
L8mg2krstPvtqzzij17L2YW9Vlge5oxzpW5yNfs2VQBUgEHA8zylpbOCzZIH4mtU
A2lJGXY5slT/izGkLZqbbqAjT67od14YWwpB616hnKfgs3a9N/o54SC90MywsXRW
RURM2wIs+T95P+QwTu5PkJ5/1+8LTSH/0VEOkU828QdjzBD/Xy3tKuMt8UUTUeT4
QBriojpMeIzg2SLxCmpZdbG6ERo5D96xltCUEdDtCI3aEc4pum9YcE993mBRNbSn
+mdUJoK2Ob0Di9XhY+ldAcBUyuv0btoydpgpEwcJlf/zkP3fbHLQmzIDKL7HoTCY
qn31sed5AGTHpAoCkacos6Te8nCZzdTvvm3kLUs8O09HfPCdi+KhuVeULUyXeZQL
V4uqHL6CQn3FdAb0v4kHF+1WWnjco1IbSpsqKokPSZhOH2c1JKNGuzkHiqOuUwL4
4fHCWjz2Nrqt8gU/+cQye+x3cW4jcKi+nA3fZmwIY7xwMzTJp40ka1T5VB4T9XE+
qvQfnaQ5n/iZzgoqYbBB2GkQuh/e/9hTp6KlVbkAOp1Hhsc+2xOu8a5dwpO5zQtq
DrbcxccML498qWXTLWFPAKaA65acZKL6C+gkH0bYiGCRBTHOYKkk/G0SoTtQxx88
EiJ8Xh7Hg3FvqDAcYbC8ujVgm3uJDVmO24anaerIEH+LqbGBHw+OO5E/6LxkjZ+7
aWG/pOKaBT6jci5eLr5dw9lrPo01TFfEBhUTmn0GdfltNXJMFz2eorjqYdEw/Dj2
nTMTa+0Idru7WCOp+DnG69TI6TZ8FiJCGtI55Y6vnHJGgo8OouEYGGqTKHD/Dgpe
q7QY9SJZ6HVJRBejT93NEUO9dukDfETnqwZ5MfzJlvzik5kx03WVQUBeOOUoLEij
MOODGldWu14GNl7W64/glI1vMrK09tMtgPly21cMwzz9CGREMRBFlTFqHHV0kEAS
RXnR61+/N199FvMtCyIrvDpwIVNdcsR3f/qB0vWJzVUOwpDLMAc+2sXInXtabMbS
OyB7tYZ/2HEl+wyKqAHDAfi+4PZIP4vluufVdm6w54513ja9LxHMv+s+GFFbYJdd
0c/D3b4a9ZRSwPOMfQkmlR9cKMD5/2jyWIpBHfPzB/JiPxywZlB3HOjT3+HAxGtg
GW5+uxpFkDxZFNiGHJ249UFYq+looPCJdz3g6qHboSwl37HycQ44i5PoaxtK3b43
30CuCZbsFKfBWzezArEyt1xO1RPZGP3aOjqmSE1dxV9bV088wI049/D/rv2+wiCW
pfohxWQX6tBrqonwomlDRo5ckhVgwLGiDGLzLDXJU0Fdw+rZ6LAmsjy8B77Ytc9e
NzAiuuJKoywnrQkoq/zpyWXH8ABu8TQBUxuvn5I5JIdhXDH0itDTHDJmDLyT5qp+
oxFabX+oU+Y6eruJmc58GwQWcX330A9l2gHGFstRiIGau02NKoMehRN+Gxg6El5s
utvMeVETTEgXpilVyoGOkBkzv191J39aEcHgIYwF53i543bT49/XkecQaUOqgUb2
VXtAZRueq/0KPgA6AkQ4tm24nPybf9B9XLj0Mqkfgj39QhCo7OY4GXMSpcQjGiTF
dQpJYaIFAcWDmJ6WZYeg//9q8tzISrkmFjoKqunPDqwIPXjd3YQeriFu9DUHLZAK
eQf62ODQBL1mQN+ooHOoCKlHLDJyIxCjnmYrHIcTwsGUzKonA49KQQkQGya0Ulke
/tMQYmWKBck+tpmL+EXrSnRb6bogpXrQqKhbQP2uxzOaPthbTX3kCPxzO6sbPn/g
6syc8Nxqy+Jq6M4Wa8mHlM4hBeTYSrgNLAkJWAoxntlW+mwExEzHUO+ttd0sEmRj
tQpTG6nuKC0ygsFee2WmMhcy4dG+LJcKMKojfj5EYhWEvVuZKj+fsGDJSEgQW5C2
vLINf82C8tAM/ivdFlD9Nnb6WoP1sa1V2kH0ChFUxFpQResP6NGAoxUjEu+xL2ci
wEzRZvgZ1x4nwoN/bwqSAR6Q2cyVSMwEcc5Hqc3ycINHdyK+u8Gjc4LDKW4BWOUz
fzdFVLJ40tODEHNSBMn6oqexsfYJ0FkjuYwynEsGk9abj/E5wi+al34kVIVMmNCi
cF0/kbzwFAAOntKQqhYnJp9JSkUh6d6PTyv/dyUSyp6UD/exH/qKeLhJBW/Yvjhv
3IgiHq+6LuP1lQFG4y/c4TGiQW3B5vDijz2+uqp3/E/YIM8z5cZQ17zVDteddZZ8
AEn0K7yqRPOHmdZwmob9Fi97X52kMqA2M0Sg7jqwYKz1bi7uRRfUnehMVtd8PKRf
ZFFrMoL0+2wE5Y8XEuldAxg+18BnVvPc+LwRwGVrZF+jr4gtgmtKWGayOlmHNfiE
fWB9vpzj1HtUQnsP9xA7QHvx9/ck538AHGJr39vyQeFwyOoOEGOdiR7nBA2J0u4w
OgAH8PZTCBUJJtp4buV4b6l6Q1TJjSuMPlk0BB32dooQx47Sgq71g0O6+akMuByi
ywq7Sm5mn+JHJkmnxJppjA6QaxW6CsjjC9cTEJUSXucb3HaSdc8uOHfT9LOZU4Gp
77x/HDJRPH4xl3pDnww4z+PAstNcdQqPzTCOtF4LgRxlo0zaJInnt77dKB5d5+Cu
oMlNl+UF2TDuZn+K/j+CyAlu/A05o6O3qYFwb00uGLPWNVFpnZ0VZF15hzcqKRc5
DO57P9XEJ1F0EMEJilcGXcwQONDp0voWR+VbEIDbIL4RkHYqboFnsMG3NA5N6dEC
DHyPMapCRwcP2gutEUE/sxhRluSQJ1ZLAD7IZkCaToxEMVNMQXvt8BofBxSVGdcz
LAvTV0oknGx40yULXM4x+Ssy2y31ybvi4zXBVxhvws+o16OmBl3yqwTmzFpm7+nH
Sb7423GDSDaYcog5JzWUp00A5h4w0Y3ZF9ksZODES46r+jsehtI0QdfnnotLyEwp
51Qxahp7X9yUSjKJ/xQLrIc/3Sn2g4o/o7uCNi1ZmucuUGGDM7mS8qugFL7PCejc
iqN6O6aCtpGkTf4UzIyZDStylKFBQK/2rqpfYxHz/2SPHzsDKRh09kaVEBfC7qpI
NqlAzf4NnYQFMqQ3sSPDbKFzJwp8BywFFg3DeYnB+IYZ2DvozGPMGf3TfEqz9ZgO
61lYfGUQ56RKkqST2a5WkURZvNYuURj2rUBWl18rc2Wkikk+OzTDwWKOcaeEmste
hoIm1EpvJSsN0uGQjhh8zp0RQMoZZQ4XZYSjiEC/fXS4XzYGfDGlaLQl/KsBucYo
Tto/Jb7kbz4FzxX9LGbqktRXk0F15Ao4/DMQaWTO8FnnOQaYjuk/MQM7cHhVIJdG
S0SVLGWlQvNMGuxyyzivPGw+ca8jN3RIR+ewg7y+1a3c89kQqkWsiVQoIY0ceWhk
CH3dSVO02s1pvFdE6YnXTgWRDCsUBqsxaDSIYTD/WfUSZKGE3XMEX4XJQQNUZ8TJ
G14v0cuk+VD4A6lQn3i866nQFDNQqIy24aqwtXAUCb4tzsy0Z9XEUvusjpr2DwbA
Bs/tjVcYbl7c4SnimPg72fx3qS49/+o2NmIo/vI3yq+ZGiMNngbQ42BbG2GDqP93
z/HqkLu1bixfU9eteCVaGGy6nKzOlMKYCOUiFrMxDrxH4dHv0xb2CFtKdeNo4cKu
pJbcG5zn0lB8XfZF2DWwSfOw9R5nyN/mtTRSNBZIa1uYPBT21+Pj7Td7vqexNfd6
rrFE6vsQPnh+kx+JTLDeiIbQ/kZDl2gCem0y/nIe2ucayq7PVzLgTKRGv6yYXlZp
eq1I0kCgvug/B0JoxDGgEde/nZmT/K2chOAYY2wD0tMQ1sISbKJcsicUKgCDeuTL
WIJfySELQlJM2Zdre6N9xoFkWRNTscPHF7YkJ+HKAX+u3ggVLU+OJb0fsH3BY5gK
gGaSkqZApYRKdDUIunG9ZtCd9Dbqdy4LixUuiXF/MVQ1Aty8ZBiEOKkh/VPd2ZIV
th22iWpe2QLGaj3179xrVgE2iXTd09b52d0Sjyy5Wm2ug6T2Lf6XPD4G+Be9zFZ4
5KJR7FB/qvJmvxkW4U5H8P747A0DxMFZNPL3LUTHaqJ15A8r8Ml2RvCtkfwSwEqM
rM3ynTvmaw9MS8lShtLXXwaihX/Rts7B1hreAPtUaF/TRvDQwTNghcOa1cnqgUbI
38YrLJMZnoEqGEXY0Ow/wHbXGLnFOtXBW7HmAyOFnQBGupaE4xQoO3GPwS6wPE+w
D8pAByL/mhQ/zUp0WkHGcX79NKm1uMXrWHoXTtoRbhrapFaJLD3C2ik5USAUM0kc
lZ8/FO6YTiKLhvGr+Thpykxo94jfpGSwsUxneLNSB1ZbBZv6AkY8KE8I2yhZnIWE
DmZzR3oigTQD4yYvE7cqCHNXRYWgMQDOzwaUMA7pYeLibZjWV8eJKvWiEIB1CCNG
GDcnCotkDJ8IRBcUPrW2dGuBwU/MaZRUgLYXfHBZiixSDlHd6RNgvN8v+6eeSPth
l7jBqzMviF+GB6A3nLdsrC+HgcWOIHBj20M8KoLDjEdLEpJOZn+BDNHfCHsAVCC7
MPNdK8l7in/G4zKa3tXtnYWjTzGNw9wh5H3yOI+DDriNk+SPpYrJJmdmWfNojiL+
+tjWpAvqPvWDIJSAVh80J/NyU+tACoUa5S1wtrWHYXtrm1HhqtSQh3gYfer6mZpx
SSECD+z4qRlx83SyNgssljIixV6CqJGP2pgmUPjCVK2HQ9aRdlgBaoAfHuRaCYDt
LFFgNmCOojE9b516SPvBh6h29xxw6aBqkWdZOgwuAjcZeH71XlTrk1e8uqnPqGXg
eqIiaAwsBzy07b5JASApw63Sv1OGCsbdwCq/pUJ+jcnFOa/4Fh9QjMisPeSZgPCZ
53YcWTNjco+Ym2RIq8MRFzaQbmEoxMsnKythKbzwdaIRIoGDJum/Sy8wFzIlJrH4
ZgL8T0vKwgnrZ2PV9JcadUTIJcBFegKE65x3tgdujMMGkUir5BDL5ZZPZBvUW+Rg
nFMogxwCNwicvMDFutycT6Ww7TSmLWnKRiD3GjkIS8KZ8kNSC3vXl47N43zgJnG0
S8mKTRGg9O+mJZSwlqQtt37kW9AG8yuj7Ai8oev2KTq4DTIU6erCAcCzOOfW4mCf
yVkLEcQrkTeQ6s/I4daTB0rLj7iSDcBJQvCSgS+VCrVpWKAUAOudmO57y15q21wE
RLGmwX2JJJ82q9gcX43cKFwTcQnWBAwW+A6ASxE2pclR+lj3hV4YfnGq65Cgj4Iu
Ovwm+xb8UYEpAsOEa7latGKi/pW/c7GKcJzoD4WOd+uFwq/6fbpq3415hLNlOeg0
4p4HE5YCPtzDjtsBXW9fmR18AeIxx7rPQm+kVbxOqEIEWybo6AfT7yuXLfLX1GaJ
lG+wEl4Y1gl67CU66ILJZ0uuV/SAEPvZ0sDrssk1TFYij2YhW2LUWKmmOhNckS5g
y6lbDQC4vXRQ3mSrQ9GdTteDgll81y0OQpzRYVW9+TjzC1Fl6WdLKh1zPJmHlap7
kLlT56HKIrnlPRSo0GE6kiqTkQbEi9Y9LFAzdr4R5f9qYaOA7izmAr857MKMEjxL
RlKK9PIhY8t4Y/Mj9CFYlhc2lJSMGVzhC/2MUeDlLv2DvWHyhlsG6sfSSgjJRv8N
lbOUHzTSGzTMS8637YkXXpsZ4I7dc5/d3AQ90iou7dq0NIPis7npNnhSfVzlgMFF
H98QPtNtEYf/9plnvutROcaIWCF6JhUFdECWlnOi0SG6RrV/LJuJEKinopKrgCMw
+jROYsXGWjk9X/2wkw8TE2UAsYlttfu0MBQmsVFPQcAvHjlDt2KNS/+cwwF8pubz
yF9ydrCA79pdvpBEt6sYq45jrGrxKpJdOzdolrfwjoOomAEb2/bpVcDG2f3/wCuo
hGHUevwgwihZt9CueYQoLgwMLlEwCwQwEZ3WaYfIYAIlC+8rulQ34OQQv5FAdoSd
j5Vujg53GAJk1mdb0AkEou6Cm9yCIxg9SJX46EOOiFfpgz3vg+Y7f4YkObuJ6c/K
Qr1hNy/TfYAfW9Wn54dAyt6zVfXGidH1pRgP804zjZHA59ED4gTwPdUlI3UqckbS
zNXMCx/rxqw2PxB7QrrM8MLOcIH4xlKpwqOrQYOv/ScXdIrIp3F3CaeX5CAww5Ov
r3FvHTj9l9xTTni4FZPvGXF1IpOWeLX7QUG2FMgRlni7aY9mwfmOyLnPEu8EOgk0
qMEtfPjLqvbw21FkZtmHhgDkM/pB/DeDdxZjg90x+aVGjzRoRGahZkynSXGSPCc0
esNsM3IKAekiE/TIfBgjo5r6lzMtORQFik7tJlHilrXNHdfWwbehrhqfAq+QIT+R
Omv2ylGajwlAeHMyw4HkQb6/EYFiXqwSfeXcFsZb9W/R41QS5PU049sODkxAOu3k
k5HnWrma1nXWSza1o5uaM5Imp1Ic35crb6LREbtTy9btFWAQITq/QyJoDSoeOYfC
tc9sYz0EO3YoCVqrPFUs+7MATIEt9Zf8o1/i6+M6lEmybCdTX4uI9rJ1qzDXMvfu
pQOamCStV8dQvE7bEvEX93wFpo59at1wj91eNMyl0DRKq7iK0QMHn9ineyxQjKaK
XU5puJ1d4AVJEU1lL3q17mbxrJUSQp5QXLyRo1Ky3IkjKwT9FicPmGpeHMOVsWtt
dJEMkoSBVey19yjXgPACBiqc0lG6S8KhDjl2DIgXoQrKMp44ai1fpPLl7+BlDSyj
mUah4TcPlMDKSAe8dBR6BJxRQ6qxzCucbRvjvZhW1QDuojg/LOzyZgeXH+unag9F
dehRjTkoFu5LURYo5TicU+9lO2i+txd+5WHnKFUTdO20VpxTZraJC9GkGpSnH72w
peEvlzig9+k6/mqAFWs1/aGhbsqEUW5icj147eFj6w7+XKOIWyl3NFEUOo7VzpZA
5mYo9wSkRNJRT0hY8vc6Mqux8kebM377UYQ2L5mVWxLBhGsNmL8gwi0U0wWdYZCj
bixTyiR3pvtyFkHpbJ99Q1kw6llZtYB050WycIGZXVY/IQhlZOdPhowcETp45642
lv5osg6of0PWzXvCIhWo7zp90mTdxINyxRgIr339tB1XHPfKOrlulToHfWSSdHGr
xmdIIlFOQbOcaNFDMfE32QVzMZtaxZ+sn66yGHzHodGf39uMbSgfzRUsQpnV/h4e
FNlkgT9D/PTibC4/tuOqymvZLsSOws8rK9EBPaPd0KF2aTELuXQo8ummeKgwQ/Nq
c3YXgMD8yfFjqda1Pdkt4ZNJIXtU5gjtexMxluZRpFajFVSYU4hVn3vyKXKxNhUP
3EP5L+tHZjy8fRII5wKa0bgojTG9EVMBtbkN9fmL1r3U0Q9enDZ7IS6rL7cUH4Qg
S9iSkc9KbIvUTgvY5dRV9P8y8axK/nKf5G3ewIqwG2CG7Aj3enjirCL/RpNcr5R4
d+rQaTA5xqxaYCKRhzLxvlOgL7SXN5S0bXiz03OO7nkRsL5UH3ozBnWU/vjTRWbg
nkAT/LGg0IcETI+tR06O0hHRpAFq2Z5q/QHz+NP9kaT9A1W9IhRWZChnwGcInPXF
Vf1lYyGV46aKILtw/Uihoc5tdmJbpiNFcf3Q34GyF+EGVOZHzoN6OcBiR5SsoMoa
k1Ih8UOi+VkwYCHbgCnR3D8axzgV6hZH9n6BgT4gqq+npqs8V84lAp7XSAoJDXAc
0pU5ik2EPI7iFHpxdXYmG3tx4XhKSuSh/x3C47YcxpcERZZ+fQS+nEL1djR91hlX
QnHpbP45/GlTfl8eozwyYsoGyTc4k4CHHlMXbnceqq+WnKKIsrLcN4GeF1x78djC
ouTCtQHifh6P9360GnS+A7Ld1SUULEQqv7oC0JhQqfTDhk1mHUdh4zTB4srfL5YI
mdhxYgKB5Ma5UTnFo1JtzkaLCPB7Bhq45fZZWVhY65EfDtUAYZWQBd4n99vungRr
NOjeJdx9axja1oqjpUIeAi3janMF/hyk9a1UwoQKPWcY2Fw2zCIbraS2dBN4fzyJ
azvsyvrZilW9xjfLDwemK97PF7IEwSerwrDAH5QP0qTthVkmQ5Yeref+HTvlBG6+
j5vOSSgxodpwKEsraync6NxQ3PpU859gQoRYfNlt+0VJxvdX1kCqbVgr3SZKXS5q
WJwS5q/Ly4wGwxHe8hsjqVxrfwsePYFHA7Y9D47iq71HlZ5xtatEzoS/D3HUtKki
HNzbWLhcPJSqKhNsyhv97uKrHa6tk3D4DL3Q32EdqvH9kwdWc9HXkJuUMVuN5xlF
GLteLl11QBMUGnFxBKViFuw4Oiq55EviM8PzCuhXmrmgQWjIUvWn7OZS9uKYgt0N
/fOPET0P5ICYxceoAKOTON9v675BcuaaLroKTG6w4PUDCzu82UbpxWyL1NMGP3/z
p0M0TjSgVKLD8WMic+YUseIfUjDAVejaAbduSkwyjkqdP+V+yJIZjKaYydQ49lwp
oXxhkaoZiJCBdHlTolcKltLnAR2eFuUELIjljjc5E1RzzpE2iGNRaKuFptXphAKL
IJcCZYWNv//rrr6ZD+SK3oySkPepyldrr94RvAhW46KIj4WxmBp388W+tQC3Ri1S
ml7aGmw/ZxBi9+hhxcpbAVkeb6t8/86nPfIjApCoTbUQFTJh6jy4G07XHvv2TeaS
WT/CkYM1BRA12u+P9fPaOTobhUCD+OKFhPnRBDANqM/A7duGjmE4youAkK1RcN8R
m/kY1i+GsQN/LKIWo36xSqSwiZcXbroh13Azcd+enviOEY5K00kutJ/oNdGGLDa0
DVV/GKBdAf53LXIjMCIOybcRSQeMOfl3/A3rHKTfpgHStZoZd7QuCiRSEKB44kS3
I8YOIlyOOO3eA4cSaVXORYvtsLIXYpQ/gFbkmovlDwO1If5v/7JuZcjf6mlh64bR
OjUYqFmmomuAb8kkDL1n3ylUhwHhZkNt5apxImHNWmv1Zxuv/HXIErWLUV+6bJuB
+4bpnt53u96qUuKliuUGPI36nkpYWPcBNK+BbjYeRe4gQBWdJ2sTzEWrznxw2gnV
6nvZ48JdbbQdMDwTyEC1GzzSyN0f2SUaXCwc2qNe0n1fPK1GOEbtE0Cj+Lw4A5GF
7roS13K+LjLX09WrZV2kkpD7cxRqi1Bg131/r77uzIpnsBrWzM2jxqZyxPvp+jZo
kHrbJBhVl4F9IJUtMyxQR+S75l3Hy47RJJoqVC1QLNjA1NmDOXFHwIOhIikWOCE8
D95NYv0ea9OFdyA1pyFrfX076G3cv1RHC/uaNHTlIXGffwhPF/WI+pkPLqeEM6Wv
rQwPVjYElT/qzY5p+8HgsNWZ3yNczYAtmLeG7LJiGr3KMEhr+vJtHZDS+Z1+Tw2b
MuOtXP0+IAN+fggXgahkp5tJQH2QKfMEjy4Ryp2CxMuL5Ar7dNpCB6Zu99q/p6v6
BsxlSgrGJHRrEaVl64UNimbn10r6xTgnxtrwIE9IDW4wkX/5KqLSEO+MlM35ntJL
AMBQkXCrtz+ANw6RPPbk9rl0RcyMjiBjRWiGeuojp0eR20b0FwfgRErV10CaRaRu
J5QskfJI4qzOpfF7qWiWjHs/iOYxbe5bCs7HZjxENcIPT8bzJPLsdp8GxopJZKdv
huokTqxlkuNhTzALOdAEYvL+qEXXNGCa9VhBu2kGVowKcqSoTtVsxiIXQQnWecO5
sm7/e+tOLPffzqZnRsEYP1XKdpyAbbB3oou0qqemk25FF6PViZ44iz0gizSsTrPv
Y5JVwr4fkmn/j6dL4ifSS9Bapx+DDPBxMgnqDyT5T70fr6QixCkGZ2rQR0wwOQTX
LrLZnwmjkGbBgmWUuOPXfjkNxTABMqeL2m4vJ3wSAJN9gKokVtUUpGR8R9GX9qsA
MolTMZHc5cY27p8eJt8JwvX/wHsHlg2fyLf4tt/vTEsqYKD6/EGO0JVXQ6tNKIyw
aaX/NjPi25YffzBgcUTnfeYG7+t/boFw2yst8ru+lAOW7ZunOI8t2VRydstPHMSW
Nd58OfElhh7lfy6VjIz796HRc3N3syHEVoJ4+KNozQlcx3mfoWayRzkK5FC71t8n
flFbperSshOG0X01IeXN1l+CGeFiOe3P7kGazPru6l9kBrSzS4IJjbDGVdTBox0I
CaZ78/4jXWHst9SemFig+7Yj4hmXqU/TfR/usotV7s/+ZioIyMZxdkLPOy77H7U2
vaje3LQlmXHss8Us4TzPXigwl7Z79jbj/y/GSsnKOjYJ8fs/L1AxALkyZwiU/CrD
yauKhYxl1/H7CHeiX361JDhPJgco8RttueSsyyXzqVcGwqrK2yhx1Q8U6xqeofZ5
b3icPafgIdeZ+MvpweC7NnumSWnr9OXfQ95z7Zth2mdBcft1Iny+nvjtAbDIkJuh
5miXaepCYu627kqN7Fd9U2UXUHXn8d9Y0RqINaTGE1SvLmcMLLQoVJvBX6yuKC+G
LcQfh1+0P7HkUStwiUfYdnIkhI2+wIVqariemMfH/tFOYT0A1bsOXz0iUXhxOyDT
Ia6ghb/jRKYKzMWRJGk/GUmYwV6t1nK4oyXoAf/MXWNE6wb4xjuuzNa2s5Zx8CDO
qbL+NfOMiEj7heqcIX0c6ou15UbT51IM5o4Mw4gtG07HQKiZNHrsLyOWETIxhWFN
3iQqYgyIL0D/b4t49olYTm+lbQ4vcI4IQ7W8+OmNmruF1X4TKn4Bwt3B27S5a/pj
8fGPrhI0LFYhTWGpHU2Y76NX2IskXmx+BcOFwi7sMfHodqcsubUJgX8DhEe2XQze
1CBmCxDtdu2QiaDuCdq3zWqMFBSAyXsicgL07UnKMmowFzFOrjoDxqvqwAfvsReh
5tFWnK/tvHuecMANnZVcNurm98T6Eh49bEHYqO6G0abnYp7P1SqBlXPMJWnED1+k
IW8URqvgRpytwFpMc0MpjypxprLRZJq5on2wMtkL1l8DsVWzwCZ+cLjZYvIurcQs
RcLpgzGvylKY9LY5iec/PhcMfgcELtfwge1V6ZFQbi6L04fGOR2klkHS2WugyrC/
uLEwII2OPZhdVssbdHEbJtyrR0kTNcIIJVRTAbyeyW2WnglJy1QMJJeGdDKcQxaO
+WdfiwNqSmh60KKrAgoq87Boq8n9S7HYc5FiCYSVJd6alIDqDGiIdOY/2tgvQlkN
hhTmtLham4kL2svKdQ76UHn2PBTtdKNCc29XzszkZInRuf2yf7c72ehFU4R54a4z
QRfDK6VvRbca3c853zLfn5LlX3oP17abwNHt99p9gu3hHde7Ivw8XT7Sg6TJuAgO
27KD8XbfQpmv9VX5iMYj6+rc7ndODjtTyk/W+gPANBTytIkAxtz/1Xz8tuGXogg5
+pvLfjRUooOdqaWAf981aFH911dRceZmmMcdcZSO2SN9SyGw/ldn3pM5QjJVDCQ7
0w8DQjrTw7zR300ZdjtLc474p9PIqaW3XejF/5ac+wWjyZ8RmTaEFvl/b5jyUebJ
ZiZII9+nb1MCCU6V/eshnIOKFa1aLpcJoN+rz9V9SlMjgZ96vfnnFUopaGkPWZkK
YIltGhbf+13luVPJh88D2ONVXqnl1jmMOJWtcM6OWkJJOI32ch6nzKG3+fwPHW2i
oT3Y+PjyByvUWZGh3LSu1UERAzdK859Rpv6IsftVTOybhCKPEP/x5R9PXEzUvejC
rM2FA+ET1JIsWG04jorf7julJRE6gLmyy3rxsugMAGPgSp0x1XK0QJLn669aHAlR
TZNDiOjcixVLC1/IigfrRx+IdqbHtcmZl6lcZTm9Eeg8DMkj6SAg7JIo/64PZgkd
9AYzA83OLUiuSKcU/RWjfWIH+BCmRyHPCn4vxkvCugzH8FRkNdWx+Pf7Ort1wO00
LqxqRQ47YKnAIa3KkGns3l9xJxNBxydORT9vbLSVwcOanbgH65VGA8QNjnG68FnX
ARQIiGy363OzTGRG30HZVlnI2YCW3mv87YAgX+WdNVcC8aThaap82CRglxL4bQ8s
4T22dOv4a0fNRIjXbS/PBAEesP49DBUZRe/LHf+YOdaEmBpUXLedyJHz9KyTGf1o
y60ZXhpuHNeD/T3GSCJdvCa15pjaKfBcJi+mfO0k9b41ieKjEqIBdeSxWvbJZa9s
V+f6Y94P/pyVdyOFHw4pkiY8diiUzCdKrAdBa1pX0ht487ABogHOWOGZu1CQ8+r1
HvbzNEFqMPKHZ5ydYyyLtKca8m+0JOIUHUjkWZ7rP0HYW5EAo82liSTBM10O0MIF
UHNWHQ535t2vL2TLoNqKPTegT+I6hX81B8VAMXUobPieL+p/H1GLnefjMI7ZcxVu
WuFR3xiBpUOX566kfxNmUCocfFM1iF2WbNoQ4lUEGhHOafqUm9ZeNn0wXluGqM6e
5DNZ/Z16qwRTIuUnnsB7A4odrw/vE93z9t1iaAJYav27YoLkuC8RZGQ2b0SxasV4
P/oMBEVz87jcckvDhByzjxl8RUH7+D2+3SYHIMk768BE4kgJFgkzz4TKTDuYJbPb
EKGnsOXs2/iXdwMWwi280vZYZ0BaflubMXxlL8/IRh9U86SAnkH3dpA/B+E6Jl3j
5abEp+NgImMOU+UeNb60B9ULUWrmIb/jyxc82nF9HA1J3rvlnW7VzO+YQEgjGHLV
KWNjOYlGh5W6gktYOK+AFxsXM+BOAWJK5LtbI7eunpTMc9P8omDjs9a6gtmhDbtg
xaVqfrRNBtgAf/T2ocqSYKbPFsJh28i70DuwNQ8WSyfj2uydTQHIpRVrPPs2tmDz
mH+1Shsze+WKFkRvjivJoma4pWuhV1K77goHKgAllIwITx38b83dU98RhfBb0ovB
HJwa4IhWigOiDQu3MLdARSh0JN3G0lkA8wDRebyzPqCslKtw56TRb+gHEnnDR/It
AfUEOcr/98IjAhjda0b6AG4uRtdpyMNZmdA9uayOH5HgrldCA+IP3Xef61m9UzHD
x4p0DBjtUoMvODyNCLej67r+/00z4DSa6OxJ3lJi1/TCf8K35VJDCPbE51Y6hEn/
AlG/+Z/rfZRj+z7cf+5TIhj/uKGaK6AcucZmsvUgJ/54kUMHH4N5aj+kFDq4wGTI
YyklfiOYWMhvkRDAbtAFIGQQqpFvuTkNa6Iy0Xy9NQQ1YLdQI8OUQZ+WrMnPLHa3
H0k3jbWK0dndip7kaNqu448HOMQ6faELOTIYZ0v1hPX1e2PSGbkPkfwft2zDdrcb
mqk4Npw8QC4/kT5huoFbEcFqhK5/cuUZhqvIpSi+31LvwoSPaVXodEH2Ge969R8a
N96rXhvTCrujHYQ4a8coGEdtHWL/mtOlI5iKmCINtZLvAtxGxXqujjlYsxr8A3m1
OXPAhCSS/vhWLDWqxoIANIWWfa7llMK36TgfI5boLEnPCHiI51dJWu6L2flBhRjv
3eFZZS71ciJaGidrxSzEbmBvuelm5gRyRZfLHZCw9PHCneTZqRdFgdDQb2NGa+SD
tG5N5zxDSgyWqY4Wdt665tceIs7RkBbdbBfWiOm+hXU6tB3Nr2aBZKHaAYXDVsS0
MM3o8SBR50pW5fV0f+H+py6cpw+ImIA4aI0k+7uuArEtfxgUs/DC6dTuHImuBRb8
yKDhdynx7guGihmTQaUP3f2lgoMppguOUSFvdtyTkxFyuangqoUmSnZWauwrCUHu
nN5/BSwnJjrOJfXDuM264quM0LhS5Jio11XWtzmmrCr9ZZ5ZCypQszV5IDlTQ5mX
L5OjToy8h8W3KMXOXen7D3cDOMbvMLKhSbJBcNffR8/PPIgd9IfPccwlXVVAm4wW
qF0YyE9Ggdefe7TXF9rgig==
--pragma protect end_data_block
--pragma protect digest_block
7kSVv3Hbqi3I0x7C3JeKTaIte/w=
--pragma protect end_digest_block
--pragma protect end_protected
