-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
CI1M3JzO1kdJkS7sugCpLb25XDCTG4HznzOj9ZJkY3W2zTPQHGPIvVfuStS6F8Pt
+pCHMvgDIEo7t+3+NjPt4nsjJLVVwcJmhpKXIlmmyU/fszyiJomlmSLNDxcUkBQg
dUeaMNQJz7p4Ue47qPJiB7hOmzUb0Sn782xLuIck2Ac=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 41984)
`protect data_block
YEiggcGB0IslcIcLoXYflC37sRuhK+i/V4gKdVpIQ8OkID5mtAPRWaeOIU1VihU1
NYfb0f1S/xeUCyY7ZLopZYolHRB2xXKP0T7RdK2heB3O9c/nyXCP1w/02Vzr8jY4
v0HELlqBayssMUzjx5kck88BzLlogNGDFn2SPAHykggsWxfE4mwLWMsHJ78R/W6y
h9Jp4N6PIg2UEyPjjSRjtparEsc1cf0ep/QsKZKLm7n549d/6Jjlmk8dUJfDGuYv
AcOBGmQ3/G7VaLdZlaERi8vsXF9Hz4ycA4sSqK5ervme9JAizbBgpfDxPebZjgs8
xe87ssykd25BCOQ/8xRYZnal5PnGBccZvPyWRQt4NWwJO+fqP/F15EOQsr1HRbZE
0czIY0w7z0IKLKU2+eUqw/nlLKoUSsfefYgjKZ+qCVCjN0caFhCcLVLsehbqSegE
IamrOoUiFZr4PaVEY8zWcAzkuqo/tSWUeLEmWYPPZ9lx1V+0kf/A8e9dr8ve0J0i
0WT7RoAB2hu7K0bX9TgeWK63kFYxAr0hhIWNVYuXT9VRsxKlo6RVo2a5QPCZrYVt
N2PYrtHiDtxVXfx1yIqo97bAIwjtQ3sjUWPzSBpJ4sLbOO8QNfUgase9874wPrSl
0MepmU5vEqtlVlzE5kLkEdjA1lINSAHTFiUCaipUSISHBfyGtCAb14ydipy9HxPb
ZyOh9sp48aiO6gdnV62g6yWbaHsgE8xDGQeJl2JdeyTVtFp6n5BDNgI1a+aG+VnJ
2T//oxmxwSqCh1hHZr/FuaCgFHQESZs/hW8msSPpZNV6tcy6BOjgztZ+Erplxqr4
SNzqZ2ENw/W4UcBkaAINTPb6gm3CW1dv976HShd3/1ze1QjDsjx7nx5MTdbWiwfj
QF6euOWPJFEOrbDBaux9jeFoCN8uWdz68epsCmyt4Mgn/tJKQ1fYLte320FFqzIl
Irk9nUz+zhrXRFiBGyaOvkJc/gpr9dKe7OgEA/QphWUt0To2aHlbFWy1/rLM1O22
FatGAVle64QdOrLgi0vd8rL170yxzRMMDgzFwbU6iFvcWLPSlGqJ+fNcyiWBbtNJ
bbpicyNKYEkPUBuKhJEJ+Qcfy8vYnQEyBaGGvCW49h4Y6+eZ5Kl4W5vMnw8eKX1Y
sGbw6W1yDYY+qOi2WBGfkKQ1k68jQHVHbtdFyWOdWPRrBOxrkBsVW1977sFHS/2I
8atqhbhuGZBTRm6BZSyigR9kSGX04dQVsJI0sjxzfCAYKCcys9GQ4Uol2s2B96Oh
pVtIv47gtMRhj3meh4/53V4JV+MR9Cbp6vv14dDUq5C/g11W/J8Nsk6EKf0Zg+3Z
3x2+dXRf2VxylxP79f2YVu33+6pI2UWpJYGlwdeURaUQyN9ZVyMgNiP1GvgzRoZ2
Z4PX2NUxee3kFtiDNcu4FZEj1FYOiyyVNTrN3KfixCEHDNoSwqABLlcp1Z1yQ8ph
b47uSG1dNSmE1YGahC/RKwDxQakqmNnZoKENadXt+SisZKL1zb/+Vme9k+B8S5/R
wFwnym9gMeK09fiDneBMnTJ2JD9xdAsZeZzL/FdknicU7tAtG0ttx4KEehQ79g/s
0Cq/gMPth/xUoVxC08oPCHO32SY3yhL1ZF5cZqhKbrYndPj2F4TrmgkEHXdIhjC9
2HtqCI3lNxRwaZCWzGmGYpWYGdDj2v2wO6jtE7QTOjj6V9UsH36r1CxJcLYhxloG
vgQqxvvcdAbjieEYyLYM2VVW2fVc5yeiOEzILYcxFJv5mD3uS6Avv0jKSdFruIYp
7BH/+7BqijIbrtG+SYylOPWcIvJP16lwrWyr7xBmohuFzXQdvoOSuTbWI0nmT3Sd
pne7yOpaSVxHrx7b7HgqHgTx9avIjHjDN3MWFpOg+YPBS5yfuYk47Piltgvej9ze
65S2w5KjOlCGBwueKaa28aueejgjzPn4e8tjLoCJfr+QoRNa1TJtDRnw/NjmDGJz
spK1tN2o+Tzx1VF7rUcCH2BG7K7pOH0sbl3ledU1kvs6OAH+LG5zSwIT5FDN6J4X
vpcFrogtwoz3Pkj5JhE4r+adRIQfnI43io9Tr2NCWNxN1HfpesSVsned+zeBTLwZ
8qA2EK6fVhX1udXDFf7YOqNBl5rkwnbe+dnujSMuQKS3EmgTprphb5SUYpxzXS1n
qRI97COQGKIfVjQxMr/gpWFXodjZ5pf8HtPgVLJQGgDjVp0ESBpsP/2rQllnWs8M
rjOrg5ybsSqBtFyTYUgoF7oHHPHsl7CXx9dL/sPjpbIMluByXHMgBcDzllDxASPT
Oh1Y457m/iWAEH7penkTs3Rh4UejKajpCfbFSO0dThONkWiYxTxkIS4UW6iRIZVk
Yb93aladEF+Q8Gk9RMkXCue6A1gJIPNjj3ozUoeqbx8EWaIbTom3fegbXx5EVOYb
g8Gg7oSnuN3XvtCI75CnLJ4CWoOfbVB3YRLOHXwblnfnUu0o27nQHJOxh01uGLlB
/QLUx143zJFrEP+xi/ZdRc8DarFcPGg8deKc44WjG0LhZ2ZdcfQIInbkjAOBJvm9
qICiIyexUeosB6T34yy1q8NHCvujaizIuWHWvqkkSqqxbeTq0ep3qpvzRKvBYVh/
IO0oQ3YvddTE4XKx2HJWmo3HClCZ3qyCRoo4RiGLgkDWZwxdgsxdgpxq0FG/3+4S
kYR0XoD7iVps6Y6up3I0wG3Vg0zVIEr6Ez9ONE+LMIZXcCT9Tvb/CetUpKqlZSvt
2sgJIELXB/Rh6lCS508hCejPqB8Z7el4J4HqOVtIl+y/4WSXeL/6FZW7+eB51GXN
JxTta3BSEC7zfbYlPCyNhkTF6EVUuneAJRQoBt52Ml+qNlvmD+gmXEfiqrj/fTjq
+tUZDiXi2nRMr7ojmF+WQAPtFxWOTabNtRfTzOTL1idO3yAiWf22RDRO0bGdS4WA
/l/rvsqNOZHYCRwn+ZBNK5z6bhuyCTUCq1hFklVGAAL0WtHroIL2uU9Wcgf6i2qt
eYzVZWcHyuvczmwu8PNrRPAWcHOheGs4/w5Uc4XIila/MShZgEnYLVDs5r9cj7TO
7aefZfdFvbivQ5Z9dMSxUSagWKi7moDaqVFh2kbMyiNLZP/vMLsiWaCqX//hTIbB
hrqytF4ObAdxz7QFY3DViu/PoSI+TaLlmVbyERhTnBkjYxq+qRskm6RZSVNuV/mx
aV4W0GH/UGCHgMPSP7vzNmDBJJLOqGggsIDMyWqtAxroUQxQlmJW7KqlmOWcD4LI
IA7IX5AgQpYfHZS40LMKzyWz/ARz4hBRrbXTez8jpe5rffV2tLNFGGIYCs/krdKm
XbD4S+QAdAslF5DFgV6YUcxf6YPVTpzdgLdqj7JuxUiHOmcshwPNr+cGA0M4nLxY
vULZeFGPvNkhjByA9aA+HymipyW0/aTAZvAAMjvdqHn/y1pV0493bPcUTG6ZwPrD
1wmTbkJpwDEPyeze+a4MpfzteaGKerIGJxADokhsckukPS5eC6YuZC4O8nrVSjf9
HOL1JwufzLb4hcclOHq4UQa4/bV5Xxw3DY0T3p0fdKSaqF/yfbVpmiNVq3e5LOc4
Y9FgmKbE52Brc2IDRBXiCYPPwiHnxKDObqa9hKetomJF5ZVTV3sgQVxU6ZcCdD04
oyJCWILFp0bJlU3Q9gl/ccO4EH43KwZ/CyTTP+P3ui02XjbVFM0KAcrRwnWHpDho
FDeyeqCcij0zVJ2Ssw2rtu0/SHi3uJhG+Ex4qLDfa6lHGqSBRuviTmggEUwv62Dv
e9v5gsIzzlr6UH8Wg8oOccqykNydiOgmKe40UNJIkfStaAFx733VJxwi5LPTRINn
dr4ze/v6duYiiCam83TLY0mIFFgEG0kXO7aObH5STDTr9nGXiCJAi22PGm96Ypa5
+OoWXh32vigN3fmqlEL2Ksnr2D7yV5Qizi8BFyaJjLb+l5xuxL3VX4PCW2+lwdtc
/6DUBdWaMDJ+Xq4rUEDxlz/hlAc0e0G3yKH1YptlIGEMMTQKJOK2iToat/kcXHnh
DpxDRPU21U+xlB+JbOmiV8FXn7jH/yyFwaObTDCnL/SH1n8ChHVIIJAm2ex1TtMK
EAfdxUtFvJjwpGISZu2Wq3qNS2fpFmp64AL72DlhzUjq/FHoy1oyaUemBBXaBlvo
huJ0B2lNEiO7hksVucP1q6aTwEjG0i2SIKZb+kPEgoYixLlMJaV498lFjKLSWfCc
8SrN904oi3Cc+sDnroxt7zw/0UPjonroYIrz/4kGS09XIcxxvfLNAoOdQFIhNZAJ
dFUQGcVKH7SzUdPFT6LdJFyD0CPk6IIMuDUOWnh6vyPk3wCIzxpFH/ROvbklrNLG
JpO3M8bfCd0gez/sekvVzFe0sMbzWNBur647S8Ku8i953lRLw0ziOPfUP1CpIYSm
UXOcWM7hIgF7vq0P8EaCHtR/dTsXVzku0qTFj4x7Ff6mH05cM3axv7/zJqX40bWo
8NZXUZATYX9SdwMwIqabrSu7TK9eFx0OyEgbBsAmjwXKogV6Obius80ZV9uEiiIZ
vFd2x4hxHXVFrYU7CNVL2vQQRQj/Ny1UDqFU0exVaO4auoHo6OW92annwErfdPoI
Y7UXr24vb7lt58JSx4BHKK1eLxSEx9ooYKoiSNbVzx7C6c+yW2Inap+GocJSYlkJ
qzgCjChCi0KM+4pTMFCDEF0BfGXxqL/YazIUNClrMgMICp8YEprHNY4y2UOeWdpZ
WKsaEFqLWdD9jKfs1aRIOMroulifj/mpAc8+uoBneiDHCaBk8P6J9IPSp7nZPU2M
QWqusAb6INlaxRY2o2SqDRdmG3B1NXFcdLv8Z96v1iezDEft5jsbPcACugP2Vepr
yN4xoqt+UM/F7hz4sdJ3Ym5/Fe0bGTxm6fXTsiQWqTrzblg9udq9NLg3IW/Icyx8
DIFYFMRnI5btVjoBcolK+elD05vwkLxyZxPChJt653NYIGSmLgvjGaVHyjAu1PtZ
hdUvnZXXAIQmP5BrcB0n9NoSyLZbe4SGM1XcTH2ftYMJ86lJ8AkiUMi9qWNu4dJB
I8nEwYPzc5jzU40O/SlDwX1VjqXn3ETvrJ9jo0emf3XTFz6LbS7iw4EhixS99qCS
WzMMcTBAxKU+okgpkUxfOohrDnm5byse6LGYm5B8nwJRP1JXZU7W1HlOJIT9jP97
ICCPj6Xxw9F41qCcxbgP6ZLKbfRo6fihMlK5DvojZntNxNqGacktpj/FQZw6EdDu
5b8yz6YazKGZFmWDeHHmPNsUTzCfef5o1E2buQ7/VNtGIOrveC8XQsI2/w6waV/P
nD0Lv7c7CvDWNk5WAwEqub6VCqJDgoMVi8SkCK61e60XPRnWq89vtYTySTXu/izg
SkZ8BppkgXXAVDTnpID8VY/59uMghTX3EUishwTEBAteqHvVxIQYs7C4DXFQmSY9
RkG+d5abkY2QbjhA1nHAI/R7t9iciWZJx6e652euveFvAScpommqYsB2/XeFmVie
ZU/VzeJtQF/PM+TTi6iC3RaNFSk3ypRGHSujPpBWsJ1Lq1zxZwpFfVwNbxAZqGGh
MLNOrEwERQOvD83GcDNVLdoe8ggi4i4kaH1750s/x+fGqihZbfrQ/V3u6PgMC4eq
nbE/oVSN87HInEZB3zSiLpZz3jtR+PHUN3X3ckyHKifiYoXEuRzf1T4Zdi8ur+m6
7lSw/Uk0aQUeQFrVRwPj/HJYgqPYjqX1LtsJv6dURCh4Cw0HaxDsNRbTxiexzuZk
+wMUgmy93WvMgnTYWOf/dtDy9RRRj3NdqHv8I3KzVvEtoQX/Jl7AKK97M5kwky/t
GvPPuudvNhNLwbLUaD76DZlAbLR08EALJWhc1DmVSmKBxdRGF8mssLG6BruznxcP
Io3eG7ZU4uWAmQLYhCnGzLJ7bD34k4KEBcudYlvGS5ObwxBoLn2IaQdrAz3uWxZA
Kyxkl1PiyaTX4C8eRcGm+TS+FCA0eqSH8lqCWiRfn2zV7tKncBY2QWoqD8n6HQ6/
U61AhA1y3HB8xozhU1tIhscm2FzlMDssoSV3j6+/S0kOTWWTGBOZ2dow4jx4CChP
4Csj4i2dajmCP5M2UgAv2j8KttQWP3LOJqHkiAUUgzD2cgJ+DrpOiei35sJp086r
ZvnusawAOsz/53pssS9jSvrPk1ps3M5HASTOmuMv+bi20JJMWtSTQwUnNmRISDFH
0haeOIEFFPJoWKkhoAnFHOYL3afb/8xcmnX9omDBv6EqGLaAgJ7/cCsJhHs8DVCe
+rO/VCz2PkAdtbijpe0C2pUf2v8gAGeTa61UgGSItWmkQHqlabr0XR3Fwa/DUiHH
kPGZGUwXRo2CPXP9ZqIzwxjnWVd5IWeQ6peFc2jEvuoqvIrA3Qtt1Dlj8mlloOko
9EvX/XBm2EqnzWo9Hy3xh9mPvAcJzPYgM/JZaJIAZuOtMD6EiRIrz3QIq3x/J1tc
EmiVhCWqp4xVUdrnygHtlAc8GBsb9USrl6pAdK8oDTI//qhLG7tTtzq1XvUFNLK2
2W+KAf5niBwTlp7C17YR1gSLWhaeNuR36+urtGHpLVrKrh51jq4fEJqr07BffjiF
2reTAXUy6GATxKWGdVuJKKq3A2ZMjct+2AZkO4a+A8ncffeH/70TiGRL/Vx3nuTu
bUUXKkRgMlAPg++SFBeknkEbcFcCcZy6CrwEB7jCJ6FRpa0xZGFS4zurz6pq5Te8
odMbLKTp1EuPhSNmniXjXRTGWRu+d7vB3Y63qCUFDA0hacxcs4NgDkn1eUC0kJjG
xJryz/PPCUuZ9AcoHvf6T1FHnwywUX+t6L953BGsFYpn4jfpaBWzZAhUkZjh9a+W
X6Y82TWsKQOkOAYoiZloF0djpeCho583ABqvuRTVgqn/cHrYHmjjh2wQOoU5gH2d
nMZBo6hrSCUiGX2d8rJ/lF0spsGq3XO7+a5mWoM1zyGZtSWD7pfnL0j9BgrPpaU8
VqM5dci2e/4b+FuO/mzUWAydjT4XV3MjbpwQtgjT5zHh2wvfVTjOZD7yPjjz1ECY
wCBK2HDWytWFk3+3j86M1K+b8cRjxb4wlSgX/pEoXTQ6G+DcrmwDZk5AfY/a8M1n
6L0X59AwuHP0AxPJ/DeUcIvC2FNucYULDMV+p6yP3ho4PRIz7rcMdIBYmVX4dBCq
3MMor4K1fnhcOGM2KQkrYChjy+kycUurNo+iXJ9t5cRv0q4qbwrDKVxE11v7mY0j
acQreRaZdqb7KPfef7tjylg+VebbfsTZ8fA9+K87YSqCUQI9X24JvFXEO9ALqzYH
vGelf9RbT9iZE+YpKq8mzbLIBbVIXnanI8MMrp19TY2oC8Y0fuj1r15bmDkakkx3
mCksP5FDpCV+4dho4A7nYGL2khbIgCYhRBW5TYgvDoQwYp89+fxbBcyFzgPBrVOH
bu9xngnBwo+d3p/SmAEvj5V9gjcYg6ZM+iRa2rqDmJBYw3wzgWJCkl3FUnj1u8eS
wM/ByHMffQkmpcIjofOiD6UL73lJWvHsnMOl7Uuzr6p4p+AOC/+PR1yeggsXzeAq
Apdx5wrl5AHqrjsj0uJrPrBThMUv2q3YSQXjyk2zjXkF03x4k06nMey2HFOhz7i2
9rtwsKPbKCbdgm0PMKKMuHPdkMbnM3JR5cEfaReaepQ4LcxFJJidXk/GPft0wOuK
Ox5Vn3hwQHIV3WfOFPIEBoiDz41UxXub7V3u8sS+vUyJ/Gr8nixH8UiOeabqeu2g
ncJiANwZYHrv8i+aHAlcJKEEv/JoqJi9yLcynlYT4KILGKMaiJRsyD3LWyLzfERa
soP79DY18jJGmvyEUuPvJLo+VEV/RELZK/lbSqBjE1DUssf99zIsI/ef6yXBu3A3
mefVdGPq5s828OKRZnSBBWWrZ6DjWzxaNnE3S4oEGr0cAS0jw8Sbdpep0MrWx7iW
x4hY7pCF8rjCRsWr2dihaGDyyZK78B/NWsOi1JoBxByfTiZsGl9qd49clBlrCDmB
yGCZl3WxI3fqhojKWNOrX7SzgMzpt/W7srgbp8yX/SKcgC1j0tY8V8w87dG4U/Yy
ybKGajHMbi9Hgl6jkOlmbmwqtkt6ex8vG5WJFwIa8YI1N93gXadTl0gyPzmsMX5J
xDO5pLucP/+EWFZ55MZfOjybpCJnTZF5AycUOkYoSCmTLnIRHk6boe5xT2vpzz05
ARjn0te/xMCzPbhqzvTlG/pz5cuulKx7YbKusqObd2I4BU5N88l/bQMrcSZSOENE
5fvQTM5mu7lOiW+ABamTxtNtcsk6VnKHIHCKcX713yJf+Nq3Zj/7V+0O1DXDg0ui
xgeej7J4KCItnPwd451QgNN4VD1ia5yFJ41Sxb64J26lkDk/UybUtRbDzPCVbR24
G6iZbBTuU53uCHvTyl9N/lYulsraMNkIjzo2AA2EbiHzcEsu4Nts7d7kCpPNuJza
DyVjb5DDk5no6q2AvXYtGum4tBnwLczhhoy+M2RppkOUBMavgiNSZjrOw3FVt+I/
vNtSwcuEgrM636TDQ6PmC6ns+reE89RPvl0GzNPr29D9bq0E6kb9g4q1VZTc3Dd+
VAN5cvX/DD+ciSbbZUeSoIwPIv8e7DJFvD5Os/aTdhlbkTC2FoRU0lIiDAgy140T
3SuEXrpR80PjY6/FDuTWIsImNZLmvtE2F9tfwp2/Dmh6jEwVgNcfu6sBLPUq6Wfk
iCG22oTgkWDuOAVMsjUtjoDJvlrZNb5R1vE0OLFEjEwzPGNB+eNQhG4orzgdlat2
HsHhlx2Pt42PyLG2Xn/DDy+vpg5tE74DJyLhNIWI+Ls7C09fv/V42QTRDjQO6H9s
uBN0vw0PiAud2ZmXvSqC+l7qkD9E/IjWLAEwNFTYZoY4/yGmb47EjprCmlaAx3kW
cQlpFJ/xElFiu+z8PpmlelXtQBqaBtrqO1fsyp1ODESit2VUToWmqIMu3IqTcUZB
2LHZ8ElJbEqkwnBcdb9/+S716GfgZBZYAPMVRFJOWTCNJFl1MVrLiU/A9U/QIUPL
yCrf15N8Fa9svcYyKYOGMHUOUY4XL1P8LqnSq+b7M9i2ACHtgODp//czyuLRjDvz
S390eYul58CrKqIHFOpDhixjOt50pgHmSCU05h7DlM0k8OVSxTcLM6y+nEDJeFa4
J5V3Zvu6b1uUEbJwFpzIFUCdOW7P6ztmU3I11syKmZbBivnEnhvEcVeJq092LXrp
2SBgvgD7ub9ebPdKGIjS6anQvhLgjc36y+QytAnuD9xMz7s2tCNShY3zn9EQPlS4
CDNh6dSYm2jk8Ts31sZeldoxIWaI79l4CEPW96iuk9P5TT/5B2vT84KbfY2vrSIT
J2SPlXK+LNak+5qsG8MIXyw0Lh+8lCgxf7ag/XnZBMT0aP75uYoYfmwLd6Q+rmHr
FSmrT+VNd8aKZ+7bO4ngKVmP+q/+8k3nJsLQKu/i7ldmnB58oRSPeGVSLHgAjyA8
V1ntTOgAacfaDhICsVwdtYVAAoNXcSOweZoqH1MGp6aQyBGtbzg6pzitvvJOpj4m
wq6b64Q6NXO6h+HFVMAvXY8gv5ev5LmuraznFcGg75y7B1vr0JiEwID70Ppim6Ka
qf2nllsXH5HqfYuXLFhCjXvKoac+gERw/PFJkCKKD+uKPwuvPtPpCRln5mImqC83
Ltf+KHuH32UNDE4NQIOrGjIjQpvQaZ5tCcSqOWC7Z0K9fw6QWjuE2PDUGajOVH73
MMZJEcl7xP0odZ2soEggsLGhJSSaIjdukG2Ch3uodj7JlRcS0+DHGoG0Fw9SIqpq
ZWhcr88lKtq6ptcwLM6+lWKPWbRBeHDI6lRTdiQYtbvA4H8m0fZMgo3pDIFszHJ6
AwEsaOXQ7dahI78Y4hsz2l2hAvvSu17VxkwgaU/jhJcayvbLGwt9As2I8K1iZOVU
dcCNUZgV5PiFOjBNX53dWuRkex+/vljPqgbPrI6prvaOws08cAZgoboFJqPTbByV
aAYGUVHJuZlmzSoeO2B+wSfP2324Xi++rZ2dBW5t21jTsvXh38UhvkHanTA1vvsz
jSmJ6995YqxegQ4HTdy335ZGMbQeCV89trbd5cFD3Lp9rhh2Y1uj4SEg1tNniY7/
5fivvdW9TMVSxVCKvdjmgBC9uGP1jcpWWqJ2AB1D5LjCbZCfeH+TSzWvSFPjM27+
omGogV4WzaI3jf04GCH08ChXqGuvXyo6NVKm7PkX0kZvGWNoPI0s262YHMSLpmEf
DeY1wQxuZ9/sit05GVmJ+Q6lYaoq7Kupwhwh1eSRGXXoiWSW6lP+gSJTAz7+LbLg
1v516afpnBsEXQW+e9fWeWBYHg3h08um4lS0WE4T0hC73Kh73cN5XLFaTt0RZxdW
4EEaeSl87K1GrJfeypOYyLHNcm7DJRJgG7eSKN86WubmlA5quJ/MsyhaWWVljIjm
+uS7slqtbxc0/PIp/HXe6WiQDm2fqr7JnS+1D8cxpVVFwGXb0ao5dTSExaD6bhT0
mLvzUDpPdwH7teMsra7N6cdaWcjQu+OhscgkvqpoYRDXMP99M2gKHSP9Vqsi4vHh
N6Z/Co6l7KHK6AWw/Q+HGI4nrAAeXfritk5ShEr0m4d6BnPl4VeR0AkfhDUf6k1w
huEPxOyRks0anooad2kx2cPmQGsYKCyaoCjwuBeE4MeUwsVDRYcYhm6FJOBAvXO8
VGr+Mi0Ev1tNmPBYL5DcdaIVDf/3ccPWylSiHSKyegm5EygHxVrMVv8964JALYb7
BsPL20lokMSt63I9BFxsvuJew77Cq6lxhYApnmMoUwagUZn2olguDchrNccuzEKX
9Fx8H4ngWCAJ3gHL88c2XassMkPzd5k4cSEwFGEftIEGUvzQKfcB2cdPOw48BP4o
nMOQu46oxxG+Di9uPMSxgKTa9H74v2dJbojWnW/IRRajnAsH8Z3DuYIXup9a41mR
ewW47r2sC6ctw9FtQ3xkdYDdK68gEQ/MQPoZEUTDaN+EvYzXzSd8rv8s8ENXaS86
wRjCb3BGSQmNp7TuM6xCYxHSJ9nJdHACD34A6NtrGlzDjoiFuFqeqm1MrCMzh142
rEirHYWUhR8k6aun8xc4z5UO+UBuiRTEcgIMlviqLBYt5R/A0i2Bl3KCBgulvjpB
8knGCftW+uhLg4MyVEbF7c2Vrkzr0LyG1IFDawaTKNua37pqjFZbhg41GOxRBxx+
Q34B28QrziRNcMLOGGKp5EqqUYBZGnoayayQaLUHZ5+YwrLpmQuMT5tYoEURhx2K
O9xmgOkWNaXIhCKnLljalQZ41TiS0tVpu7I86Crh/NT8KKEdqLYGQCh8iYOtfsSu
ABJdk61hKOj1Gi131BAVBmu8nyPL55Y0dAjukTGMopPlccWSPHmYAz3P0n9H9qDc
Yc7JPvbC9+KGXw4m4QIK5BGegfxRVA09edJLoOyPfgZA7Q/VsjCywSh/G5FSNYbE
ITy+KFYJcLzysy9EOkq5M6/ytxlbtWYWSSZbnZuCu+mHCQvT+3KMDkZLzHbLND+v
LcKGDVOEHpnDS86KBJ7q5HfsBSdU5ZF7rKbdKP84bmeFmY5ciIQn8A1wAXVXoOY/
ZFHlN5Ra2mlmLkhSOROMvDFdvY4KK7wsSNQp8V2IMiYOLDh34545frEV9nwxhr8I
qUB1aKg3Mgju3pVjelYZGzneRdCwwOfuhIJD6KVU3vcFyFVyI2PQ2pvrLADjAOnK
5pBTpZBFfAby08C1373I/jylpba//42r61oaoVkBdodJO1rpqZEOShMCP7f4tTPy
UrIr+IlK2z77tECBe+FlhxBXgg2PIz9jYAZiy1AEkyhVBZrP/0qb/9ftDOlhJ5+j
pjf1kjw3EqgMKWHCbNpB8NAGL+gJGowmbZm1cHFJrenrs0vlh67Wh5y6mz+2CsaH
6wuf3gMhBx4z5vxe7vYXfK3ZFr2Nvf4vw33Atc0u96ylG05PnzFpC53WK/9CDcWz
rCdUBrbbJv2yNPOtJAqHRQWnvLVYJZDA6CBCdFNt2yo0vzY2iKP9XmXeyI5pHQSp
hLoqpNSRUuCgG8cgy8smpmLg5+E9yVFL1oixqQ1S1/Dq3VL+5aAShKvskNWfTurk
+FcY1b4TPGB3AvUFPEu976VGn00NY0RoHe6PTxC5GBzXa/+OMk0u4UyvFSkqE+Hs
JHQaTqJfBGhvTIF3uBTzIjXyMkPjsq4NpBFl5hFwXbRWhQ26hbiXblw42zW4qRr3
BV8cRtPGJoOh7C+42Ut33amirf5mF7+FDO7FnTiueiOMTD485Zu/f5+9wQj2pCt4
imWQ7vM43gE3drHQ+e5NswEYUc8D0LM34aqek12jMO4/ppDwusDMzW/JZwiY99IT
a5OaA7xFhVokbhOwDmbkDo6/vfpRwA+HoABtgsGA4+n7EIcGky9bjRI32Ip2DMJq
cd9B+oa87Vhk6Ea0SzUJzsEGQQnkAe9nARedP+waxxI4makzAU25oMya0/VzP14H
Pkl3FiTGY9G39hY4KnUcxu8Zj4ic3C89MIqKXEfExn12bfZs3yy1q3NOoAvr79qm
RSHETTOPZNVJj7km8tJ+c49TfV6z8cPBbSnCvLLf7I3UQ2eiCWdzMeaEiaJNnHWm
AAFuvYNX1AdBihGuzPJSH895z73wiMYkvAPMpoR7V7VDTlcfPyW2i1c8iSKmQtv3
qQafz2YJCuy4swFxUR0eaORBBIXeTNyQvgCeQJwOLIJgB3G7yxFXbljBUoJAUX1X
t7gPNEFWRiYYJ9DhGoUcQRu28Hx//4RdBvqw0/2GabQyZJp1fL72606zR4b5mHI8
B8oeOGwd5P2J8LNMUZxmowZx5sjuVfC+WhWEaXjF/D8yKqG4H/RaoQbIOjEJF/U1
x7LZBsk4ByVae644n+vYcRuEqR3fIAh9l0BrRDD3AsT11E/K9Ktm049/B6/pc+aX
z5llbOh82tzCWJ8YrbaTfERJZOWMfeK0eVkG1nEAIgo5vYCPpIZiq058Etg+tsXi
jRAJty08lN4U1t/+uBoxyoeROssqvmbzliNUogyWneUqd9JAddSmnNAGmfpo00CB
jifyKN+yBImgFBpDvFvoZ3XBAfI/8hoLLG0/P1CPXWdC63oohQTZ7o0RsAs0W/Yp
E5SVyBUaDr5HJcJzqm1xO32wJb8atcCytgyQzjhOnI5wWncrZ+pVGaWH2T0XySpi
OdkxjXP5KY+9zEo49hefytxNNg0fBQ/BLrTOGICGA+2WHlgMwrAHm4kXn5930fvY
1odlmo6iPrd8w9hd+FJZStdYagHjV8cwyJVg073Yp20Sa3Jb+QGqYbuZtvtrcWiU
0/5T3lQGT9W+GTG02ZqPJsnOGQ/SKQWCL4cRxOl0UdVLlqdE57c4B0MMEcjh3NFp
cp3LVl3iglyEaJ24hITEVv1XAJjqws6LwopIDziURNXke8h7dkl4t2Zci0ORNSjb
cnQGxNXRJm/jMBRjgc+n4PZIVS3tfMOedhIErAFqPwf0pVBVF9JgIsZnvUvPs+Uv
bf2KDHHMRnW9diUW+xNkl+D0wK3V0a4dV38kjUnasx/YYllJW4qgXEEk8hoslu1U
1NYGe/DJxAfmlD2bIcFfA+pn7Knio92ksTYsGgG2A0zjWa+CAiGfI08LHlZmEzBH
ao4cBpY2ATQ9Q6UTr8v1nFNgybE4w3ugT5gIhuflVV/4sdhn894zHt++jKc7AfJa
IWm5UeX+hQLo/RBVWWuGbZUv9EkWCDCIIDRzd4E9PgjBmJiD7h86fDg2gdcg3NYV
vN6rrZ0Sz346td5QkTKcMyHvRXsdBEHOV9dvW4GkyUYup+8mfATyQ5c4l1eIKh4R
TtQegFiUsD1uLmggua2XKNEcyCmHvBlFjXNDHNHvb5Tic9N1xe0lhYD92GwP2qWA
mU8uyLRuHXm/LC1v9vbzRRnUj7qQW5UFdJFwHdNK2xO9TkZKADu/rxEjWc9LSDZI
SDlrt9Xa2YfYbVf4L+1frLuNQTZUhVUegKh83RIJycLcd+MaqsZpAqwT/4i5+mq7
XVugMSdQskPScwHWNWhZxW4RiyLyW89FMyAqgu/XNuys05gLKoN4WNYe9FXDXTzb
boB5TQtydgejjikDPh7D16rcHfFancHJfx9G8Y14ZP2WlBOVdpO0Ddpd2HoigeBU
hjbIjkZ3+bXYAZQAubDC67H7uCkZ0+Kx3vO92oXy3Bw1sB2KIkm1tBTaCs6U2veD
yuGTNDvBTIFrTCCHFNGw9S4+ibqfu4poBlCN0ujHcsvXI1jlhjb/5K0a8hMMjTgj
Tsjmn06UgmtgTeSSockladFYPILkPK+0y3ZIuDVTRI1PgivWEXEm1JqQLtuQlmkC
QCXqy+kX/jpGCkhGeXQo0rD+dIwDXgSlWDbidbQPuNxHYCaQfHmpWxlSrppqxOzx
u5qzWYeS/gopCNeO0+k2z60EcWtfBxOHuizvdNKBqiiRsgHZBX2Z1zHufVWF+STM
jbBX3vVfDZdgVUI6YGkKxGJ0ubvnO6Avg26DByV+D10YJxuv+/sYMWlWwFavrH8P
LxohBFi5wiUR8DBHRTQKqizFHF4lqP6sNz4RrbpBvyyAUA0RHHF2ic67SdrPfRMs
S+awCfFJHiSYY+z1iJg02ZkMcg0HVTvYiCCMtQBWV100rq3MXjoCJuz7fEsi3W22
7vc+/o3qpuIFMAe2zH9tAqZthZUaxwbUtLNwJJ3TmOHcp92l2b6YRQIQNYIUAaOB
YUf/VNZNkf3Aw8LLhIpVt94gZXnq5YAbvY4UPo/wCOYDJPLsO+t31zOBA5J89g2T
vGw3u78XYdHXcD51C7/1RfAjhMWfjOE35z2ma7oaeQXCSPjgYDvZJ+xjJpxBhbP4
4u809fjhkcQaG/dI7Z/ZOZ697tupa+KHLP1TMNDEmxsub/KYTDsUte+l+31MpZ2v
OLWsXfT3pn/hSBTDzPRwJiix3Ng+8wjFUYdIPZ/Y+VPxgYhL5S20C28HcA0gzO85
/80TNrBFN8C6FAPtEpWiLBZyGm9JU+IABqngsoUcwQUfZnW/IsYKX44mkh+CjK+P
iUYg+3GNmEv8XBRv+1NftiHzpyTlYD75HogGecbAqNgmMmt4t8aatxYK3OHvn8B7
fuOH0L7/78wofRWtKLUi6ZEJxeVFPlF+Ygb9HrJWt8x4rCIvSa5uZocIqEC/wYIY
9mX9tpd+HWYwmjz3YjErgI7KrRRghPu5CSVNdybLKa2pTdSw1lk6c2pWaacxjNX3
kbK/Yi8olLwtqJFZQ/vC2eR5PnMrOrvcdDev2XQ85zDdHmKBbbBkqmerlYb11+Tb
XuLHUT5kEh23u9vFEla3zEGomSYwfiEqAg/4ACPafBIV6VzvTbyeXh3r8DARgfeN
vETCZsc1YNZSw7NUub+EbOfFN64cMnPy1By1Eez663KjH0DSVfapowbRAKX+XFM9
JtIXwRbB/o38Rsc4qxeNpzJZKgFgjdPLQU7Juoctas9jVPHNUEUT7UxuOmKJFppH
voR9wpO2S4bz4T39wyEpsCHYY7Qb1Q42q4kcDHNWE3bxED1RdbeYuHxG+tWn3Bo4
F/pR7GDtd610eSHD6ueRhcQGqGNoq4YEePpCUnhXO0C1yK1qfPuS1mcwIOz6F22P
soCK2oUCSLVRdnPbjB11CVqPsHwBbGj2byO/UcV4/HLpF/vUGwts+HwSHvXXy12p
ACxqyzwVMdMWJOl6morCAAWS23fTkJwd6Ut0qZFAztrka7M6VnLS+PSfFC39PrDN
XBlsFb+uD2BVmp1xjih0lX5p0PH77kS+5PTfXs7hMUj5JvXlCeM7x7VGjZ/hwtQ7
rk+q2Bx8IGUqhNXD8azpov7iq8msZ6SVNHpSYElTBqa3nkEF6RkCPL5gDETqnwnT
tI1VlzuwxOCGmZy5C9OZRD1HiaO5tP4JTRIAmhmsJQT3PVCwBvefBU9hTTt1fevR
pA6x8GPe7DVLASwhcyUrLFemKehMbkfALLqD13AzfMAKQXp5SBLBEPtkkb+lKNEL
ILMldqe/WOACr60TrRHjZ9Y703yvAmuys4DCTKVlidzAU4U4yBNWO/eHvnEaU4GZ
HkvYndQl/gaHcqgFy7Fdj+0oBO0xv8dh34tlG5YZ2S+8qo0AMYFdGW6aKGcFVnHY
REVQomkhFTqrqR6IDiyMcLNxrZTMo/PX6GGpcmy3MbmR6a7YJWv895zZOkOvJXLi
VUOAS4nTHfJK33tcEJzMgZVkGv+W/bNCaUfYTTRI2CwHLH5k+Looipw+uZtOZAhT
QmgHjeCxJSO90tixT399i51eEXd9XxI3H1Y1BFHmTXSnGr8D9s/aLawBwpGrZUQO
PMOUc8edny/ZOqfeQe8cHIFmed6hX+f+tr8gClJdAIiHVyV4WlmGMMZUDRlcn6x1
WEYlAIyIrwXol13N0IF/TLk86g/NHirjN6nkzpa+42KXkK6HmEijyeUislqZEO0d
QxuZ1rOYvLoMQmuLrhO4iZa1r5V+oGkZJjjNi+JUxywtcwdQpfklnnuH7G5gpT5G
H1B5t1HBnKDYdXR3A5uEN6jN0NJuEn8FQnuNvrgxT3zOQhGANa5BI1MHjxetdOTy
L59C5UbwLuFAcBoCkWZ/q+Hj1xguB+S/4d0hfjuXlOY59MCZsQbEaI1CpiTYKiQ7
dcxWYXsLhIeOETCikb3lWt/4EJgsHhVsaZVK+nyiWfjNSRXmfbHRwZE+Rrf8cYR6
Qhwu8Hzv4fq0OP0TZD/D25KvgpBzJrZJUVSiIpvkga9CF/QbiaaYXKoNRiWsXsjY
P+gsj4SxkOS0B1Mk9uZMXyfOKE59/1BR+/R3MPl6iJqqAE7iQLkrbHcTYcP0anYw
/sM2A41kvypLKb8c3XTYuowpLJOY/mcrvKffurM1O/Y4iSpYBLEglxt+2aL4JJu5
vqAJZX9VVrQAh5/DgplxbUABA98r8uTOWZVTZfuxyEEcsmN+79EnrpV+IS4TxMfM
euC5QbJ7OUsGVl31/VRm+1U04px1D8TH/c9d0ivkYmgjGIiv0xfwejPsF/oVru6L
3zOuoUu5kKbUwiuSqhaPtqPBrHPyUWMchPkR7R7+4bLkoIHdEWysr5r7ZNoFVxBa
6fPzkTjno/kPyKauzPaoEFeqJEaNFeImLBzi+ZwRVIEdiihreZYXrEpRAE9hlac2
RC3RL4r2VNyuZKJIz1NJTmGGqMftUkJb50AoVeDQQhZ3tY3c02AtWMe8ikQKT0qF
L/C5R1/LA6H4cLpj52+NiJ69BN+D+E/yVaRWI4wQxjIq21DdIQaHdcDqDkGZuT/P
GF5NIiXnSV4F7BOuxsB9No4VD6M7xyw4jZCblYDWnxr++vjEfyHL49MgG+1CvU4i
EcTw3eP4vcQLC+p4T7U1jEHr6dSXILJFQg7XDF9UUN/w36+hNSGlJSoOrUCViW7A
lV9KKD+08BBMmNm1lcTTc7dnpOnB6S7eG8fSqjxltZKtXnvzqNcD/roIQExexfGZ
x6I/SO9Eb7aedQ/gF8tBQ1UMiM5vBOrqplo4+7QRytPFmPEcrQidZfesAa4DaiEj
O+NuBv+0laYa3HT2S9JvGijPjL8kCVO7sdNd4iycrg8H7getbfMfQ+wEe8UbZZdu
NbrXZ6xUwpZ1wE9gH5riMk8Svp5bSFEsU6JbGJvU83zOQZaL/uoX2gmyVi2rN4aK
Hu81LnPIgxmxzOcipt6MzTwwdLgZLwtkJeHTzwRR8ps9zhoJKz4yUHL07OnOQP9I
ft94BP5eYfVAL6Ku+f1aRxG+F2mM8/wpKQ5kkelVLFJTUz4Gs1FW68CmfA+v009w
uOKnPd6EdCQRMCvA0Pia9OlT+oxOMsZ+enL2kfV5OvsmxGTNzRPJVRQ3Bg1WGL1n
Iz4gIwV+9dc89JncXxiDrjsY6VmbOg0P6p12HjzebpGQyDLY/7T+1R5dJ57PPae3
hONxpkWYufbLqr0Nzgi6Tfg2Jwcm6zx0Ddl30TD0etk36DG79PK9rKDhrvr9qEOA
Ygxix4OsYzfpR9ha2z5Ojb7MuUd9TYR2dQji5PKzIHaS235ol/YxZrtBGRnf5AjW
O164IkZFvGiWIG4tI4cIVG0b5XS0p6vAy6YReBvufqUAW2y2i/2OdgHCdeSLXRkQ
oDisK9uQSE66b9OkwPUxNMLAyVJEkjPqYLGSQKA7sbIEailnGO4Y4GhXHzlsCye2
6ybwL3xcwiM8KgTwYfPfJThHw4Nz4zk163za1+pLAVyLgYT3+XbbAvceCVbQyj+y
LIovzMH31BqdwOXvk2hR5NmJdo9/22ZHrTQqL7R+y1/t7ZC2Xh1CMaZvPNRiDZ2z
V39Qle5uo0j0k/PIPSkzap0SM22c/n/xVYZGIPGs/TGKMHJkMH8JtJ/PgFmLi80c
xjckJxyK/pAKtPVmu2AONB+9sffBXGCdOrMMf2dercBn7DiW0jkeehsUUeZPqddK
m3Qh4A7cB62pxdcCKfsP2u9Bysev9D5fz1yQclQqZtyBvdRrMS/YSSocqMrnkNUy
Ezt5Zxmq7y5fieihKjE6HgisnBw9AGACY4E0ubarXRxQp17L15//GIdYCXY+YeL/
uL8A5Z2NAeNw6SFeP489YUqQ3VgfI3GYdoXKl6YtXE/c9BPIKktTsm36vU+0zgiz
7RrGlTE1bVJK1qrA7kS0/deQFW17NUHbgc0r9F794V+9UVY+SB8SBypjSfsgSnpd
Uskfb5jDmy72hQj6OL6n7yYo+7LAcp8WKPUx0SKf1mYpXOqPMRnfnmLAihNRMruN
6RkDSJT8BHf6DsV5T4UTUONniRhDMKVNmsIdgODJjyr9rw6ihsXB2N2gG/YVGR2N
dfNbMe2x2iSR3xVdvHTb6uVTFpJmqk1PZzZ0KGGgCFRQFxUgeOlpXo/AFFxM4axI
1ui9J90YbgG+FIZcvc9ra2IAfZoUrN422cOgHdnkot8FzKGrdzx+jD5rnNv5NbsU
pMfmVRZxmC7LMIruB1Mdcv6sriTB5/+k19xc54yefE++uhB+ugP+oMpqZe3Syogf
R6d177Xr9DFZUl0IUNw/MvsmLthwgqxr/NzXfzjOe0iqLTBmHk2P5O0GX2G+EVt1
6JcrJM+wU6B74+JzZYiWyEFkxTDxW4p3wLUN9l+tvLk2X+mfEvsa48ve6nLUyM1k
J9zumqCeBQyR63esomWvhs+3MAPHzHDq2jflpYESIP/veoODoTfzDzhlO9uA/a3F
l0EB/N3k59KcFBSfowz2AAgapmIgszOgmiWA5oQOdvFZ8ReR4LSjZqPqGPfh/Npo
6dvuEA6eyikyrqqlfcD9bS6Oe0JxTq2gREH0iU5kAnigzwnYuaEpIpMOcXHinven
0RtVTND5e9+c+bHV7XA0shp9qzCnYaVCZWSmEmZG05zS3rfvCjR6PSHujOoBtktK
9e2oK/+Y/59WqOzlcpC+EzGCje4KhQdDPLQ1UJtJ8GZWsO93TuWofeaFsuF1DdIl
qw54KpezYdwGR288eqspnnlkVAVHu1m0nhhetzXmKVJnCzYACoHswYaCho+kUIcO
EaxHL3l/X7g1XmGTtABD67x/QI21YYP5ObVN7bVbl9ztl+pt50Kd8a/cP+yWz3CF
1F/SqpqVyi89iHdJN18IvDyvbFowIElC0nhQzKDU3TK2BH9Gn/NCZH6uluQOOit9
GKUedPC5vF11Dj65WJ21aI/7xJt8MzaazkDu5QL2C84oq5hgW/IwjSGgipHGvboc
1zHfqbldNAqCrndViDVHHhHweVqV4jdGaTEsIMYLVf++Z7MeOagYHJpHlFhFaIXz
KEcnIKG2VJoASWhd7EvbQg+ALRT9PBIdpROWLfutK7pqBDkBTmdTH9nizNwzehPO
LrQHZ7Zwim//p+rgPnfncTe9GTSlEPNB+dh3g0G/bolBJmjQPJ+b0UxTYLiIHexj
p72YR+o83K0Ki+9+CUSSSP3nv07PnjeAAyOxA7qTVlBUxkGFGVD/PcznQj3jii6g
bO7aqt4GqTLwzpEmUV029KE/HXsZlxam2xAgZAyoK3rMFi3/Uno98/PNd3KYaLrP
2nBnw3pehYyoFqmxO6rVS33DJx35F26eZ15NkxtKy6vGFG1lppVfDRiGPerlv7Os
eBYhbBoRbJE5GG1gaERsx1dtqPzQU/oQMor+zw7I+YU6J5EZ2JuqkOLk2Xso6xb0
dCZoJpfkH5n+nB6HPbzpcGB9qL90QXZbtjhJtn+ZbINQRseCEWuaofXwfKF4ydFz
rsKg3dDSjjLW2qz1Qa5Hqd4PaldGOQqsrZCCIqbcyjaRAXfyYTjfRA4m6iMK+/Zk
D4Xcc2LaAjVX/jhX3lf2mZDnAmQKhe7IzWpWnV3fODZFBvlPXdMLCcfTjZC3a4g4
T1aLxHStwPViAcABOXQbHA8ZaIr531BOrDpSCs70tFusEUU3eNNCkqT3iJXuvOcA
kBjz7zEv5l8GTC3NettD5Bt1GljWo3n+PuKYhALelc3CH76h68SfDrN/KL2lqb9V
nH0h8F5GMOJqCMEAxIyLv8acgAjm0afB36CGK8l/GrQrFtlahZQtWMJ5/g5Ir3m5
yIK04b3OjffpPsd3/mdU4DRkMroLO4WQwge8ls3u+RNQ9AA2PBlR2PvFI90Md1UZ
Dgobvw8I+4P4OHrbuw19lMTPFk90sOAYI3vnNtMdRgZClU8oPUZCBdQN4GttUWtO
pk1S92lZbadk+Pl6od68QZ6fsTs2ldg+5ldxo6AP3ELO+1fJNlHy4h2HeuD20++P
thRDchdeOT3FSqmjVGjhVsNghIRyKUfmmUmkiw+yQPhMHkceDNEanBl1p8JKQR0D
2tO9qe2Y+A4DHm2eczQWVE6ExQpAsmfPm6xtRgRqfL+dv3lRXz9qFskVXqrwyqv7
mlEo0jJz7UjVExFL7UiCKAs21F8rSWtumDRqkXqDKPkHzOEACGv5VWcycF+wylkV
VSyn4Tn+mLsPNdm/QYNfg7jlUdNGkNc9eYWqxyZd1LOd+aTBrDM97tecU/n93cP8
kxcGxTk8Q/y39Q+D7tFkm/hZbAz1YL8lcbzxp5uM3YdxBJy3Rr9PBd9Gx3PMph8L
COZXzkgg588K8DJGcqAWJrSizLbDFVq7MaU02czJFCcqgd9e/KRcf+Owpj2ROpFj
PKQKGWPrzzJLNKn5qxov6wy7eojbqoNtLQbB1tF9a0UmmYVfK8T1k+9T1QVh6Twn
SZX6E4hYeOgCPTJ7Q6eKvLVA38PWD39Qm5t2fWa2GVjWZWY5GM0EwjcGA/Y280yC
poByoqre2PPYtSFCQW1bGpyCaBWcDcqxgOO/pP8ySWo7syQBRutS+Sy/fVGY8tg7
t+lX5oWeM8CJ08gWttabSEfeEGdI/w6ZVADQBfHCQS4NGqaaug18Ut/MDjzoQR2s
Se3MSuOMgjzz1TJG19N9DXsy4Og62L57KwtqlnNyqTh/n6yLr04JZ8HMTk+67rvS
KPBDbQqw4v3ZbLSdDDNyDEOY8VP69pHIajroZ6vlrOsBYsg2SszKnZBnmXeRdxqm
AAr7xXVqwUZLuaqb/tqgPg0/clTLbiBVD780V4ARS54Q3yVPRHLJgL8NOO6QSTEc
+QiWhGtwk5OxCa+hjr6Fekf63G3w6K8EppRs3VHdbOigZzAbnIxbp4noCdYeN/hU
5+1culyPPuPNYUs9U7UkWGwucnPNwF5y5f7JhNyFGgKILrAcxGD/cPZqYZDtqOz4
gaDnv+JE959CRPy9/uJ+Zh6oQ2OnsiX1TIGQLJq4v+Fvc0XbAzM/EGbO7sd9JZjA
H2ERKX7RAJ4E3BnqBIQGTwQx7tv1ohG/Gn93HGynYLf7uHjfeSjDGXFmUL7cnUAd
fqM8hQmOhbrTPnsY7uJF4SjxSVhn8ANsmarhS0bG5nbz3LXJYlTYGoVYA+8p48+Q
n3dHIteILlTX/7O2IZM5D+S7UbVTFbQJdY2k2E7grVqankNFAomaMbNiFGNNwAUj
DKnD3v90j56bAL5acp2DSkNEJfccAyNc2aoqezsxOV6G69qpxbfmPbXKJxK45dRV
3Nb6aHGFDwTMUwPHqZyXJR1Y9VvJDhQbQEN/9TaZ5qPHWP2UfkIxFFrs/Y3ko/y9
4lh3UsKRkY5rZTO+Q/qDVYgNh8xuSy0QfswhVSps+4d9ozSFofOPiMDMseTpSR7M
rjKQ6j4023xXAF5/S446HAVibB0hCTLF9gA93MwdV7Evl+jP5CAwlPgWSW85MaUH
RlXc6fwVUCaMK1MmsC6OmxWeYVfa03Mu1jiK7y+MQSezX6SXd+qcP62iXS9ju2jO
w2drzzUBabAIGfDjoUn/+OGVjFvHxglR3RGA1AidzixofD+rf9BUTp9m9cTDpVRx
cG819UAEdCLKX2kCm3SgGpKoXJ8Fg5zGH00XTeVzWSBmnxBT8BAYp1XCTT+GIAoT
48tO1lw+IIUO8AMVpZVWf/xmhahjffiNysk4SvYwRtgfuBzR8qcxEAmPVOKD81OJ
HL2K3K5+3foJl3F12T/hYYfzJ6Ds3SKxDMesSdlgblBX84IavtRRofN06CFLQnYt
JAzAId3VYcdPxnsUGTDk8GI24stS7h1pbGv9qNZKtbgfTg/pljAD8B7SRMBU80Nw
guk9L9T7Vpu4VQ+LbHbz7mH8kWXaPN6xskUVQ6hUrKTulrpplI2+2IOPK5zCSyEe
mm0gpnPfl/xCgOA6c2LBPnXZhkuhHsgmwaRrpdZ8bQotXtsXLhqewHvVQPiDfSAD
H4A9lwp4tDEumJwRzbXDdsWqJCttNeshlCzWBbPjeAc55M1Z2vpqGGjKPA+9xVa6
W2RBZ1wDAwkCe2884YMfQ4yWDCrmNLeKYWvrg+GW/Jc+yKPVIw8UlrQ+8eEQdbZp
RwPJes+8GnhrArsabDiC442NyK8VKOTMxgcY1JBrIFjga4R2rf0jBojPjfM4J+pV
/ZQIeKySOlQgy3/WgX8ug0yRVfELZITDoayWFj8lwbbaa7es4E6gf8vR3LrHRSdx
NLMBl2VfN/zVVeEEwmEJlnlaDp6S4Ye0lca3vC5HqTefpe/rooGEHXUwUh7xTJ5N
yrsylHU9xYwD4p3pNT93cAv+E0kC0YEPtks927l3Z5jZ1e3dC4cv3l3cPPk7iMgi
joQOchbmKdFZbhDH7nnXNwX5UOQ2KSJBqz4IQdwCvOpClXOfc4Ht2BtoqJrLWyXB
sQ8s/4hiBp0lolIvZXbF75yIs9l8PP59K0uJTBV9nCoBlaHV9Jp8NsgM9DfvHdry
lNTujwbupgg1BQ8mWiZpHQfJELasaiM4z1njAT7ZMpvqttQT4YlDul1yR/e1difq
eJdaQiGOIdpkLa0sN/2ggG3tbHZq/akrwGtV0J+r6KBoEfND67KPbcXF3+AvxBKt
DtKBRnoZzGfr6tcI7eiRqQ+RHduQ9VIDfuXpu6C13t6vdRGpptclfAAm1erioBn3
xq6BurJYdsJWEQPR6HEdOSHjHSHhDuDMwkXQ+600ZpY/pzu8k96Bq3HYLf0pXZr7
d5GnqLTN6VFqsvbG94HltkVclPM7dTK7oUOOC3WK8SU1k9QXB+8+0Hp3HPu8tCCX
awRiS79nArNChJpe2GOJFokw5NSWJvE/0z4y0MKfYf0hbH+/wRegTWfPRDwE+6Px
h4EX0Q5rq32bHA4XpLUCr5CuBlF2hgyly0Kitd+vdKtLMauG8dFRVuARIyLT3u4p
CkAeVyVrx785rOPEQMB/SN3NmjRuOblhD9i6uwcH8EkTuR3wQRvMLGiGOQdwgz5t
AvZywsBeQm98p8S703xfc/VV+fNciwHuL3G3o7Vxldp9noRWJQqS/PqciPDwGo2H
P0/bCIO4tfubiL3DLp2/itQi/oZvy0mkOEbYNKrJVkoMSu0uA2TBvkqQR7bTMDGq
KD8FXwG/P+jtIfX5ttpS71D5znxdCixrppfvuYEXJRr1S7ycSazu8R7f7dQYqOXb
lTNMDJTggk/sqd7snpqs6zdurcaJ0EcjWs+Nl+6+v/u+JwOK0SOG0HaxWDtwG4Sw
+UvGpMUQKReuI6MSCOtfnUUKmmunYCnDn+PYtRa9F/3tFcXxhzuedPGGAXkSCxc9
PvEw6Vsw+FTlQmFqg0JJg1cgIzWpNGEX2L0IBYknMN4wd3xYOTVWqdDXjuHe8dIC
vbP7nsbsFaE09cYTyaeisdGEDwz5/pYYAFoyW/9Bfg5uDUhe32aZvIEFlyHm9xxp
WOprpIVx6RuSQXxC87Vt0p/Ru/1GXVKOh6ASXKuqGK7oPWsL2IBVOhT31wWU/bGk
OBYwGeKFxM0HcFUF4vWrGdiPor+lBAysdakHacGPIE6la7GEal/J3xlj3D77OvIs
Fb84opP4zeBcmMesQJgVzQ1gwx+WYCfuREjVv4rayfzhk76qZwjR0v2+86A6YCki
NBsm5mWkgGkXs+lXZvna9YFVDCtFmLUDrPSea2/C6YfqG+9GloSEcSBUruifI36q
K5QoBBXIDdRfzgggpEtJOoeeaOfR00qrmGViblV8c0rsg7JgHevvnQF+JlXjtSIt
llisx5Ynk61NfIBpJhb5sTnAG1O8gz51zLXnSMfwniyOQysgZfWrmHNNRufs484e
yGGzX/mQYu2iRLB0o+BHeA/VG19MkL0jW83WMi1BeQXKYwHEIWmf63QVLEyTCVEq
x7hJM2ZTx2g27VTL9sU2+tEQ1/LbvPPvZs18rZHoJVwgMoWU8xokXZvyBuzDTyMm
Y+zMFWYFfaHIp6K0jZMIXU7/pYcbyVRmR+J8iR5XIJZKxekLaU2RwBsLS3yC4QrQ
GnZljp1yWQb0kHE5Cu4sUIWMokof23hrzzVhWGHD4IP2hCoFEQl0L/7i66g2TDGc
oeAK4goy0MPhKEjMvQ6517aZrsmSU4Tag152cIS7vafLEj3eoEhod6Y2xxx3QSSC
D1Q0D7DUcbkSPYiJ+xvA4YQ/uHjisutHI0/mFQWyA4wpl3vX5htnHLNLLjsbjEsF
DbIdGwXbYpakQ5/c+nfzeejVk+uEA88NDv3dojd61bazGI2jrP+FbIpNh1NPRphZ
akVvfbClCzYIaNtFWcoVKkBOQH2ch6WEQmpevxETV2t1PjZbSn5QYxtVYkniH8OO
gClx5hJ1LU8r4kIchCaGewbXoJsBDkdYS8rGuGW+KgEvKur7CiWdgxnM8AWwtAXu
8WNVrBhr6vbi2QNvb1vCvCTdA4+xuWe40X8CIdDFdoZIVMeJK3lQWB2ufFnfJCIE
7CErchHRn+uqyRNHvZTKjW2pkKQt5T1n4w+VEtoQg3pbKnpEORIer6XpbxhIEz/N
EH1n+6Tu710FT3P+Csv0UykF1r19ulgcsaVq8e345Imu+QYPAeHtD2t6j8e8DRKh
t5Y4wObXUu2kWbOqf9jUZQQnPUjrMxdDHxVG+AzNYkhadGLF+JYqs10o/8XH7alr
rW0a3dsNWOY4wSeRsCKgpLDgW4GaKTa8Ql2OMXQqZb+4FBEKSCtILKl6fOI5c61C
OzoSJTu+q6eLlUv6dUpPF9m9DDkZpkmXe/QP+7SMNSggcFYMABYuvdnPGK9OREy+
H/o8Raj+5CZKj+SCNbmWS+1MmbWbsCF7EqQCG7P2ZS746v4JwUr5yQRv11UX2xyv
sCmKERw9P6uWmyNlJjn3NPnRymxIiqzT1ceY+sROIXczTerbX65gdsEuP/pSUg0m
IH7UOBkVWjOzGq3V/CYI4J2tKHmqrua9V1nPw+IbMsQOwYIr7a/oudmWuN6tzt3P
AAqK9DMrwJ2ppgL4iBgy5V3jSVmDEOlTdsZ2cwcXP8S28YRxgxEf/yLeG3DhIQlR
DRafwt8VZEz61Ehj4VwQTHmSVEqIlH6l1ogW0LlNO+aSbtQ1XO9Dt5Wsup7qTn8w
tM7sW+59RyYZW28czB2qx7JwtA42mYNmx7FuW+CCRxKjlUgk4Uzcax2lILds4dFj
MXyTW0l1iyEiVsafK6g5oz3Z/ro9BtQmk5e9zfpHbGVhiFX0DPKhXG6cXcrGOr8Z
WQ05xcJPJD859Md97z+wJaz160FCXfkhQ8gIXXi3uwVXd1HswLeOPDk8dzJgoru4
GvaHAZ69r2aynJt/WHNs9PR7EsOKc7Umc6zSkpZXmkRn7U+69t7bYn5HWCT6KmjF
Uv0D7nclgTZjatrR3y53TiNJopvZfcZfL39ih0ftD08/2Vx8mRX7/WuEBN4XXTNh
py/gR4Cc2chynHv6bXjU6EpFB6nzpS48P5TNGO2lx6uaA3qWnKm7KGjKePDmccjn
YtLrI50ZZ5AnlwdisXto0U6l0YLFj/5ZfU8kO5UeLEVk8BdJpV71ZUw2IeXZvmRy
ImDRFIwQSOWgNLNylcywd84+KSlib2eRYL8jSzlqNLwLexT/D/BRrkgGom1NJvPC
L4S+AboOGdJujSnILphfoZo+EryWfGwWUru8HQJuxJqgzxeEG3GJAHmiQZ8Zx3X7
Bm6l8lPVcF517b97QFpzfyg4yrEd6ZCrkN0fg2HC2l5y3G8n4Yla+r73jcBv3sRa
kMBSojYIQUTOelLxNg4eB+d+e5Mc7BGrhYuDJhvgA9l/huSPHo13VsLYGJ9LljpU
DA6W1r2g5dsXnz4Nvr0Aa9e9KN+GKlcvre/erbhS7Aqy5ZzJAcZQjvNFpiqeCmQr
Ar7f9G0qmcPZJrC5+JAuCG5c+8DvqQ0SNwM3Wv0kQciWw5ENP3XvKoPYYT3cUbd+
4X/CTz0Gy42K8mCY0Tz/UqMLtmBiolAtO6IDUQsXabu4UQmy42mbkGXflazzo16m
xncSQs+4aUhLBNuHVTdE8eGrtMyJeIKoRWjUqC3luokp2XpsWzv1OpVoD7aHaUZ7
iezv7+ycQAOmDqZggXQyRQAo/HUdVcj3jgiGr6FkVQL1BDsVQkyFpFeA4XG4ETUP
eJNJNP3HBVax0Vv0qFz0nkbvEzJnYpX9lxLtTyvsv4R57DYjEj4V5gjHNQ4Jdhw1
HHmpE1ZQRD1p43BDqqVs1m3X9yoYpSCHTeOPkuqkpos6Y3AwOSONBkV+Yv0DUHTY
vdDCScscFwBYNAuEvmzY6eP8xlm03wlTCm1FTk+WaVyP9AuSSTFFwM0F6HfwPyo/
UxNNdl9w/hEsyf9FE1D/E79JZyDs/DRKopzBF3Jkk/9bQM6q/rLXyoqh1LYQCPsy
8CLUsWpFuqA/9hN9qbSdjLbuTOENo01AqMr3ETFq9Oy5tPP8xL7YOyv/p2cN667U
AcCAeqkL2Eb5U8cxz+7DSoDXqsk7gI3j8QpIOKvj/E5aOSNIZ/qNdbwgwtBJA9W7
/q4kka9E9XlO+w0S1uiwiU9VA4lRZ2TlriXIhUtUgybpnTqCC8+r53ZPcDUC0zWs
RalaWCl7+Yxux8LsyTmCjHSfqpbQybcVS0lLUnaCGWmcJaqFniSqfdUNnaETweK4
oOQAfq9slRUs+ra3j13phYB4/OvK78IU8Ht1b2pZqL4zvLqdjcrmsT54pCCfUOj2
8J/31oxdgQJzlrgDHwkCs8gdtE/gBkqFcykOPD0ue9HMN2Stle6r8wfCSgjuK7th
HA9X/gJkCdT06C+RslOTbcK8rn70tbcYLlsiUOmSohtWZFDn6tclQU3QiqUC95Gm
bHq++lJ+mg9A1p6CBLwovVIY7sJRDqm7kKR1FCmb8+kKk15ggiIYA+KhOHgUu7ot
Ap86L1c6KPugBsiv2tt9sJupNh36PGtpi6fpO78BBqU9IcqyysHmnqR6oE/cIoaR
X27RDGt+4qqmgxGzHlf5qsBq6HTzrwPKiwfE5nuT4uyVh8+OkTBy5QdOpBKfNVPR
8G+RrIrTBPXzhFoL2w8J0mSc7b/JkJIdhMT8cvtpoJWhJpALs92WumELXFO+ceNz
T7EzadvSa+EKoAdySNZOaQNsvOZwupWNyMel+nWIdsmTXvu9GryaNkCJ2G31BYXC
6gV5jYVrVjpjJZLvH/qd9XYjhYKjVzL2w8kECZAK4wXoVHIRhEqjoTVljTBXKk2C
yiG/bv6z/S6UtcUS4kDXmWrgaAjy+gqGjrUMQ5X/QsF8GSTXFYmU2jg2I3GpZpaW
zOf+gqSQnENkwk+Vk5CX40enH7x0sWR/GsDd0YtHW6H+UdOrRsE2HV8jOpfw+UPA
CQzm+YUqFBbPasaRbjIQrGDs38gfOGXuI++WA8tCAG5My5lquLX7vp+JchPmhONa
c/htZx4bPwOFWpZdgbe4ndYD/hu4FEh1woeMidzaHYIy8aiaF6KW4tya+bSjwxPN
qC3iU2uQB5EjNkl7UdBz4QEQIo1ILgEWrJJf762LCfSC3USjsNUyv2QW7o4askG6
PdMRBnT8Be7IstreC89drBIAQVAyssbzQTUJR+/4SEMcA032g54KqqzNM+LN7oTH
bvHgDT5RO9pOQG2QEmGdD77Rghu4d2XhvIeSWCiuFQrXe1UD4CJwk7kMLumE+41d
CqjwlLPumnMedhGU73NjIor5DZq1AzSgWbVrZjQpudaPqlrVuOF4lhqi1Q6dm3QE
rsC7xod5y7qpwEepUD03Jq90PPDh4dQoGeNPOClwywo3KIhHq3yS2N7C2dePY9w8
m/f0YXb80TW1nPOI9fT+HTR1HahW9kdmKWxSiGL54rwO7MnSeExEBdKpaqmprZ+q
79VmbAugwQZhr0qkSZcW+VeJma5E1bkITFoEIMSaUkjEdm7JVLX9LCWE2cgIvwId
StWnP+7H4DZDzPfXPrEcJJEknuaWI1C+AKp2OH51nv+eJPcg5DPbH5+HT3XOJTW7
qnu5/Y9/ZljmXtktNNTDpONgkeEFjKO1WjxH7M/WBUQH+GKYClzFN3tu2otQB60C
63Q4s3xrxbu7FmcwUdUk4rii6O0Xk9KC2KRxUoRojdBwb+PYuif57M2zwD2QbQvt
mMwpe4t6MW64bMZDJv2riHMHZ0H6N8faNWCdRduZJly6v3EKBQTWtYGYRu7a/3gu
4ImKnAXI3ynwgTkfv8XS5o64xHHnyznWX0eJsQMSAPpdWDiZd4j7cIJ+W/Prt0S2
f/GIHSDi9VNtB8LcQI6d0eij2259QZDGhucvoHMPD0D6IhRsa4/oR+nKgRBHB3Vi
BaALojsJ9oVIS5JrcFp7Z2bKpbMjoi+hgjIjnuUGXRmH5GEQBMp0+i/yKWqhjpc3
fevEv8GRlc9TXrvzdGanb1Ia1pXeoDt/+KkJx07CkFQfzBYyIvj108jYb58B85d4
720OwuefWZKKCMafQoBnUA9xeDgBSFTG3ZXaCVvSxNXkFnf5Z4IDX8XW73YqmEHQ
yO3GUo0GSSPua1CY063Eq2eHkbWboWMDxJdPukiB22IfIZO4CeN1tsyJGW5mbb57
Iu+/LRNf50uhLowk9apoRBSqvkk5No0+HOOP0rhRyq56yOEWvo7o+R90AXv1rNGd
T0h4o3TFh3apKzgHLaHYhg21vQ8L7hcxEG1y2osjJ00MvthotEnkC79XYXgNR/o1
zg85d50O8NmvCXqWh0eSK6UtOGlPZeYdSOyboZ7bY7BhLjbiYSesf6AmOupxkzAU
I9CNO1YD3JlV3ZHPpQJbhHpWYPwasw3w3BDFN/1W1qcmO9dfwwb5ixQbGwc7DYux
3cFmfeAAsAu3ZQKl5Wa4DZPRkpiP3B7wd9oiAPFmNQPww8rTuo1irPtyq1gM9PZL
Xdf84iY82dzCNJVs4+IiVi/9sVFQYB3s0mDET1wzxvefM/dS5SW8DtMkRNmu094+
q6L6Upt6eRENi9iySDP0100QDfQJfJ4akyOUooC07eXLPFCdvZUDt7BNhpAYvoFb
39ODRKdK/iqaADeo1ATXWBkaVeJYjffIwJrrf0E8JRDvWv4XEu2Zo3sa1F2PXd7j
8lYccRkgq1ZeEIEgCY9DudTqcMSXHesX6wI/2QSmb9AvH5SPzX7Qi7CYXONAbPWi
ow0sJFYHbRTNGqQLgRmsDmbAcFF6CtwUiCP64J6j4visLCFbBfOOpTMs8dsRlvXz
tL4mIwp6sADFamcJr4hlX6wl2BpXsyLJ4wrjFwK5XRNJ+KbIGiu5YHwoie6AR8/6
DUmRCvPOYcoQhDB/cgmCiIpNf2FtXtT9umlnggVwiz7ItWx3Eu6/0fH898DWxsF8
6SJvUmW5xD0cJTZ9AdLuJudStFrnHuMddSL0rvK7Ss9acveGJ/W6IHpxFpuiIc+V
pfHnqw1p5ExBEBVgd9r4TaYdskKVhsoNMm8j2pzwgOEmtTZvWZKbasSjFajSm9qC
K1zB8GHt0sQ3GBNRwDuyJfi1VS/glbUbdv7nS3TAF8JpVGbcsd5mmq0gb6rEenQM
nE10FJmZ+rNh5cL6kwt7ld8h0fGrcwq8Kxg2Sfg5hbU0vzJiCl2Ar9RVTm0xlyB6
/vMWz0otSgiiTKhA1zkmoi3KHqbDxuGZ63KfVbutix9VBgFFOVEtGqT4hnV7EWjU
gsBGOK9M+zjSqNTJf947rHqyhiCHYw3nvdWeDTjONrpaTPLk/OdC4fzN1sEwIu8n
pLLA+FgeA9vqvi62sfGgcfKOtYjN/ci9BJ9dOutVvPo5+XOhl8Al+t8SCQy3naKA
ExuPl/GrPm5qDyHQkbgHhZj1k+RfddV3H1TwKHpWBY5BFHB5nLgO28p8iBr5+e0b
ACOGacGSnrqOyCXez/cxInOmlJIjlSRFvUCWJVGURa99mC3bLyi4g0dZP7/Ppk08
ImQNamYGPb9HP7Dtir9Ge1RrWJxpw+7UotPXnJ1gWuSJIyEe6muVpZeBdunH7hfC
7bDtJbdC6gFxYE2uyC0QERBSJZK/j8dyobBIsIz94s+jQ2GH76ECEBjdbIPQ2D0d
ECW3VS9dKvkdeefwb86wTVUoY3kTfcC1Kv1MVcgBrdRqqRY45FYDjLTbXVSAA/7d
FTzBFlW2G38fQ5mh+7F74BctzobOHAS6b0j74j9an5+GnCYTIdhPOyWEarFTsiws
0oJwW5Ymx+DD1/74JkoTx286APE6GpgjcORPI4knqXP6aIxdVWULk3hyBK3q4w/8
UCHmLvYan7S2wSLbioj2w9eCb918aofJHcYPwQ4z6j8GZ9iuh3OXk/0hgQvuKvVs
1aXji5qvFLaknCKn+QtnjowSqnblm6gheG8zuJt2uZaSzktCaO660fukdBslRqvK
SoEJ48i/tBYf1YOLFWUlr5b88jLEQ7cg6jrmdumHxxJO/XEiNgAMtpu3e2anj3J1
BZ4Y8Z6aNVkzikaM2emZqeXg6N7td1+iS121KFXcMpypxxx7aTaoc8bbgWrMwALV
RFlqYOwLjzW1hUrlHO6ScenJIAlgqdnM3baGYBD40gpNtjjIQCvExsFo0PLImsuG
TNocR/kqUj2MEax02STtkTZPjgC/TIZEpmY22FpWQnHLhX2RSkrTg5lSfSdC9DUv
zalhv+QLDxaDP5srb5fR+ak46I5RadYKhWmvmSg1nX/CqV8mYl63l6La8/FQZHSd
rl0Iv/0Az743jHrOMzQyn6BcKRpCaSQ0JX/WZPF25OhhFEsVwbahRNI9hzxIeMhN
Nx3Ch7Fg0PPZOiJCPgSmRCkSeFQ5cLmtQuU002cdgJ8GwBnt1LxszJEX/b9ToOkR
9jblfIJuI3Ab8icAbePs2nr28C5dTn1i/ZTBqa4kMHzkj1uSkn2CC10eyaPzmxz+
P0PiqtanGzCqDguHFIe40UNrvwI29vN3aG6D73UxuRzrS9aR/BFTIikaOkMxtui8
pABO+vpeq6eBYtnhQTuEAQ6uWkIvPOK9lCcj7p657OhbDwBbwdb7SdYJeLGSIeF0
6BBJjA+cYwoyRoHAwQG3w6xy2xXbuRqsEUyjK/RNdazXJoKY/ye6xPJcuYfvk3t4
qFi+0enh91rFmyHqea1bb6p4pgRgH/IfaE77CXeE7KhmabqmMwb6OoII/Guh50TO
qQfMR2N7jMuwU7QurKqoUMjEIiLu28W73d6OEpm1fdMLRo2i0sdQ5gAK0xTbUN0g
3Fnjb8DPdjX5mEDpAuODwqZN0IBznY0O1KkA2I9b0GcaJgTGYGSiDaXLN3sNewGm
823/aEHXraII6RdZWTCTwvxSglR6ndBGQtTcRtGwcUenHramWQqHT864aBQhg+SU
yEJvCeyGHUuVdJmHf9Yf1mIc8oTn9yAfPaWFKwUc/e4gazDypz+MrmyBkkEkeUV6
EQn6JOdVR/51qjmPWqEFS5kiAT0iItls5wyv288gka4NKm7SXB3PwvJn/bddGm+E
CP6MODii9ynzYdAdcOu2b16UDjnTTCge9kDFemix2N9SrLCOW5QgHbZgUNQmlh9L
hPnu+a4frgugOJrgdwWrOLaXo7V9WzvldDOZXjwx5LZ6N/wnmoV1/sYSy5Y+O6aO
7Cph4VglnBrlyw82O5xkh9wPA9wylr3tAD//UgcDNuOhgYzFXC8Bmq3MeSkT+NOB
ux+Ut8/sJq1hVKvLS3QJ/hj8mHCJTEzapQRlIKuwaHxPw7kbzEDJk0pfc0RmG2sG
PFJiDgCAYKmNtXbjSJ0jN2kfFWfUOb6ML3hob2hfvc7ocI9COFG4BAxsNETics4k
1WqSOmvkMXPQ3CCdWuRC++mjTfnx3o2Us2VovwrRT9C93SndToWv8BX0rRnzRmi4
KOVOXBjpt5Dm1RDGDyFX8h1ItkQ0WWUvPKd9iobc/zqlbbq0/tyconDbm5sC7rYl
p5CmfTqmtaFC9ba/6GXBEuKNBTKgBexRvZ/cs4xVNpZro7JUBRQADyS9jlZIuFsD
Ev95NF15o03skP7x1i+ZLsenhnsRq+xhz5L8nREVxeWXVIBNLgw24ZtTgogS7cXW
KfAhcDlfR4Yui+oyz3IyBitRxZGMiUfcC8f70388hwOKnEMtcqdYR/z8TnFuTi/X
vfxgGXH7VJbxb6BKSuOKJNB+OPMAWMfWMT+LMDaZ6SdX9cyNKaDQaS/1KQKPBxPJ
fcEsjSChiCzZXHC1QizOy6vaPYzIrIY/3ga2ZnYIrwvg9yBR89KQ0vCsV3Er4sIS
06xgxbP5wRhnn43MQM718cKvkW9fT08hzKTneCeEd1ZUSTHRTLBjSrHr+y4Dc3yH
eZZsJ0xlyriaJEj1U/HLVroz1q4K0bb2CJviqnQFpB1azfQ24ALYI1UQCJWlObTD
GqbmLOpoiKF2Jv0gTw5CJn4Io0QM4lJxI/PfAuu6Cfts7ATxOtVNK5sLLqWs90J7
ybhPAaOALPJ/XTvaMVzP5S/PgCraXbudoGtXcK/OTnritPycDqUmSrlnipDTx3Ua
7nxEFZLjsM8PhT1fWwqytqXw5iG9+wQLwe2J6AUNo9BeH5j3q2UfIPyG+RKsr9J2
ehFMW5BNkZ7TrG2kX4zmNdZVpL6dZDkmEjJEeFXIgfvacAN33l6LIWhpgywU8y3z
59olv45mbWefd9SO3xkINUTuzMo0an5mv5grf53pvfLz6DoOOrTngTENcQsp6WIo
iioIjjYIc5S67Vv+mMemotEL/bQRybZ7/6k+WNyA0/sYGN5IBLyGfGBF4ZV8D6To
byepMHpZJ5v1zPJvkfIYk2ySgrOP/w69fN/w1hZjvXS0B3PBgdrE33OuDcRx7vw7
W0W1irjSCQ4ndlCDTlm6WjiJHnGrUhkctHVcD0uSosRcEq8zLmVpCLR5KcRXyWOp
NYUS1Zk23t/sRuWEBfyjoVO22Fyy3DBUnlZDEXGvi7HQ4gfKiATtO5nwXNF5ZJpf
+BJD3OneH+iiNQCilbPBvSmbMZC0FwLEf5YyU+tqRubg11vtYLSVh5/uH1bIqm4L
Jmp00aCAtDyW6hElTIRNMKzTogDIXZtzEo7xrvLFRL3A3XAGp6aJok1i/xepqgv+
g1w92tbZBQmerERs/UyOZvc3TEqO1wzB4QsG7FNuvo4GHFTxTmfkE52pFi3Ocx5i
z+oCWd/3DviruyCnjX/1KFY9F5JsRCUaZCfY9qFqMtotTiTsVmNwVHcpiLJM3gGb
Crp1zWqEZif2X+gJfTCyvtErOpQcHD9GqCRwOYgT/8xt+2YOa655u+u3Cnlc2cCD
/uo5BfujR4VDen9V4Ku2KtnvjNRT+VIP8+bIwXZLvRcHRUUzrvYHoW+VpDboWGu1
uK+Uq4sS+eckFddItOhXL/OIxqgdC24IMpYYOm9zLyCdM8UGLT2oDqGGu78PNbWH
Ugy9YsKtv7DHygNswYerg5FFYNEAFpt9bmt9xsRVJ/J2+7s8+aj6b74Hz4pnC3CW
IxxBBqWzjNqCcfO9NSRi4uDNs5c3BSo1906MUpBPq4b0uzckKY36Cl08m6zeaumA
Ig3tr71DcC0b47v4A5ahMkskSpK61Ih5ItGhnT7XHwzd5za6O81cJhtNb+qwzObW
UEE57okhYNCH39b0F6z3mgluB871abqeP+7PUHyCgG74nN/Or/G+iJ+y8XBvTgtx
hzhAjACXlGL27i2D4E3Qg/+b2xux9RTc0VRUTcyzdWRVfCoHMu7h5o1vsPno/ryQ
QwQiGT0KVi8DLCk726ISuMIIsylXG9XjcWd4mUWaMFVIYAauZcbvKqP783bi82vn
XiqCoOMN/8StT+CV1EryR/WFRtYqIz1VPOyN6ELp4JY1l6mHDXfD9SdAtA2c/pSy
ekOUEEoAyAMX1T67+3NjlVxVAHwkkEngnWs/5ER8qHGWXBh/RUGAsBzX5B00s4zP
U1YAo80FYDFdOGIZ/m4eEzFX9cFQD23ExoyMrNlbLAYI0PLL/JvXgOfurjRh7z6L
H8VMpSanfgcwWsnCLYwUC/oT/etpzCTkr/vKOoz5hI+6ag0YqtfnXCn4T8REqe+V
C9W7CtBGedALdf9Q54OHeABpjBBShJid4/OeONgtaB2elCD1v055zchaPorCG4qa
jPLS9C9TtJlC/SvSxnTuSASJQvfvG7hhZcZcoXJqqIHMIBUdQrMZs9H3IhbnKYeJ
PboleXN759bkK7WIYPXZtGg+yyLq7GAbao50sGjUnLzVb46w9HtCZvkwTRI77tnj
rQ1Ysw309raEirpyrYHU9KSNWAscb/bJomqmJq1f8qPmoex5iLDUJrhl0Mtu9JPu
EGOQ0bo/7Z8BoFM9vMOkLxDyAgOWnaslg1hjGuCzU9Uv1uKtZD1/9wMUX3KQlIAg
dPz/PZVohiV7Ews/2b+S0gfo8DJfWm/ejjOpLmvwznka7stqaLbgv/nVXi2gFPlv
GIXZmdBEKHreK4Vpy+rj8+eKOBA8lyj2gE3BJu5oDz+bh/E/IIKTlq17kq7RtUdJ
wwYxSgAja4b12U0rLXqdFrH287cKesMUQ2cM8SXlZ/BFJi9M2dAB6G4gQwl7TmDR
Y9obxWzSpzLdebpTZo4HKKUte7CW0NmWprhcK78M4dYmQ4SzoczECRW+gDCvmjpg
XuD48M6bLQDyeirUS1Vmz7z9ZI0U5NvDTl2RxOMScFp4zniCOSLXZAQmC9/t1diJ
hSU1xd6zirfjIs6tdyBTytB33vAnr5Pbaq3FS5Nl0iUPTNnB40x98MlRj1dwRQ2O
dAX6nDBOQ8Z0Js/WdFVSjOnsCERHqqg8J7fOZEwt1hexBlumVNtRxSAqrUWHgTnm
ifFlw30clDqhtReMrf2tBMKEZwNTpm1KmSIbADwl8Qu8JwT2LhaUvELCR51WCZuh
vVM113f+b8QZdcQG1W3ahYpZHz5B0I4uJEYUsJF76DAizqQfTjGDlnMBQYX5awZT
XPagsD9AsqLZErQsP9eA3cHvMWUATXcUCtDwjG2YNy7bsCNmXfZl7F2nHp6eWc0Z
IDOKJzzITXPXtQhmUhUySqozDBzIBDlx+3p2Xm80KcALE7A6TPh+FHsLyv+NrMuF
J9Cxf6tZbDzAdycG0QpqcqQo1xn8Ja5bsP1L8uO8NwOmmBDo98EYOZ8I/SGgpsVg
cjyoEqSwUizKFhyiZV9YBMjkj4YV7AsGOrWExWNewiMomV6gRSKiKgz2YnM6NgTf
44y6otStbeRclpsTusJl9gBQeWv/RCZdTHnrPNbxtdqcz0oulpj5CICRBH7BK2nC
SCKTgm6lZ3AjBw3pvp5D11j6BOFK9kYxRjGide0O33DGEX9HHlnHH5YzLzbXBbPi
Cw51jMO3JLsHJcJexlT6eYdP7uMHTJ6SPV/vDefawVf6BG1Y/Q9s4PUNaCkBxnYL
uX4THkiVGvD/thSyhS7ummdxqqUoksgq1LD58UYe62Ip9jkFNdMshclGozi0fcD6
coY91LZY8imuiY7tNE/rRn7jDGqLIjFwC6cctQFT2VcDfnOICWXh5YOWmGHq0Hm1
/LcPjxF4TA/iyGN3LO+0jzXqZAYJnoEyabZWbJMUa1LkOmW5ht/yVKj6UalhDzMP
RQljUGbREXtIN/aER0SNXZmKzmn9SK8g0x4vabm6w44Ux8o1YUcXPEWFO9aDtHsb
v/RsfELpID9JzGTmWpdJoP42Jx+jvfxGB4iQO4AE4DcyWtpu/C+C6s/moKaFhhlY
5w4/7nh6EdeDMXmk4ZJ3BOwmOPAgDj37VEP/VzngV5CpSpCUIL/H1oId6dUHW5GT
u0QjbGaLATdRMS0idK0jH8U3DBsyaHbzYU/b376Clan3yytLShAp3saO15KBLvqC
KKbU64wCIZGqAKL2asMZ1JSripBhj3JLABmpv3iih40qtr6ZXigQdBRZhiXUrUxq
V+63P4VrCuZkrM1sbKqBPL8Tkrz0UTsgBi1E7aEmglckr8FDwEIwspJdzWxi85LM
bgYjWYaIm08/crcOqB7D8f3WidPFutJVVo9kQxkMuJajW+KKXaFUB5zGwJgwsAkq
JtVtaSdUL/PgDwzrAhyaY8KZ4uX3LTSeUxsu353oQnDb8mrBm43Ql8GSuMOVivD5
Vt7fK22xCWfBaF0QqpTqTxJAKaRqnvAqxqjlmNnknITFkSOzaJZjpNrm253recDT
NgrBxVVvNTVh7/cpuM2oZXMKhc3UksOShTSDT2spw7Y1D+TLC8YF5ZaDrPeX9WhS
KFGvlDp4/nDQa+RM5705QW9O5TrRG51uHQaF/I1RlQjcLgNLnfvNGFQ9Jtn1Wc6b
I+8Ohq3aa7RMXcUkpVMdgZ7n4WB0wpI+8u1jVqYW/Ifg0VlbXWV/YDD8jMi9x+Pm
wgnwxQY7VtbFISIliUvPpIc0zNR1DTwOYNx2yL03B6B4jhWPNp9BzWxh7AdhBqzt
rpwjh3GJBP0cBNEuK735cUb4uSMubTBVLRHqlyYXGR/OURsyJnvPJX1EdH1anVWa
pgf+ry8YtiqaQTk4SyZBvL/Vg8h9zrWFzyakDSBYGD985ITUW1vcnxYh8wF7jA3F
qOU3fteuIXSCgj29Kke9oodjR7sJzxKc7DDylyTWkBZDcT6FlvjNq6WxMH+dpaC+
H3vHzpcGjK2ciBjeTlxODkpz8dxlBvb/3Fw97KzwvyzyV1moRAG+70TC+/DvdGaE
+vMOG3GalwRdN/RvVafdVOR1aZvVbeMwHsKCNN5z+OIT9szBMFRephPVWoILgnOn
0Agrf/CQZ+FTc/C/ogp4huEPZDXoa5t89H/nre3FAYkj5tDToAjLd0SXW2FYnR7A
GfvYbuthUoZjqUgdOcHMJs0+S+Dv1KzB58WGETsDZ9mvRE0wR5RqE4ivioQqa/AP
9+fsu/DW4bw5buyCkw43JW2Eq63GL9x/cgJfQPWWEaGE3ush2/V3b7RCr0Nz25AS
qQY6SbK4kk7L/4xaA9yctQpZP5iAFB6Dyknh1XkX/DL4BJwWnQJ1Wo/jDXk66Teg
Ny1nHazCO8gZ9lYwIIqCPyw90NtNOrLnOIFbGZs8eQZL0PdXrQo8ZnD4lzCwUvvD
2cAHVXRKojMaoMqjiDyhn2/woqY56LiVCrJxfPL2crCkW9ImYPFSVIX9S8p4mlr2
H5cM8WPoSZOZRZR6hro02qFvVdVQInncQx3U669rRJ1kvzG82grRlS5PKh/92yP+
Ga82UzsyxA46fXLOJ32LqRaIp7ARkR+QjsKfyNKRmaH251izbdE84+sqdJnMc+n8
8KKzDG0ky6i33sPKkGu0ETtsDaSAqi4aJP5FStPrN6Vf9dnH8/x+oo70ztUw6tUh
/LchDnwSHBrI291+k541savP+FQVyTy6wvfFE4r4FPahST54T1MgzjyG6j/VkwSJ
XyRFsZZZHRkTt+FnJ/ONae7AgG94hS3rd1/iBrVFQaa9DGeSvBh0AAxt1hDjDy7M
SuA/qm3h6m7qhVWSxHNZ4nioWD6a3BpQS8ReNvkkUrRPrcwi12tlMbm/2STR1Sp6
y84XKAYazjSdzWuihYs4uWweKwdqJNoOukZxDIuTVqUV93TcmhDLrbKWwJwwAOax
cAxcuBRxNMXgEQygVX6HibdTxpj+iyTI52lV4EE8FuHHm6waxUD3CDLV+pw67rbj
XXIH89rpBqup0518Lu/vu2jEfRGJ5icyEiXUCqFvrnCrkaA6MsSIbRKhzs5G772J
Mr1DUfYhqWVXBQoAEWjqkMtyi3wVJauz6rMPo7fcbATmHTgS1cAHvbca2c8jGrE1
vexC0CPNUgsnvgzXs/l5CzZMrBVpYtPcL7kpC6BN0gsyZ5zDI4Fzx4POcS1iHa1k
Z+OcfFciUp3HdQfp4+aMXDF83sPF8lpEfQhNxtVXZry7IZAc+gc81Ikp7+T4v2Hd
+aK5G7VCX8fI8e4OVHmVs2Q6weDwya/wahnJH/+2m1SrGI4wLKdWLQocdjgDP0rv
G1bIT6aw6JWioLJoJn5JQkmCU2rmEAVAgI+Bd69MuE9WBNIu6Nuarpca/ggHxV5N
lAz73gfQ3B3CU/RUZC38DfYWR+WVsREO9clpySKhpPqLaBiSAEJ9iRS/oCseaEdh
mAGMEiaB0GcB6JW0Kh/17kTlZrFTMKMMoFhWJuM9WTs/OucyrVks3Z47yiUASrO3
5VOqGVdIsXundT2kzk5qHSPQXBHUYdA6R3rB9ViI+HUfWt4BOPGKrg27bjwLIpB6
oDY5i+voHRV//Rg0FZuz2xdl/Nw8IWOoxMHzggwqrm9cQbXioYHFo+EcO8EJoQrB
5yFYB/CUJsUH13w3OAQeew1/FbS26ieTyz2c+f4tkrscfIm/wylMNfQuSXBYA3ow
oQW2QxHNlVbiXLfTHd13lPvH3uiWjHfEP8jC0LfZVbRtD5yjN8jmKrCM4kPkfdGE
j7MtwVGH8eYaiBWpiDPpCSbVr/AlSLh5PstAM2SiiUGMMv+iSXfNGRDW8cTAfjBb
BuzUWTTOQnQvvJdTL+FtaDkEntieYfxfGUFuXGN9TYD3jMyRTrzC3/sdMXM8iJJB
lxphVSb40Ebf9QloQQGL4kQ9LekVnerWtRaeTBqiUEEIPF6+dfOB3OLFIYGG669l
FRc82bOuyM2w4QesBFWUdDXB8oVbHVdylcLfaoYD3+rnu3gqphmyfHaKo1s7NtJx
8avUE89MLXEU7qlqimJR8d+est9D1/4Q3d+O5ItYyAA5Vr6FJImgoGS4VjwIWGE5
x4IWtAKH9AjyrxkdAnHMVSa+XeiDGkBghe67l73S0SJnPjVbUOEiml0Nh2Mg+3Qg
/yHZUvH3gMFped0W2V+ptxXtX67FkEjGEAWTW6BsAqRdljO9T3Nb6lkIwOkYRZyg
5lXpbfZ8yHh0CiVCrPS6Lk9/WEOYwrl8jeZQgxSSN/JTSzuWJzf8EqmdJaH2GDTh
PwdWzMiw61AXhfHFXSUi8J6hP3/S27AubqUE9sVfFPxMcw6l4Oi8SF1IQ2n4OKrf
N3QqnN1+uf119S1H8Iu8ABDSudmQkr6yQASVdeJ8dWPlvXSOiCdMyA/JvyEuyrZ8
htabwuV9klevdKuyiB4qkzM+gMLrrSyiNIyq2IpF7F8y6pl0RrS65oac9qqeIOx8
UIqVZq5QgQ0cZC/pizmqqdLJcnC8mekvslx27j2tRdW7UaZ/M6gPEh4ANSG81u/u
bBPpjjk6bSqkvMgj3P0aMVh9JApleg5PQ7q7M4saOXYDiNgMkgTcTEIK42sVUjZV
1tEAWB25R6qu/qStxHxxIFXctYgL4zcdflV9b3R25FPSRZCgCCyoBLNuhm1KJp4g
Apre59e/T6K3pBcnxy6PyocQtDtER6GTty2+VBa4iklV6HOL4Dyv+9jm+UvIu1tp
2uXqWcgAyYMfEvs+T6eMtJAlTHh5Bdh5shSqSrJexB58dAc9lwuIV/jhwy3bmV2/
biYq3vXBU9/7qEAbURMCd1aNkzYnpzUucZkqMi3Uf6wn1Hu9zDtac8ekAn366Plx
ytsVp338mkZp9SkMNBFuh5WwPPHIyEQRsetGRwOxe35CBunUV8sxIkAcdbA6jfqh
YWRuIbUzgsIkPpzUYsOavo3HHvsHtYXXje8Qu0OLsd7777pjkXolFV0/fV7nhBAn
qJdAH+BT75nr33UKrzWAeP5Ap0FF2W2LKIlWkC5GDAfHr6BDJo7tQrmpspSYLTEh
zJqpBAvgRkEPciWUkjsXmFD1/q/NxluXeAD0+GYYSYbTPb1Ivo3YNHUzH8IsC6QL
C8Fw3GCF/E7hRppXQwemtIX2vV6ADgTVVvIjWivXwJzOV+ywgpdq/keHNxPWpDl5
YUj/rhIoAYoSGAMPQM4S5kyw483taYT3jVqVAkGynBZq75tv9wNYSzFTALZkm08o
qSyJlW/hzuv4TTnBUlEfC8s4aGB1EImBt1U+5Zk60fFmP3/7yyLv/K0kyhCN4zs8
inkLztOjidKEL0iOSk5Nh+U3d2oEeWTV7wGwtqPLZ4czno4vSf06kDYbqzU8O1dr
3U4/yraJs9zKmqsZNii7R5bvyrtJfogW9E9cQrezMyrxN40aggeI7y8/H95pkF9M
jAC875XUj9jneG8zxXw0CtziLxPz8qULrARaamSANbFyMljwiOcnqT9aOTUfb1Pp
r0HxPdSZbUzkTXlaSs8oaB6htw7+bqJgGm6a31K8TH+685mMv3ogO1dBs6JedTrc
3EhmXGq+MCIrgqxPCInTG+U8c1tGmklTc0hzz6P6BAxaesgWdQ3K1eIpR9Fq5wb5
l1FiLmZ0rLYzblduvAv17sCEC13qp+mE4M22gFWx9Zb98NIv+YK55jfMcGmt7VPG
hQPGnz/E8L9qKNzN0p44GpKktChvMlnDEMzLSYJIlHVKWhLO0oyjChYpZwMRPo2U
Ki5GaaPRGgTc7BLCDMWcStUkZWsamH5zOum+2z4yQtnUgXAMp/0odguycaldkAWK
C98OdP9d3ljY/9KY8R4/iK23b/NdbrYXIbkfneupdZfpeR4SLMcMVmYsctNC1Eg6
rRENXi4k1icrE9iuc56ViqDQTjfgK0Ca+3Nc8LQQdGq0bkjsrdG1Ngt4flpUCEHc
IotHp3N06khv3n9P7Fjw7TJuK6M04NAOUn0qjMllGliWOLbj4vH2DnVqhLrOoT1c
PoLM2jHFsMQ66BzKkmeU8yiS3exphiVFzzv9ClI2xmh3+7hLRxvqH/pahPkeo8u/
viEVV/n2xhLKJE0FfOOLnzLu+fC6ZQgj54D1Y09MpvhxAulJr+MVpgqBjXoRggEF
V5Q3+EPeS4tYFNni/axWmvv7Usmt3qWL9HJ7W3PHYGkIwI197jSbVaGHyYSW6oM3
9CpahAvFfIhfqNo4UlZNr++iNj54E2DeO2g0S5o51qnMJ2UEo5fuEQEV/mZkf1GA
WK3EnjebLSLb4NSIry4KorEAvq41g2KdHJRpX3I0yOyVxmFfxcz58VRtplabJ0HD
XpDz3IqDQk4o6mkM4i+i1vsiGqW5FU9nyJKedAtiNsXvI8+rStdLbPTC8NvezX7m
CrZLCVehZnE+4+9PfV39/OzLm/TuWTccIcLX+dslm01uAex/pHRofRA3GxzdUrF6
0U3jdGRneqiRbHqqm3CssGE1YpqEafc3CeAmlcO/6P6uXFPUM25L4Z/6YOHeOhVY
yWjZ+exVqvUQd3L3I5Sjd8L/YpHL1IlBwXPzsgzMck5s7rerd6KOkoTwgs9IVcPT
Hf9/z5+nKwd/FxTFQklwfJHa8qn5lkNzIPOfZOUI11eT8b0tVImuPDLZvY5D87Yy
eTVjqUHGrdql9Zo8fLNUTZHZwICqkTb3QihTOKxRiZ55Bqx6MB7sQLpuBptLAO9L
L3NZHqBAE1Bq5xB0F3ipR1tOGZoME6KrqB1NjKM7ebBWYt4rz60EhLR5waAyL1Ai
xiTpIMLN8rln9IstNjp1TOuxoso8xvXF8Wmh7R8u3XmFgopZk2gDI4GYREYS9nXi
2Zmoj20M+CaLyvk9NTxBRyR1mhjgyxOa4j0d5hxNSgxS6DUfu1IjBw9d+lRxXl1x
QcXJ1MgcT/D0Kin5+2DFKhdCO1GF1XS5sxPUQ68trA62SpA6IckEoNReYPZdOkwp
77SexxPukvjM+TD0lWM0zr5Zkf8OQzbzLKNOgh77C7bob8VWXqtwaTRLEJkRRfzv
fzUVX7hJbCHYAMMXr1NACA/1kTO2S6ozbSioSJweiSxPgJq2ZZLuGL7jdzCuEHQH
iQQmVcJUi0WbQRvcqaW+J6RV3Gpz4JBDLsfViUq2miytsW5PeYgRMlgRzQftsB2Y
u8sPe34HQX6jZzuC7Z+HNsTURrdg5b8z+PYX0vZDKKCpdLcgKneni9yyR4+eT9aB
Ooi2T1PoESlFK4sJAIBTOcAoXr9/mPyBNuE1K0nGvP1SvqzLWO/xlP6JbfNPGIY4
whK1JJym6Bk6DWKqKz2chQv3jP3CM/pLaE7GhcyNfk0Jw1Qz+6W2Mc1e481Vz8Y6
6HWvUnlEIe3ikZhcYhr/kcBaoC9Ipgf9CgJQTdaaczHKRS4uaFWvIIo2U9RgrqID
Ig+CCzQn9iM0OLymJh2OVJavwXSllvdxIzVRQQ+N0goGk8FSeSZAL8yR2uH39sYj
Gk6Rxg2G1gn5eqWNlitT5yDl18W5QgqgVJj2q0NDtpwZWYrzP1nMPPCGIV92TEpE
LZZSXWvuHvKv3IM6utEcHrLRzQDlOfQfWPAn3xdRLxBUizSrT7KLQrMlevqHqtMT
WdD3SDZt5j/q2m8bUnGScYTFv9KdhkeCInYtomRK8rjfERL7TLa+T63qfZhHk9ge
ovTBFf8qX+yeRIYJaEnPNz61PLbn4TpoFupTXr6+AsfSlRzXN9gTseNKmqZsGC+H
6SCNL5/xOloeXXxbIsmQu2pN6iWoHDPCnA8ISRmO3R6P5pGjmWPYUuoWEQX9zboZ
yWRTGUHqm/72rQBRzPvrmkX/xDebHbJVmETW8+oze1pGZXT7a5M2AnsvxHg1dW4x
j2XIJ81wq0pe3BeqF7SL8R7jXIUue31IKZ3RWzeOyioVrAvXB9Y8gNJLT7AgzSJX
zkMjFehPNZsgLddqY7JKqq0Bi4wapfG5G8NE/WpH3JRIEF/E+sKKwfxzhwwOm9oO
pdr4DXlSeJZMAOYwksHtBELu6koHCuxq2RUWprFjaEAKK95x4NA5BhMNCXl6qWlo
s4q0dZVIdarv8MTITF9QdUHEuN0JfFhDxEux6+5iQNtiKe9RfpLT3Gv/l2dDb5Qo
1ko769O0XgoDe1crNLXPXFVB4zJr7yeDv9nCTx5G8FMtN1pQztixeyg1ORGGf5Po
iRHnVWzpP0F+EArZfHhin6jI/PQGb8QW7rpmJuJ0NftEppTRyv6BWfADZ5v+ZQDJ
CB0ewMbdlPuIr/tNXH0AF4TWXDr+/l1Hanm9aHxsVm2FgaLB0OlzaiYFx0k3q3gq
Rm1C2FZqh6y/ajYCCRJLwImk9IiTi5kVWjjOyWVDQwGdSEajFxPwCecbumVGT0h/
2whEQy1/WgNeXXpjfbK3AtEWW7mgd5U48GpEw+7SgYe9zO9xtZKXz/iQRgL5Ge8f
MVGUD11PtLY+J996OEyrpROjSJufUNwNUdb64pICe3r7SjWwaZUyUgOmhlTuHgF5
rcafxomHDrxuQR5scRCHHPnwTtea2131PjhDC+3DsW8w4vN/R+UXmQCu06LWr6kG
inAI6uSSHQRNcWKwHHHyvP8QbY3B7LMu5nLhpedxDOoCCUl4b6zhHJiEo8UxuaqS
JXguU8AZ7MxCs7ydNfs6Y+XbBFr+rvJv99+7F9VsFI1w2FUOgWbl9O9/LDeG/cSj
y+u3sjtKvAiv6Ff/IIu4TAnDW/jSUdRKKgk9OyvG4Pf/Az/mTDx92M6zaX0plB/O
70CeDH/qaaBGOxSr4AwW5SKvacxJAu6qc4AKGQr5SNZxcktLabf6g3SDhyNhA8iW
fDAI0XUQ1guzLentHG1+z170uRoDzRybZDWs02orbjOl5WKN04mtw5LrB+WmEKFW
dZpxiqJos1oIOl/KNgOeBWBNG4T6W0onA066+W3O4zoSkE8IiYzyrZasdeLq9DF1
I6U8nYN/NKUCJ2Mz66Ai/vSHZ6EbEI2wYpikzOjOa7+Np2+2JmxILyjl16E2jv0Y
y67aVaYPWm4jWby05NpX22MV0rod7IO61MybmDDDYa2j5Z/FLkIKCCCThfEN8jk/
k0EgLI7ky5gSr8dAeimZqWhPoAEB74TBfluwMqcM8Bk1GH9U1wdCEUMoUctNq0lD
9R5EiljP8b9O9nbc1L+AyJnUvgaAHUeIsYWtPE5+rCdqUEswrqJ/UXQfGQYWBH76
S8emtDhqiGJykvo44FZ1E9FBHyGUmD0J+xTPlBRrUYl9D50kdAGxYzhLgSKXAD1E
Mjt9YJ3tRpuFEePNNKd4en+WySZ9pprCDZNP4j3xMFPtz/NPbLp2C48QhQgEXdkG
tH/JUiYQlWBGF3PcTDAVJQFHKpxvcTz0SkvYj6yj8QtIKhbWiVR2DT6VYi8SaY6K
4J44GotZwdatfD8JrYIefAYU9QKAF9GtZhXeJYN0TOFStqVh3lwV9HLzFIeP2NeH
/pzemlD3m43m47mw7knJ3YpGLbwn83ugihXILWgx9tKnHLqHfQdkiFupoY7kezto
267CSJmP+hpjPk8jXfrIcJAzUv5CkhWM8F6kXFwTQHnS++4tYKaBB2EONczqnpMm
NuoCj28tGlQItMO4oRE+/bp9CxB6ouCnHIhvMgsYZIZI7Ic5ZnE9o0QSO2LPVXvZ
vUkHwFLR3+rj0E7CQklXsQ3smNE+ZP7FJiiwUTJw06F/+inZqe0th+Z/W0TBSdyT
2ROcactpPu3kJ+/riMaDKy3PdbmbnSa9CcAejAZwLptl9mwuEbs+A/XVhQqB10pp
s1z0YNTL3Aj6OdPcXo4BY22gT9XdPo1dpheBBDLKXqI2qzzXwjLEBC5oH3QSGjB7
VOH4cmSiw7PVKQ0019eolncbkaDphZ4KH4A06c/XaZAvqX21Eg+3GkefhWTpxqaY
QzZvBOcE4Bqzv252M2RyT174h1MRO0SrulfofHkzHJe/mff6TiwXBP0rt0IK1FBY
E2ZgfSyrenU4II85oGeeOZQ9c2lCpwHU2Eb3NW1YkrCMCaMh7AWFl4dfh3CTS7Cg
lv4kBOu/uv+8tRnLo9m0ENO2GXmQgCOYtbfxWaqtjIQblr8Mvo0EoKYdVhfP9FUN
+XasQFuJmylGzzfbmYgamPW/yjD40znsavotCEMJOeu8VWlrIkk185fq6a/p6O8b
m1DUhLBY/o8SUmCZBH7I/DJKPNkESaRLPwCDysX6X4MX2A0TIN+3aCNoC3MeXtk/
4z0s454+CJGiKf8xrvb4ZgUjvxvCTC3dCU0rADBz4aLgYcOTTNN0ANoo64DzHfWl
Jcg+2BOZTqByPiAmzxgTeSZRSAu5rIiukkqhBMGFh01w+6rKG0fzHO52Bj9fzCfc
8JxDml4UDk4LdBH010T9X7X9/+cfm2zSl2QHlItMCpmVIXVPVqyQZSZBSolhJNoV
gqxsKuIj2aSzRfvIbG+K3atSDQUhYgRTz0FPl/eFwK7Mkr23M/yVa6maWh5PbrjX
9wZTDIj+7PI3NhkaAUkfRSkS9bS4ocUdbnzj+PhJ6kxVCwkNeqYbEuU3PL/9BgAR
WfigltiM0kM0NGHX5+mD2CE44gTo8pVSb6+1dbq+SJRIMVA55TZKrfj1Kbkw0wEv
FQzUYyIl/B6bg8C7qYG6wF7U8ec8QLXgi2dpOEXxLcCpVR8LQtHtH7aHOtOCO2/S
1Ysswz8kdMQtWuwW5cOOjjN69fKDnLRgp/A0iKZYDCbvIghpi7vHYGYnoUeX5P/b
pXAUQmKd1/ywXjU4Roo4JgBmk6BN7kKgvSokzeS+PVfVo3aUN4oNZV6h26lHDLTk
hvCCXXwLolReiiOs5S5Wo/uBvwykTON4Z34rN/xzngUJzEu+VFjwXZ3Ak2nJW7Jc
aJvQejvzF590Pw9wfQrVqBtvJt/KN11X4Jy6GaO/NEbdqImVCgTkoCf38zo/koq5
dW56JP0j8hMnGJ41w8S72UcE3S4M19PYk0Jd7e5BjiqBapnVMtlDV+HRC2ZtO+jx
TEWaIhDOQqG3ThPFqj70GTbT939vKa0lZZgxlkuYrDZdc6eapKJj7GcfoZ4Josf+
KrVx4j4nECfAD+I9THsYs1IQIW9e7Ydg6Dg60HUQpulC7jtAKEAF+PrrAzkC401J
6iADJ9WBAG79TZwuYvXukzYpd/yte7I/gHEcw9v/rz80wgieiv77XNC+DCgA7tuh
Pk7yU7JjhEdsIzEU/+Lrls8Ejc614cvPw0YSPOYEtSHpLpcC3u5TZckDcud7TS1Q
4vtka3VSn/IPTyN/gPP6b0bTB7OnP+N1WxC4OR9A2XeN6wZ2utVdxXnX18Fibx44
0FJH4uHBeQ12VoKD2ghbka2mp8uqwOfpUgIjc9Ons/yAKvyFgUVc7m8B23BUnkE0
YmCyV0mznKh1kR4R2yf0dN8rcrE1S36WIYYoMxnR7vMFbiYlBUNSIoxtsCYV84Fa
aa5BDgp9inn3Zks935xAk5sjB3gkYDsjVWXwuc2ZFPRVfX47IKef+eh2cJzQxJ5J
d5V6Cp2Zq4Z+MuMWR88n+/C7+V/dvTVTLeNOjizzwR9dOGO2/xMKzVC0uf1Ub4ye
EDWA9qQJxZWvoqMlvYagNTAxkFVQJqBQrL8MGHVzi6Pb6g+d5pY9A3Vn86B6v4h3
n61Yp8Xt9OIWWDGBW+rvPsa9jML0CyEMn9/q9c1USqQtg5f+lilsoxSoJVFVeUww
MpfhpbRQ75x0Cr8JIa4TsMFQ8XOkNhPB08zU0LxYDm1C+u9ZwH4MhO7asPmg9q3M
4hqHHyJiKY1vXX599nsBi2nIHW234ak1Tak65M533dNas88RYDkGIDPMcUD6sBjg
QF9Y1HKBvdg3tLBj5xEy8I7YtXECUKHaW21mjpRKE2CFBzLe6kpDQje+9XoJnCwT
KR5OkFoTG+YIYtwMoCnqMYwPa5r4L3c8VFvREaPV3SIyJe+q+/0ZxplbwaVmDJJZ
bwQCGeHLA0ZexBwQONqTxfZGlBQK71Os9Hp1LIETa/w78AF/iGE/qI6mL+YbNq6+
/CCZZEwqnlEjUHsvUwrtJMeWVv4/eQWOpjwK4246BmaFVzdT11epPiDMXuYx3AlS
qzN16WsvAmyoWUE3xiiDrYkk2zFMeCtlTFI8od/mo0SJGiv9+tv4+nhsKqwb2zgu
y+xn+sCqFAQnan8URZKXwsmThTCd9eEBGnf6itcMKHmIw21Ja/FedazepAO+M2bI
bqUi0ospePmv8I1ynXlkwDwBsF3HEgZttlVniTscTWNTAhEO/yWjfxapv8GEq9gp
pP71UZhXCkSX7Jl8sodzNR+iKCHhZHzyzci4hVlbxsuoA6uAmkZ0hQu1YMLF0veq
2UfNafcApNWkWaHlnO3rAD1A8RmERLbRuLXPY5MWNWXunURFUxbXZ7N81w++OkLa
tyzWRUkrlAFTVh2lrjuc4LVdYXE7p2PtUlZkhEUhxhfZOwMmy/M4FJbDmGXcUJM+
6IkWb6ZH/6cDxHCjKvhbamkh1rGK4ifU6F50pVbazSQE1vbwEqjJhcVoHnPqw0xJ
7O8O8AE4d1bt6BwD2befjhyPPxZByhP2OsuVuqWgPDMxE/+C8axILQ00xVbSB96d
DIpJfrHAVNmrxDiFNDEGUaes8RvM4y85UY0S20cAvFIVQ5FanfrLTyWreLVB3sRB
No/ARj/mH9JCxXy+ngy4MPo/iN/Xw9JUVUDLwUJt+2z8O2I5K4UqLj9vgn6Jd0WP
uCiEYjTutNXX1nW1a76hA7lvK/Ktti6/KELBw0pluy2UfkqfqvVGA6Xa67mCrqo5
d1reX4Y8e7J+OVp3ZExeqM4TMoVremBpZRlRwhPB1u62URU2J4d3Wm1Um190IgjB
EdYNSBLlzBU51c3kSHMXwFOsJIwTkNSoHx3SDoImzSGWLNCVp+GjEK1HAmS432x0
f/mNpRLaVL0P5egB1gccTVyIar7vpy2rK7ahhRYEWoYZtjvmzRPcqUw5MK8YBc2Q
YH6k/FefIjWAtGQkGoSsysJmWcZoU/2hdMSZxBywb78Xbsby158BF2mU6HPl4zgD
e7lkJVHI4+8v2Q67qyu5M4QEqQfx9fuJZsJjACidO1+Rk0ObtrKe/OOMLrHKKTeH
1gGw6RfUn1YBp5oVmfR1RsWwyfReTq81sprEpT36JQ+A3gmTlcDw+UUaQyZSGnLu
7oJzhTErgomRUDUhY0kVa0IaW7jtxUfafNXl417UGiPom0yYNrZuS/URmLdqjkyL
ZbYrudAztsoiQxjiwT1NWlmj7k+PrJOOi5TiqVqCv1EWOzd0bcsEWrVgP7BuhP1W
DQ0nyzUOlrfk9KIXkr6qDMasoJLCS2udJ/3cWERJUMGl0ZUdL31pQGggs7jN7WXW
EbR9ioRywtHLoIpNdY95gDdO1GhAMGX879ojvtq459aL3cBB66ZQd9CyfqnLGee4
Enss81CsgI6rNXSsGjGDkPkxBpbgf1ImB/4Jo6V2mu047ADuBu6Q7CflAmx6RS0f
kQhJAGNhIGk+ieIcnHRgkk7q5OOp9O2k8EIgrUsEmCNowiGDomM/LSnDqnhcbzPQ
Mkh3ox/Uz8xvLmKl19e+PW7B6pQPO3GPtkOWaoXKQ/b8+pQmW8AiopGS4JgddQhK
wfx8XDdt0VRd0FYI5pmpzpa6txncBTwH6oMj6QszICSkJUgDnGhgXfSZHSeX6Ecp
R4gCQzFt34nt9PUyaQpsSeL8ICyghfyVc5auTUd2beMMsQmK74QWuTbQm/UKN5n7
eLFxppBwHiiPT88vV6NkGgRT987p6vRd0J1rij6VD1siG8rqDed/8hH7g2XXhXQk
Hmq91JW0EoQDm5b0l+tay9jGiLXUIoVz5PoZQT+vaSdnbnnAUABjSe2cRqLSx407
nxJgrUQdg8ELOMENRduT/m4GroEgCmdpPUV7Ex8/thzN7d1+nJTy7XUDRPLUh+zh
+AGRI9j7uCojeo18MZQHcBpsNpEj12RylizZ8xdcN/5ol1j3IwlbT3MoO1HRwxx9
MyRVyj/vSyScoY3eEnx35izewWV8D2dOXpPAn//OujeGj21INz26oVi1VZPRNGBK
n8ZcOB95rU7/kF1ZNh+iO2FlqQb0ht8hyXjTxzEd6tsM9gcDtn44UX+EaWGE7P5j
QBpFzRoHzf2w/zK2F0yOSJzRQKhoKff/qU2UmD2BehNcVNtn3FEFo7Kvss76vGKR
meZr3G80sOPPmj28FmR0rfqFA86k61bLyETehYNjWYuB0AZM8y1xZ7vM/k/nyEWh
xvxgKEYONdON1DdOB8EcoyofrhoUvClG/Meuph2BUH383eRtluTHaTxSC3HYqXXC
sVsuXT5eyosL2y8kEeN7sJtrmuTCJQrSJFmWIUG6f/E7sMEDxZADzVYxyMu4VMO1
Xn/ZCblmCGCZJh4m8JN9/sQjeueMHtw0rQPbBzna2VNE0AC7TxwCOihhAouyaK1V
a3OenVY8NWN5XudWP0EKpgfE+DVuOUbZxKT8hRvRb4XihaCOQuo2KVBe7o0AKOil
8znIJjV8XdFeWPZ9iVESBANuetNwYJKIIODS5NgxRseKFbruCo06LiavsskUnTB5
p/qDEiZcw4txCnWYDXZ0sMlIlj/bK+kflZy+xpN4fy+A5UKWm/jman2mV1I1bv+I
WQl3oTkI2kFYu8KkKZozYd/ZaonQMkZ8P+A7tU2x9lKrJnN+Pxps/qcQlUQFXXkQ
3vOP6l9+n+1kyA45/TDrYHTwt4lZZ9YH+GJNT1xm0DcOjEtCJAgSM3n7amobMWgp
cWFziK1wp+oFr0uc4Uygk9imFXoxoEEyOveK/foz9jzKU4f1G6i1oyYQfvMW4KA8
zlrovrPq+y58UYa+KTf/zSMhLxwuQfsbJWp/sfshKRi16H/FDeT3wblGhtF9v2yK
2I1HdVoKjE8b2wO4f/bHs9SekKXZb04iGd4RT0YIO7lcBYRCtw63UbaiFH4SJL6K
0j+9M4vgQvtFL9g25ptFNo32eKL/q/O3XXTrwXOSatNIJegpbSlIOMtgtTUv3hMg
9clNpn4CHhjPfRdHfadzNxy59jdv1AqORvX2KczyvFs8cGyw0yd7h6d+xLKSdazG
Of9oSRdJ77fYmCyBeehu0cw7AVvY1NOwRkANRlCzeyB58yWtJn0goJ6Cn8rXNOF4
xYOkcBsdMn7AFhMoXc7eU35vuvZR3kjfQoetCJFgZZJebuv+ywxyPx0b49XZ5cnv
AQ0Ss9UH8paEXgnrOqFv41ERINDsWguIQRe9/DDKmYB/rRKD2hqde8B403jsC1eQ
Ww1mtTRhRUgRZDIE+GRMXUGE8mEdRIjREZXnndDT3XNRLsyixsehA+dFaUdr8VEf
7nInJkECC0tBQerhfVlJkOJLdM/viyG1mEZ6jtGXXr5M8Cua5+4fHtqOJBOJRnM+
kuAjB5Ig8gZPak9PBBOy6cNtcXI9zXpfHUEwYN+kdhElej32Al4EMDL61fOiMuKp
pA3z7EFVtYykUJxBUMuV5CjpEkoOLz9jcwxkRZkHL9uJkfs97eXpoZxw4aOqDhoB
NmSB6sX2i2YsBk4f0L4COnUJMWUjyecEZztLRq+fY9karz5Ll8A4xOkwrd/lZ4B+
1b/jSrSkZno7ew4tj++t6SP80VMP9yL6bQbX94YBbVnJzsqHa3wq+6GF/dLgNOSi
KskVLc+S01wk/I/v7sb2S2WGRoetY2Rf0opWGGWuCTrOccGqMCny3KMjZ4wGUx7Z
EdROK0n5UtefzUUZWnCIqOCcdC4vbcq2IjaAdlipXbF6sBbi/C69J0ktGU8Wx5mg
Rainr11zKEzZSMP1gimKlWxBRrHe5wLfqGleEzt8UcfZ5suQS8LFeKfLva95btRY
00AyrWZXZsugg49sHK3vFEIp5D1mvFj8b7dpfg8/kHcCkNf/jJFGNyR/0KEU3GOD
RLpSSj0hLG5YSgzPrGECPWahuQwrvsgrdi+cpL/ZZWeaJlFC+FoZl8wveo/lsq4w
S0cKlVOmLPDM9EyekRuUisV59HuG3RLGjaZ4/w2NlsFxhgng3xIBnoC/0FVK+/Zb
uw9JmnZvUkd4bh9E7XmE6VEvz/d8HFZUmwa8J4iH63zHUlEA0zmLTpg3HA6qboXe
iYJkLkojhxbY1j9YdYp1ZeiuA1cRJjrwHqwruQfW81/qpGIg+8ys+tyZklfRJaZ1
MWAe47ilJWGm3UWawIj+WRecrgX2P5+7p7kq07gSzEotZ7jQ7VA9Te7IShjumXFx
S1OYmgIkwUEcWKdUCsVBgdtaYwKPTRdesk31dkOgexZPRk73K8WGek1INpQSq0Gt
8PyCq/KDjESm4Y6lRYDNG10LAC0iDuoWIiUr53T4+/3IsqW9PWY7n/XYMEw6IHPE
zuc6fDXLA7OMiCKtVFwMdhtIOv9GXOH7qjdSUcuGhpXfdgRWOIA9ayJeLJw8H1bi
6Zp/DilXzs3q0mCLGAjrp9RNahwTV9KQNfZpG1fT9DL1Pv5lA2DqOOzar/yXTQWx
lvgUnSc+NxqAMR5xf/Q1PikzciDwmkrRIDuLk5mYxdhAnsuC+KNwV1bb+33/T0ZD
kEC8IyOX5s2E3+WrK1JIfa6+XEwSQ7sHqAfYCdSNXviY28DSIqM8LVZOixIxTGS5
IMWjoVPDOl0/3lAIXydKKJzcrnZNmRPgI+e1/G9JCNU2yytjz+s8sAYllxZWNx2D
tO6Zl4pC+5gXMFsNWOVGGgd+f1B1hbkfx/JItmtEEkJaG5AbSvZl+bYcIHZh9XFV
ErIz09GnA3IvHWsl3/paLid7PEEBkwtVjNVLaGJUiXqdP9g2Qcova4Y0CUuiKlKz
KkAvC3/y2NGohII0ZWAPoS4Jxzhuc2yv9sHepqTrO/enTKJe1koWG8ZFl6HE6oKC
nPv8DdxBoyrRNwfa89zgjNLrQjtJwEzL9KUn9o6od1r8MtPUdtG3o+EoMifesM5v
jSotV3sDmNHFVm1CLeh9Vh7xDnUgU5Ba7RzG5yWFusz2ufu2cXp7Ll0Zy5I96ah5
QHH/80S8Q+Dyuj907iR8ldJF78ynyV/TSgFBA8x6XRNdCaxpTfCvOEpUY8No7b6+
54KhT05DPFx+iWzwIGNE8NWnNmszZinicfkvfAbkzGjFlCS5QX0o7EMxeVMrlBms
7JrzRDtb6z8QluuM9HMbdw09Gh++lVUEFF6ThVAb5wzO56UI1bTcqZJq4p45KwCt
siPFQvPpVaU5JRJvqvEN5zWRf2pIcYsWPOtIYBBPUbtchN/PdUgLRj7VU/8xk62M
XVPICG8igimz8EKbzbVxSTZUCiVNBXZg9nB3eBuJVJnv3yUA12wxZBY+avDoi3LT
e6DXxsF3o6qXkbVCy+zjj+Xyt8mG8EJeig99BfDbLs8igwFa4xwsVUDKgoQTREak
WXp/J5BkzoMPsb+3o1r72jz7w8UYROkn/6JXjXNM2obYNn/TkNwBWysvpwOmU4k8
rWW0rGRVlj2cO7x8MWbyFrBXtNLITceD7FQRXJfcyCm1RILhL5FVu1dcbCAS+EFo
nG7H2Wh2/wHXUKJo5JHMLut7fbTqtzz2BfingZrRpJan2kT7YVwEAFuql9AjX3y/
dtQLoe65RJ0gf/uaDu0IGpwSC/OozSQStpsGnPja8izmrewLb27NVBftSVYH221k
mySc4oBjVwnbVaJvVeK21s5ZVOoKyFWF9myh2utQiNTLiqqlhWZfuiqQlFXAmWIi
oDNIFE/tu/CMC5SbhntnUFnva2YYwReXEfLo5TXzS4ZUjVpubU1AWIYeebw09yKt
g8T3WoEdl8Pm42J5ciMZz8DHHYz3/cA/hkrwfuVOaHgYQbXWh3KHrcrkT8EvyKm+
q2h/+98tLJuFl5s7EAz2Alw02OOTENgAly8RW8h6Tuxxe/BoGTmJq1Gd1dYMjojE
1xMEfyANIdDfUeU+ZOIBO+NlS4Iys0LhV/dlxzuOWtzjIBr3/jRk/TOgG+Is4Cz9
GIRoCXJ9BV9zZ32K0dBTU0+2RIia0wMizJtYanQTY97dJWVPKJ0Mx73Ad1ZH32V+
hWmjxJbtZLEOFsDC/CCu0PFylYzC/TTcLOQdeFJybYuZ88856j17e0pcBnbuOhY0
5L4mExlAJBOAtRv6uxmUTBOy2C4gnULOce5Ht/EIrMpnfwi9XV4yZRc4zUaa0nYN
+HtrDJrnXrdFW5XJFYeQR3F0vv51O41mfH6SZzsu/JeKyEkoSn8jpP8Ga7oeiuXS
218+mu6edbEE+MXbhirqxD4/MRVqXYXWSU3CZjnTW2ji9l7aFwe71laCC5dCEBob
UtFVG7z6yQwO2aU0f/NP7sJeA5ySZpYBx6X12xX3062mei+nQ0sEjI+4yOEMS04v
hpgQTP+4D+Ns2W86v6cbUo8jM8D3b701P1rpFIqKV8FSTuX/FJ1ImiJJT0M8L1B5
IVEENB1UItdjKkUsWaBO55HmRvzoxXro6LCe0PYFNb8lodbP4yekFvAPGCVr+VM4
JgPZY+Xl+99RFTOzzfEv6RhfIHNveGC7BoHMT10dd+lLAGOhXGuALze4S3VVJIJw
sO8kHi0vbpG5LxEHREzWRD17ffuIXwbBeA9Vxik5kgvIcvkii83hQgU4l2495hsz
2li28GcNygdl5Jc2gPEnOpM80RHY6o8d1eahL65Ko4iQjagSQ2/qUEnsFayffdZk
sbDavJpkroRmTQK1poCnWFkcO67gQGDpRbmmfNbsM3z/iJTnHakfgRhAHYALtWMi
ZLHUbIjPSFvFRPX+aABvNvMdQiyNAV54yGZsLdXTRqhWAwFrMi9oKTW0XcKPHKaL
L2Uy9vCSfyBwHbOlOLORsrUVi3vwBrjJaODY1cO3odOroY+IejHRrdWeisl8bTif
6/2iQPf+mTd0jOjnGZ83WkqFMVdANBzLqvLfPM/QVAHB/3ujUgK8xILevo1TZOkL
kSg9XOK1tloUeprs2qrfvFnbWJyvCWFf+3Q7P2X+VunbR+DS45pMo/jnGRoG0sU8
h+aV8g2Jdy+ZsfP2aW9D+euCMfLKDs94srI96BnBm0djIDgWj0oOzoB9Q5F9anMn
gK/XpvTGbBbvHhSD+ldFnIf72/kTS69zNvP8RTleO2rxJ5bWvanbcw6hQDn5oALS
8NYU+MHkqLSRBXsy6O6mKN56EGYHnu2EY9WKonoRoU+9nucAx0I06PIvYKl5K7s1
v+BYmVlM0abJQ/MGr3Mn31Ei6k502/MmwcjvP04m4fpcur3Nq3LG7EyRUZ6lE+dT
4PMS+aeNP84D3Z4pQ4+sHPi1FZgtX/LrQANwPS4OEwkwhLFOI3EgaYeEdfTuk9Ln
UVbeRGtjSFVz2Mi5SsCpzJuGWN53Y3fvuaZhMmFVzy1MdXxy6ebyHf/vtnb+Xtcu
yCXAQKjS5WQ+EXSuPpR2Cq19XsDPkiYEt0INm4TTJFbqQnTCsBits1I3PTQ4kwGX
huQTs6JTkcZezSAI8Y2RuKXSmvE0gUl9U1lw+GjSD860Chy9JFfyZqL9tWNRbnwd
AzTF7gSfViWzE0hpnr8j1qVOZGhkP9/dyU25koRGkAHpMtGlf8dcg5Z0wlEYDeRp
zC6VdLoHVr4gC/RqLfRwlgwN25iNkFiwwOJin3d/GHamqbb6ajxn4lvp00AAg0T9
2Xw0q37pJj02b+FiV/CA1SVnajaZf7SpJTBR2Y2unCk2WGyFRXijpu9hx9j8uRgD
0lTQTZykJmtKdZ7ksH8GSMC3BIEQsT10IBD3wuJ5P2Nst7GlW9XMAi37BL+BbMMU
djiqUYJnALEdBymkb8corAUObKvF1QjTS7OBCctK/AqjMB0I1YmRvwagtkD2rHtg
hWEwb7popr2Z+X++Qnu6XYAOiDE1uefi1H+awtM5nsbASzDiBsaaMEyyRBBK6Vn8
ViUa85SY22eBIATyK22wxznlrK7NxUoqIRM2ViHNJLjJva56hNuwk2GvlwLJvxbL
2ONcSUBj9kDsUzk6A7Buz4P9rUzWHkJ+P/DhDo6QW6tN6XMQn8m0gBRMH1R+Zsue
Sqtel8t0PQrqpFovamd3C9jD3+ZokcQOn++hzUgNHQTVBI0D1Lx/BRRNQo3kZwWs
9cMGc+JpOQzhak7Xm/a13v/GuH32lDK5PrkuEix6OeJi+nfRRH2O7zctv49WOvoI
6J7+Xz9ZdcB0JEW8SNo4n4vNJ6L9LOD97gdfr0DNFdXElQ0aZK3oRYhISdTrQ2JC
EXg/DI1JBq0fE00Pzo7V9mVpjrjU5GECU1viIg3zwWpHM21ojppW9aNl04FMZwcP
yLOx8PKbd4syi2WFzJCnG8EeTV+/qKzeVQi5X13PbklOfPH0gZtbrm6sImj+QFV7
UzyBaL5TmVx0713wh1dPlV5TqE/ComNfOWwyMQBnfXP/HfsQeB/EahQIvhckmPGO
u33B2TcGJQchssL/M1JBtl9P+ljdFCQqFjhEXweyRpXDD4yhN2UNjgz8zv9Tdt6C
45f4vzQsnsfUQBYyibIAeKlctjZ6xFMBl8OjVEUgQybIGmwQ1ua9Uj2qqbmhMOt+
VLFu+Tgh09Xz7+wd57W4TcWLygZUbq/DZghgWEFYIBfM4Be/fKobuiEQXW/Qdi62
eF88TJma2I/UWRZMs1YV0PbOGbTV/2Z1t0xkRwee6DM=
`protect end_protected
