-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
hQK+7f6427tzi+4mIgTvkZQr9GFHklwoISAIkUmYta9RxFDwEzk+6tNOwTpyhBQ7
FtZpo70lFGaA34M1aCiju3fVQCM3XMwQ7xOzGcWV5sb4hfDW3VJzw1fRMVa8I4bB
7XJt6B+d9ESZNQdRPEW1luI9B7C9nHar0hG8ORWuxSw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1040)
`protect data_block
jZOuHdmQUjBcoojTHulxeexuZuRvUJX8qZBmQ2xFSdzRfVBtejNqFv6q4+neQ8nC
l9vlvNkJ0UA62+AXxn19clis543U7BJM2X2aLBbpEUCZPupmGzTxcZBmXspmPDvv
aw++qUywfLk9Oa212YPXSdwswcJmFXu0uniiH6sGi6gE7sG4Y4/n1D9d1WVkltI7
mKU3GkV2iycfJqHfjDR6OYhFTvaOPWWUpz47oO6ihPL7Uf39S9bUkUaykH2NdFp7
+33lnnbBw3DCY7u530/GGFWJVp+2guOlm5nE0I2EFHhhOdcSKqQwD1Pb6WD2kysi
JrMednCqu9oA9ThU2ulw39m8AtYP8lRpbcyHyQfEWbTQmtoRQv46vCTmdwhP4/Lu
fPOs7nJJDzF5SIa7/pFsFqjpIuQOP3np//ZzxxWLbiJbQHGsxbmSxC/AZbhYhgpQ
k0Pq+bSiZelY0jTZSnlND9QqENvq0c7lb3Fiv7Zm98BkhpFWhvjdi8kiVOnUoBVV
4HrhfgynStb64jqGV+gI/SWTEL2FF2IEtWqX197ZVtHNj1SGMiXq0dM/X6uS447G
u5NOsZ16sZyeAWP7V9cIUlr0Z/7q7lRcQd4dtaLZXTg3E7T+M+G90wCLccG3EI0t
KOQzz55LSrDIHR6ZtVaFBOVNpT5sGZwKFamuXkvxksmDR1w3cihUO5U/r9CDd/Kj
X1tA7zaPy6lypPvxAezVXXrMCr0zLnWn/3QwfrzFmO5K6M98jKDVC4YTMUF591Cm
74t6g0SgJW8VPJShTycbnUEb2aPn6I02cwCkOw6j/H+Kp/WgnGT24IIbK9D1OQ1/
9BK6KB2sLDeKtrVZLIy69MOE/A0a7o+Y6VRboVmZiRDzrjcohtKk2dypuqECoHdh
UCMZGPnieiZY8H5/wO/ig+v42RYO56lqL2CsK5LiT9chg0Dd5ATqkdR2o87HtqBq
1FowP+dG4sov7W1xyayxCcWHNz5S1PoMI8OLM58f8h85I6d+ont4M9G3SLEQt4mr
7gelofL6ZALdXSH0XCczuG58MuYnmZA9zCIBpAje5P9jgq1RiCP97stk7Rr4yboD
qibQFliLWVkxQ4D47XmyqkKfGvxMXdw+NKTVYRVmE3OjVKq9Dv4zYfL99kJbyC0n
CwdgKViW4JoEu4oulWY8cZcUYIGciT2yPfF2/bA5FlPomz8mESckefXkqYCrcZa0
UHJGSrZssOG3CzpNnBBa5Wa2md4s74dAmKDxcVckyfOo3xVD7cMrn2tfa/2yKoQi
x6OAjK817yzgJwWzHgjFnMeyaOeXl06Kmo/Ix9IB3ggXEoT5Qm4aue7AiJyHWV6E
FKdCqDqGWOnphoV+828avDIDU1j1zdNSdWHzXpGIHi8=
`protect end_protected
