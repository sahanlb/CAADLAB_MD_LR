module resetRelease (
		output wire  user_reset,   //   user_reset.user_reset
		output wire  user_clkgate  // user_clkgate.user_clkgate
	);
endmodule

