-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
3rdbX5lZQ/Rmq69vW17iCwKAd6IIokrgCcgVH2VmsmXusA2+SVV3pDuWzbkErV8e
ZyNR4P3Q+rTG7vSA868kUR9J0fbPN8WhHLUpnK5R7uzEgjVRGEdyGFwChIKCD97C
xz8hW/SOqoYHXaty8vCH6NeD5jAVB/U/82XJI2yR8xg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24944)
`protect data_block
jQHX/idWEaHk1iyGxbhiiultVOlCZIoKrIoVq8UdX5nRzEx4A9L4PKyorSZGqtb8
SCiRz1o8HCvpNXPOeUi6J+QxDKtVL0w9SCC0MdfRohFppVt9d3xCtfhYsncI6j9U
aqfhwvoAEaTATo20akXkIz2GqVyZt2PuILBO+S0F8CExjHGRsan45L9ZXox3RfXV
uDzwioHdcuB1teempbe2X9gD4oGkAn5Ypt8maqlC/SGrlfjixPvOfSIRzQe83DU8
Vi6CrbMU03NjYQLgAvawBC74wpzRVwRX55rSCy+AQaLx/rqvXXBCUKg53tNw2OsD
IAaNzKTkQb/kc7Y7vRToOWuynbN9ayzyGGyekpDG/xUxF/sqUnaeuU7XeRUWe35n
/L86OADt3eylWW50rcQXxksg5rf4iPNCc85C8pdUQn3yZenUnVSHrTEIjJ6ku1qG
V/OW3e3yKf0KNE+EahBBhoASc2AjRXiMDewSHyevuff/EsDqmpszLUu70oLQYNSF
xVmBD0Bn1KMIY2lgdRdEpp/A2dY6xK/E/WEIni4lPRJrffIPg/G/9bMoiEyrqEes
ItK5vBdfm+Ga81IlZPPPUnXB8w6sDKzC10LtUrJOsYuFgjS6FnPVqjQxPdqZi//F
VZTdGYE+RaYZt95J/WbEfLhzLTblzDpSqGtouDJAW2GdGwJxP0FTw89Z/ZavEuTx
sPS5l2zWjgxL/zif8EDcHF9z8cR/fEhYb4VNe9QmBjAKu+MbnZQvyFnYBYBS+Lqi
KuYsryv4qpi3q9EKiWe/pTW7dUs7U73KNDR8zKcLiF5LVxVOK4iG15sElp9M403d
GSRcU59FZC7U0MkeW9cmHPE3U70unspr41jfuoZbBYPB1io/AMcsDPOBxURwMQ8u
rOm2BS6qqIyNBw0Wp0qo6UaAdGWPnnyNf2WDk9/LPVA/WzfQnAAiG8YKoRchVHWn
IrUKrNwu4fe3OCtSMZkCVqIm5tCFlBFE6AFEYHdH3EIVCSYIddObhNaufyLlPPPF
fd98mlr9plbBzFwyNqQhrEAGt4tOr37DpZSbP3jKbd41hH1imnp/r42g0pq0xOTY
meTrK/qrhC4ZcfEGyXyhQQbkXhP86EvQgfMc+ztgTSbmhxaELApx6QAxWQG9h2mo
G8WLH9LIWby4c1bHBXDrlgPJnFL0EotwFheqUbXIvo4zKpMhwKb/1KpGuHkXVwKm
ja5nkNcfERs0ENlcaiU9qIIW6GK4Dkkl7a8oNw11fWgLrDAvdgakrZzZfKMUvqLd
Sqzn3qgcyrRbafsSh1x3EhncIPA8LUl5Go7+i/m+NjjLz5VfuahOtA0yTzf8DjRy
k3B38uUt68s0neGJjwlVXEdcAZC/k39iAFt9wOr22yvbLz/vwSjMpDrlpEz4+NFG
3C0mgqDtBnFb6CcwXIaa3r0Poz6SgX41msmFQqbeFm3uE43/YEEnqAaTXqZzQLYd
5vBhaX3tN7aOUOrEDbfDMUTsjYFK86hMRiUamf6dXGeFjFT0IP3pKkWkBqYG4W8g
ETka8gXyMnxbCDgyk8wImimb0j9QnnalT57Cz0A36YKPdrZMB5cydj6sJnD8nGh7
UvTtXFxmRofvLGichKAXaUqG1ZMV+P+CcOyM2ZErWASYTylhLRU9AsWpeXdLENPo
iOCF6xMV38aQYlPXhBVRGqtKQqaikymEXQFq1R4+PPBwNFWhhq9l6SCasbXb8nqc
4j9dSLL87da95k4Eh/vXeAPjeNrNo/UoNQa+zLYs0JLxzFmB7G53B7R4g/b7KYAJ
C0m1Ek+u/L0EaFqTPAUE5JbOAp7ifvjtUZEzp8asMBwKQKzMO25mkXoVsN60hi9E
u7/n98RrYRh9oG6pF4GIxICnbngsLu1pTVDjwJ8A8c5IoByiLhEPJ5ulmONmz+6f
J2MAUCGQELdqsuFK7No/3A51+AOliFZU4Fgphba3B0yDWh6a898N5dWlvXZtHv79
jfvjHEKNGaiTrtXqcNDhFi83D3Hhszkq2tf/YzZuP17MNT+5eoii+0amFxZynHkV
f00CYTfqY5E9E4XDMcYLhcCVJzBZdPy3a/KRcN2XI9xgMrtto2DhX1vrbLBRQONb
Jd/8eLJWMkoCXyUX8ZzTRqBDsN+R9iWosqEAlD/80pFDOlK02pGZpWf3gOIUvlz9
/FjN7on2Bg53msDc/hkBqbMqpUvRy6/U+0BaLLum+QIYprES1hB1UJKm7RSoSWm1
tzH3P0qQKo/bhvmTXLZEhih3f0DY6tqd0du++JVqEmD4iVX5nSDH9S8IoZeiXAYH
jW4g03SWohX6f/E5qkSWjWcD9vRAN5Tucv9wYoGkkxePiYL07boOYw/AFR1RcILV
6CXJrQFcADUfzq9kQg/HhjG+lMndw3ak79Y20ipcSTpRGtIPY7G1asS3WIKPyUT7
yCrrkwU3Qz+ABJjazatGMRuLda6gReGSrg0/SlTUz+Z27Pu/CK/KEGqYG4hsPowh
lPqLkOt3dxA8NKHfhQHOtcc6MQAMvMAzU1vxYTlo9aTX6txL/FcF+0w5Zp94qnVh
01mt/MnTdlailRS/H1R/JqRwxQ07c1rXXNofy6Eldy8fJQgnWsrHDZfaX2K5TM1v
1NLHKSyo86+mfuvGcTchABRkzbDbuS9IurkwHEht0wX2W6xWG4zeREtNK+n/RyDD
UWAB3+jBKPU+8SVzR0Pkld0m12PwYqX8ca5n861BhcYhtjCuOEqeSmm5lOFoj+ql
t/o4z3BsjCIx07erzwg7uSNH6g5I3Z+7LxyhdwYP0GhC444y6CcCXtgEDr1TzzwB
k1IoHJCLxldjyJOGeQA+L1681fmb56ierBeOmDanM7RSXQivZa+VpLgla73Ss0Ya
1a9bPu3APS7EYYwdf0p451UppWKPteaTQmgR1QAju/wdLXZEoBJ0sfsf3aDDkaJb
1LqQhcvOHcrKfiXS/H7Icv1wfyYi8W14Ufo6mpHGqZvkiYL77K+Al8fgcjJY1CY6
966P7rGxpfjPvJxcIMkEpH831FB0jENJKS5+U8zYgCOhK+YONQy6BDmXhc20hmAA
bx8EY87tf5K+9nzDsbkmoKh63LmQfWAOxYrSo96JcYfXHNLdfWhKCKd3f4StvlPo
RUYcgsrqRXgwRaTFwY+fBtxOW6W1RZnZlDMnvfaG1wDxLwGygvLOhU+99P0PdHUF
4HJtkLAIzp957WgzDQPHeJ9wR8J3PnLDkD9AdYQQB7fur440XfXPCQuZcxvYPo2e
M1ycAsopGhgNZU2qd8Bhvx3gOffBi3oxAZCCpkgGThpEF9NR04uGx2y7r5NYnpVo
FCLVPJ3Qnw9yHKJPlBuA29ruaok2gLXvDZmyYVlRvTDRWYb9oNtcD9L+yl5dzxKg
e7uXI5zqSMd+gPZP0JG0AziKKDJI9wuROcIzCvkAEnU9gaXuPJ76T+sJhlP60CSU
CN+IMJJOfibuWsyd38M3a+n6boqHtMFRjkvyzp83SOwE0QET8nHXWeVN+cLBWehH
QuZ+s7SF6Pz2Yi8aXnOgxHeAOWq7bvZ5UtjFGlGXK0000LrmlwxBlDauwrkPtyfJ
ke86ljIDVPprM3D1TwAIuP5t3LNVVy1sfUDDBAU0pg32gVJ1piF3OgNHDqDXVTMr
LA85yeNXJIttwW8FVhot8iD+cJhAfKnXMkmhMM5rPUHubbHOrpN1NhIzGZOfVIVh
151Ro4EDU3SYtTy407AXA1s5zg0IdY9qlzFM0uxHS/GCARrLfQVzZMfvgPNYsDhd
NW8rOsx0iD5PyENfGTNeaWSpdid0Tc6SlQmkWo1fRDV+FpPpGDJrUqBjwIT03ZTl
JHp4SRz8LGdperyvPf1E4s5HUeCpaHkoy3v62L6i3YsvcwB1lZ7rGXpNJ46OFz5O
UekEiDvMnDxS7sceX5btWXZ8lS0PliuxONfsWNzDG6a0aBm5kpe9a/BQ0pKnuwan
8oMLxmSEHTgJa/+fvb+S/l1lTwGNAHfTMDQ9wrZ6WPvJt2Q2kPorFeIhCgaWKTHj
npM+yerqo7MMhXSjHRh5+++tLhLvflrG0ZaKpMaN1xsNcG240A8yUYNhicPG1asR
Fk6aUQdaJ+185tAXO6hlaaLtXUSgBRLTrSjq8hChbtRQh5jCdr4kTdyIlcBtiHWK
jYXmwTQI//X4Cb6hF2r3JkaeYEyaldxBPP9yefMc7nvljzVkYxkd/Ga3YxSOmqM6
FSZVgwwHZctFBP8YUDFjQJU5NLCrPH4DqT9jSktKth2Xp6KEbZOltWl5C3acd4/a
NC8Am+tBTwrVQ9TeyY8lPDqNDiby1/5jMFYkn1TsJbLAzRqV/47jlfe9aZKARpXl
ibirqCYNqO8JqXLoy7Vew4yroolakkbGTI4Lc8kGGr4bokR/3k+0qprMcWeV5oNG
NxriTSv+rXVYg5fhkZqYK4G0i3h2j3kZa/k66crGBk6LinejLZXHwECVbKQ8wu0L
8JiD3hDqWWJvMGw7zG/iy6NKYx0ztSDLZn9gO9/fZ1wTDizUWKhgLPUvt861mHIh
d68L88EKleLx1i0SepRhroqCG9R7cE83W0JOl7tfvCyFKtjZpQG5c72h/GBgp3uT
0Q6Yd7qP5wf2d8fCeks0ikAkD4PceJDmKEQc2/yu0MnxGfn2B5czoTV8GICRm3DA
xoVvYidekHx4FTx4FU9SxKBsZ/BozRvt8UPKXzBeSMuDVipxLOySGYCnf2mquUUx
AapBMeozCDBgYlNMAGGEqb4Jzr6CUKa42CAUay6tzvtyTUYnHvgimVbzMWk1uSEv
JzZmIApFF9yLhFpLMlhiwOaMpuhtZjW3u2c3sMEHdL5hkktZgqkr7H+k7CkC/L4m
XiRd9jLPFe9YsjSHyi/YIaRZDTTqNZe7JniIODyWUA3vbqZOwHZB7cSiV1J8mbKv
3CJj01XDmF1ByErNDLUXtxdcEDKoBPEudNn56uy+ukDExcwWMO5zS0T1/eUYmgTw
dkjGOkyIkqNwporpt28/MHmVxFp3J3TbR4inkiwY1tRXOe9B+B8fAKt1crlz8UvY
8hzu/eIA4DAe5y0v9ynoQ0Vzvm2nGED24DJzbR7erm2GbKG4GGtGw2tkPfqMgpY6
iOPnKh3n435qXHRAPA6PUVYpDr1ww6niLm0j1/2zlBFsXfSi1UwgekrhPTM7dHDS
mv5b0wTtM9VAHxU3aSsXZ6fAqGeIy1fO3ufPbLNmYPbzFTLdhVPahImnKHWjwhZY
DIIwWnFsCfRv8BXDKLT4yqQSwAyGoho5Cuaq5h1BdDhyv/mEAkA0oLITY2TLuzSm
OSqzM+ijPVqym+xUi5MBYXcjHJI8JFJ0uFIuy+S8NwbEcqO4t6qR/bv/417Jaq20
fmWXwCu/QVNKbrDMWepkEPshN40cZwXfwG9eyISAnlVsWtE/DMm38a9kcrahLy3T
DwLJ1xN3iZGNctmepQBOfs/L/WXGFU/FUzKuyv+cZi+QRAIu1h8YYsEwadVzJzFF
iJLqUNJzYCQJXFv2EC8X6nOXHpWtze16a81hDto5YhbcUbyQuBhOnynHgOpzQ/oI
NfcghzNJ6mRlikFYjytkC6K95jx7kxSMLsp/nBtR1ZdIF0VSzK31Oai6irk5wDE/
SJGQYy43x1ELI2/Fk5oX5mmKznZruyWzCf999PbwHguiSnBjDtWEnls3Wpasas3G
fGvkGwPUk6gn2SKcDn9TmcSOohzlrTg4Hs9vCIzMF5tslMvOQCDzJ/Oqe8HfLOld
lNq/Broaptey7R85mUX63zVzq7PGGO/v7pMiYO8Y6WLOIwfeX75sCBEJ3jJLCnqw
1yNKYpCU24SmH3kZe8p1KG6Z6HScsXHQXe/KQWDXwJcpQ/Efz5brBtB/0B7xl9ko
kSjPOLENO1W6Q7s469GSN4gutzwzkksxlsxWd1vm14CEOw5UHfTkh6lkg77esoVy
nWmaXmMPTnnbSq5OGNTNT6QLUYyLw5xGicTQMtZJnhYhSjgHWs4wXZq6ldBUqbBR
hp58TsKU6FbI68xTLV0YsWWGOYQmVRimXfQLsF/bj4L3/wFNCGExmB+r2ufavAcQ
Ce/Q2k4+JiLWPSENczjAr5EEa0YpvSi7SdbLc8ZXb6SU9+yo44uQ5yapUgoFXpNA
vpYz3EEda7jkhsxfyJwGHUlfzvg3V6py5Ku1mlIKZHjEnTRXzvvBqQ/6xvJ8em1k
Ybwa2qsQ3banWgnXBuW16DXTQYQlGbpB5/Ty+7PmrvNqRjGnOmszdkrMQxnEXhRE
2Kt5raSVRlt5gDRnrqcUVQhTs2E/xHlqE0u9psYEPAikREYI5F0KX+JUPqVzUYbd
gZkVYsuObBASUMb3PYwEb6BwjUjweFzSbgyU64pIKP9GPdgxW6gWivJ3oi4zsoVw
Ur/jc19BD3SzdoVHDX5Ywr6twTazsgrSukTFTg1uwRL+O6dxq13lgx/n6ou41gKV
fZyoQPqE+/MD1modinbyyNLwnrNqyKz7fbymw9qNHsobuxLlJoXQcxdFYIvDlk+O
gwA6DC3U6RlYd+zFCfnyWnogarbtT9eLICm0cTtGi7WNrCNXplO8wLxVH+qxGk9V
55RM9jby5V/alNp4JEY/8Zs4Tc9BUD+nLmsLyAk+e5+SF6ejsRH1NqVOYFkDVXEF
s5qdAR0hM3oHGW97f1Z9pdjXIdIxqsMk09rDW4P7E3fhJsk/NflTS5bw8nUk2vGa
wiidjEkU+B8y+aI5bUGuubLJh0R60Y22NI0Ztid2r8IANmCSnrGouYYzTJDkjQwc
8+gyKFlufVxIhmmVfhWTzMJc//2Aa8kQPc8Zh7SuNlwI4N2bFww6d66r7ZMwf2p9
grEpbWXcOPSFs3drmRNZnrIBYBA35qT86iQ7xQJisedCejxtMUsJ/ZH6CTbIg9Ve
+7CdWzczvJgwY9FtcNXvzDmS6eSvZxSd5nkE3Q4HTIUYoGMPxkkS57R/F0Zp+BaR
BscMCTq/+/pmszS+xBfEkCZ7ObuyWhYs221tFNb4OTY0QQwFapbx4UDeog+OWEZI
rNXi9jxSGyKa7pRsAeM/i8vMMYNrzsDY5wUOHx1E19iy85YxTcAHiNBbjbr3LoBI
xXNwdKXV9dWs+eacuARUqnDLwrTOwKRoWI/XEgdoHJp5QjVqvd6hSi2A+yYq0m9I
IPIboMgdTamM9uIMaz0r1d/RO5AoGZfBCQ9+21nG8ZspPZ3vACFVJmiK7ZLOwkdO
kYeSTBmnpSc+4gp/Ji1yMwplIwvSqwfsJZqUuLm9KzP+Sgbk0IIh+kmViD+RGOGS
SvTMZ6R51y/oExhnPPj3NdIHvEYKS6l5chB1p8WwJa2m53QIous+9jg2vAEzCIdO
FpdVNBQvRTVuRsk/ArQ5/+sYdsOk7b2x090HImZXP2y7NED6O/bs+bOIIKKQ1zRi
MEIGaP3mAZEjyPuBJiG5RYuI1RxuHtDOCK7HxA/wC+42Y+JXzBemD9LzI5/capZs
fkiElwK9ueUukHQYzyt85oUi646vMEpwfKVBpo3+vumkcKlPtRynOIZztI4FimEO
6YBhHCirk2gvVsfMpnvVT8tvg+sUHOPtYqEwxqlaMXEzp0pMR22I83Dw15K/qdVk
6VsddYb3gXVscdYx+9JY7N0yp49lxgmSAZ6Hk64/xnU+fH0iGxHFefwktRQJ/ujj
YfHW8jIfbaCflgYvurz33FPJWJQrxC9bHrWHGsLuR8w4T1ej9bzB20RP6EUcp4Ja
EVXwmDffVQ9UP6Rpa9wGt54JBWOE6kXBmlZNPqcVomw+aUHLOWmcdHgW2AC12ROJ
vapIj7jSRlT3WIH2jvMOVlVhgekDQXg79XhUmZYLuWFuatvsybfsOK/L3gvDfOXM
WkYtpbl2wrnIBTOEwhd6cNNCiaRsryIJA6Cw4qI22LaFYUA27dXZIHo6pRL1PAEf
KWojIhs7g4JAcVNrK9MaQN9kFlK9GTzwgRqqk5IXwE9aaFVP61PUSmofzhzU9Ukm
K1DZESFFrvlh8GYDE82HApo6075jfMrGVn0yJ0nozopcBCkspCHHaWBT1aC6Au0L
fhHPVRoKWF5nl2nOTx/FmNn+/UHtdJg4YPcDiPt+4X/nqx4huHwTGmLfYwHIAO5r
QHNHJImEdDZFD6V+/YXBP/bsiJb+25L36yjpSf+clTRu3w0d7qnWOHzNx9i9womK
na95h20Gpnk11TM+BYfNSQtOqM9y7o0Ic2TJ1GXRuwF6ww3bBBKXtObT+EI/8YON
C1E0C0kb70M2O83ryXt5fH+aFXAE/sgES3NFAWJeSkS98LJb0T+em1olHrilxX21
XSmxdifd3FeqN5dIy2k2W+wqfeknNnZiRbJqLptq6QAomt9a+xOpy1KILu/+5JA1
VEWPCj01thpbFqbvdhdkUgpTDP/+2L6YMDu6jWq+koUqzovC8GucsI95Vlocm69h
jKHpuusJAVp8IT0Anm3ACQoWAZ+FzchB683fZ0AFfnRYsD1hqRO6XNMnZrMzL+8I
LSHJwMNOMeiexAca2uBNvOfb8CM91Qb8IuQu5LaHtFpGnnIimsIetheahxBUHyQQ
zzqxrBaDe6MaicRG3sB6r7vIy1LpS3RYdAApO7/4rJctT9wW4JXFJXcyiZENytxs
uJsk+vCm6OUbwHeHoRKIdnLOrTDCUUz2XYkf/FCKgkH3r70k2flIt2F+sUYvxFf7
9hHIYp6Xy9C9whm5gtFPvMxvXp31YJ2mvXTk30zAPsYAmoW6eUC27yRBTOlE8y/R
cYBjQKXoXQetio0sQW3IDSb0Xe/KwM5TJkBVNBiqj1I2KMUKOndgDLvRwDTI4gMp
smkAEUmiFWTJkn1aPKDg4/qPSbNrRQtQXmmEOcjXUmFUbDaUvmO5OdFEfT7lNL9K
DCFPu5EwP5BzCGLwwbQN/ouzKc7YlgB2egomRyFv+atXjoVP87oAMtx1uctESOJX
oVPIGT9xDT6KlWV0iq1IKpfvTDA6y35NbNvHpYhvxeVFC56q88MYCGaufepzAjvU
niAQSXpILuv8QNOnD9JXi7b2pIHtVCyc+VGT5uZFryNSlFGLONW2etpZ3JLARYur
tixqD4hJKTlYdtflz6a2VPLCdxW+6VxdKCSXkQGtz3WjYg4yaBoUgJi+OXl8oc8O
Qqd9Tbh0dUbHk8gXVIjlbiGHPMfIOjKHr/wxuJ20CYjzEnNWEf/R/ZxnxfTC3vNo
r5IV6du7yhhv5o7eVmKhBlvF/4iXQrJs39FUttCNSVg9GNes0oISHF52XukWVxMP
rbMZf/OzVFzqTj2VVOqWwiHB4tCguzsS/oJOB+zkdZUwl4dXFiqi/e4oRpNWu3Uk
T0EYBG2+92F/OYlOEovpTNptvJJ8w4/FMDiKqoAR7Tf2ZveuAt3Ba2qEkGz74dw5
YogevMPE/yx+p6lSWIlCp8zQ75MRQMjnqeCans+NGkw+EgOQShEDwfRHS0aEVAQs
UShkzIHXHOL4c7v+eDtVHM6ZRgHJ77NeYpGiXP4/QKMpuZD560rmJMVTBrsvyCxW
Dr6vJWwe+XKJhWggQPF5vj220x/3sPzk/ibX+ZMo8L7Sd+RF9Z3Yw1u4xpJmY1nE
B3hbUmUsPe4OfvVHEl7tOZT/ssXahBIotNwuQhGQbFb1B66SpQynEjPdYQmHxq6g
ym2njArF0D0nyUII+0BH2vfa+o8qqN4ENrp+HH/C8hvSP9mel0osTTLTLH6+o6zu
2grdnNA5Ctc8x7Bn3tpImKoA0pAUkw433jhdEQ6S41By1f7GCzpQKDmc/WzACech
/9ejy+ijdsMe0F1Y7JKZrHi2MeiuIcKvm2TOSu+NaWQNHTV90+lame5P9qBICNca
ECfnIxzZhiL5dWKjqgsnjncy8YpTLuvweWwVafsKnHF/rMpqBBeSFSqlFs0aXdxq
NtY46NJiOCoNNcqbvCAazg1Rm30TA5SB1HCvLQ0ctX4qrxGK0lMswAD/6Uu3p6Ri
KZwPPvb9Ud+yp9Zz8+hr6k+0d+qO5q6SwiqPcPg1OQlUTtDAh8aXCRzSi2wbreJE
Q2lDDcschyayuXg3WqjYcPeQ8dHFK4JMZzp+n6muSI1CQKanhh2ACR+Ucrza6XrF
nSQsJONgVrE2yBq/msfNlEP3Uyi6FwiLwRVWC84hH4Vh2R+nw/qvQKHFkvdFX/b6
XunK3N+plozaBUSRBeHEo1S5AQfOj1Zlr4Lg9NLiUcRBX25r/jmOn0jC6LcirqvG
92TTWIjgi+5u8dGu/OYE6eQIUwfZA90TM2MheqJrRMbbQE9/ChGv4P3xJA34hf9C
gNnKAzwV2F5QhrslokXZBuZy8aJz8HFIs0gh4lDhAemdHEuawiXdRiyR9eDC8BgP
dPNXISZkrvQAZWxFrS//gUj9HJZc6Z1ZD3KNxIj8bnHnHgxW+PzLn1jnJv6+SnUq
/TCPatu9mYnOT+I6Ibc3CbqB3Cw/YjNta5QEtN6IoMPTQFB6OQFtwGgxW4u74fKM
2nnoxX6UammczR7fZS7s6rs6Dm4iVTEltFtnSafDid5zSSEoPsTnDFeJmdJs0nGN
XOycbc0eYGRK6kdVXZaZcRppcQoDTEzKIBMujBTm7r4JljyYfWDwz/VJzzd2RoJa
+qIpb6nipliNWIV52sNhFk2Y7S19MVirvvwHNpQr+5mXUuL01BeZIpmsJSqNaK2w
gnKlyMFNfMWgVJ4jFNLUiSiHKRomcVlMHHXb/ciBtPZkiF24zFhs7JTym/SiETu3
eAsKL3Q5kmZ+zQ83OqWLInNv39WmYnMq/h9S/uXPpwIBluJWP2L7uz1joiDzJMWQ
ggwU24ECwgJlTzdGX3kdKfOBZ/ZKkPDQX5eo7ETBvjJLPQot9nUAdgmqGmhqxPnJ
ALdm/yxnFIRS5/AdIWUlR0hrhWSeXV04q3NXd5gVREzkykMB/LeuqG6bfOc08KWw
KGBAmTMGLTlsUznsq5FStpxrazeKvnl/ZdfxNoUjvni+AWETRITDgrRRFjebEAMt
z7YjbpdpiHnBKwyPiJqIJ5kY6c0EfCW92SyXd/qSPL0+6JOibyedjREIFF09Z1Qd
5ChTU8qXLCM6Yw+1B3dQH791KE9/2bJb37iLCveLEckeGHkMyfyKZH/E0HvlKyyD
ivhmtluengbOQiALl3aSxGOliriK5szGN2Hr6EWgHbkn9aCrCYFRtTmOrXtG+cWq
Fj96ZQkrnDBTp4FxyEK6Gnk8tWxpHdgC/lzsvzLD2F5P5aHmFce5Y3q0xNj/Nv/h
ZdboTBJAuIyGFIO0BOl4gSVVpcX/DNjnoaczFluADRCa7jDWu4LY65/DTZKq2vrA
uWOuB3ebqN2rEKpWhh8b1i/ftfU8GvwO36/gmRDnlw/ISmDTlpljUfrlU7MVtQ2g
VKkQPmjKai8MyvLymE4qHErzs6jjN53SywToWpZEHmzKsrc1eOd8gjktZuVRYLfz
DXF8H5fo8pHXBbfdSikC04Vv5FrPQSLDigOZ2IsG9hvSvzdykUrPCwV/Hm6xOcgY
JvsutTh07BLxBVgEeENtFR4Ii0DSPMzDILnp8+M2NIocO4hYPywjvFO3XRi8PmrG
mzeWwaFzsse/Yy+OKDmqLGr5QcKv0WvYPkOq7+RQMPt/qWA3gd6Ji8rG8r60xhvu
yk4i21ZES/B6Le9vzqSFFvKnujliP1vtCgbVd+QKhO8K2RVrONwmBvhS1sLg+POU
RcjXuEoUY/CTM+YkwF8ly2fyqm2xxf/OyecbhqfJMgSdT8imxmkF67RC9yv/orR+
CSpX+pQW4hwNUlzEtAHwF7iknV+Mf4A5MjNeDHA8HpZ8nxlm+7lxrcALCBhSxny1
0fvwePkvrfCB0jJPbcGKSm4wi2e2M+3tkQYrh+7hJ40ogJsyzs4RL6SUjOPIxdhI
aiz80kpV7xpP2/99lHp6Hxgve3jt0m5/B9KQ8HKGRIrN2NYpoBj6sTClESGZyzbG
tgyplr55KKw+nHcBJSSqMjk0MgcwJuqraLAyqYN1zKCspAQ7HIrxSapVO3MXKmXj
Jio3/i+ut72qjeCPVg4p6HBGMkJlU3/2f+vV4zR12+YK7WJK4BWQNlYJ8h0/UBZ/
Af4wdZDHGt2DTr5CK1wee0QeRdy15aj/mY65WLfRCeLuUKLTjzeKeOIDCQw5V46R
3o+39bfLqFXPLRHhtWtPcDzVjADsN7O871cisurb2C2mmu7QDY1c+z/VB8QMVr3k
4t9xil3BvxiMMq8ukz+P075BJjnG/ycVUm4L+QkiYl5a1+wFfElWe+pk4xXD35hx
bI5j4S9NFypi08SAKKc7WDBYxUuK0g+N5nqTaOcHMN9bhKeAfJhQVSGub/Ll8bnx
2Zhy3Pfrt5Eku5rwTZqGw/9Mxyt+TgJIp4llH1PbGJ1sZa0tsAzVyDnHgmLXKjZn
xUkEpEIhCI59ylDFrr5T15BTWeiVAHByiDt8RoK+pgNyxZf4iLj4Qr75RsFH/bcu
HPfb+tFZm1hS2o19F32VRCtae2FEjh78C3E95fm9yOtX9+LTrPY+SmKdYzUwmzoj
uLSfNofHkRQfnoxpbxSgSBOl5hvd06SC5cmvm5s1pX64W14Mfhz306zFddeGjMvo
VU/iOMqpFLBdtdMrj9W6OVOeCDN0IUhqoNa1DVbkcINCaK1zGJg5DxF6qQ5NmHlA
4PYkzd2yC2EPk5C7SRs5dV7Nift+bFZ151kWC1Edzncg+OsDSY2HXo1hcM2D9L7m
XcTY707vZVnoYgM7DJ+EZPC57i3i0TpvGrsHxYTw9yxSaK7+xoiIG1ri8UJtF1Tx
uDR571xSvDFg4uH64OuqrqkxepvDozzCRUkDvo3WDLPPluTdmXmKBXPnxmHd76g1
m6EnP5qL9JM+fWv8q/y099cXH/HXWM4WKgavKEd6wsOyACDNer87PekNX5ff3hKJ
y2vy0PmOOQ13evuoHOk0bez8IlPcszhoTmO/sh5q5tuDp3QuihvJnIljjsXZJRfL
h8q1dhSLZ6FiBzoHKNvvcB7HYYy+PVEiA6+B5I/j2vQfXsR0lAyI8sUNxZuXWLQ1
3vC9kg2WrMdDLQz69agihORaGPtQ7Wsf7GazTHRYWsR5SzxzeDLvLH+W/7llJWhV
gE+iZT0sLWKfMyWLBbj0/VU8IwjfA2p9lq4dkTRkxc6zFVmyihFmdYLnZ9ZQuDDN
V7IIj16BqqQPZeJIbFRPBZDRAsnaZlJaMMWLoBNXD/AgistBoVLLLNktSVzPwFQi
p4oc+MpY3PlE5O3SvDbMGRpWT7Hag4IxLGf/GYqbmSXyJKdHr9JfqL/qcVA8XYSg
U8HngWxJEfHgXcdhiv5Gf0cXrmg/te1yVISSXFQ/PwweBGehYp+aeR/NrQEzQeEy
2Mgs1Q8prQdlhuMIeoy0Ftsz6yuq95wgfNrvTImoMVWU/4+sykNShOA7uEyzi6iD
MspyJW7/GaWs0owZGLoPRT8Zpxr6gPsMiVXi4n+N3LijNFFb/wf4WY3HqJVeLS9T
HNbh6EsiVUdz0ygUdtPco+7IKyB2EqBRjI4G6UnnKuS5dVi/3iYU3t7lBkk/kAVs
rL6JZRSM08XKwp0XrOhMcKzPvsHgAUqHkaxoxM78EI7WHz56DGj+4rLitdR9K9Ho
tbXAFQ5ATnCmZOgUnzK6SW7Ir/1HOY/O8KiQ76cKVqgFtDdbqwrF0Zh2s+4sTZUx
Ny7hZTscpkwdHqBnNMEDYkjImd87b/T1WNKhKxu4JtknxIkqDQmw/nFIbTpbuWKW
UN+uba5ww//ExUvpqWP/C4WLq5CKe8nzoVn1i57N9x/Fo6O/c7TwRvdLgS6DxjaR
eoKPHjM9yQVXgU9vFTkAxxytkkAHGgRjr7Ug/Ywd3eHtiJa6lG/2ZzEzsbZRyhIz
pXxupgLJIFDzRlPEfuA4UlTnTEVM7//hUePkuzXjxjvWjbvktHss2UpJ9ceVWtG6
ZKp77Fuj2IlEEwL9cX+Efif7VeRcFhi1MAT1YPdK0BwksgEO5EaLBNZnq5r2R1Xv
wuqzFK7yAJqKAvMRAZ15zHE0mMS4VUXHC6SJ8VuWSD0g0a5SPLUk3ZvsU7+ixiwO
UBAD72Q2HavOUdyCEzY1JmDeASNbiW182u153dGrgV1xcv7DGPm1IZSAVbioV+0i
1daBWfHBelZbliUYkIP1W65ZyX3qwV/M/fYvQboEn+SmIH0JfeqWS8BgwNjJYGpK
EZCORVyZ1a7iDNx+focMcLgKuPHcwyHaErFj498JKr83Oh4EDom5OEyIjaKfFh33
Cw7zeWTjAj7Wrxmn+irOr41dWk9aKicNU0TNkTxcafJ+VJIe5MaUkNT9EpJ8Vf5b
m4n+809DlTODTcHQ7loAM+XmkVJEr5e/bLWKhNQtO6sbWE0E4hWkNvx7+iOSuse3
lViU+LpMMWmjB9c+GoODXqKWtOqI0vHTgyESzkSYRFjfvQfvdvfPQG48wE5cYk11
OmY1ELcZ4xwziP/eM17WVdr4K8ZPU9Ew2+QTfemfd5sCmROUSeWEBeGrBqPzHNXv
ScoKX3Xjg8IxdJjjhkNEqnv0qJKqGmdtai5SkPww5kmTIr/Y93p2YMmg0xRQl/Ax
q434N/kywHPsIo98t1mOhfKu0GGeh8cNJfc+1hdDz5R/AK6UXhopogSPPvLdln0T
kcTbbb5dYMgmMFqUib+xW91qVFlIuZ2UN3yu8RHMhhQKF6yf6ReCv/lJ9jXw7ezE
FXandbst9K2wW1o5IzLiJFQ+Z5Ew5K5x9A9W3EDfEgwejDWT24WzBwUXt+ygn4ml
ziw/SfgVjAKWlJ39p8EnK6PjtbWTYKQBLtVR/tgRsogW/KfyVZVNKTTkYWQUaYZF
ilSLW+S6TYZdCV7TSKD4YVMU9OaqMNqeDCTlQpJfFFnwoLQ2nS6ioC0NotRfegWf
6XAPM9KKiXtQQigKPXEOnVWSsdDd858cTW7Jo0qTX+K7BGI3b5rVmKOTPbBiWjI6
GeZGB7Ji+D+XFAKWUPCq7eON7aRW8DvamiJEU/PvlZ9gTXM4MTyDbz4oBecoNaHL
+ARSC6203OlBSRn2NBf4mA1+zaxYomK0se61OYCIkflIdMHCvNiQiUi2ccxzO4rg
T0fglz17cCWNJR1ZgGdug7ak8cAoC5NL5uFW6kYmzKg5Tm/9K5CR219IcgELIlkt
tRXvA4u1EnWP+jzy9I3xnPAGX0b+zfIOzl0rWH+NEmP0ranfWkeUq6xTLltaLXS6
QltHa0xctABl+V8dQPINei9hTkNEI7Js86dRV3f2fNRJtRc0GW4BfAspPUwqF1s0
tFYqRef2QPq5M7gvqGABLOV9alZckgnMyNRYu2tD2oG79gia1tWdJfLd/7BTHq3g
GazexsJlOf7etoDXNK2LBrfeapdIzzsmvOrQouyE4L99RzoRBBC8RtCsvwINY6gb
5Ica/iAMzyCGomcC/QR3Ln9nwcmlU8pqfpw9jQwU6VeorCNhBG9ijZgIIG5HiY2U
wlBb03t472NGVhAwrnQD5uuedNrvvEkp6aM7Rn2GS8I7lhaFTYnwPkipGAr8pAtG
zhLAq0ExIP9GUmP1qCSMPDiGiIANncUat/DRGF9+wLNABIY/gBVGkowow7Lm3V25
q6khH621zoWmMqyf5j5bFyGQCAjGODm4mFWaXmIGfpBD6HoSBeyDl+lm5w3eSYwF
3EVHD1mEc3YhPkNBd1/Ec6QBUBoIXtryWRwfglTewXZoqRz7kDKYKMilsY1hgO0H
n/EnwVwt6ItDuoCxl8+Mir4Tpi+McXvKbmpe+AKp+2C28gfx/vib0ojbbE7ckK0q
zhw+RPBNljc+CCXA4QemD/AN6QqyfjC2SIDoh3P7i6MxIycC3CS7fq0AygHwcd9Q
Z9DFn0Z2MfS5HSSP5Ilhs9SxLZUos1J9jArOfVtTXZhj3Az9ImygxKvCRfiEYi4c
QiyCaiEstq3oQPzFasgg6UySuLA+D/wZAfn4v6J17LoLwOSFYT/LoWSIHPqk56SQ
s//cI/6FVUbczH0MPXae9/0HW3fTI/N6s+5zzea+gGPv5mLQCupqwV2GYjioPPyo
I5tujox7MIFy3mdEeJgBGeX6qIc/R65uiY6CcfoOXeNhHq9/ItQBk+7bEOg2eifV
JEWxbF3nfh/c3bagVnxetP0BoKZ1WsQStIpIWzVf4FPmMf/vbk4TR4yIxbYXSV7m
ECPXFRoMVH4vLRN4TlnnxQ9LM66TBBWe3cYy+TdFOqK5NyRdJ+uduQWM8WxkKH5N
2ZYlTsfFf2maMxsBLsPpEPh7c+xv7j5y2Z0zFGBV5v4kAB6bOiIfWJwh+swQUz7E
sGhH1WNc6DgNnrBKD1ge/rMsUq402cvdKb6BholWxEUWEDgcLECcdgekHqVdUlAq
JCNlhnXFqzROP2D8J03EeFF7V3dFhoXXHPpnXiT0xFecgbL0MJVch5Gu4Tfvc/Gg
9w3p+T1CJ9Aclt1OFrvLIlQa1qIP3cJ0uvc2dyDMIO/EPUQ3TPwzdXp4MBpKR9Lu
+FZR1FnyMXUdULygTiDRfKUszh8H3toTWHI8TZuKC+2kNyRSQdxGCmRzbcmmMYV9
ijD5kNxwdlvwDRxvQyK47g89LWvpMai2T9XIiXnWmawootG9ioXRYy1k+UJud4rQ
MNEpGhLGCQYb8lgCMMNscxAuGGHniEK5TTgbtV8dTTooGrAX45qjtR+gbZ3xCAI/
fuyFsDub9ykMAIa939lZqvCL9I9ZTF9al2kYn8wIyABr7jXwM74oZiGJ0rO2EMrG
UYxBePf+7E29tm3BOvfdmaeCTv5rsf3C6UqiGRHeZPdCbKm8NR/3fmLrTa+Hf7oX
rvRKYaGvXpgNqJnh4JvXIoGO5vshHQEJrqdXdGSPlBtdB6B3xL/rrXJ6WpibtXdv
X3y4FqEt3XTouM2yonGlJQiXhA1BbU5VCgxJ6xwOYW447eV+h25LuKj0Xz7MSPRw
AJNxC59M4kFj7R+YQObJ6vW5YV/Z21o4pxaOTlnu97TCaVhVB1iWhOCVti231Kt7
AG4w/z8QRLdqv+5KwiaFJGpEdF9AuDQ7desIc1nCdDIJbyX+EiZ20LC/a4KRwugO
DmckdofyrBmJLiytQiKvWkVlo7rMcYr3+rBDaqtHL0MXtBK7+WMqpumRrsf9Ag6G
t16ixAP0mVMTR2ewD4X+SOeSQH5yFM3UkNdPNu4GMfR2rg6+fAaG9CEgAuEEdcg+
SOK3NsJFiLGWXaM2ypuHcResbYAAuKU1IAaOzE8+Ta8hSC43l67LtHrg2VmD5Y3L
AIfi7+ZNFTcB4zwVRTWfPfRP4BnBOFAPEeDoIQYRBEJbZg3D3QcyuREcgGwIz/W1
OIqHTLcIZGET8haRnaHqvPNmi9FDmYllQW2Jc3w9EOuB2h3O1f1T4/l+Gpf/SzSK
LfEdOqYkfBs5utaLGqCjPx2t+us0tG5Zypts11tXoy2ofKD3iSFS93KA/Dv+xxY/
VvpFreVw1ILdeYzOA+W4ydBwSg3TCxyB1eKpAI8ALpFgwytD7QzRPrxfdcs9SeXd
BsrekU4WJ1+ODaRyT3jbuLk+AK+potmJ0q7ljiO84R0zSMZEPiWqBaqoY8AlPpYZ
kLUNkfybuFTJ9y8gK3f30mXYjzua52UgLxkP6cFZbedorKiG5/FwjtS1bL3iQ+sY
1UJEMgRKONQoZVhACmgAuR7UHSeenBvd0cJgsoTQPyCoiqbrhzXEqbqJxGuUbPu1
K3GQk2KiLDR//pneQus4tCnTSTweBsJGfYGKyHRS5yl9tlbaRGcr5njffV0yKtJe
e/7V0dVaObhBoRc8r5DQv8DM7QUISMMFhbF3a2nq4MerE1w9YdE8cGAvFjzBTWiJ
LGtLb4IZu8fYDPYYYLbVUlfcEdNHO5I4VoBHA8jStDWvGmCapHMrBk8XM+YvK5oZ
R6G0XwO6EWxJQvtlDghifFtdXWDVDR4JQuqcsgO1OmZRs55/KyupI+6IeuXMM4VA
7iTDtR33w7D7vKYs42YBLfpOTX6eOtFbw0mnk4j5QGu+JvCh4qeLOnm4Q+e9U9Z0
XdQlMr9rhV8brHO9mqodEaDcYj74iWCGX9eoIYoHDiLlsnYxtWrF9Zw165eioFDc
QXQOtckFIf+x8kmOFfOHxBEflRT2luz6TjwI/hIh2JeHl227wzkLlRGYOTUGOEjy
3e3m1KaDD5g/pysY6CyEwWopLbUTGJar+3CL5az3213BWHufYt1xn0e4zl6tGT+y
JMLlCcYsEIu5tCRQWDbVsBTZO52IYINaEkNYRR15BJ/nQx63kZ7acdMd/cyaQ99D
o+tM5kUUKqbqgJgKdP9T255UZKOBDauG51ufOsEgImoUKxwEDDuFrNKKOciEi8Ld
5OTehIrXyOhziPzIXraMI3Ldz5Ww+Vn4pvusZ27zj0UqQL8tyyH89WFGZMYpdpsR
xt73xGrQqYIBjKEmEJnfTPGSz0m3IJsOFTy6TNAB6L3vcO3I/TgKtW1bdFxZTSrV
kNPSjPWTuTiNzWPHJrJi+m+gU17AO0+djzr5B4bbCapLHmpI9ryhxaEQLipM5GIe
3+BpMC37LsSJwUa4ZvRrNHE2hQDcYAj91l7Pvjz34Xldp7oal/Z/uK1eKtPaqUqK
gr52H6qOyUaCihwaBhZS/APGHCnjhEC76eapgNahsZQstv8RbCZudqhUss/Z5d6s
ybGskLOmSFPdBK+ht3jW23tH8EyxPE4z/I/FDKwLUdy4WF/JRRJvjxrnxwiD3f+H
GufCb4Dbx1elnkHmQ4TLo11KQAEMULaq94Dzb71HVrRQyva3w4r9oyiTyAfdFo4u
e/+PfL/rmjpQZ4XQdUvk0e0iFHTOeGkyEPToS2qEQUfLomcTqbXF70PQJGVHnrb2
fCm+4gGMZE7e34fIidP9ZMy9zyAfPAOmAuXft9/rMbM2QKboNgAH+H/cNIrbEXUP
UQ7HhPZNTLOu35STEOM8VXZE6+SQtJ/1I1yWeyV0QzZ232h5BLp5aCUHat9tacvg
6FEnTR30pbHSFu4LF6F6idPbPbtqUoP6yLpZt41m65nPPWHKa3oXSDowpuVSxS7P
ovD5CaDKl3x2t1VMTPj2U2GXE9tZp7BRG6zwsbwWjMWMLk2JWtaR0Ckqu7vpLcNw
+PE95BbCE2QHrLS54QD4uC/Agf6mA8MK/XSTA30XaaSKuIhJE5Grex6BymJ9c1ri
MQ8jjP5OGWMaEHRnQ1k0i0ZSH6VVFKxT1aje/1A6Sv2jwyfV/PGzi0WQT8SLoWIT
RJEXJTBahuC73RPEUzJlPNL3GvnS6ma0jtiIb91ay559U8B4J7jxgYDUMklsoQEe
+CLPM/2bxfm6589EpX9rMsmB7p0GH+TDBXqgTT3WaVvrm9Bar9kixn5y67E0Z/OO
gbB7U3DbvGhOMmeR2C5GJU9+/apwlLIikY/ismL9YdVNOfEZX5l7wb3C9VklQW+V
jnJQ7shmJgL4r3kAGy4G4JSlZ+gpirWURlZfN0o8YQc1nD/I5ZGWxyBt/yTg9HU0
BQA67XMyIW+n5PvlhFx7dqKnHozoLxWo2IxHULjgJET1QupcFrExytlsNZ2wu6NU
ZjR0tYNMTGY1gj4w2poj3P4A7d0JD6gHRuUIncNSeUqfAD+FwnGwo69ezx/cVMTg
7xaxQGta3lJwM9yi4WU/LaP531qG/JUODCbVhcP1j3GMpIeKPR2BL5HD6kiPyy5/
4jRCct5QNl8ibxBUttzcBrYEMryhIWWcSnHAbJskHhZaeWhBZbKh833mQHd7hrMA
AZeGkF4NJ0EVWBSv5LvlcPrA7Sdj3vVy1fdTswOyeaos9V1Rt7j3AvIhVOpKqt4X
nzmLrDfknn+sdY8pAOwtorA/WI8OiMGSKJ4YRjvzpy/2IWUm8gY3UU4OwioyhbRH
rOi2Xb2PhUQZbSzUIq9ZN22UYgkB0tAQR1NVJKQNi2gUjCDxWYN+MI6caYrgATC7
eR/NDoddb0QJ3Inzw/RSU5jkw/xdWUjVj0BF//QjNM4CL2ZoQayYZBIQtKjUf1o2
phv2hd3hymlncipb/YQJy91jEYNs87Qa3eLAo6DwqhrS2QY9lT0EtZunrpeXtNx8
onp5AOvmSQNbMy4KxqWuNTP2umHh5gbKdTIGG6fhrBxR1NiTUPpog4e+xSN3AKvn
Ek0rfJAOv/4+jyTa6zcVBdGyW9h3a8kDnD5M1Gk5HLDfx0Wr1pEpxsk86mHdX7pC
3Jqwj0GGMs0uZgHhhsVqLADJp4HenhGwqS027yfA5UOQ/Ei+yrAdISCJlbZTapsN
rmkuorFjCFpZ66GdqiulAGE4uUJ69/EsMoUDIBYcS4qV6Vu8kXxpBS7+TY4lWP3I
bJ9zN/tw9oUDlb0rAAOdiANBohaCI/Ddn+NropdXboLZAJz75Kt42qcZXPmhKkEE
sdbFd+A7p3dYQvzq4mM1h9KzByQCQwjbI0KggTYj7yKP6AskwLH0rvI0u18yysW0
zHn45W/rRotKMK7s5kKqE8MfqnORAfLPuVAGGLW94sGZpmNpjbglJP1nRQtJkK2l
2WlNivn0eUoaFrhElbluk88fEXpL6J9oDJjg70dDP6QmHbM4kZE0QQ8z/WGD2JL+
++wQPluTtPDg/xZHsdFcDvKQbNe6KiOXJXKfY69J6gVZRtwl+Em2X+gIjFuuGhW0
h6MGXUrKfaXcle8d4Zd6NXG48vlVDnY0BkahrArRh2dcSraF0U1iIFtCNjvXm7zn
agTpxscPBUA5/+YnsMlFcMUnP771QPtYT7MNCqDkdSPnEvAPMHg4FgLyrp+1CHb9
P2soFVbLMU4RwJvTL9LjAxada1rXO9juCfvGNDsZ+vsgvwriGv35ua+09zO+wmZG
QkjlhdBjgdP9zw3Ic3xrofGT4VMgIhm6xDs4/0k5zN6eXhogxC4hqDnB1ezfatIC
pMuRuQ831Sr8XWvf/57+L83vbkJA3TNG1EzbOPZdqBAVLG2rEpadZ+Tnm93SZO9Z
WMiRlQHcoef63PrfRZmkRarW3qb+w44gFDzFa7qiq1oKLWAuroXHPxJB2XIF2b8l
E58boZts2iFK78lfiQBc4EzW+XNAdBLoqjqiI+7V8H+DpfNBHItdfijCmgbgWro+
Mcf0daVLEUUVwsNjtWg0WYAbhq2kqvYeoH1t1CINfIc41GVz76y/yopOdtwmMhSH
c+WQ7lHuYhra2ohkW8RbToKuNcuGiubgOvxM+a2REKwgXFml83d0hGnSPRj64Aw4
6H71vf8/jo3DwBdMDI8VaNl44uded1nf2wvNHm9zGEgUr3Ewwj1bEYxuYIM2Kll9
8Dyip9n4SpsTdXfKryK9n+wGQEHMoVwbp5JJ8XCqtxG3zSzF18Nhn45BH+o2Vfbm
wXegogOsciyMPwduA2eZvnxzyUctSu47QDaPSxOs6UUUITCed5D43fRaLUXPoQAy
bF9HtqAJi7cTaMd3q4wVyEmEHAkBpufFNV+fmlA2UwRdC3m1in8WOBUdfKWoE/nC
FNb44HHmtqXd8zQerNSA4BASntWPNnk7wQPZhd1jEX6gKE6hR2L/q8n8OWZqp09p
JNfcDaJQBvWHFxZEMi9xbuCKC/tUJ60NENk8dEw3KoA3SVynjS1ARU+hyCw46BhK
BFfG8fOWcIlO3D7Ou2tevBXQwOEhkPTCpKnEHtIA+DZ+t/Jw+2JZmKReo/g3MDmO
ZE4n+pXl4a8kOmMGA9sPC8BjX7yKL9Zbli666jWhQo5aTPGZH0SHw52jUvKl8gSa
DDhL3FEtvWrFEzKOybdiWYnS/+gBiFp7+2CzsF9Fa8ihcS5SKpSvcHtawAiFGjhi
ViEHkQcZ+DsGMF7X4YePj55Yym9jFRnmrktbi8/ANr8M+gUBRSyQ+j1+YXpCnBmZ
Sw696ezS/WszClQsnC4nUBqKslFA+bu8WCKqpmSZUDwpm+IfO3W72a5lV+WLhOK5
Aj8VIzNhmwV9QPZCeyXVahYiV+4nDqtYyZ/vDIlnFmRlvHkxD6l79Vvrdy8MXnw0
rcEgrvi/ASEbT7hUQ9khrTY6YrXZzLFL8d1G1reU/L/qxcADjBXjqpYpZ7w15ciZ
vHkauzVkM/xgZrpeeu2R0484+UrEDbno8GmTXJMbHilgYd8wP1w4cMN+phTA+pq+
cYVPo1Trz3sugfu1Tv0qKLXTw3bGWzlSzjp33FREGzfJAZ4Ke4tAVUeL9K0rYHDH
WOgs3T6LxoeUhm3pALsRIsVK6c/4eAm2WdqfyrKYnJxArdEjwGsV6tXqsHayCjMG
GqLPzA75OUmUbB9nAEaNqFjgMJSMHVHx7nT3+HCUTKdUU+8BHXOS5/w9MAcWdd/Y
x8hFnGSUPKcUjrWHfhWxya/8inktzhRlz0sT2V45dib7RLmvEI3b/wko3tcGogFy
7GI9Q9pbEJky749D9FTPQ1iXKBzeloAa0SLfOTjzZDqjzMzD7blThIlsnJcLG8r0
t1RTvg5ArCQ047I9c3UJ/XLjaVeYOjyKFcUXJTnmXZlXIUGVStphA+qZhuDltrAH
QUMBiEsmLU/SEoY1YM9NZFCRJI6X81z5rU60EZsxngqi++t+jy18ASFm6JGNVzkT
5/MJRte9D9bFHxlostz+2WOYVOVy/V8NUxLte/SsYH7UjxJr7VIY5VmABE6ojJlM
GzjEg0ukBmI61z7CtQ7Njl7WWZbpDZfLvv1WLiqK70MTA2Pr3XnJfjjCPs/mniKu
H0ldHAX/mjGQdTwTa31maXMeMDBfZ2W2O1/DfXobm6dHF0aBTY+p2sUGGPLZQd2E
CJ061XqFOxhrCv7QjpBeKBCafhYTph5y4FUB0wrNkaGPHZuzzjeHnstLmWt5F7xG
NbwTL3zE0kmjbcAq/ThauqG4a6i67gsJ9Y1XIsfqhnj9iDOUcHhb9Y2vtfK97+h9
+FisQxiIJwJ3SAjllsk5b645Ea5DUYywCH5DdFljpyuzLgxjayFNQRIsM9uYhwDp
Vg2klk9TbhoP73uy5Cebo7isil6Makq9EXGQ7I2n6ZL3u1zPcUM6VVbuL1AkasJT
oWO2WiZpZK2uM14q1AzaqaR7MZq+IsgIfYS5iFjso2CBI8LRkesaAOTL33jiqElT
+8Fn5p+/UE47tbnMydHUYoUSSYkeNy8EEMvvi7IaJK95Vt+ah0x6jZWpwCqENz8G
cHax3jotzrFzsfccIhJTeuqPQh1poLbFvEy+8OzV3V4Zz/Z7+W2JByYBIB+ldori
tF0F/A8WqaB0BZ4/Evr6Q5S/QfUUgR96ofZzESNF6M1lKUBB66JHI+bc/Af+RiMm
mEyOszBluC8r0KRR/CVVYOYhStvJyTLILnq95gaflm6ep9v16OxSLxwgQcUxtlE9
/y2PtUcSSEawI+nH8i4KQFhy4KnMZRqaEIA6Axatm7Hl37ppk7am7lD2D8nrRnHz
dfM4LHuXnCFM1A8/jOPZG5nmWM+S1ze1W8fCUa8NmtgGWi8qRg+lmiJOaMbLhRhh
nTYi01ILO5933t+zRfB1QBhRyR/zdCRathx8L8jvRgBiclidhydGxvhCSyVvQ3Fm
OSrbcrl6WMLQ/T5ZSUoq76bmoA6u4Wrr4gLoZtwNtYORU2JnfVryZqZHF0t63H5k
3vZPCjZib9LI2dB1jL2LK9NuZbbG/bAjEm3IMEnCdhHb6msaBfFoUGz6Zmwj5tI+
06tPxLg/R68dPvYVpufMDiSyrxAt2OZTQOEz+TKoQEnrBaaO1iET6fXqU/pL3Xv2
kWyfa5Inqp1tDBguWr1yLWOoXAvTUyF84OdRUETIQKssiTL/pT0P5AHjxdoLvKXx
/ta+2mA16a0p66GwP8HTM0rw6kDRxx5jMOoxzMOo/NWn3WxwVsBD8X+M1TfGvmSq
YkF/g1skHYIP6vgHSfYwp+T65uO1Lc8b81itKAlvEyy65Din9UCXWP0cDKS8Gf9W
1PPqQtnNUwc4fPsiUI6IobFDfusA1/0Oc/LQUe3xLPWW/fUwT1iaw/ozFu1kqWCS
YOJV7GfDPVOaNMmsmBFDCodbnzOet7aM/2NfYx3xN+x8tVXPnMnvG+mTvjGgrPnM
/BxVpXCy+YrBG9QeOzR5dBgcVsdZMXgjT0rYisWd/yO13bXgoSOgRr9yBEE7MI+T
CjDSHRo9VVdp5YHuuRilSVFKSNXvzjA67wEnz7LrDNJT8qBysCn+t0zfp/nShqX7
b67QZWTTMwMgPgw9xrGoaJP4Ys8rzE0xCw/SfO+wTwAOFDYdXis9nprECPsfBN7l
XzAENtDobe5Sjb64T+9OVEIjuQdlwgRzVnlBqLlK+PzE4u1XK3nnsRWHoiKkdenC
Pwxi0QXyGn81KO/lhstp6+Z0lXBm7qnKh+hm6S4EJUjquCCx1ZhL49I+LYr7DVIA
8f0tkavfFI078RyMsj94hS1ob61E1dqsqqnBYRP7zbkJrzGOvk1jCh0HxBRqh8z7
qTlX2PthKh2oMw0QHZvI2MTmQ0cpRFBkVzNl3DfNtBunufueHBkrXmSijyE7XNHN
8MdORjuD+oi55lzzfXM5eMh32+3kDxeR3QHuMBT945ZZa/LJkcsrWENwvzAgITYs
foKjqTuAW2Ha5znJREXQWZEffKGASGClZen/oJVNDuT8Vb6O2GHu4W22YD/STA7h
toN6U2pPhMIJbqtFlX4t088gqcnn1xXBrIn6fhPpx/9gj+zvuwupqXEVPXayi5Us
jh0BP6CARTyI9Z/U1hNqwJmgbFsVpxBiTSvIywYDMANg/4iFiuF5uZJ2nhln/1M1
62grwRZ/+j0A60eiIRD9g8jz9tL4EKxc9lRb5wQrOIf1M3JGm6pMIQzPnCK11OcG
KXQHDcwCxI/L5NPJNWBsQEME9o6OMBP6AihS9wje4R3sRI9KuTpYAhKmiA+cCfZr
/2mb170wa6b9CyM6nmwmj+JxcQVgVFvSDJWsMd2rgaZpjfCkg6rqGBZvb/Rn7X8T
174FJrwiQIchlrRoHoFDA3dvWuIbbNv7fX/rh7hxfkoH6+jyABgsT3JAmLypbrxJ
zW1w6HyghrfAt52hhWC9ZFSCm0ArsJq9PXb75EbFQVe0eyKfMUMCZRUDsz8wox27
vzlVxWU83BvKuvAcgX3YUvcX1JV24563AR5lINEuQ+rzzcVU254ivZB53Jnium3V
6/E8eDO/iJPLL6sgk3PZg5FPljmCG91bp6SCqb1iexBjz9pn+L1XrXkkxBAYjKfY
PAvI1p4E9o4W3pjQ9tgjHc7nzEYD2W9YAz/JTD6dGJrg7Du4c4tgPpUXhVy0G/Av
hSMuXDT5aw8FPsDxpF/neTtle1FAh70uMXWBcwutHt38Ep3SlP+rU3uU95hhtskm
+mu3Odxe8DQ6rl+4BW1m5y3uZcqsTaBgxNE1ChMxpbatmJpPHd7soLuXpIC8yNPE
6SVtzOdLF9wbM9oVOTDhMBJ3fax4COtav5kvnI3aOmtW06o1A6zDkOO5c4cLO6vy
nfKVkXoabhUmsxUM9kLcxfC9V4AYeHSW2gJjNkVTrj8zxndF9Dets3q8wFuB7y+F
He1dMo1ePnEvKvrxOx+DEtUcqnw16l4kHZ/f8Ws3ZOVj25DxwQ7cHFZGEibNQ7DM
iaOUmqjs7T6hjBgeeyZVbxaTyH5I/K/vUkBBvPyAL1gISc01/B/2fscHKFOpxJUi
xqED5eVnLzn1aNYVwvjVqsav3eY4a4+CB1L8/s2c0QKsz+HKF/1XUV7eGMFMDFTL
DvUt9cZdLTT+8aNQCESgn7ghIagIEhJklL2CtPiJCM6LB4YeGA4d3TqGxBxIl9LD
18dJqq6jRuWo9JqAtMMHxcHF67De/buS+wpB+c2zeGj9Zc9Wr67CEhCLdW43IZH9
7zT9S0WmMyzQIGKtKK1S5rdge/bMaL58aVICoZ4qzrVBlmr2UFkatmscCwTpA/a9
s04gJOZLxbhF0xVG4svp6xiteO3+UTxXxu47iKu8oKvvjOtg0l124qObRglH5bZt
j7HgSp7avI51BRycyAL8qE70EWPaT+5/ULPvjl70b97gbeML7GgWScY3iPe4/yKG
LioKIMkG+VK4BOaoqb6steNTiEcfQOQUctcatchMR2O5SBECI0Tk3zKFnzRgKi34
nHhnXpmDCzN62Oumz0YLc7Soyt+fvIqyL2J7vibqvUaSRZYHMg8vwDQnfQzUUoHc
3FzZWhfVQzeB6dXAOI7c/KCzj8SCewi9G8EpD/34rm9CgQ2ioaa33lNxHkgc/LhF
zZLi5mdQxH1TsuBFAMQaoSQSzgB/0uFfTN2SPTFp0tQgDPgi2empBwWPpsA7jEWL
J7onm9s69+IF5aeLqZpjIrRodArMI7sFnrHj3Ld2jcfnC1BZo+8WpteE5A9kAgwq
fdOYJBfbmzcVYF6dVY5Eew6jBy8AqL9pUlLivbXsoDAuJZr3qQJUJ65lpnKULFcG
U14CQtTRmZNEa2bai3uqZ75qn5djy6sVutz8XBjEOnHKx4lXUPjPW98Ck+C1av/q
bmZkAC+beo5+JI4EF+L9mQsxP+E7RTHS9CGn8xqGu3m+STH723GvETcPbPydWyAu
L9OJKT5bOxbyOcSxbQbbZ7fab/g1YQd8xBMvcBTj9i9MUssN6FZR5TSFOCXJZFdd
70IVyp0C6M2hiDBO5KhbBIaYjfKNCdWvjv+O2krM0OKcWwJ16Cr43hTdekdiySkO
kHlOhMvaY1mmy+k8cBEQA05Fge6FYWVS8h2zYhq02LwN5/rVgTamEQiWAeALKk4b
lWuLsELHdj09T8ETVIZ7dBpgUSnKYQO2vqDanSnPqxo3H7OdkvvYGIbC5SEat7Uu
nQzyyjdNh6H4+2f22IgqVNVOnYm3o6nbYVbGcEfJ3ijsL/Kvb0RFryxDFBOOUw49
F9tQE8GDHhshB2clDJ1tVdZrTjYOxtKEYPGze6DPJLkbby094Hqafqs7FBdLky3P
AsR5+RICGRWw9spDCBQ1WzXk4dlqmHdjR0KOLhbOp2OkSfW7wDqxshzo/xVCD9Ia
RFCoOVkKPGQnsARWbUKbs76fw0Nb2wdSzetHtio5uDvUtevdSmfpaI7jmEO8TFpK
qGsw++VkiJfGad5fYLYWnvlgnxLdMP6koHygQTINcaf4vp4q55zjcd485JWOBbpd
ClzD9AJn8JEOzuHnD0fZ+3mluNEARgTdhWp4pae7FU5a8YaOVr9pbKjdIyJmoo/Z
ytyvTNi6G0kAAlum/URWkh0vy3WAGOWKamy6cIK6tpzZvpd5yCCRqySzNNT59F+H
amw5nFQgNyqktpr5ktQCqPZ/AJn9ZrlfDJUhdjzzMLncwXEDsbYLunfDfNy+vKLk
deFzgZJ7o9GRBcHDqmn56B/q7Y5dFHVLK34sCk8p23KU3GpJyYWe7aHqmEIxctin
zPi9Qj1/RshI1V0AkFuEhtAko5lFszoH4PAfSHB+P5ALgVmVaVvsCd1SHZ+edrGg
Td8YBkseGjtEAN6Vig8ksR5L3ccMJE10RdZVTMKPP5ITB0wO1Kc6yG0pMBvTNqxp
DobCJgK+nzBGP5x0eJMh9gZT+T6/lAWyXFTbRlGTsSjRBBs929HO/gbyCW/d/0yk
6z+bcmJVIl98mQMWiG5kW9vjzy0vgGKW57VGMyrPeyQdD6H6X/vroZPq1gKZ5Tic
X1VuOxoEeJ4yAp/tVXdF61mCecBEQmJH/pc1MNDACo20oFyxe48/ayl4Vvd3IaK6
xwLFrhG2e+tus7Fbf1XfiZ0r+CKDRIYAb1ZmPsT5NRS9f7U0QnYM22gJSPSpJCo9
7Mk9vmWMUAO52ELJLwmbqFNnwRo+NXea6qNv0KIijtVmhyRJuTuBakAwlWbRqBJB
8ZReWREku5pF/Oq84DOA00BSfG5g4eX82KgQ/6+t8r/64LNJ099Q81yHZlZpPlj3
tZl6CEMk2CHR8tQA2zqZtJnnNah0QjDI2s87DCmFrn1jGAplWwCdm61ruX6jItBM
J4HIAhIgVarWu7byLnENnThkTaNzfv3AELRFQY4wuqdEYUhOyvPC8qwU6aKihHL3
Jlbi5WAsCdhy9yPvTaTsylgouElGs8I9pHbm2fpDbkta8SkbJYk62qmWutOvt0io
ZDqG5r48ATczksI882psOainFT4FGUxPYxgFe9Q7DrZfAps1fPSJlSqiG+zGMrvs
xLalHwVC1187NxjpQ3wjKtOd6wMwQahatV8cwey+o78W+dbph1XcIehzqlmJLY2U
4XXZno9wxOYIRsCtgMofbnrdPuY3WG6VFV7i1cj6JMSgGCt0oAq2PdKcYStJ0JAQ
PS7AVeakm01+MPTUJ0uVwJ5LEQOjsOZSxQpy4HcDS/coAYdICnXKUU7CKIBIGoSC
dTH/o15iDgBBtNDqr0Iluf7dFcoKF0P9iWTyee4rRPW3VHzhiqC/gUbx99sUpKP+
e52EDMiGd+DdRHk9775S94SV0a6I5YQm2zLcT5hY+ufvGAKlBml1/1zhDE3aAqSt
1AGH7ZxP3NS5TUTfFHOqUfkv+KGE3OPunAiq6ys0+J5p2YgHypc6jO733+Tw4om4
dDtdrxen/JqgcZCwNgHYd/l4wMZqDf8rQ8Q1yXRUzFJQZuX0I16xoFywuQWwsUEF
poNrL+o1KNlNgMp5w8sT2SrQVHW2mHzBLph5o/CRgvGOPWfLPF5mxiJl7VkAn7wS
KD1KBz8rfPUCO/9ULXjcHUcp8WtEqEBs1AwnwTWoxYW5f+RtV8Qbt+Qw9dFATzh/
rycMPiZlj+RgwqymT+R2YYwVfgcsN5QU0JoSdbLiCXDriur5BfvIAc4+ES/FtiIt
wIr93V6iqbO3swiFj149ndXel+MMneG8J8SR/hhZLVYSdu5mhoJEGdDj49WnepB+
fEKP7edUea4kfU5yJ2BrQIPIuuUXHiDakYNIy+0mfWvw764K3RtLrPc3ejKsYKjC
gcQN8vEMXh8TJhYdG7T8kPUDsaWTvK9Nzv+F1GcJ9sBgz0Zgdqh9OxvzrxdlCcJn
iejmH4PD2frZWE0Cb8Ddp3mPGe1V6+ZF/Is/suTTNosAigzSv+fDzq9WNQ1zjQ+d
4Nc9Tew2yFr4YfOtqf5JpQNw0+9l/VjAkKCK0OifVVyItcwbjyD4t7YTrsOX82zP
kUlnUOdofFBojDGfx5P7ewPtdgyENoJMG/m/+eVEAqDIU6R6KsjXKiH1XuqRTVKi
0pljt6s8JuBRarlqilh+wuN0F5kv39VCNrhvdzMzorUDpb4gNKmnHzf7nMnCLOMc
XP1TZeTR1ILggxtdQpDwISpyVhnpUeBdmgJ9FbsDcmu5QvboIs8dA9PnPks/V5OX
FkZ95b3qItHxeLKsZFTLub2yCvh5j8LLK5PLVGEBHXFMov9t+d/IE0FGhLnepjv1
7pUFGk6lw3HrXQIGAqCsBFF9fZT2uZIsSuTZ8DhpyKkaOu9VFjAwFt+GJHo+ElNj
WgcaAZNj8js4evHED4eYFWfx1Clp6gcuIRYIWMGfGsr0BUCPkZRCNCvPrdjXPcEY
d/s/hMmh/5ICU7TTmsqj8tzUkFcrjjFseTEmsFTEyW5yHi+JSA83xI5WoHy/zs+a
Vqde2gJbKJsiaihU0cWRDwkwZDqeALMWQ7bzrIBCsU7fN+cwAWRZyY2bQ7Qxqzyx
UObE3K1gJYqDm4yV0Z1JAOoKxCD0/bNolF1m/JfBU8yzvDske3Imtq34Ri8kxEV/
Jws5fUG2alEPMDrzplb8BfEANBaguy6pg0uvdrl+5qPsWjsBHini5qFacPue2Hlo
8hO3OWEs6M59KAlLxHtq548veXB7gTDqFVQENneFliiGRnRMfoz5Q5nGmNQgAnOV
Bk1P6wPGd6S+M2/WXm3OFkOeGCZuv4UexVEKHmrJCaDxYboTaHeoS5KnoG6JQD0R
7pAOYd+k+eLUnd5/QwTxW5o9/WWAQBCntAhPt5j+ivo15AuKuiYJZ+lPfIUG0UIW
gpBFbCbydw/yPxzRE9HtgAG9eXE13EgQfkTbk13UvoyuMhJiw/ksA4TYwPB3+Lvw
9xgrnDTXinoIH0YmVwk+Ofd1lD/JVNe4+nmN4uCU61hw+mGbIHWXmkJYcPODUWT2
6FJQSYYzsLsp/SghAI9H2XDejUYTN2WCrTghy+hDbfV7U37wTYVSPqpm2QSNa6yX
eG8maIJSOOXVmLEbaWvhLi2Qub5LgE6sjaPPQoyPG/dstBTLD/trMXD7qtIbQEG+
1blzD7fKFqlobyJuzfd+SehnAhErhc/Lw+TpAK4DE6hX42RTvzxBCSiEuo6NXzQY
bkekpsBGRGhoedl7gxyQK78h/jBnVmh6/CejlOxmE00uBWVwSeXle/pg8mkshVC3
1PZxWaXX2iM9ZJTxUG9Ebbg8TvtKElpaTY8fsVD8qhZeu8SdGlpWFKKbp5U22M+Z
P58mRoB+IXAUAy+migv93+pbIFLEosLE5WuZWjeQrHr1jrcI69N+gFNepSQmPBhQ
ZZI66r6oaNZpoy5wg7mcTB5lvOAknwHzh/8ahW3Meom0ysR7cJ12nzAzItT9lBAH
TTU5sH7k2411ePbtWDeZzsCFZtjoPIA01lWYBislFZR9OfKYbmOSDDBNjfqE1hsF
UPuloNhI9n0phvado34WdRDMH5gUPruRlxK1bgcIFat7J/Qfdk1CpLcnpphmf5ex
Mj+PfFTLQrSYQ+jv1c0oGpYUVAM3FJct5yg30/Tvv0yThVYdcRcoIa9VJKHV2pB/
9JseyK+mm1+hH6FuCbqskKF0KVfLrTCCBvNTKXpfusO4jjAup8EzVC9p1tLAJg4U
IhrO3LroMeWSnJW35SDcuwyNj3GEDs+qoe7HLQDfSdYHw+VuixbwbY8RWUY5TWEU
BwKeSxWHN7ZP+c9p4ktniaWqAjcic8BoKDlrwT83ebyYYazE6w7Nc0QAfbkzlG5W
RZXX1fTS+H5cTzqX4mxLUTIn9TaAJrPjuaeBlR/g5Ov4mwQ3OxusumK8Btmpiyr/
GWGSFsDEUQfJugDK9tOw3tZvjxr6t4NptKtKGHVW/foeuRecgcFkQfIuiRwcn+K3
LezZTDcVuGk//j+L28Hr0blDWdaYE4Fkyuf3GioT5fH/0fA77/N7vB8vAdfHRrh4
2F3YPnPODcs4zEdjiwvUS3d9sQ7whf4RIqynRv0VAALK9mKBsASWKXsAiwbVmo7r
29JDUFcuf3dmdsyIlgTXRDWXyhNSK8DD7qyX2GF6yTbrQ21hUKS+zSRcrR7FuILZ
Qb+AVKyCCTm/qk0yhG45MaSGRpoKZVn/GNrvs7I0jOlazFORDC2lULVos2JME9dN
e5Nw20uu4BOQUzXRT/yJKCchtK94BzVWIhYYDZefokHMrB/TZeuy4HIK3p0nOyqD
bICP5zHOlz3ummEa2PMdAXChkdfh8C677pdPtDvZZUDPTIgE7MyK287/5wmGFpnW
t9joWxrlI0ccCs+81xUKJpuD0A1uUpZxT15Lj3LAEJVbp6dgABu2lcOf2yj5NEZ9
f5ZwGPk1HMJWJ8YCdF6PiOwA7yl6tQCznnSHCIp3CEQcr0ct3LCk/ToOFKjF40Cr
s5Gk5QQux6CQgdkSgzE08CgkSaePx8bA5aXFlp+T8LAuTddpgpxl20VzprEWv6hi
MoigWQ0BjE7uYOm4+eTMpIMjJ+xby1goq1aihX8UX2iyZnBkl8nboL3MGPSO8YBg
6W3hxD3FZAtuyGve7IL0xH+PhQTEQ+a9I4kkHwof5atgSu8vI/HCdj/MuQJQrhdx
/F7fFPLnu3xjgjsQm8ceBKdKDx1Jl+a6tMUc4ektVTCab4cj2qbAQvAlU+rDAEI5
wMcBa6jX8+CyXzGWupX9mHVrHCcddpOnZxuNJjZ37rwQzKO/uH6o4Zqfl5M3Ue/R
cINg4M/2vEXtf1o8lwtSiziYr8aTGNbQk+W+igmlmSZE9Xg6llxlI3bkIrzFt9wP
sTP6JzhndcGMXlWI7cf5M2UleVeGv+3J7PKEXsbFmabuNPaq7P9/9PYjN8h3QHAY
hb+K2AungH9L/t8KfZmCUznan1rxm3oljjXMGK96Kfs3UJ8yrjyVpzkmSn67ln7I
63gCe4s6il17yItFWkI6tKbfwyZbX/X8fX/xuyd9R8o0KE+K4u4qpQ4EyolCvGzr
mNxGSVqDU/x7hPm9/DBjU/RYNtky51mjJ4lvb0xRrZVqHmW2IblkwO9qx/mdiqt3
Ww2UZciQG/r4UfQux9v3aRo6fAkWuEe07aS4GvnjCOoyV9wi4SS/Wot5VocygPRp
27tAK7MGc/WxFY+Lz7WLKsy5df5kTx0dHJTu4g6Pf2i83VKY94GfoZsStmmhVqbq
rVUJ6qI3VjgMKbEP7hvnXHk/m2sbNjo6IWMC4HoIJB9pY/vJ77PtIR4BVU8CuGxG
4kDt/gQPZRjKjk5hjhhbWgE8hejsDyBn/bebMsJp9RqAzoWysoOQtd8G9Y4AXvKG
mSZSKkQOqJcfx0sVU4pJCx4nqSWUZH00TAHOnDJrvzVNJLGksFWP5CSQt5qDSPIM
ztwflWxraprijLxtJgu3xx94xNBFtfs855cAcu2jRCd0HIVwBIV7QF0grQ0jPTs8
3qGvICADERWHVCSJe8mQIZXHmPxsqT/gVZiiIe/90Mbo4kp3tuHHs8Y3wIfkPPh4
H9cn0iOP+3baB9xU373EclAoqFgMHMy2m39TXa8P1Vx7z21w+EX7wfJF4mEsCf4W
g3G/O8S9BcZzawU+nhYfy9iF7dVIU/gto4NI4mWt7nIfCeyPytsWGGfgPAmG4TO7
H+nEen/51/tTqASWWdLwoe8JGMIOKK8k7nEDWg5fui0w8iWzYYLmkCmOnNB55jiH
VDaaFyi0A37+XeSgdf4wZgkh6YoALVmOWhmFBqjGJU+jBVeoTcXipdvulDCYjaqS
iZLTYmtwJ5IEL8RvgF4KxupJAVl2zFN69Cm3z5MHYvm0K8q5higpBkHuRN3JwQdK
HF25Wr6rNUXQKq3YtqAl69iz/lmMWZmTdrlDTZSWXg36yOe/Dv0iLUys/1T9BvPk
m6u4F9CH9q5JekbwUtX9cXQCB8RxJYH7kgHcyo3glT2rFGwOQ55dI4ZyqRh1FEet
kxgQMxv1DawPAfEoqFhC7jeLs1sDpXVbDbqEj+Oe+pQknAGYLf72Mw+zBg3L8Bp/
tujQwTI8BiPtEdeCgHGB/GEOG0gnZKCJ6g+mYAuXnGWaqhF/2QGHuYGlARx90Mvs
fUAxsx1wU+7GwJO8Aqjhwuvfb74SAI5wBVgZztQNRGI=
`protect end_protected
