localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTZ_CHK = {
  {32'hc3419a3f, 32'h00000000} /* (15, 15, 15) {real, imag} */,
  {32'hc285f0fe, 32'h00000000} /* (15, 15, 14) {real, imag} */,
  {32'h4358d1ac, 32'h00000000} /* (15, 15, 13) {real, imag} */,
  {32'h42dc3078, 32'h00000000} /* (15, 15, 12) {real, imag} */,
  {32'h42ae2544, 32'h00000000} /* (15, 15, 11) {real, imag} */,
  {32'h439ab249, 32'h00000000} /* (15, 15, 10) {real, imag} */,
  {32'hc29b067a, 32'h00000000} /* (15, 15, 9) {real, imag} */,
  {32'hc4034353, 32'h00000000} /* (15, 15, 8) {real, imag} */,
  {32'hc389def8, 32'h00000000} /* (15, 15, 7) {real, imag} */,
  {32'hc3fffc3a, 32'h00000000} /* (15, 15, 6) {real, imag} */,
  {32'hc46fa05d, 32'h00000000} /* (15, 15, 5) {real, imag} */,
  {32'hc4493ad3, 32'h00000000} /* (15, 15, 4) {real, imag} */,
  {32'hc43f7b6e, 32'h00000000} /* (15, 15, 3) {real, imag} */,
  {32'hc46fa5dc, 32'h00000000} /* (15, 15, 2) {real, imag} */,
  {32'hc3d3cf50, 32'h00000000} /* (15, 15, 1) {real, imag} */,
  {32'hc322b1e4, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hc2cd1b9e, 32'h00000000} /* (15, 14, 15) {real, imag} */,
  {32'hc3fff3fd, 32'h00000000} /* (15, 14, 14) {real, imag} */,
  {32'hc2bc0a68, 32'h00000000} /* (15, 14, 13) {real, imag} */,
  {32'h435a7a35, 32'h00000000} /* (15, 14, 12) {real, imag} */,
  {32'hc3059775, 32'h00000000} /* (15, 14, 11) {real, imag} */,
  {32'hc1f91e10, 32'h00000000} /* (15, 14, 10) {real, imag} */,
  {32'h431c1d29, 32'h00000000} /* (15, 14, 9) {real, imag} */,
  {32'hc2f57166, 32'h00000000} /* (15, 14, 8) {real, imag} */,
  {32'hc321e1f1, 32'h00000000} /* (15, 14, 7) {real, imag} */,
  {32'hc3b5ca77, 32'h00000000} /* (15, 14, 6) {real, imag} */,
  {32'hc48cc096, 32'h00000000} /* (15, 14, 5) {real, imag} */,
  {32'hc3ae4a6e, 32'h00000000} /* (15, 14, 4) {real, imag} */,
  {32'hc41ac87b, 32'h00000000} /* (15, 14, 3) {real, imag} */,
  {32'hc3a73e42, 32'h00000000} /* (15, 14, 2) {real, imag} */,
  {32'hc39588ca, 32'h00000000} /* (15, 14, 1) {real, imag} */,
  {32'hc3b31176, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'h4380ba40, 32'h00000000} /* (15, 13, 15) {real, imag} */,
  {32'h4319e4f2, 32'h00000000} /* (15, 13, 14) {real, imag} */,
  {32'hc343d7d7, 32'h00000000} /* (15, 13, 13) {real, imag} */,
  {32'hc3ef1496, 32'h00000000} /* (15, 13, 12) {real, imag} */,
  {32'hc2942f3c, 32'h00000000} /* (15, 13, 11) {real, imag} */,
  {32'hc37d4197, 32'h00000000} /* (15, 13, 10) {real, imag} */,
  {32'hc45e6e94, 32'h00000000} /* (15, 13, 9) {real, imag} */,
  {32'h4351a120, 32'h00000000} /* (15, 13, 8) {real, imag} */,
  {32'hc2fe48a2, 32'h00000000} /* (15, 13, 7) {real, imag} */,
  {32'h438a3dd9, 32'h00000000} /* (15, 13, 6) {real, imag} */,
  {32'hc22c6c04, 32'h00000000} /* (15, 13, 5) {real, imag} */,
  {32'hc3d5dfce, 32'h00000000} /* (15, 13, 4) {real, imag} */,
  {32'hc3b4dca6, 32'h00000000} /* (15, 13, 3) {real, imag} */,
  {32'hc39945ca, 32'h00000000} /* (15, 13, 2) {real, imag} */,
  {32'h44137830, 32'h00000000} /* (15, 13, 1) {real, imag} */,
  {32'h441cd426, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'h44016f5a, 32'h00000000} /* (15, 12, 15) {real, imag} */,
  {32'h44330924, 32'h00000000} /* (15, 12, 14) {real, imag} */,
  {32'hc19411c8, 32'h00000000} /* (15, 12, 13) {real, imag} */,
  {32'hc33a8ef0, 32'h00000000} /* (15, 12, 12) {real, imag} */,
  {32'hc3ae788e, 32'h00000000} /* (15, 12, 11) {real, imag} */,
  {32'hc393c3de, 32'h00000000} /* (15, 12, 10) {real, imag} */,
  {32'hc2830aee, 32'h00000000} /* (15, 12, 9) {real, imag} */,
  {32'h4159db90, 32'h00000000} /* (15, 12, 8) {real, imag} */,
  {32'hc31c4d86, 32'h00000000} /* (15, 12, 7) {real, imag} */,
  {32'h42400208, 32'h00000000} /* (15, 12, 6) {real, imag} */,
  {32'h4363ab3f, 32'h00000000} /* (15, 12, 5) {real, imag} */,
  {32'hc33107c0, 32'h00000000} /* (15, 12, 4) {real, imag} */,
  {32'hc41a8343, 32'h00000000} /* (15, 12, 3) {real, imag} */,
  {32'hc2f4dd16, 32'h00000000} /* (15, 12, 2) {real, imag} */,
  {32'h436b1c59, 32'h00000000} /* (15, 12, 1) {real, imag} */,
  {32'h4343f2d3, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'h4457a892, 32'h00000000} /* (15, 11, 15) {real, imag} */,
  {32'h441f684e, 32'h00000000} /* (15, 11, 14) {real, imag} */,
  {32'h43891cdd, 32'h00000000} /* (15, 11, 13) {real, imag} */,
  {32'h4401dfa6, 32'h00000000} /* (15, 11, 12) {real, imag} */,
  {32'hc3d8aeb0, 32'h00000000} /* (15, 11, 11) {real, imag} */,
  {32'hc3994e74, 32'h00000000} /* (15, 11, 10) {real, imag} */,
  {32'hc2c725cd, 32'h00000000} /* (15, 11, 9) {real, imag} */,
  {32'hc34995b4, 32'h00000000} /* (15, 11, 8) {real, imag} */,
  {32'hc341d736, 32'h00000000} /* (15, 11, 7) {real, imag} */,
  {32'h4354e052, 32'h00000000} /* (15, 11, 6) {real, imag} */,
  {32'hc31735a6, 32'h00000000} /* (15, 11, 5) {real, imag} */,
  {32'hc3dee575, 32'h00000000} /* (15, 11, 4) {real, imag} */,
  {32'hc35a3503, 32'h00000000} /* (15, 11, 3) {real, imag} */,
  {32'h4392c598, 32'h00000000} /* (15, 11, 2) {real, imag} */,
  {32'h42733a66, 32'h00000000} /* (15, 11, 1) {real, imag} */,
  {32'h429e35b9, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h440c958c, 32'h00000000} /* (15, 10, 15) {real, imag} */,
  {32'h44376b42, 32'h00000000} /* (15, 10, 14) {real, imag} */,
  {32'hc1643a38, 32'h00000000} /* (15, 10, 13) {real, imag} */,
  {32'h428646b8, 32'h00000000} /* (15, 10, 12) {real, imag} */,
  {32'h4422e408, 32'h00000000} /* (15, 10, 11) {real, imag} */,
  {32'h43d3bfd4, 32'h00000000} /* (15, 10, 10) {real, imag} */,
  {32'hc41bec56, 32'h00000000} /* (15, 10, 9) {real, imag} */,
  {32'hc4207b42, 32'h00000000} /* (15, 10, 8) {real, imag} */,
  {32'hc294ae3c, 32'h00000000} /* (15, 10, 7) {real, imag} */,
  {32'h4292d34c, 32'h00000000} /* (15, 10, 6) {real, imag} */,
  {32'hc3139cb4, 32'h00000000} /* (15, 10, 5) {real, imag} */,
  {32'hc2a168b0, 32'h00000000} /* (15, 10, 4) {real, imag} */,
  {32'hc33b3c2e, 32'h00000000} /* (15, 10, 3) {real, imag} */,
  {32'h43b06634, 32'h00000000} /* (15, 10, 2) {real, imag} */,
  {32'h43ad609e, 32'h00000000} /* (15, 10, 1) {real, imag} */,
  {32'h439971ab, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'h428de9be, 32'h00000000} /* (15, 9, 15) {real, imag} */,
  {32'hc42168bc, 32'h00000000} /* (15, 9, 14) {real, imag} */,
  {32'h43c804ae, 32'h00000000} /* (15, 9, 13) {real, imag} */,
  {32'h413ee128, 32'h00000000} /* (15, 9, 12) {real, imag} */,
  {32'h43643450, 32'h00000000} /* (15, 9, 11) {real, imag} */,
  {32'h43b5c5dd, 32'h00000000} /* (15, 9, 10) {real, imag} */,
  {32'hc4412b86, 32'h00000000} /* (15, 9, 9) {real, imag} */,
  {32'hc40689fe, 32'h00000000} /* (15, 9, 8) {real, imag} */,
  {32'hc25d3c2b, 32'h00000000} /* (15, 9, 7) {real, imag} */,
  {32'hc40020b0, 32'h00000000} /* (15, 9, 6) {real, imag} */,
  {32'hc42246ad, 32'h00000000} /* (15, 9, 5) {real, imag} */,
  {32'hc30caf0a, 32'h00000000} /* (15, 9, 4) {real, imag} */,
  {32'h42dc9a69, 32'h00000000} /* (15, 9, 3) {real, imag} */,
  {32'h4384b3d9, 32'h00000000} /* (15, 9, 2) {real, imag} */,
  {32'h435f7ed0, 32'h00000000} /* (15, 9, 1) {real, imag} */,
  {32'h436d553e, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'h42b566e6, 32'h00000000} /* (15, 8, 15) {real, imag} */,
  {32'hc427161e, 32'h00000000} /* (15, 8, 14) {real, imag} */,
  {32'hc2a99c54, 32'h00000000} /* (15, 8, 13) {real, imag} */,
  {32'hc1a3172a, 32'h00000000} /* (15, 8, 12) {real, imag} */,
  {32'h431f22be, 32'h00000000} /* (15, 8, 11) {real, imag} */,
  {32'h437a4a0c, 32'h00000000} /* (15, 8, 10) {real, imag} */,
  {32'h4320391f, 32'h00000000} /* (15, 8, 9) {real, imag} */,
  {32'hc46cabea, 32'h00000000} /* (15, 8, 8) {real, imag} */,
  {32'hc4088501, 32'h00000000} /* (15, 8, 7) {real, imag} */,
  {32'hc36d9202, 32'h00000000} /* (15, 8, 6) {real, imag} */,
  {32'hc3c1c901, 32'h00000000} /* (15, 8, 5) {real, imag} */,
  {32'h41a621ca, 32'h00000000} /* (15, 8, 4) {real, imag} */,
  {32'h43948efe, 32'h00000000} /* (15, 8, 3) {real, imag} */,
  {32'h42e78410, 32'h00000000} /* (15, 8, 2) {real, imag} */,
  {32'h439c3900, 32'h00000000} /* (15, 8, 1) {real, imag} */,
  {32'h41ed7e60, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h432800e4, 32'h00000000} /* (15, 7, 15) {real, imag} */,
  {32'h43183174, 32'h00000000} /* (15, 7, 14) {real, imag} */,
  {32'hc317ef5a, 32'h00000000} /* (15, 7, 13) {real, imag} */,
  {32'hc3978aa3, 32'h00000000} /* (15, 7, 12) {real, imag} */,
  {32'hc3f9871e, 32'h00000000} /* (15, 7, 11) {real, imag} */,
  {32'h4224be9e, 32'h00000000} /* (15, 7, 10) {real, imag} */,
  {32'hc192c994, 32'h00000000} /* (15, 7, 9) {real, imag} */,
  {32'hc3b25ee2, 32'h00000000} /* (15, 7, 8) {real, imag} */,
  {32'h408b2ef0, 32'h00000000} /* (15, 7, 7) {real, imag} */,
  {32'h43022fc8, 32'h00000000} /* (15, 7, 6) {real, imag} */,
  {32'hc3191f9e, 32'h00000000} /* (15, 7, 5) {real, imag} */,
  {32'h43154a76, 32'h00000000} /* (15, 7, 4) {real, imag} */,
  {32'hc2da4b32, 32'h00000000} /* (15, 7, 3) {real, imag} */,
  {32'hc3799644, 32'h00000000} /* (15, 7, 2) {real, imag} */,
  {32'hc37335a6, 32'h00000000} /* (15, 7, 1) {real, imag} */,
  {32'h42bd96d0, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'hc329afd4, 32'h00000000} /* (15, 6, 15) {real, imag} */,
  {32'hc2802be9, 32'h00000000} /* (15, 6, 14) {real, imag} */,
  {32'hc4035954, 32'h00000000} /* (15, 6, 13) {real, imag} */,
  {32'h4297db3a, 32'h00000000} /* (15, 6, 12) {real, imag} */,
  {32'hc198dc42, 32'h00000000} /* (15, 6, 11) {real, imag} */,
  {32'h43e6a19f, 32'h00000000} /* (15, 6, 10) {real, imag} */,
  {32'h43b14d28, 32'h00000000} /* (15, 6, 9) {real, imag} */,
  {32'h4383c546, 32'h00000000} /* (15, 6, 8) {real, imag} */,
  {32'h438bb2aa, 32'h00000000} /* (15, 6, 7) {real, imag} */,
  {32'h43504994, 32'h00000000} /* (15, 6, 6) {real, imag} */,
  {32'hc34c264e, 32'h00000000} /* (15, 6, 5) {real, imag} */,
  {32'hc28eb6c6, 32'h00000000} /* (15, 6, 4) {real, imag} */,
  {32'hc2ec6f02, 32'h00000000} /* (15, 6, 3) {real, imag} */,
  {32'hc3ffae79, 32'h00000000} /* (15, 6, 2) {real, imag} */,
  {32'hc4019e97, 32'h00000000} /* (15, 6, 1) {real, imag} */,
  {32'h4240912c, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h43607b70, 32'h00000000} /* (15, 5, 15) {real, imag} */,
  {32'h4366b4b0, 32'h00000000} /* (15, 5, 14) {real, imag} */,
  {32'h423fec28, 32'h00000000} /* (15, 5, 13) {real, imag} */,
  {32'h43da6f1d, 32'h00000000} /* (15, 5, 12) {real, imag} */,
  {32'h431615b4, 32'h00000000} /* (15, 5, 11) {real, imag} */,
  {32'h42148a74, 32'h00000000} /* (15, 5, 10) {real, imag} */,
  {32'h4384f662, 32'h00000000} /* (15, 5, 9) {real, imag} */,
  {32'hc1f64d7c, 32'h00000000} /* (15, 5, 8) {real, imag} */,
  {32'hc255ddc2, 32'h00000000} /* (15, 5, 7) {real, imag} */,
  {32'hc3d7f83e, 32'h00000000} /* (15, 5, 6) {real, imag} */,
  {32'hc3d9a3f3, 32'h00000000} /* (15, 5, 5) {real, imag} */,
  {32'hc416e43c, 32'h00000000} /* (15, 5, 4) {real, imag} */,
  {32'hc3beed40, 32'h00000000} /* (15, 5, 3) {real, imag} */,
  {32'h43b84b2a, 32'h00000000} /* (15, 5, 2) {real, imag} */,
  {32'h43925ea6, 32'h00000000} /* (15, 5, 1) {real, imag} */,
  {32'h4210904a, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'h4335d140, 32'h00000000} /* (15, 4, 15) {real, imag} */,
  {32'h40996e80, 32'h00000000} /* (15, 4, 14) {real, imag} */,
  {32'hc36ff34e, 32'h00000000} /* (15, 4, 13) {real, imag} */,
  {32'h43880a11, 32'h00000000} /* (15, 4, 12) {real, imag} */,
  {32'hc1ffad6a, 32'h00000000} /* (15, 4, 11) {real, imag} */,
  {32'h439e30cf, 32'h00000000} /* (15, 4, 10) {real, imag} */,
  {32'hc2de8c76, 32'h00000000} /* (15, 4, 9) {real, imag} */,
  {32'hc1ee1ae0, 32'h00000000} /* (15, 4, 8) {real, imag} */,
  {32'hc32497a6, 32'h00000000} /* (15, 4, 7) {real, imag} */,
  {32'hc38d5845, 32'h00000000} /* (15, 4, 6) {real, imag} */,
  {32'hc444fe74, 32'h00000000} /* (15, 4, 5) {real, imag} */,
  {32'hc2e4f730, 32'h00000000} /* (15, 4, 4) {real, imag} */,
  {32'hc312b8e9, 32'h00000000} /* (15, 4, 3) {real, imag} */,
  {32'h43756b72, 32'h00000000} /* (15, 4, 2) {real, imag} */,
  {32'hc397acb2, 32'h00000000} /* (15, 4, 1) {real, imag} */,
  {32'hc3a3bb25, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'hc34e2a20, 32'h00000000} /* (15, 3, 15) {real, imag} */,
  {32'h43637332, 32'h00000000} /* (15, 3, 14) {real, imag} */,
  {32'h4356f640, 32'h00000000} /* (15, 3, 13) {real, imag} */,
  {32'h43da6562, 32'h00000000} /* (15, 3, 12) {real, imag} */,
  {32'h434d1452, 32'h00000000} /* (15, 3, 11) {real, imag} */,
  {32'h44737b7e, 32'h00000000} /* (15, 3, 10) {real, imag} */,
  {32'h42ee1d5a, 32'h00000000} /* (15, 3, 9) {real, imag} */,
  {32'h4215954c, 32'h00000000} /* (15, 3, 8) {real, imag} */,
  {32'hc400b741, 32'h00000000} /* (15, 3, 7) {real, imag} */,
  {32'h41c8bf0c, 32'h00000000} /* (15, 3, 6) {real, imag} */,
  {32'hc45adca2, 32'h00000000} /* (15, 3, 5) {real, imag} */,
  {32'hc3e4bae2, 32'h00000000} /* (15, 3, 4) {real, imag} */,
  {32'hc3203e82, 32'h00000000} /* (15, 3, 3) {real, imag} */,
  {32'hc425243a, 32'h00000000} /* (15, 3, 2) {real, imag} */,
  {32'hc345b0f9, 32'h00000000} /* (15, 3, 1) {real, imag} */,
  {32'h43b725e0, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'hbe69f400, 32'h00000000} /* (15, 2, 15) {real, imag} */,
  {32'h42946f80, 32'h00000000} /* (15, 2, 14) {real, imag} */,
  {32'h4461249c, 32'h00000000} /* (15, 2, 13) {real, imag} */,
  {32'h44242026, 32'h00000000} /* (15, 2, 12) {real, imag} */,
  {32'h430c4eaa, 32'h00000000} /* (15, 2, 11) {real, imag} */,
  {32'h42efbb48, 32'h00000000} /* (15, 2, 10) {real, imag} */,
  {32'h43b5b6fa, 32'h00000000} /* (15, 2, 9) {real, imag} */,
  {32'h437ca09d, 32'h00000000} /* (15, 2, 8) {real, imag} */,
  {32'hc3fa8618, 32'h00000000} /* (15, 2, 7) {real, imag} */,
  {32'hc4884625, 32'h00000000} /* (15, 2, 6) {real, imag} */,
  {32'hc4387a04, 32'h00000000} /* (15, 2, 5) {real, imag} */,
  {32'hc48aeee6, 32'h00000000} /* (15, 2, 4) {real, imag} */,
  {32'hc4258408, 32'h00000000} /* (15, 2, 3) {real, imag} */,
  {32'hc466668f, 32'h00000000} /* (15, 2, 2) {real, imag} */,
  {32'hc4386333, 32'h00000000} /* (15, 2, 1) {real, imag} */,
  {32'h438d43e5, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'h422b1c40, 32'h00000000} /* (15, 1, 15) {real, imag} */,
  {32'hc357766c, 32'h00000000} /* (15, 1, 14) {real, imag} */,
  {32'h42279ff0, 32'h00000000} /* (15, 1, 13) {real, imag} */,
  {32'h43b25bc2, 32'h00000000} /* (15, 1, 12) {real, imag} */,
  {32'h43d9689c, 32'h00000000} /* (15, 1, 11) {real, imag} */,
  {32'h43c25c55, 32'h00000000} /* (15, 1, 10) {real, imag} */,
  {32'h4395646a, 32'h00000000} /* (15, 1, 9) {real, imag} */,
  {32'h42c1c24c, 32'h00000000} /* (15, 1, 8) {real, imag} */,
  {32'hc41ba2e1, 32'h00000000} /* (15, 1, 7) {real, imag} */,
  {32'hc4a4d312, 32'h00000000} /* (15, 1, 6) {real, imag} */,
  {32'hc4c7810a, 32'h00000000} /* (15, 1, 5) {real, imag} */,
  {32'hc45b578f, 32'h00000000} /* (15, 1, 4) {real, imag} */,
  {32'hc454da58, 32'h00000000} /* (15, 1, 3) {real, imag} */,
  {32'hc3d0c54b, 32'h00000000} /* (15, 1, 2) {real, imag} */,
  {32'hc415f7e0, 32'h00000000} /* (15, 1, 1) {real, imag} */,
  {32'hc401c918, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'hbf7ba900, 32'h00000000} /* (15, 0, 15) {real, imag} */,
  {32'h4317b628, 32'h00000000} /* (15, 0, 14) {real, imag} */,
  {32'hc34b0812, 32'h00000000} /* (15, 0, 13) {real, imag} */,
  {32'h4280c034, 32'h00000000} /* (15, 0, 12) {real, imag} */,
  {32'h43169d39, 32'h00000000} /* (15, 0, 11) {real, imag} */,
  {32'hc30bbe62, 32'h00000000} /* (15, 0, 10) {real, imag} */,
  {32'h416c3780, 32'h00000000} /* (15, 0, 9) {real, imag} */,
  {32'hc3aacb06, 32'h00000000} /* (15, 0, 8) {real, imag} */,
  {32'hc3dd5ef0, 32'h00000000} /* (15, 0, 7) {real, imag} */,
  {32'hc3b6beb0, 32'h00000000} /* (15, 0, 6) {real, imag} */,
  {32'hc432b638, 32'h00000000} /* (15, 0, 5) {real, imag} */,
  {32'hc41d2880, 32'h00000000} /* (15, 0, 4) {real, imag} */,
  {32'hc405ec70, 32'h00000000} /* (15, 0, 3) {real, imag} */,
  {32'hc407062e, 32'h00000000} /* (15, 0, 2) {real, imag} */,
  {32'hc3af12f3, 32'h00000000} /* (15, 0, 1) {real, imag} */,
  {32'hc372dcb5, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h43cf75ee, 32'h00000000} /* (14, 15, 15) {real, imag} */,
  {32'hc3c293a2, 32'h00000000} /* (14, 15, 14) {real, imag} */,
  {32'h4276cf89, 32'h00000000} /* (14, 15, 13) {real, imag} */,
  {32'h43145f11, 32'h00000000} /* (14, 15, 12) {real, imag} */,
  {32'hc2483cc8, 32'h00000000} /* (14, 15, 11) {real, imag} */,
  {32'hc3ff6e5b, 32'h00000000} /* (14, 15, 10) {real, imag} */,
  {32'hc44e118d, 32'h00000000} /* (14, 15, 9) {real, imag} */,
  {32'hc418b642, 32'h00000000} /* (14, 15, 8) {real, imag} */,
  {32'hc3deb2fc, 32'h00000000} /* (14, 15, 7) {real, imag} */,
  {32'hc2f3ba08, 32'h00000000} /* (14, 15, 6) {real, imag} */,
  {32'h43066f12, 32'h00000000} /* (14, 15, 5) {real, imag} */,
  {32'hc410734c, 32'h00000000} /* (14, 15, 4) {real, imag} */,
  {32'hc4267986, 32'h00000000} /* (14, 15, 3) {real, imag} */,
  {32'hc3b035b9, 32'h00000000} /* (14, 15, 2) {real, imag} */,
  {32'hc4857e26, 32'h00000000} /* (14, 15, 1) {real, imag} */,
  {32'hc38e21ec, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'h430f6054, 32'h00000000} /* (14, 14, 15) {real, imag} */,
  {32'hc413ef92, 32'h00000000} /* (14, 14, 14) {real, imag} */,
  {32'hc0aeb260, 32'h00000000} /* (14, 14, 13) {real, imag} */,
  {32'hc39fa5d1, 32'h00000000} /* (14, 14, 12) {real, imag} */,
  {32'h438dc9d2, 32'h00000000} /* (14, 14, 11) {real, imag} */,
  {32'h436fc894, 32'h00000000} /* (14, 14, 10) {real, imag} */,
  {32'hc429b060, 32'h00000000} /* (14, 14, 9) {real, imag} */,
  {32'hc4054c66, 32'h00000000} /* (14, 14, 8) {real, imag} */,
  {32'h42db7813, 32'h00000000} /* (14, 14, 7) {real, imag} */,
  {32'hc3a241f3, 32'h00000000} /* (14, 14, 6) {real, imag} */,
  {32'hc3feb63a, 32'h00000000} /* (14, 14, 5) {real, imag} */,
  {32'hc3b0a9d3, 32'h00000000} /* (14, 14, 4) {real, imag} */,
  {32'hc4045eeb, 32'h00000000} /* (14, 14, 3) {real, imag} */,
  {32'hc4273155, 32'h00000000} /* (14, 14, 2) {real, imag} */,
  {32'hc444598a, 32'h00000000} /* (14, 14, 1) {real, imag} */,
  {32'hc281589c, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'h43d44672, 32'h00000000} /* (14, 13, 15) {real, imag} */,
  {32'h43d4eb2d, 32'h00000000} /* (14, 13, 14) {real, imag} */,
  {32'hc3860387, 32'h00000000} /* (14, 13, 13) {real, imag} */,
  {32'hc47edf70, 32'h00000000} /* (14, 13, 12) {real, imag} */,
  {32'hc3d9e84d, 32'h00000000} /* (14, 13, 11) {real, imag} */,
  {32'hc2999c64, 32'h00000000} /* (14, 13, 10) {real, imag} */,
  {32'h43592560, 32'h00000000} /* (14, 13, 9) {real, imag} */,
  {32'hc2e9e614, 32'h00000000} /* (14, 13, 8) {real, imag} */,
  {32'hc404dff5, 32'h00000000} /* (14, 13, 7) {real, imag} */,
  {32'h43abe8e1, 32'h00000000} /* (14, 13, 6) {real, imag} */,
  {32'hc3a4bba5, 32'h00000000} /* (14, 13, 5) {real, imag} */,
  {32'h42c1b104, 32'h00000000} /* (14, 13, 4) {real, imag} */,
  {32'hc3d8349b, 32'h00000000} /* (14, 13, 3) {real, imag} */,
  {32'hc4310732, 32'h00000000} /* (14, 13, 2) {real, imag} */,
  {32'h42cb2f14, 32'h00000000} /* (14, 13, 1) {real, imag} */,
  {32'h440bd9b6, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'h43ad2878, 32'h00000000} /* (14, 12, 15) {real, imag} */,
  {32'h431819bc, 32'h00000000} /* (14, 12, 14) {real, imag} */,
  {32'h423a66d4, 32'h00000000} /* (14, 12, 13) {real, imag} */,
  {32'hc304d73a, 32'h00000000} /* (14, 12, 12) {real, imag} */,
  {32'hc4b07f20, 32'h00000000} /* (14, 12, 11) {real, imag} */,
  {32'h42640558, 32'h00000000} /* (14, 12, 10) {real, imag} */,
  {32'hc410a01e, 32'h00000000} /* (14, 12, 9) {real, imag} */,
  {32'hc418a2b1, 32'h00000000} /* (14, 12, 8) {real, imag} */,
  {32'hc40b4e3f, 32'h00000000} /* (14, 12, 7) {real, imag} */,
  {32'hc410600f, 32'h00000000} /* (14, 12, 6) {real, imag} */,
  {32'hc3af0188, 32'h00000000} /* (14, 12, 5) {real, imag} */,
  {32'hc44421fe, 32'h00000000} /* (14, 12, 4) {real, imag} */,
  {32'hc3b9253e, 32'h00000000} /* (14, 12, 3) {real, imag} */,
  {32'hc3ecd1a3, 32'h00000000} /* (14, 12, 2) {real, imag} */,
  {32'h44160570, 32'h00000000} /* (14, 12, 1) {real, imag} */,
  {32'h43a7d3a2, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'h43c2dc5c, 32'h00000000} /* (14, 11, 15) {real, imag} */,
  {32'h443476dd, 32'h00000000} /* (14, 11, 14) {real, imag} */,
  {32'h43e5ddd8, 32'h00000000} /* (14, 11, 13) {real, imag} */,
  {32'h43a72544, 32'h00000000} /* (14, 11, 12) {real, imag} */,
  {32'h43eab9e7, 32'h00000000} /* (14, 11, 11) {real, imag} */,
  {32'hc4496ef4, 32'h00000000} /* (14, 11, 10) {real, imag} */,
  {32'hc210afaa, 32'h00000000} /* (14, 11, 9) {real, imag} */,
  {32'h43c90eb4, 32'h00000000} /* (14, 11, 8) {real, imag} */,
  {32'hc397c470, 32'h00000000} /* (14, 11, 7) {real, imag} */,
  {32'hc3f56986, 32'h00000000} /* (14, 11, 6) {real, imag} */,
  {32'hc3860c30, 32'h00000000} /* (14, 11, 5) {real, imag} */,
  {32'h4447bc86, 32'h00000000} /* (14, 11, 4) {real, imag} */,
  {32'h4326ae82, 32'h00000000} /* (14, 11, 3) {real, imag} */,
  {32'hc34f41a2, 32'h00000000} /* (14, 11, 2) {real, imag} */,
  {32'h4386cbed, 32'h00000000} /* (14, 11, 1) {real, imag} */,
  {32'hc245f674, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h42e62069, 32'h00000000} /* (14, 10, 15) {real, imag} */,
  {32'h44835170, 32'h00000000} /* (14, 10, 14) {real, imag} */,
  {32'h4299799d, 32'h00000000} /* (14, 10, 13) {real, imag} */,
  {32'hc371bf66, 32'h00000000} /* (14, 10, 12) {real, imag} */,
  {32'h4350f0db, 32'h00000000} /* (14, 10, 11) {real, imag} */,
  {32'hc3806305, 32'h00000000} /* (14, 10, 10) {real, imag} */,
  {32'hc395474f, 32'h00000000} /* (14, 10, 9) {real, imag} */,
  {32'h42fd9a70, 32'h00000000} /* (14, 10, 8) {real, imag} */,
  {32'h43b31aa6, 32'h00000000} /* (14, 10, 7) {real, imag} */,
  {32'hc38212da, 32'h00000000} /* (14, 10, 6) {real, imag} */,
  {32'hc33812b2, 32'h00000000} /* (14, 10, 5) {real, imag} */,
  {32'h4401be7c, 32'h00000000} /* (14, 10, 4) {real, imag} */,
  {32'h433a89f5, 32'h00000000} /* (14, 10, 3) {real, imag} */,
  {32'hc3ff8ad7, 32'h00000000} /* (14, 10, 2) {real, imag} */,
  {32'h43ca7471, 32'h00000000} /* (14, 10, 1) {real, imag} */,
  {32'h440679ff, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'hc22f0a00, 32'h00000000} /* (14, 9, 15) {real, imag} */,
  {32'hc3334946, 32'h00000000} /* (14, 9, 14) {real, imag} */,
  {32'hc39185ee, 32'h00000000} /* (14, 9, 13) {real, imag} */,
  {32'h44877c55, 32'h00000000} /* (14, 9, 12) {real, imag} */,
  {32'h448f9597, 32'h00000000} /* (14, 9, 11) {real, imag} */,
  {32'h440eafb3, 32'h00000000} /* (14, 9, 10) {real, imag} */,
  {32'hc4b5b81e, 32'h00000000} /* (14, 9, 9) {real, imag} */,
  {32'hc31751d0, 32'h00000000} /* (14, 9, 8) {real, imag} */,
  {32'hc391f2b6, 32'h00000000} /* (14, 9, 7) {real, imag} */,
  {32'hc45040b2, 32'h00000000} /* (14, 9, 6) {real, imag} */,
  {32'h4329a587, 32'h00000000} /* (14, 9, 5) {real, imag} */,
  {32'hc40b38dc, 32'h00000000} /* (14, 9, 4) {real, imag} */,
  {32'h4324b536, 32'h00000000} /* (14, 9, 3) {real, imag} */,
  {32'hc3a15a4c, 32'h00000000} /* (14, 9, 2) {real, imag} */,
  {32'hc3cbfb26, 32'h00000000} /* (14, 9, 1) {real, imag} */,
  {32'h4486f088, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'hc3487f71, 32'h00000000} /* (14, 8, 15) {real, imag} */,
  {32'hc44815d6, 32'h00000000} /* (14, 8, 14) {real, imag} */,
  {32'h4246663b, 32'h00000000} /* (14, 8, 13) {real, imag} */,
  {32'hc3dd5079, 32'h00000000} /* (14, 8, 12) {real, imag} */,
  {32'h44202718, 32'h00000000} /* (14, 8, 11) {real, imag} */,
  {32'h447aba1b, 32'h00000000} /* (14, 8, 10) {real, imag} */,
  {32'hc32c076b, 32'h00000000} /* (14, 8, 9) {real, imag} */,
  {32'h43aa898e, 32'h00000000} /* (14, 8, 8) {real, imag} */,
  {32'hc3c51524, 32'h00000000} /* (14, 8, 7) {real, imag} */,
  {32'hc44dc8a8, 32'h00000000} /* (14, 8, 6) {real, imag} */,
  {32'hc2872124, 32'h00000000} /* (14, 8, 5) {real, imag} */,
  {32'h44311590, 32'h00000000} /* (14, 8, 4) {real, imag} */,
  {32'h4313e97f, 32'h00000000} /* (14, 8, 3) {real, imag} */,
  {32'h42246fb0, 32'h00000000} /* (14, 8, 2) {real, imag} */,
  {32'h42f6b9f6, 32'h00000000} /* (14, 8, 1) {real, imag} */,
  {32'hc075ce40, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'h408fb7a0, 32'h00000000} /* (14, 7, 15) {real, imag} */,
  {32'hc42998d9, 32'h00000000} /* (14, 7, 14) {real, imag} */,
  {32'hc449bed8, 32'h00000000} /* (14, 7, 13) {real, imag} */,
  {32'hc499b09e, 32'h00000000} /* (14, 7, 12) {real, imag} */,
  {32'h43c4e308, 32'h00000000} /* (14, 7, 11) {real, imag} */,
  {32'h445fca10, 32'h00000000} /* (14, 7, 10) {real, imag} */,
  {32'h4454c07e, 32'h00000000} /* (14, 7, 9) {real, imag} */,
  {32'h437152ef, 32'h00000000} /* (14, 7, 8) {real, imag} */,
  {32'hc3665d50, 32'h00000000} /* (14, 7, 7) {real, imag} */,
  {32'h431a7f2c, 32'h00000000} /* (14, 7, 6) {real, imag} */,
  {32'h438ffc5d, 32'h00000000} /* (14, 7, 5) {real, imag} */,
  {32'hc3899eaa, 32'h00000000} /* (14, 7, 4) {real, imag} */,
  {32'hc41de54a, 32'h00000000} /* (14, 7, 3) {real, imag} */,
  {32'hc3539290, 32'h00000000} /* (14, 7, 2) {real, imag} */,
  {32'hc2c09fb8, 32'h00000000} /* (14, 7, 1) {real, imag} */,
  {32'hc350dfb7, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'hc2baa866, 32'h00000000} /* (14, 6, 15) {real, imag} */,
  {32'h429a6698, 32'h00000000} /* (14, 6, 14) {real, imag} */,
  {32'hc3bbdede, 32'h00000000} /* (14, 6, 13) {real, imag} */,
  {32'h43d38843, 32'h00000000} /* (14, 6, 12) {real, imag} */,
  {32'h44a88592, 32'h00000000} /* (14, 6, 11) {real, imag} */,
  {32'h43b088c4, 32'h00000000} /* (14, 6, 10) {real, imag} */,
  {32'h44acf4fd, 32'h00000000} /* (14, 6, 9) {real, imag} */,
  {32'h43a38e34, 32'h00000000} /* (14, 6, 8) {real, imag} */,
  {32'h43ba7de2, 32'h00000000} /* (14, 6, 7) {real, imag} */,
  {32'h42d55cac, 32'h00000000} /* (14, 6, 6) {real, imag} */,
  {32'hc42524b1, 32'h00000000} /* (14, 6, 5) {real, imag} */,
  {32'hc334d10a, 32'h00000000} /* (14, 6, 4) {real, imag} */,
  {32'h43f0a23e, 32'h00000000} /* (14, 6, 3) {real, imag} */,
  {32'hc42543ad, 32'h00000000} /* (14, 6, 2) {real, imag} */,
  {32'hc21129a0, 32'h00000000} /* (14, 6, 1) {real, imag} */,
  {32'h43c40420, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h427cace2, 32'h00000000} /* (14, 5, 15) {real, imag} */,
  {32'h446f5e22, 32'h00000000} /* (14, 5, 14) {real, imag} */,
  {32'hc3fed396, 32'h00000000} /* (14, 5, 13) {real, imag} */,
  {32'hc409fd8c, 32'h00000000} /* (14, 5, 12) {real, imag} */,
  {32'h43f1b5d7, 32'h00000000} /* (14, 5, 11) {real, imag} */,
  {32'h440576db, 32'h00000000} /* (14, 5, 10) {real, imag} */,
  {32'h4417f197, 32'h00000000} /* (14, 5, 9) {real, imag} */,
  {32'h413dbfc0, 32'h00000000} /* (14, 5, 8) {real, imag} */,
  {32'h41f0ba2d, 32'h00000000} /* (14, 5, 7) {real, imag} */,
  {32'hc3b747b1, 32'h00000000} /* (14, 5, 6) {real, imag} */,
  {32'hc4522339, 32'h00000000} /* (14, 5, 5) {real, imag} */,
  {32'hc35d8f5f, 32'h00000000} /* (14, 5, 4) {real, imag} */,
  {32'h43c6495d, 32'h00000000} /* (14, 5, 3) {real, imag} */,
  {32'h426963c0, 32'h00000000} /* (14, 5, 2) {real, imag} */,
  {32'h447174a1, 32'h00000000} /* (14, 5, 1) {real, imag} */,
  {32'h4221e068, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'h42a25340, 32'h00000000} /* (14, 4, 15) {real, imag} */,
  {32'h42dd4750, 32'h00000000} /* (14, 4, 14) {real, imag} */,
  {32'hc3f8aac1, 32'h00000000} /* (14, 4, 13) {real, imag} */,
  {32'h43c170ef, 32'h00000000} /* (14, 4, 12) {real, imag} */,
  {32'h43be61a2, 32'h00000000} /* (14, 4, 11) {real, imag} */,
  {32'h43b9f5f1, 32'h00000000} /* (14, 4, 10) {real, imag} */,
  {32'h43184e46, 32'h00000000} /* (14, 4, 9) {real, imag} */,
  {32'h44260526, 32'h00000000} /* (14, 4, 8) {real, imag} */,
  {32'h42fa146c, 32'h00000000} /* (14, 4, 7) {real, imag} */,
  {32'hc3e959fc, 32'h00000000} /* (14, 4, 6) {real, imag} */,
  {32'hc4afd7e6, 32'h00000000} /* (14, 4, 5) {real, imag} */,
  {32'hc254e928, 32'h00000000} /* (14, 4, 4) {real, imag} */,
  {32'hc3bc677a, 32'h00000000} /* (14, 4, 3) {real, imag} */,
  {32'hc3f0dc81, 32'h00000000} /* (14, 4, 2) {real, imag} */,
  {32'h43d8a4a5, 32'h00000000} /* (14, 4, 1) {real, imag} */,
  {32'h4326b4c4, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'hc2c0f66c, 32'h00000000} /* (14, 3, 15) {real, imag} */,
  {32'h443039da, 32'h00000000} /* (14, 3, 14) {real, imag} */,
  {32'h44497428, 32'h00000000} /* (14, 3, 13) {real, imag} */,
  {32'h44952fae, 32'h00000000} /* (14, 3, 12) {real, imag} */,
  {32'h44866418, 32'h00000000} /* (14, 3, 11) {real, imag} */,
  {32'hc237c190, 32'h00000000} /* (14, 3, 10) {real, imag} */,
  {32'h438b0b81, 32'h00000000} /* (14, 3, 9) {real, imag} */,
  {32'hc38d69f5, 32'h00000000} /* (14, 3, 8) {real, imag} */,
  {32'hc44fa6f8, 32'h00000000} /* (14, 3, 7) {real, imag} */,
  {32'hc405c4dc, 32'h00000000} /* (14, 3, 6) {real, imag} */,
  {32'hc4467eda, 32'h00000000} /* (14, 3, 5) {real, imag} */,
  {32'hc4d5e42a, 32'h00000000} /* (14, 3, 4) {real, imag} */,
  {32'h4370a5cc, 32'h00000000} /* (14, 3, 3) {real, imag} */,
  {32'h42809048, 32'h00000000} /* (14, 3, 2) {real, imag} */,
  {32'hc2376610, 32'h00000000} /* (14, 3, 1) {real, imag} */,
  {32'h44a2e26d, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h445b0168, 32'h00000000} /* (14, 2, 15) {real, imag} */,
  {32'h447ec286, 32'h00000000} /* (14, 2, 14) {real, imag} */,
  {32'h447d6dfc, 32'h00000000} /* (14, 2, 13) {real, imag} */,
  {32'h449f4544, 32'h00000000} /* (14, 2, 12) {real, imag} */,
  {32'hc3949eb7, 32'h00000000} /* (14, 2, 11) {real, imag} */,
  {32'h44b88e15, 32'h00000000} /* (14, 2, 10) {real, imag} */,
  {32'hc3aff5ab, 32'h00000000} /* (14, 2, 9) {real, imag} */,
  {32'hc3e0890e, 32'h00000000} /* (14, 2, 8) {real, imag} */,
  {32'hc44a773a, 32'h00000000} /* (14, 2, 7) {real, imag} */,
  {32'hc483919d, 32'h00000000} /* (14, 2, 6) {real, imag} */,
  {32'hc5035d80, 32'h00000000} /* (14, 2, 5) {real, imag} */,
  {32'hc49b09c0, 32'h00000000} /* (14, 2, 4) {real, imag} */,
  {32'hc43dce1c, 32'h00000000} /* (14, 2, 3) {real, imag} */,
  {32'hc40bd9dc, 32'h00000000} /* (14, 2, 2) {real, imag} */,
  {32'hc40f5596, 32'h00000000} /* (14, 2, 1) {real, imag} */,
  {32'h43033cac, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h4388f88c, 32'h00000000} /* (14, 1, 15) {real, imag} */,
  {32'h43f2db60, 32'h00000000} /* (14, 1, 14) {real, imag} */,
  {32'h44063386, 32'h00000000} /* (14, 1, 13) {real, imag} */,
  {32'h44527dc9, 32'h00000000} /* (14, 1, 12) {real, imag} */,
  {32'hc3b0a96a, 32'h00000000} /* (14, 1, 11) {real, imag} */,
  {32'h430434d2, 32'h00000000} /* (14, 1, 10) {real, imag} */,
  {32'h4498547a, 32'h00000000} /* (14, 1, 9) {real, imag} */,
  {32'hc0bae120, 32'h00000000} /* (14, 1, 8) {real, imag} */,
  {32'hc49bb88b, 32'h00000000} /* (14, 1, 7) {real, imag} */,
  {32'hc4e1589a, 32'h00000000} /* (14, 1, 6) {real, imag} */,
  {32'hc4f3bd87, 32'h00000000} /* (14, 1, 5) {real, imag} */,
  {32'hc4be4008, 32'h00000000} /* (14, 1, 4) {real, imag} */,
  {32'hc453eaeb, 32'h00000000} /* (14, 1, 3) {real, imag} */,
  {32'hc3d77279, 32'h00000000} /* (14, 1, 2) {real, imag} */,
  {32'hc498004a, 32'h00000000} /* (14, 1, 1) {real, imag} */,
  {32'hc3c39e8e, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h41acc1e0, 32'h00000000} /* (14, 0, 15) {real, imag} */,
  {32'h43d9f2db, 32'h00000000} /* (14, 0, 14) {real, imag} */,
  {32'h43ecb58b, 32'h00000000} /* (14, 0, 13) {real, imag} */,
  {32'h441e7fbd, 32'h00000000} /* (14, 0, 12) {real, imag} */,
  {32'h4383d16c, 32'h00000000} /* (14, 0, 11) {real, imag} */,
  {32'hc4428386, 32'h00000000} /* (14, 0, 10) {real, imag} */,
  {32'hc32e4d60, 32'h00000000} /* (14, 0, 9) {real, imag} */,
  {32'h43aea49b, 32'h00000000} /* (14, 0, 8) {real, imag} */,
  {32'hc4972690, 32'h00000000} /* (14, 0, 7) {real, imag} */,
  {32'hc48bb3f1, 32'h00000000} /* (14, 0, 6) {real, imag} */,
  {32'hc435a9fb, 32'h00000000} /* (14, 0, 5) {real, imag} */,
  {32'hc3e63bae, 32'h00000000} /* (14, 0, 4) {real, imag} */,
  {32'hc3a830c4, 32'h00000000} /* (14, 0, 3) {real, imag} */,
  {32'hc32fbc8a, 32'h00000000} /* (14, 0, 2) {real, imag} */,
  {32'hc32c619c, 32'h00000000} /* (14, 0, 1) {real, imag} */,
  {32'h415824a0, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h42f6cf33, 32'h00000000} /* (13, 15, 15) {real, imag} */,
  {32'h434ed171, 32'h00000000} /* (13, 15, 14) {real, imag} */,
  {32'hc336fa1c, 32'h00000000} /* (13, 15, 13) {real, imag} */,
  {32'hc31f6fb0, 32'h00000000} /* (13, 15, 12) {real, imag} */,
  {32'h42dd1adb, 32'h00000000} /* (13, 15, 11) {real, imag} */,
  {32'hc485f62a, 32'h00000000} /* (13, 15, 10) {real, imag} */,
  {32'hc44f892f, 32'h00000000} /* (13, 15, 9) {real, imag} */,
  {32'hc40989f6, 32'h00000000} /* (13, 15, 8) {real, imag} */,
  {32'h4302eff0, 32'h00000000} /* (13, 15, 7) {real, imag} */,
  {32'hc40ccdec, 32'h00000000} /* (13, 15, 6) {real, imag} */,
  {32'hc35a0552, 32'h00000000} /* (13, 15, 5) {real, imag} */,
  {32'h40faa570, 32'h00000000} /* (13, 15, 4) {real, imag} */,
  {32'h427039ba, 32'h00000000} /* (13, 15, 3) {real, imag} */,
  {32'h4382023e, 32'h00000000} /* (13, 15, 2) {real, imag} */,
  {32'h43f9848e, 32'h00000000} /* (13, 15, 1) {real, imag} */,
  {32'h4480a779, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'h4394956a, 32'h00000000} /* (13, 14, 15) {real, imag} */,
  {32'hc3089b1c, 32'h00000000} /* (13, 14, 14) {real, imag} */,
  {32'hc40c4c5a, 32'h00000000} /* (13, 14, 13) {real, imag} */,
  {32'hc365e8dc, 32'h00000000} /* (13, 14, 12) {real, imag} */,
  {32'hc35d7644, 32'h00000000} /* (13, 14, 11) {real, imag} */,
  {32'hc4ab2a52, 32'h00000000} /* (13, 14, 10) {real, imag} */,
  {32'hc48dc80a, 32'h00000000} /* (13, 14, 9) {real, imag} */,
  {32'hc41996bd, 32'h00000000} /* (13, 14, 8) {real, imag} */,
  {32'h43811a82, 32'h00000000} /* (13, 14, 7) {real, imag} */,
  {32'hc2f8dfa8, 32'h00000000} /* (13, 14, 6) {real, imag} */,
  {32'hc39d036c, 32'h00000000} /* (13, 14, 5) {real, imag} */,
  {32'hc391963e, 32'h00000000} /* (13, 14, 4) {real, imag} */,
  {32'hc3a50cd6, 32'h00000000} /* (13, 14, 3) {real, imag} */,
  {32'hc48352be, 32'h00000000} /* (13, 14, 2) {real, imag} */,
  {32'hc3d43177, 32'h00000000} /* (13, 14, 1) {real, imag} */,
  {32'h444afc47, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'h43af3492, 32'h00000000} /* (13, 13, 15) {real, imag} */,
  {32'hc3e1857a, 32'h00000000} /* (13, 13, 14) {real, imag} */,
  {32'hc3db182a, 32'h00000000} /* (13, 13, 13) {real, imag} */,
  {32'hc3d22b52, 32'h00000000} /* (13, 13, 12) {real, imag} */,
  {32'hc2f5d926, 32'h00000000} /* (13, 13, 11) {real, imag} */,
  {32'hc3c9c100, 32'h00000000} /* (13, 13, 10) {real, imag} */,
  {32'h42b20734, 32'h00000000} /* (13, 13, 9) {real, imag} */,
  {32'hc40a69fc, 32'h00000000} /* (13, 13, 8) {real, imag} */,
  {32'hc41dd1cf, 32'h00000000} /* (13, 13, 7) {real, imag} */,
  {32'h440cc859, 32'h00000000} /* (13, 13, 6) {real, imag} */,
  {32'hc40b157a, 32'h00000000} /* (13, 13, 5) {real, imag} */,
  {32'hc3a1daa6, 32'h00000000} /* (13, 13, 4) {real, imag} */,
  {32'hc3d5cb8c, 32'h00000000} /* (13, 13, 3) {real, imag} */,
  {32'h4292704e, 32'h00000000} /* (13, 13, 2) {real, imag} */,
  {32'hc432fa24, 32'h00000000} /* (13, 13, 1) {real, imag} */,
  {32'hc2c8072c, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'h43f0f728, 32'h00000000} /* (13, 12, 15) {real, imag} */,
  {32'hc2f1dfc0, 32'h00000000} /* (13, 12, 14) {real, imag} */,
  {32'h4383b98e, 32'h00000000} /* (13, 12, 13) {real, imag} */,
  {32'h43d35fcf, 32'h00000000} /* (13, 12, 12) {real, imag} */,
  {32'hc280c634, 32'h00000000} /* (13, 12, 11) {real, imag} */,
  {32'h42d289f8, 32'h00000000} /* (13, 12, 10) {real, imag} */,
  {32'h448f69a6, 32'h00000000} /* (13, 12, 9) {real, imag} */,
  {32'h42efac96, 32'h00000000} /* (13, 12, 8) {real, imag} */,
  {32'hc4472812, 32'h00000000} /* (13, 12, 7) {real, imag} */,
  {32'hc3eb2590, 32'h00000000} /* (13, 12, 6) {real, imag} */,
  {32'h42852686, 32'h00000000} /* (13, 12, 5) {real, imag} */,
  {32'h41926480, 32'h00000000} /* (13, 12, 4) {real, imag} */,
  {32'hc385be2c, 32'h00000000} /* (13, 12, 3) {real, imag} */,
  {32'hc4761a17, 32'h00000000} /* (13, 12, 2) {real, imag} */,
  {32'h42d652f8, 32'h00000000} /* (13, 12, 1) {real, imag} */,
  {32'hc3b17796, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'h42a56966, 32'h00000000} /* (13, 11, 15) {real, imag} */,
  {32'h42887f50, 32'h00000000} /* (13, 11, 14) {real, imag} */,
  {32'h4394752c, 32'h00000000} /* (13, 11, 13) {real, imag} */,
  {32'h41923e18, 32'h00000000} /* (13, 11, 12) {real, imag} */,
  {32'h44290f99, 32'h00000000} /* (13, 11, 11) {real, imag} */,
  {32'hc181a7a0, 32'h00000000} /* (13, 11, 10) {real, imag} */,
  {32'h43a990bc, 32'h00000000} /* (13, 11, 9) {real, imag} */,
  {32'h4456e00c, 32'h00000000} /* (13, 11, 8) {real, imag} */,
  {32'hc3734a4d, 32'h00000000} /* (13, 11, 7) {real, imag} */,
  {32'hc4a3f718, 32'h00000000} /* (13, 11, 6) {real, imag} */,
  {32'hc4076483, 32'h00000000} /* (13, 11, 5) {real, imag} */,
  {32'h4269398c, 32'h00000000} /* (13, 11, 4) {real, imag} */,
  {32'hc3c1d0b6, 32'h00000000} /* (13, 11, 3) {real, imag} */,
  {32'hc46e38e9, 32'h00000000} /* (13, 11, 2) {real, imag} */,
  {32'h40af8400, 32'h00000000} /* (13, 11, 1) {real, imag} */,
  {32'h41068d80, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'hc1c687a0, 32'h00000000} /* (13, 10, 15) {real, imag} */,
  {32'hc3a4f27e, 32'h00000000} /* (13, 10, 14) {real, imag} */,
  {32'h440c7578, 32'h00000000} /* (13, 10, 13) {real, imag} */,
  {32'h448d8d7a, 32'h00000000} /* (13, 10, 12) {real, imag} */,
  {32'h4449b74b, 32'h00000000} /* (13, 10, 11) {real, imag} */,
  {32'hc3c8e171, 32'h00000000} /* (13, 10, 10) {real, imag} */,
  {32'h43b42ada, 32'h00000000} /* (13, 10, 9) {real, imag} */,
  {32'hc3b0a4ec, 32'h00000000} /* (13, 10, 8) {real, imag} */,
  {32'h431bdcd4, 32'h00000000} /* (13, 10, 7) {real, imag} */,
  {32'h43c451a4, 32'h00000000} /* (13, 10, 6) {real, imag} */,
  {32'hc40c53da, 32'h00000000} /* (13, 10, 5) {real, imag} */,
  {32'hc3c3a7aa, 32'h00000000} /* (13, 10, 4) {real, imag} */,
  {32'h442925dd, 32'h00000000} /* (13, 10, 3) {real, imag} */,
  {32'hc3dbf967, 32'h00000000} /* (13, 10, 2) {real, imag} */,
  {32'h42bc976e, 32'h00000000} /* (13, 10, 1) {real, imag} */,
  {32'h443ed7dc, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h448787b2, 32'h00000000} /* (13, 9, 15) {real, imag} */,
  {32'h44c0628c, 32'h00000000} /* (13, 9, 14) {real, imag} */,
  {32'h4306dd2e, 32'h00000000} /* (13, 9, 13) {real, imag} */,
  {32'h444391fe, 32'h00000000} /* (13, 9, 12) {real, imag} */,
  {32'h437c0540, 32'h00000000} /* (13, 9, 11) {real, imag} */,
  {32'h441d5fb1, 32'h00000000} /* (13, 9, 10) {real, imag} */,
  {32'hc38bcae3, 32'h00000000} /* (13, 9, 9) {real, imag} */,
  {32'hc3acf6ac, 32'h00000000} /* (13, 9, 8) {real, imag} */,
  {32'hc3aa5132, 32'h00000000} /* (13, 9, 7) {real, imag} */,
  {32'hc39ae912, 32'h00000000} /* (13, 9, 6) {real, imag} */,
  {32'h43b96eb9, 32'h00000000} /* (13, 9, 5) {real, imag} */,
  {32'hc3571760, 32'h00000000} /* (13, 9, 4) {real, imag} */,
  {32'hc1462e00, 32'h00000000} /* (13, 9, 3) {real, imag} */,
  {32'h43a86ec0, 32'h00000000} /* (13, 9, 2) {real, imag} */,
  {32'hc35be1c2, 32'h00000000} /* (13, 9, 1) {real, imag} */,
  {32'h4326dee9, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'hc328808e, 32'h00000000} /* (13, 8, 15) {real, imag} */,
  {32'h414a88c0, 32'h00000000} /* (13, 8, 14) {real, imag} */,
  {32'h4359d507, 32'h00000000} /* (13, 8, 13) {real, imag} */,
  {32'h43d1828a, 32'h00000000} /* (13, 8, 12) {real, imag} */,
  {32'h4429fe0b, 32'h00000000} /* (13, 8, 11) {real, imag} */,
  {32'h435bfaaa, 32'h00000000} /* (13, 8, 10) {real, imag} */,
  {32'h439b079a, 32'h00000000} /* (13, 8, 9) {real, imag} */,
  {32'h435aa30f, 32'h00000000} /* (13, 8, 8) {real, imag} */,
  {32'hc270b486, 32'h00000000} /* (13, 8, 7) {real, imag} */,
  {32'hc44ce737, 32'h00000000} /* (13, 8, 6) {real, imag} */,
  {32'hc3aa8c12, 32'h00000000} /* (13, 8, 5) {real, imag} */,
  {32'hc34b692f, 32'h00000000} /* (13, 8, 4) {real, imag} */,
  {32'hc447d0e5, 32'h00000000} /* (13, 8, 3) {real, imag} */,
  {32'h43cbae4f, 32'h00000000} /* (13, 8, 2) {real, imag} */,
  {32'hc3932da2, 32'h00000000} /* (13, 8, 1) {real, imag} */,
  {32'hc4250cad, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'hc3f02076, 32'h00000000} /* (13, 7, 15) {real, imag} */,
  {32'hc4338aba, 32'h00000000} /* (13, 7, 14) {real, imag} */,
  {32'hc40379d6, 32'h00000000} /* (13, 7, 13) {real, imag} */,
  {32'h449390af, 32'h00000000} /* (13, 7, 12) {real, imag} */,
  {32'h44818e70, 32'h00000000} /* (13, 7, 11) {real, imag} */,
  {32'h4398bbfc, 32'h00000000} /* (13, 7, 10) {real, imag} */,
  {32'h441ac6de, 32'h00000000} /* (13, 7, 9) {real, imag} */,
  {32'h443b3516, 32'h00000000} /* (13, 7, 8) {real, imag} */,
  {32'hc221bed4, 32'h00000000} /* (13, 7, 7) {real, imag} */,
  {32'h44300f76, 32'h00000000} /* (13, 7, 6) {real, imag} */,
  {32'hc3978180, 32'h00000000} /* (13, 7, 5) {real, imag} */,
  {32'h42d382b0, 32'h00000000} /* (13, 7, 4) {real, imag} */,
  {32'h444c17cd, 32'h00000000} /* (13, 7, 3) {real, imag} */,
  {32'h43f216aa, 32'h00000000} /* (13, 7, 2) {real, imag} */,
  {32'h440bede6, 32'h00000000} /* (13, 7, 1) {real, imag} */,
  {32'hc478fa6a, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'hc36f9c50, 32'h00000000} /* (13, 6, 15) {real, imag} */,
  {32'hc33f96ce, 32'h00000000} /* (13, 6, 14) {real, imag} */,
  {32'hc3642d9a, 32'h00000000} /* (13, 6, 13) {real, imag} */,
  {32'h43b4b8e0, 32'h00000000} /* (13, 6, 12) {real, imag} */,
  {32'hc3997a30, 32'h00000000} /* (13, 6, 11) {real, imag} */,
  {32'h44c94a2a, 32'h00000000} /* (13, 6, 10) {real, imag} */,
  {32'h44a5fe80, 32'h00000000} /* (13, 6, 9) {real, imag} */,
  {32'hc34c31db, 32'h00000000} /* (13, 6, 8) {real, imag} */,
  {32'h44dbfc9c, 32'h00000000} /* (13, 6, 7) {real, imag} */,
  {32'h4393c18d, 32'h00000000} /* (13, 6, 6) {real, imag} */,
  {32'h43af9d0b, 32'h00000000} /* (13, 6, 5) {real, imag} */,
  {32'hc4395ce4, 32'h00000000} /* (13, 6, 4) {real, imag} */,
  {32'h4288ee50, 32'h00000000} /* (13, 6, 3) {real, imag} */,
  {32'h43e6ce22, 32'h00000000} /* (13, 6, 2) {real, imag} */,
  {32'hc38572aa, 32'h00000000} /* (13, 6, 1) {real, imag} */,
  {32'h438dd5c8, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'h435777da, 32'h00000000} /* (13, 5, 15) {real, imag} */,
  {32'h3e7ae000, 32'h00000000} /* (13, 5, 14) {real, imag} */,
  {32'h431ce042, 32'h00000000} /* (13, 5, 13) {real, imag} */,
  {32'hc3188984, 32'h00000000} /* (13, 5, 12) {real, imag} */,
  {32'h437172f5, 32'h00000000} /* (13, 5, 11) {real, imag} */,
  {32'h43b32886, 32'h00000000} /* (13, 5, 10) {real, imag} */,
  {32'h43ecafb4, 32'h00000000} /* (13, 5, 9) {real, imag} */,
  {32'h4358e081, 32'h00000000} /* (13, 5, 8) {real, imag} */,
  {32'h43c26bbd, 32'h00000000} /* (13, 5, 7) {real, imag} */,
  {32'h443d2001, 32'h00000000} /* (13, 5, 6) {real, imag} */,
  {32'h43802ab1, 32'h00000000} /* (13, 5, 5) {real, imag} */,
  {32'h4488cf6e, 32'h00000000} /* (13, 5, 4) {real, imag} */,
  {32'h44380936, 32'h00000000} /* (13, 5, 3) {real, imag} */,
  {32'h440f794c, 32'h00000000} /* (13, 5, 2) {real, imag} */,
  {32'hc23c8780, 32'h00000000} /* (13, 5, 1) {real, imag} */,
  {32'hc0c67220, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h43f76544, 32'h00000000} /* (13, 4, 15) {real, imag} */,
  {32'h4419a474, 32'h00000000} /* (13, 4, 14) {real, imag} */,
  {32'h43a84bf0, 32'h00000000} /* (13, 4, 13) {real, imag} */,
  {32'h445b2deb, 32'h00000000} /* (13, 4, 12) {real, imag} */,
  {32'hc3a95ef8, 32'h00000000} /* (13, 4, 11) {real, imag} */,
  {32'h4308d12b, 32'h00000000} /* (13, 4, 10) {real, imag} */,
  {32'h43a264dc, 32'h00000000} /* (13, 4, 9) {real, imag} */,
  {32'h44598575, 32'h00000000} /* (13, 4, 8) {real, imag} */,
  {32'h43873b80, 32'h00000000} /* (13, 4, 7) {real, imag} */,
  {32'h4393c1ec, 32'h00000000} /* (13, 4, 6) {real, imag} */,
  {32'hc45c928a, 32'h00000000} /* (13, 4, 5) {real, imag} */,
  {32'hc428e59d, 32'h00000000} /* (13, 4, 4) {real, imag} */,
  {32'h444caec2, 32'h00000000} /* (13, 4, 3) {real, imag} */,
  {32'hc3314721, 32'h00000000} /* (13, 4, 2) {real, imag} */,
  {32'h440fc184, 32'h00000000} /* (13, 4, 1) {real, imag} */,
  {32'h43a5420a, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'hc2a52b0c, 32'h00000000} /* (13, 3, 15) {real, imag} */,
  {32'hc41e938e, 32'h00000000} /* (13, 3, 14) {real, imag} */,
  {32'h44f710c4, 32'h00000000} /* (13, 3, 13) {real, imag} */,
  {32'h44f323c8, 32'h00000000} /* (13, 3, 12) {real, imag} */,
  {32'h444d4c5d, 32'h00000000} /* (13, 3, 11) {real, imag} */,
  {32'hc332180a, 32'h00000000} /* (13, 3, 10) {real, imag} */,
  {32'h42a9fd60, 32'h00000000} /* (13, 3, 9) {real, imag} */,
  {32'h44b59e3c, 32'h00000000} /* (13, 3, 8) {real, imag} */,
  {32'h4436f7f0, 32'h00000000} /* (13, 3, 7) {real, imag} */,
  {32'hc4930413, 32'h00000000} /* (13, 3, 6) {real, imag} */,
  {32'hc417b524, 32'h00000000} /* (13, 3, 5) {real, imag} */,
  {32'hc42cce04, 32'h00000000} /* (13, 3, 4) {real, imag} */,
  {32'h441c7661, 32'h00000000} /* (13, 3, 3) {real, imag} */,
  {32'h4380fbe1, 32'h00000000} /* (13, 3, 2) {real, imag} */,
  {32'hc3baab82, 32'h00000000} /* (13, 3, 1) {real, imag} */,
  {32'h442471c4, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h4419531f, 32'h00000000} /* (13, 2, 15) {real, imag} */,
  {32'h4481b192, 32'h00000000} /* (13, 2, 14) {real, imag} */,
  {32'h4486d5fc, 32'h00000000} /* (13, 2, 13) {real, imag} */,
  {32'h449ab81c, 32'h00000000} /* (13, 2, 12) {real, imag} */,
  {32'h43d38bfa, 32'h00000000} /* (13, 2, 11) {real, imag} */,
  {32'hc4608262, 32'h00000000} /* (13, 2, 10) {real, imag} */,
  {32'hc2f3067c, 32'h00000000} /* (13, 2, 9) {real, imag} */,
  {32'hc3e1906b, 32'h00000000} /* (13, 2, 8) {real, imag} */,
  {32'h43cc47b4, 32'h00000000} /* (13, 2, 7) {real, imag} */,
  {32'hc424822d, 32'h00000000} /* (13, 2, 6) {real, imag} */,
  {32'hc48b1782, 32'h00000000} /* (13, 2, 5) {real, imag} */,
  {32'hc3b3ff81, 32'h00000000} /* (13, 2, 4) {real, imag} */,
  {32'h42d4dcb2, 32'h00000000} /* (13, 2, 3) {real, imag} */,
  {32'h42b520dc, 32'h00000000} /* (13, 2, 2) {real, imag} */,
  {32'h42f59c14, 32'h00000000} /* (13, 2, 1) {real, imag} */,
  {32'h42d628b4, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h44222c7c, 32'h00000000} /* (13, 1, 15) {real, imag} */,
  {32'h4426662d, 32'h00000000} /* (13, 1, 14) {real, imag} */,
  {32'h44b676fc, 32'h00000000} /* (13, 1, 13) {real, imag} */,
  {32'h44721b12, 32'h00000000} /* (13, 1, 12) {real, imag} */,
  {32'hc440670a, 32'h00000000} /* (13, 1, 11) {real, imag} */,
  {32'hc3b20e50, 32'h00000000} /* (13, 1, 10) {real, imag} */,
  {32'h442d91d3, 32'h00000000} /* (13, 1, 9) {real, imag} */,
  {32'hc2ac05f2, 32'h00000000} /* (13, 1, 8) {real, imag} */,
  {32'hc4822edb, 32'h00000000} /* (13, 1, 7) {real, imag} */,
  {32'hc42c025f, 32'h00000000} /* (13, 1, 6) {real, imag} */,
  {32'hc2a46cd8, 32'h00000000} /* (13, 1, 5) {real, imag} */,
  {32'hc48ba4e1, 32'h00000000} /* (13, 1, 4) {real, imag} */,
  {32'hc4881c1b, 32'h00000000} /* (13, 1, 3) {real, imag} */,
  {32'hc2f77fce, 32'h00000000} /* (13, 1, 2) {real, imag} */,
  {32'h4292ade8, 32'h00000000} /* (13, 1, 1) {real, imag} */,
  {32'hc10f8710, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h4337e90c, 32'h00000000} /* (13, 0, 15) {real, imag} */,
  {32'h42b52bb8, 32'h00000000} /* (13, 0, 14) {real, imag} */,
  {32'h448f9d92, 32'h00000000} /* (13, 0, 13) {real, imag} */,
  {32'h4429c844, 32'h00000000} /* (13, 0, 12) {real, imag} */,
  {32'hc3b2104d, 32'h00000000} /* (13, 0, 11) {real, imag} */,
  {32'hc32d661d, 32'h00000000} /* (13, 0, 10) {real, imag} */,
  {32'h4349ba9a, 32'h00000000} /* (13, 0, 9) {real, imag} */,
  {32'h43f09c06, 32'h00000000} /* (13, 0, 8) {real, imag} */,
  {32'hc3dca6e2, 32'h00000000} /* (13, 0, 7) {real, imag} */,
  {32'hc3cb3916, 32'h00000000} /* (13, 0, 6) {real, imag} */,
  {32'h42b76400, 32'h00000000} /* (13, 0, 5) {real, imag} */,
  {32'hc23d4e28, 32'h00000000} /* (13, 0, 4) {real, imag} */,
  {32'h4308ab30, 32'h00000000} /* (13, 0, 3) {real, imag} */,
  {32'hc34c2f2f, 32'h00000000} /* (13, 0, 2) {real, imag} */,
  {32'hc15a88a0, 32'h00000000} /* (13, 0, 1) {real, imag} */,
  {32'h4337c49c, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h43e69c4c, 32'h00000000} /* (12, 15, 15) {real, imag} */,
  {32'h438192af, 32'h00000000} /* (12, 15, 14) {real, imag} */,
  {32'hc3a3df78, 32'h00000000} /* (12, 15, 13) {real, imag} */,
  {32'h4384b737, 32'h00000000} /* (12, 15, 12) {real, imag} */,
  {32'h42cb6bec, 32'h00000000} /* (12, 15, 11) {real, imag} */,
  {32'hc4492dc5, 32'h00000000} /* (12, 15, 10) {real, imag} */,
  {32'hc40032b6, 32'h00000000} /* (12, 15, 9) {real, imag} */,
  {32'hc41802cc, 32'h00000000} /* (12, 15, 8) {real, imag} */,
  {32'hc38765fc, 32'h00000000} /* (12, 15, 7) {real, imag} */,
  {32'h419f39d0, 32'h00000000} /* (12, 15, 6) {real, imag} */,
  {32'hc25fbf7c, 32'h00000000} /* (12, 15, 5) {real, imag} */,
  {32'h43f0890b, 32'h00000000} /* (12, 15, 4) {real, imag} */,
  {32'h44661d64, 32'h00000000} /* (12, 15, 3) {real, imag} */,
  {32'h43a9a976, 32'h00000000} /* (12, 15, 2) {real, imag} */,
  {32'hc33bfc51, 32'h00000000} /* (12, 15, 1) {real, imag} */,
  {32'h430235e2, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'h442546e8, 32'h00000000} /* (12, 14, 15) {real, imag} */,
  {32'hc21f58c8, 32'h00000000} /* (12, 14, 14) {real, imag} */,
  {32'hc42b5d81, 32'h00000000} /* (12, 14, 13) {real, imag} */,
  {32'hc4131f0b, 32'h00000000} /* (12, 14, 12) {real, imag} */,
  {32'hc2b0b332, 32'h00000000} /* (12, 14, 11) {real, imag} */,
  {32'hc4faaf52, 32'h00000000} /* (12, 14, 10) {real, imag} */,
  {32'hc3b8fa9f, 32'h00000000} /* (12, 14, 9) {real, imag} */,
  {32'hc4013126, 32'h00000000} /* (12, 14, 8) {real, imag} */,
  {32'h43cb721b, 32'h00000000} /* (12, 14, 7) {real, imag} */,
  {32'h4444dad0, 32'h00000000} /* (12, 14, 6) {real, imag} */,
  {32'hc32666f4, 32'h00000000} /* (12, 14, 5) {real, imag} */,
  {32'h44183671, 32'h00000000} /* (12, 14, 4) {real, imag} */,
  {32'h44074dc1, 32'h00000000} /* (12, 14, 3) {real, imag} */,
  {32'h43a28040, 32'h00000000} /* (12, 14, 2) {real, imag} */,
  {32'h4390adc1, 32'h00000000} /* (12, 14, 1) {real, imag} */,
  {32'hc37d266e, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'h44246460, 32'h00000000} /* (12, 13, 15) {real, imag} */,
  {32'h42da42b4, 32'h00000000} /* (12, 13, 14) {real, imag} */,
  {32'h43ba793b, 32'h00000000} /* (12, 13, 13) {real, imag} */,
  {32'hc4295bb2, 32'h00000000} /* (12, 13, 12) {real, imag} */,
  {32'hc1af51d0, 32'h00000000} /* (12, 13, 11) {real, imag} */,
  {32'h43a34585, 32'h00000000} /* (12, 13, 10) {real, imag} */,
  {32'hc2653da7, 32'h00000000} /* (12, 13, 9) {real, imag} */,
  {32'hc23a9fa4, 32'h00000000} /* (12, 13, 8) {real, imag} */,
  {32'hc34a5202, 32'h00000000} /* (12, 13, 7) {real, imag} */,
  {32'h43a1a779, 32'h00000000} /* (12, 13, 6) {real, imag} */,
  {32'h440c9f4c, 32'h00000000} /* (12, 13, 5) {real, imag} */,
  {32'h442f3868, 32'h00000000} /* (12, 13, 4) {real, imag} */,
  {32'hc2d1461c, 32'h00000000} /* (12, 13, 3) {real, imag} */,
  {32'hc334cc7a, 32'h00000000} /* (12, 13, 2) {real, imag} */,
  {32'h42239457, 32'h00000000} /* (12, 13, 1) {real, imag} */,
  {32'h433b059d, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'h441dd190, 32'h00000000} /* (12, 12, 15) {real, imag} */,
  {32'h44927882, 32'h00000000} /* (12, 12, 14) {real, imag} */,
  {32'hc3c9a397, 32'h00000000} /* (12, 12, 13) {real, imag} */,
  {32'h43e74191, 32'h00000000} /* (12, 12, 12) {real, imag} */,
  {32'h42fb039b, 32'h00000000} /* (12, 12, 11) {real, imag} */,
  {32'h43dbe350, 32'h00000000} /* (12, 12, 10) {real, imag} */,
  {32'h441ccd88, 32'h00000000} /* (12, 12, 9) {real, imag} */,
  {32'hc25ed5d4, 32'h00000000} /* (12, 12, 8) {real, imag} */,
  {32'hc3e9a17d, 32'h00000000} /* (12, 12, 7) {real, imag} */,
  {32'hc37ee284, 32'h00000000} /* (12, 12, 6) {real, imag} */,
  {32'h44258212, 32'h00000000} /* (12, 12, 5) {real, imag} */,
  {32'h430bc1aa, 32'h00000000} /* (12, 12, 4) {real, imag} */,
  {32'h41d6736c, 32'h00000000} /* (12, 12, 3) {real, imag} */,
  {32'hc467b318, 32'h00000000} /* (12, 12, 2) {real, imag} */,
  {32'hc3156b96, 32'h00000000} /* (12, 12, 1) {real, imag} */,
  {32'h43fd9226, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'h43b479ef, 32'h00000000} /* (12, 11, 15) {real, imag} */,
  {32'hc2d85499, 32'h00000000} /* (12, 11, 14) {real, imag} */,
  {32'h4385dd46, 32'h00000000} /* (12, 11, 13) {real, imag} */,
  {32'h447fe28f, 32'h00000000} /* (12, 11, 12) {real, imag} */,
  {32'h44654b1b, 32'h00000000} /* (12, 11, 11) {real, imag} */,
  {32'h43743001, 32'h00000000} /* (12, 11, 10) {real, imag} */,
  {32'h445b53ab, 32'h00000000} /* (12, 11, 9) {real, imag} */,
  {32'h4459e2bc, 32'h00000000} /* (12, 11, 8) {real, imag} */,
  {32'h4487f307, 32'h00000000} /* (12, 11, 7) {real, imag} */,
  {32'h4113b988, 32'h00000000} /* (12, 11, 6) {real, imag} */,
  {32'h42f4c4ce, 32'h00000000} /* (12, 11, 5) {real, imag} */,
  {32'hc3e40cd2, 32'h00000000} /* (12, 11, 4) {real, imag} */,
  {32'hc218e190, 32'h00000000} /* (12, 11, 3) {real, imag} */,
  {32'h4429ba4a, 32'h00000000} /* (12, 11, 2) {real, imag} */,
  {32'h43762ea4, 32'h00000000} /* (12, 11, 1) {real, imag} */,
  {32'h43ebd474, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'h442880e2, 32'h00000000} /* (12, 10, 15) {real, imag} */,
  {32'hc3536514, 32'h00000000} /* (12, 10, 14) {real, imag} */,
  {32'h43ac6682, 32'h00000000} /* (12, 10, 13) {real, imag} */,
  {32'h444f67bd, 32'h00000000} /* (12, 10, 12) {real, imag} */,
  {32'h447eafd9, 32'h00000000} /* (12, 10, 11) {real, imag} */,
  {32'h4480785a, 32'h00000000} /* (12, 10, 10) {real, imag} */,
  {32'h43c370d6, 32'h00000000} /* (12, 10, 9) {real, imag} */,
  {32'h441ae92e, 32'h00000000} /* (12, 10, 8) {real, imag} */,
  {32'h4371f0d1, 32'h00000000} /* (12, 10, 7) {real, imag} */,
  {32'h4403a18a, 32'h00000000} /* (12, 10, 6) {real, imag} */,
  {32'hc4831014, 32'h00000000} /* (12, 10, 5) {real, imag} */,
  {32'hc349099c, 32'h00000000} /* (12, 10, 4) {real, imag} */,
  {32'hc298a818, 32'h00000000} /* (12, 10, 3) {real, imag} */,
  {32'h4383a342, 32'h00000000} /* (12, 10, 2) {real, imag} */,
  {32'h43e50b82, 32'h00000000} /* (12, 10, 1) {real, imag} */,
  {32'h43b8f883, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h43a643c4, 32'h00000000} /* (12, 9, 15) {real, imag} */,
  {32'h41c2a350, 32'h00000000} /* (12, 9, 14) {real, imag} */,
  {32'h439ae6e5, 32'h00000000} /* (12, 9, 13) {real, imag} */,
  {32'h443e72ec, 32'h00000000} /* (12, 9, 12) {real, imag} */,
  {32'h4496cb9e, 32'h00000000} /* (12, 9, 11) {real, imag} */,
  {32'h43ecce2a, 32'h00000000} /* (12, 9, 10) {real, imag} */,
  {32'h43e4dbca, 32'h00000000} /* (12, 9, 9) {real, imag} */,
  {32'hc4845580, 32'h00000000} /* (12, 9, 8) {real, imag} */,
  {32'h43370299, 32'h00000000} /* (12, 9, 7) {real, imag} */,
  {32'hc383fdcd, 32'h00000000} /* (12, 9, 6) {real, imag} */,
  {32'hc47ce746, 32'h00000000} /* (12, 9, 5) {real, imag} */,
  {32'hc418a160, 32'h00000000} /* (12, 9, 4) {real, imag} */,
  {32'hc40fc2cb, 32'h00000000} /* (12, 9, 3) {real, imag} */,
  {32'h43cc7cfa, 32'h00000000} /* (12, 9, 2) {real, imag} */,
  {32'h446b09d7, 32'h00000000} /* (12, 9, 1) {real, imag} */,
  {32'h43d23920, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'h42c0aa5f, 32'h00000000} /* (12, 8, 15) {real, imag} */,
  {32'h43f82b9e, 32'h00000000} /* (12, 8, 14) {real, imag} */,
  {32'h431b98d4, 32'h00000000} /* (12, 8, 13) {real, imag} */,
  {32'hc334d396, 32'h00000000} /* (12, 8, 12) {real, imag} */,
  {32'h436db38d, 32'h00000000} /* (12, 8, 11) {real, imag} */,
  {32'h43167dfd, 32'h00000000} /* (12, 8, 10) {real, imag} */,
  {32'h43c0f76e, 32'h00000000} /* (12, 8, 9) {real, imag} */,
  {32'h43e6907f, 32'h00000000} /* (12, 8, 8) {real, imag} */,
  {32'hc2e1cbdb, 32'h00000000} /* (12, 8, 7) {real, imag} */,
  {32'hc24c7230, 32'h00000000} /* (12, 8, 6) {real, imag} */,
  {32'hc4ac7086, 32'h00000000} /* (12, 8, 5) {real, imag} */,
  {32'hc450d23c, 32'h00000000} /* (12, 8, 4) {real, imag} */,
  {32'hc421bd76, 32'h00000000} /* (12, 8, 3) {real, imag} */,
  {32'hc3b3822e, 32'h00000000} /* (12, 8, 2) {real, imag} */,
  {32'h43f67c3a, 32'h00000000} /* (12, 8, 1) {real, imag} */,
  {32'h4354735e, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'hc4858d14, 32'h00000000} /* (12, 7, 15) {real, imag} */,
  {32'hc469e72b, 32'h00000000} /* (12, 7, 14) {real, imag} */,
  {32'hc3026430, 32'h00000000} /* (12, 7, 13) {real, imag} */,
  {32'hc28eec34, 32'h00000000} /* (12, 7, 12) {real, imag} */,
  {32'h44329bca, 32'h00000000} /* (12, 7, 11) {real, imag} */,
  {32'h43f6422a, 32'h00000000} /* (12, 7, 10) {real, imag} */,
  {32'h43e2a3cb, 32'h00000000} /* (12, 7, 9) {real, imag} */,
  {32'h44577d2c, 32'h00000000} /* (12, 7, 8) {real, imag} */,
  {32'h4377b30c, 32'h00000000} /* (12, 7, 7) {real, imag} */,
  {32'h43c5a3a6, 32'h00000000} /* (12, 7, 6) {real, imag} */,
  {32'hc396995e, 32'h00000000} /* (12, 7, 5) {real, imag} */,
  {32'hc40e9876, 32'h00000000} /* (12, 7, 4) {real, imag} */,
  {32'hc22c61c0, 32'h00000000} /* (12, 7, 3) {real, imag} */,
  {32'h421624f0, 32'h00000000} /* (12, 7, 2) {real, imag} */,
  {32'hc385d3eb, 32'h00000000} /* (12, 7, 1) {real, imag} */,
  {32'hc2df5da8, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'hc487f4f9, 32'h00000000} /* (12, 6, 15) {real, imag} */,
  {32'hc3f3b334, 32'h00000000} /* (12, 6, 14) {real, imag} */,
  {32'hc21abc60, 32'h00000000} /* (12, 6, 13) {real, imag} */,
  {32'hc3c4eac2, 32'h00000000} /* (12, 6, 12) {real, imag} */,
  {32'h442fee15, 32'h00000000} /* (12, 6, 11) {real, imag} */,
  {32'h42cd5f96, 32'h00000000} /* (12, 6, 10) {real, imag} */,
  {32'h442dd4e6, 32'h00000000} /* (12, 6, 9) {real, imag} */,
  {32'h44227912, 32'h00000000} /* (12, 6, 8) {real, imag} */,
  {32'h449184eb, 32'h00000000} /* (12, 6, 7) {real, imag} */,
  {32'h441aca7a, 32'h00000000} /* (12, 6, 6) {real, imag} */,
  {32'h44d84519, 32'h00000000} /* (12, 6, 5) {real, imag} */,
  {32'h449b0836, 32'h00000000} /* (12, 6, 4) {real, imag} */,
  {32'h43363ec4, 32'h00000000} /* (12, 6, 3) {real, imag} */,
  {32'hc3b5fea4, 32'h00000000} /* (12, 6, 2) {real, imag} */,
  {32'hc4a95773, 32'h00000000} /* (12, 6, 1) {real, imag} */,
  {32'h42edc3e0, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'h430973fe, 32'h00000000} /* (12, 5, 15) {real, imag} */,
  {32'h440085ca, 32'h00000000} /* (12, 5, 14) {real, imag} */,
  {32'h41c26154, 32'h00000000} /* (12, 5, 13) {real, imag} */,
  {32'h42c91ce0, 32'h00000000} /* (12, 5, 12) {real, imag} */,
  {32'hc416ec08, 32'h00000000} /* (12, 5, 11) {real, imag} */,
  {32'hc332d23e, 32'h00000000} /* (12, 5, 10) {real, imag} */,
  {32'h444e1eaa, 32'h00000000} /* (12, 5, 9) {real, imag} */,
  {32'hc4355c90, 32'h00000000} /* (12, 5, 8) {real, imag} */,
  {32'h448e38d8, 32'h00000000} /* (12, 5, 7) {real, imag} */,
  {32'h44a105f5, 32'h00000000} /* (12, 5, 6) {real, imag} */,
  {32'h435bcc78, 32'h00000000} /* (12, 5, 5) {real, imag} */,
  {32'h4424b328, 32'h00000000} /* (12, 5, 4) {real, imag} */,
  {32'h443a7492, 32'h00000000} /* (12, 5, 3) {real, imag} */,
  {32'h43c0843f, 32'h00000000} /* (12, 5, 2) {real, imag} */,
  {32'hc2993e08, 32'h00000000} /* (12, 5, 1) {real, imag} */,
  {32'hc106fca0, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'h43a26f6b, 32'h00000000} /* (12, 4, 15) {real, imag} */,
  {32'h42fe4e43, 32'h00000000} /* (12, 4, 14) {real, imag} */,
  {32'h43a94322, 32'h00000000} /* (12, 4, 13) {real, imag} */,
  {32'h44a52dc8, 32'h00000000} /* (12, 4, 12) {real, imag} */,
  {32'hc2fd3bf0, 32'h00000000} /* (12, 4, 11) {real, imag} */,
  {32'hc37676b7, 32'h00000000} /* (12, 4, 10) {real, imag} */,
  {32'hc3211c3a, 32'h00000000} /* (12, 4, 9) {real, imag} */,
  {32'h43e56024, 32'h00000000} /* (12, 4, 8) {real, imag} */,
  {32'h445d58ca, 32'h00000000} /* (12, 4, 7) {real, imag} */,
  {32'h4395d3b6, 32'h00000000} /* (12, 4, 6) {real, imag} */,
  {32'h44897030, 32'h00000000} /* (12, 4, 5) {real, imag} */,
  {32'h442678a7, 32'h00000000} /* (12, 4, 4) {real, imag} */,
  {32'h44179f6d, 32'h00000000} /* (12, 4, 3) {real, imag} */,
  {32'h4419b6db, 32'h00000000} /* (12, 4, 2) {real, imag} */,
  {32'h43843005, 32'h00000000} /* (12, 4, 1) {real, imag} */,
  {32'h427edd2c, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'h43c3c3b6, 32'h00000000} /* (12, 3, 15) {real, imag} */,
  {32'h43f6d4fe, 32'h00000000} /* (12, 3, 14) {real, imag} */,
  {32'h43ea7cf2, 32'h00000000} /* (12, 3, 13) {real, imag} */,
  {32'h448a0041, 32'h00000000} /* (12, 3, 12) {real, imag} */,
  {32'h43620787, 32'h00000000} /* (12, 3, 11) {real, imag} */,
  {32'h43f7f742, 32'h00000000} /* (12, 3, 10) {real, imag} */,
  {32'h423a008c, 32'h00000000} /* (12, 3, 9) {real, imag} */,
  {32'h434cc362, 32'h00000000} /* (12, 3, 8) {real, imag} */,
  {32'h4423cb0f, 32'h00000000} /* (12, 3, 7) {real, imag} */,
  {32'h448785d0, 32'h00000000} /* (12, 3, 6) {real, imag} */,
  {32'hc38089a8, 32'h00000000} /* (12, 3, 5) {real, imag} */,
  {32'h4405b900, 32'h00000000} /* (12, 3, 4) {real, imag} */,
  {32'h430c5873, 32'h00000000} /* (12, 3, 3) {real, imag} */,
  {32'hc439f3bb, 32'h00000000} /* (12, 3, 2) {real, imag} */,
  {32'h43d9a1cc, 32'h00000000} /* (12, 3, 1) {real, imag} */,
  {32'hc30718aa, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'h4358d2ba, 32'h00000000} /* (12, 2, 15) {real, imag} */,
  {32'hc2d1753b, 32'h00000000} /* (12, 2, 14) {real, imag} */,
  {32'h43f54356, 32'h00000000} /* (12, 2, 13) {real, imag} */,
  {32'h43c99263, 32'h00000000} /* (12, 2, 12) {real, imag} */,
  {32'h430c3b4a, 32'h00000000} /* (12, 2, 11) {real, imag} */,
  {32'h43a17d2a, 32'h00000000} /* (12, 2, 10) {real, imag} */,
  {32'hc1dceb60, 32'h00000000} /* (12, 2, 9) {real, imag} */,
  {32'hc3b48244, 32'h00000000} /* (12, 2, 8) {real, imag} */,
  {32'h43c05e55, 32'h00000000} /* (12, 2, 7) {real, imag} */,
  {32'hc3059b5f, 32'h00000000} /* (12, 2, 6) {real, imag} */,
  {32'hc46e34cf, 32'h00000000} /* (12, 2, 5) {real, imag} */,
  {32'hc3d39ec1, 32'h00000000} /* (12, 2, 4) {real, imag} */,
  {32'h4368aa2a, 32'h00000000} /* (12, 2, 3) {real, imag} */,
  {32'hc35a11ac, 32'h00000000} /* (12, 2, 2) {real, imag} */,
  {32'h441ef719, 32'h00000000} /* (12, 2, 1) {real, imag} */,
  {32'hc1b22098, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'hc31cd777, 32'h00000000} /* (12, 1, 15) {real, imag} */,
  {32'hc3b74fdc, 32'h00000000} /* (12, 1, 14) {real, imag} */,
  {32'h4443d03c, 32'h00000000} /* (12, 1, 13) {real, imag} */,
  {32'h43111cd6, 32'h00000000} /* (12, 1, 12) {real, imag} */,
  {32'h4489f4bf, 32'h00000000} /* (12, 1, 11) {real, imag} */,
  {32'h43bdc9a8, 32'h00000000} /* (12, 1, 10) {real, imag} */,
  {32'hc29c5b9a, 32'h00000000} /* (12, 1, 9) {real, imag} */,
  {32'h43efd431, 32'h00000000} /* (12, 1, 8) {real, imag} */,
  {32'h4370d707, 32'h00000000} /* (12, 1, 7) {real, imag} */,
  {32'hc3cec268, 32'h00000000} /* (12, 1, 6) {real, imag} */,
  {32'hc3c4c714, 32'h00000000} /* (12, 1, 5) {real, imag} */,
  {32'h428370cc, 32'h00000000} /* (12, 1, 4) {real, imag} */,
  {32'hc394ab1b, 32'h00000000} /* (12, 1, 3) {real, imag} */,
  {32'h41e0a948, 32'h00000000} /* (12, 1, 2) {real, imag} */,
  {32'hc396aafc, 32'h00000000} /* (12, 1, 1) {real, imag} */,
  {32'h437fa5ce, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'h436857db, 32'h00000000} /* (12, 0, 15) {real, imag} */,
  {32'h435b14ac, 32'h00000000} /* (12, 0, 14) {real, imag} */,
  {32'h4334f3ca, 32'h00000000} /* (12, 0, 13) {real, imag} */,
  {32'h4334caf0, 32'h00000000} /* (12, 0, 12) {real, imag} */,
  {32'h429b7d4d, 32'h00000000} /* (12, 0, 11) {real, imag} */,
  {32'h42ad2870, 32'h00000000} /* (12, 0, 10) {real, imag} */,
  {32'h43305ac9, 32'h00000000} /* (12, 0, 9) {real, imag} */,
  {32'h438ada1c, 32'h00000000} /* (12, 0, 8) {real, imag} */,
  {32'hc331f1e7, 32'h00000000} /* (12, 0, 7) {real, imag} */,
  {32'hc39401f8, 32'h00000000} /* (12, 0, 6) {real, imag} */,
  {32'hc2e3d5b3, 32'h00000000} /* (12, 0, 5) {real, imag} */,
  {32'h43963b76, 32'h00000000} /* (12, 0, 4) {real, imag} */,
  {32'h438d1807, 32'h00000000} /* (12, 0, 3) {real, imag} */,
  {32'h439b672a, 32'h00000000} /* (12, 0, 2) {real, imag} */,
  {32'h438877d6, 32'h00000000} /* (12, 0, 1) {real, imag} */,
  {32'h43c89632, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h441bb08d, 32'h00000000} /* (11, 15, 15) {real, imag} */,
  {32'h4405c094, 32'h00000000} /* (11, 15, 14) {real, imag} */,
  {32'h4294abde, 32'h00000000} /* (11, 15, 13) {real, imag} */,
  {32'h4414053e, 32'h00000000} /* (11, 15, 12) {real, imag} */,
  {32'h43a154c0, 32'h00000000} /* (11, 15, 11) {real, imag} */,
  {32'hc2af55a0, 32'h00000000} /* (11, 15, 10) {real, imag} */,
  {32'hc3a31db6, 32'h00000000} /* (11, 15, 9) {real, imag} */,
  {32'hc4873b65, 32'h00000000} /* (11, 15, 8) {real, imag} */,
  {32'hc3513355, 32'h00000000} /* (11, 15, 7) {real, imag} */,
  {32'h4413d71e, 32'h00000000} /* (11, 15, 6) {real, imag} */,
  {32'h438495c6, 32'h00000000} /* (11, 15, 5) {real, imag} */,
  {32'h4481359b, 32'h00000000} /* (11, 15, 4) {real, imag} */,
  {32'h44265b3e, 32'h00000000} /* (11, 15, 3) {real, imag} */,
  {32'hc42861de, 32'h00000000} /* (11, 15, 2) {real, imag} */,
  {32'h4405db84, 32'h00000000} /* (11, 15, 1) {real, imag} */,
  {32'h43121a38, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'h447ae9cc, 32'h00000000} /* (11, 14, 15) {real, imag} */,
  {32'h43e52146, 32'h00000000} /* (11, 14, 14) {real, imag} */,
  {32'h44309040, 32'h00000000} /* (11, 14, 13) {real, imag} */,
  {32'hc3550d06, 32'h00000000} /* (11, 14, 12) {real, imag} */,
  {32'h442f3c06, 32'h00000000} /* (11, 14, 11) {real, imag} */,
  {32'h43889145, 32'h00000000} /* (11, 14, 10) {real, imag} */,
  {32'h43820548, 32'h00000000} /* (11, 14, 9) {real, imag} */,
  {32'hc42d9180, 32'h00000000} /* (11, 14, 8) {real, imag} */,
  {32'h442f45ce, 32'h00000000} /* (11, 14, 7) {real, imag} */,
  {32'h447812e9, 32'h00000000} /* (11, 14, 6) {real, imag} */,
  {32'h448bc5fa, 32'h00000000} /* (11, 14, 5) {real, imag} */,
  {32'h4437d666, 32'h00000000} /* (11, 14, 4) {real, imag} */,
  {32'h447968e0, 32'h00000000} /* (11, 14, 3) {real, imag} */,
  {32'h42cfd195, 32'h00000000} /* (11, 14, 2) {real, imag} */,
  {32'hc39bc60a, 32'h00000000} /* (11, 14, 1) {real, imag} */,
  {32'h4390be4e, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'h40f8a900, 32'h00000000} /* (11, 13, 15) {real, imag} */,
  {32'h44cbb4a0, 32'h00000000} /* (11, 13, 14) {real, imag} */,
  {32'h43b678b0, 32'h00000000} /* (11, 13, 13) {real, imag} */,
  {32'hc3e29407, 32'h00000000} /* (11, 13, 12) {real, imag} */,
  {32'h4158d700, 32'h00000000} /* (11, 13, 11) {real, imag} */,
  {32'h435a3e16, 32'h00000000} /* (11, 13, 10) {real, imag} */,
  {32'h445912c2, 32'h00000000} /* (11, 13, 9) {real, imag} */,
  {32'h4404b253, 32'h00000000} /* (11, 13, 8) {real, imag} */,
  {32'h4507d5ac, 32'h00000000} /* (11, 13, 7) {real, imag} */,
  {32'h43cd8b9e, 32'h00000000} /* (11, 13, 6) {real, imag} */,
  {32'h44060a84, 32'h00000000} /* (11, 13, 5) {real, imag} */,
  {32'h44b7636d, 32'h00000000} /* (11, 13, 4) {real, imag} */,
  {32'h425dc200, 32'h00000000} /* (11, 13, 3) {real, imag} */,
  {32'hc308611e, 32'h00000000} /* (11, 13, 2) {real, imag} */,
  {32'h443aecb6, 32'h00000000} /* (11, 13, 1) {real, imag} */,
  {32'h43cad7ec, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'h43c9d66a, 32'h00000000} /* (11, 12, 15) {real, imag} */,
  {32'hc3f2ec60, 32'h00000000} /* (11, 12, 14) {real, imag} */,
  {32'hc3725287, 32'h00000000} /* (11, 12, 13) {real, imag} */,
  {32'h448b462e, 32'h00000000} /* (11, 12, 12) {real, imag} */,
  {32'h447cd650, 32'h00000000} /* (11, 12, 11) {real, imag} */,
  {32'h444a2e4b, 32'h00000000} /* (11, 12, 10) {real, imag} */,
  {32'hc2c80598, 32'h00000000} /* (11, 12, 9) {real, imag} */,
  {32'h43866de1, 32'h00000000} /* (11, 12, 8) {real, imag} */,
  {32'h4471a1eb, 32'h00000000} /* (11, 12, 7) {real, imag} */,
  {32'h43ab160c, 32'h00000000} /* (11, 12, 6) {real, imag} */,
  {32'h42cdae9e, 32'h00000000} /* (11, 12, 5) {real, imag} */,
  {32'h44af795e, 32'h00000000} /* (11, 12, 4) {real, imag} */,
  {32'h44348d70, 32'h00000000} /* (11, 12, 3) {real, imag} */,
  {32'h430c0794, 32'h00000000} /* (11, 12, 2) {real, imag} */,
  {32'h4488515a, 32'h00000000} /* (11, 12, 1) {real, imag} */,
  {32'h448f20e7, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'h43dc271a, 32'h00000000} /* (11, 11, 15) {real, imag} */,
  {32'hc26a37f0, 32'h00000000} /* (11, 11, 14) {real, imag} */,
  {32'h4405a22c, 32'h00000000} /* (11, 11, 13) {real, imag} */,
  {32'h438ce914, 32'h00000000} /* (11, 11, 12) {real, imag} */,
  {32'h446f09ee, 32'h00000000} /* (11, 11, 11) {real, imag} */,
  {32'h438490a6, 32'h00000000} /* (11, 11, 10) {real, imag} */,
  {32'h437c7404, 32'h00000000} /* (11, 11, 9) {real, imag} */,
  {32'h4351c024, 32'h00000000} /* (11, 11, 8) {real, imag} */,
  {32'h4441db4d, 32'h00000000} /* (11, 11, 7) {real, imag} */,
  {32'h449bf800, 32'h00000000} /* (11, 11, 6) {real, imag} */,
  {32'h447c13fc, 32'h00000000} /* (11, 11, 5) {real, imag} */,
  {32'h4404f87e, 32'h00000000} /* (11, 11, 4) {real, imag} */,
  {32'h43ddc768, 32'h00000000} /* (11, 11, 3) {real, imag} */,
  {32'h4456f2d1, 32'h00000000} /* (11, 11, 2) {real, imag} */,
  {32'h44a48a7a, 32'h00000000} /* (11, 11, 1) {real, imag} */,
  {32'h448670f2, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'h43b6f974, 32'h00000000} /* (11, 10, 15) {real, imag} */,
  {32'h446271c1, 32'h00000000} /* (11, 10, 14) {real, imag} */,
  {32'h4279f110, 32'h00000000} /* (11, 10, 13) {real, imag} */,
  {32'h4414aae0, 32'h00000000} /* (11, 10, 12) {real, imag} */,
  {32'h438370da, 32'h00000000} /* (11, 10, 11) {real, imag} */,
  {32'h43eeef17, 32'h00000000} /* (11, 10, 10) {real, imag} */,
  {32'h440bc5a9, 32'h00000000} /* (11, 10, 9) {real, imag} */,
  {32'h4412f1aa, 32'h00000000} /* (11, 10, 8) {real, imag} */,
  {32'h4505d834, 32'h00000000} /* (11, 10, 7) {real, imag} */,
  {32'h43bc374a, 32'h00000000} /* (11, 10, 6) {real, imag} */,
  {32'h44a8333c, 32'h00000000} /* (11, 10, 5) {real, imag} */,
  {32'h4499e1ce, 32'h00000000} /* (11, 10, 4) {real, imag} */,
  {32'h44054d0b, 32'h00000000} /* (11, 10, 3) {real, imag} */,
  {32'h4480eb69, 32'h00000000} /* (11, 10, 2) {real, imag} */,
  {32'h44b6f15c, 32'h00000000} /* (11, 10, 1) {real, imag} */,
  {32'h442eeb26, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h442091b8, 32'h00000000} /* (11, 9, 15) {real, imag} */,
  {32'h433b0cc9, 32'h00000000} /* (11, 9, 14) {real, imag} */,
  {32'hc31e3eb0, 32'h00000000} /* (11, 9, 13) {real, imag} */,
  {32'h442c330e, 32'h00000000} /* (11, 9, 12) {real, imag} */,
  {32'h448a6b03, 32'h00000000} /* (11, 9, 11) {real, imag} */,
  {32'h444c19b0, 32'h00000000} /* (11, 9, 10) {real, imag} */,
  {32'h437ae8b8, 32'h00000000} /* (11, 9, 9) {real, imag} */,
  {32'h442197ba, 32'h00000000} /* (11, 9, 8) {real, imag} */,
  {32'h448be10a, 32'h00000000} /* (11, 9, 7) {real, imag} */,
  {32'hc38cdd44, 32'h00000000} /* (11, 9, 6) {real, imag} */,
  {32'hc41cf9d0, 32'h00000000} /* (11, 9, 5) {real, imag} */,
  {32'h438920f4, 32'h00000000} /* (11, 9, 4) {real, imag} */,
  {32'h43a0996b, 32'h00000000} /* (11, 9, 3) {real, imag} */,
  {32'h4353ece2, 32'h00000000} /* (11, 9, 2) {real, imag} */,
  {32'h44b72603, 32'h00000000} /* (11, 9, 1) {real, imag} */,
  {32'h43cf1ad4, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h446d72fc, 32'h00000000} /* (11, 8, 15) {real, imag} */,
  {32'h445ed76c, 32'h00000000} /* (11, 8, 14) {real, imag} */,
  {32'h43b8e864, 32'h00000000} /* (11, 8, 13) {real, imag} */,
  {32'hc447d9f4, 32'h00000000} /* (11, 8, 12) {real, imag} */,
  {32'h44190467, 32'h00000000} /* (11, 8, 11) {real, imag} */,
  {32'h436314b4, 32'h00000000} /* (11, 8, 10) {real, imag} */,
  {32'h4421a2e2, 32'h00000000} /* (11, 8, 9) {real, imag} */,
  {32'hc33b4dda, 32'h00000000} /* (11, 8, 8) {real, imag} */,
  {32'hc329b390, 32'h00000000} /* (11, 8, 7) {real, imag} */,
  {32'hc3ed1500, 32'h00000000} /* (11, 8, 6) {real, imag} */,
  {32'hc2461e54, 32'h00000000} /* (11, 8, 5) {real, imag} */,
  {32'hc2af36ec, 32'h00000000} /* (11, 8, 4) {real, imag} */,
  {32'hc44ffdc9, 32'h00000000} /* (11, 8, 3) {real, imag} */,
  {32'hc3a2a46a, 32'h00000000} /* (11, 8, 2) {real, imag} */,
  {32'h440762aa, 32'h00000000} /* (11, 8, 1) {real, imag} */,
  {32'h43a1335f, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h43f1fa04, 32'h00000000} /* (11, 7, 15) {real, imag} */,
  {32'h4447f3ac, 32'h00000000} /* (11, 7, 14) {real, imag} */,
  {32'hc4c3c094, 32'h00000000} /* (11, 7, 13) {real, imag} */,
  {32'h42c0b7ce, 32'h00000000} /* (11, 7, 12) {real, imag} */,
  {32'h44580743, 32'h00000000} /* (11, 7, 11) {real, imag} */,
  {32'h43464eca, 32'h00000000} /* (11, 7, 10) {real, imag} */,
  {32'h430f3b90, 32'h00000000} /* (11, 7, 9) {real, imag} */,
  {32'h42f7ecf4, 32'h00000000} /* (11, 7, 8) {real, imag} */,
  {32'h43ac68c6, 32'h00000000} /* (11, 7, 7) {real, imag} */,
  {32'h429e3df4, 32'h00000000} /* (11, 7, 6) {real, imag} */,
  {32'hc3cb5252, 32'h00000000} /* (11, 7, 5) {real, imag} */,
  {32'hc28001c6, 32'h00000000} /* (11, 7, 4) {real, imag} */,
  {32'h43fb3482, 32'h00000000} /* (11, 7, 3) {real, imag} */,
  {32'h4366cc5a, 32'h00000000} /* (11, 7, 2) {real, imag} */,
  {32'hc0415c00, 32'h00000000} /* (11, 7, 1) {real, imag} */,
  {32'h434a3c76, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'h419c3040, 32'h00000000} /* (11, 6, 15) {real, imag} */,
  {32'h433be582, 32'h00000000} /* (11, 6, 14) {real, imag} */,
  {32'h442d4994, 32'h00000000} /* (11, 6, 13) {real, imag} */,
  {32'h43678ff6, 32'h00000000} /* (11, 6, 12) {real, imag} */,
  {32'h44031982, 32'h00000000} /* (11, 6, 11) {real, imag} */,
  {32'hc3e3b83d, 32'h00000000} /* (11, 6, 10) {real, imag} */,
  {32'h44a6229b, 32'h00000000} /* (11, 6, 9) {real, imag} */,
  {32'h444e3d2a, 32'h00000000} /* (11, 6, 8) {real, imag} */,
  {32'h44dbc615, 32'h00000000} /* (11, 6, 7) {real, imag} */,
  {32'h44798122, 32'h00000000} /* (11, 6, 6) {real, imag} */,
  {32'hc32c285e, 32'h00000000} /* (11, 6, 5) {real, imag} */,
  {32'hc42b0222, 32'h00000000} /* (11, 6, 4) {real, imag} */,
  {32'h446dd9da, 32'h00000000} /* (11, 6, 3) {real, imag} */,
  {32'hc2556758, 32'h00000000} /* (11, 6, 2) {real, imag} */,
  {32'hc457fbea, 32'h00000000} /* (11, 6, 1) {real, imag} */,
  {32'h43851bbc, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'h439fc646, 32'h00000000} /* (11, 5, 15) {real, imag} */,
  {32'h4384dd38, 32'h00000000} /* (11, 5, 14) {real, imag} */,
  {32'h4184e7b0, 32'h00000000} /* (11, 5, 13) {real, imag} */,
  {32'hc35915d0, 32'h00000000} /* (11, 5, 12) {real, imag} */,
  {32'hc3fd7e06, 32'h00000000} /* (11, 5, 11) {real, imag} */,
  {32'hc3e5f1f3, 32'h00000000} /* (11, 5, 10) {real, imag} */,
  {32'h449d8121, 32'h00000000} /* (11, 5, 9) {real, imag} */,
  {32'h4462450a, 32'h00000000} /* (11, 5, 8) {real, imag} */,
  {32'h44d2b3fa, 32'h00000000} /* (11, 5, 7) {real, imag} */,
  {32'h442ad32b, 32'h00000000} /* (11, 5, 6) {real, imag} */,
  {32'h42ed423c, 32'h00000000} /* (11, 5, 5) {real, imag} */,
  {32'h44ab27cf, 32'h00000000} /* (11, 5, 4) {real, imag} */,
  {32'h442f3471, 32'h00000000} /* (11, 5, 3) {real, imag} */,
  {32'h443c588a, 32'h00000000} /* (11, 5, 2) {real, imag} */,
  {32'h43a159d4, 32'h00000000} /* (11, 5, 1) {real, imag} */,
  {32'h43991de8, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h4409713c, 32'h00000000} /* (11, 4, 15) {real, imag} */,
  {32'h443a7d9e, 32'h00000000} /* (11, 4, 14) {real, imag} */,
  {32'hc40dfcfe, 32'h00000000} /* (11, 4, 13) {real, imag} */,
  {32'hc41a4eea, 32'h00000000} /* (11, 4, 12) {real, imag} */,
  {32'hc3ee651c, 32'h00000000} /* (11, 4, 11) {real, imag} */,
  {32'hc3cc58fc, 32'h00000000} /* (11, 4, 10) {real, imag} */,
  {32'h4335ee3a, 32'h00000000} /* (11, 4, 9) {real, imag} */,
  {32'h43f62f3f, 32'h00000000} /* (11, 4, 8) {real, imag} */,
  {32'h4465ad44, 32'h00000000} /* (11, 4, 7) {real, imag} */,
  {32'h44064192, 32'h00000000} /* (11, 4, 6) {real, imag} */,
  {32'h41f0c250, 32'h00000000} /* (11, 4, 5) {real, imag} */,
  {32'h447aae9c, 32'h00000000} /* (11, 4, 4) {real, imag} */,
  {32'h4496a3c5, 32'h00000000} /* (11, 4, 3) {real, imag} */,
  {32'h43d7cf6a, 32'h00000000} /* (11, 4, 2) {real, imag} */,
  {32'h443906a0, 32'h00000000} /* (11, 4, 1) {real, imag} */,
  {32'h43bb5e9f, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h434bccc0, 32'h00000000} /* (11, 3, 15) {real, imag} */,
  {32'hc380ca32, 32'h00000000} /* (11, 3, 14) {real, imag} */,
  {32'hc4001aaa, 32'h00000000} /* (11, 3, 13) {real, imag} */,
  {32'hc400a42f, 32'h00000000} /* (11, 3, 12) {real, imag} */,
  {32'h42b58dc8, 32'h00000000} /* (11, 3, 11) {real, imag} */,
  {32'hc3efc950, 32'h00000000} /* (11, 3, 10) {real, imag} */,
  {32'hc42ce5c5, 32'h00000000} /* (11, 3, 9) {real, imag} */,
  {32'h4206bd3c, 32'h00000000} /* (11, 3, 8) {real, imag} */,
  {32'h437dcbb0, 32'h00000000} /* (11, 3, 7) {real, imag} */,
  {32'h420081a8, 32'h00000000} /* (11, 3, 6) {real, imag} */,
  {32'h42b68fca, 32'h00000000} /* (11, 3, 5) {real, imag} */,
  {32'hc3e5d8f2, 32'h00000000} /* (11, 3, 4) {real, imag} */,
  {32'h44b5efea, 32'h00000000} /* (11, 3, 3) {real, imag} */,
  {32'h4435b842, 32'h00000000} /* (11, 3, 2) {real, imag} */,
  {32'hc379164c, 32'h00000000} /* (11, 3, 1) {real, imag} */,
  {32'h4305758f, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'hc286ee5c, 32'h00000000} /* (11, 2, 15) {real, imag} */,
  {32'hc479732e, 32'h00000000} /* (11, 2, 14) {real, imag} */,
  {32'hc354b00c, 32'h00000000} /* (11, 2, 13) {real, imag} */,
  {32'hc2e2fda2, 32'h00000000} /* (11, 2, 12) {real, imag} */,
  {32'h447cc2b0, 32'h00000000} /* (11, 2, 11) {real, imag} */,
  {32'h4353b85c, 32'h00000000} /* (11, 2, 10) {real, imag} */,
  {32'hc3bcbcd6, 32'h00000000} /* (11, 2, 9) {real, imag} */,
  {32'h4260e23e, 32'h00000000} /* (11, 2, 8) {real, imag} */,
  {32'h4292a338, 32'h00000000} /* (11, 2, 7) {real, imag} */,
  {32'h43cabaf4, 32'h00000000} /* (11, 2, 6) {real, imag} */,
  {32'hc44f26cd, 32'h00000000} /* (11, 2, 5) {real, imag} */,
  {32'hc39210f8, 32'h00000000} /* (11, 2, 4) {real, imag} */,
  {32'hc279c000, 32'h00000000} /* (11, 2, 3) {real, imag} */,
  {32'hc44b8359, 32'h00000000} /* (11, 2, 2) {real, imag} */,
  {32'hc36ea134, 32'h00000000} /* (11, 2, 1) {real, imag} */,
  {32'hc19eacc4, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'h43a8f72f, 32'h00000000} /* (11, 1, 15) {real, imag} */,
  {32'h43a0226c, 32'h00000000} /* (11, 1, 14) {real, imag} */,
  {32'h43d2cf4b, 32'h00000000} /* (11, 1, 13) {real, imag} */,
  {32'hc24a1190, 32'h00000000} /* (11, 1, 12) {real, imag} */,
  {32'hc202a242, 32'h00000000} /* (11, 1, 11) {real, imag} */,
  {32'h44507743, 32'h00000000} /* (11, 1, 10) {real, imag} */,
  {32'h43727475, 32'h00000000} /* (11, 1, 9) {real, imag} */,
  {32'h432e76f6, 32'h00000000} /* (11, 1, 8) {real, imag} */,
  {32'h4457b30c, 32'h00000000} /* (11, 1, 7) {real, imag} */,
  {32'h4353f910, 32'h00000000} /* (11, 1, 6) {real, imag} */,
  {32'h436a3f5a, 32'h00000000} /* (11, 1, 5) {real, imag} */,
  {32'h44689ee7, 32'h00000000} /* (11, 1, 4) {real, imag} */,
  {32'h42791812, 32'h00000000} /* (11, 1, 3) {real, imag} */,
  {32'hc3956002, 32'h00000000} /* (11, 1, 2) {real, imag} */,
  {32'h42b908be, 32'h00000000} /* (11, 1, 1) {real, imag} */,
  {32'h4361fff4, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h42fde50c, 32'h00000000} /* (11, 0, 15) {real, imag} */,
  {32'h42fe9234, 32'h00000000} /* (11, 0, 14) {real, imag} */,
  {32'h428c88e8, 32'h00000000} /* (11, 0, 13) {real, imag} */,
  {32'hc38942c9, 32'h00000000} /* (11, 0, 12) {real, imag} */,
  {32'hc393a70a, 32'h00000000} /* (11, 0, 11) {real, imag} */,
  {32'h4342cb7c, 32'h00000000} /* (11, 0, 10) {real, imag} */,
  {32'hbfebca80, 32'h00000000} /* (11, 0, 9) {real, imag} */,
  {32'hc22bd7b8, 32'h00000000} /* (11, 0, 8) {real, imag} */,
  {32'h440b0b80, 32'h00000000} /* (11, 0, 7) {real, imag} */,
  {32'hc349f99a, 32'h00000000} /* (11, 0, 6) {real, imag} */,
  {32'hc3455cbe, 32'h00000000} /* (11, 0, 5) {real, imag} */,
  {32'h443a4398, 32'h00000000} /* (11, 0, 4) {real, imag} */,
  {32'h430741b1, 32'h00000000} /* (11, 0, 3) {real, imag} */,
  {32'h44512761, 32'h00000000} /* (11, 0, 2) {real, imag} */,
  {32'h432e9bc7, 32'h00000000} /* (11, 0, 1) {real, imag} */,
  {32'h4413e850, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h43cc8ce0, 32'h00000000} /* (10, 15, 15) {real, imag} */,
  {32'h4395ce4e, 32'h00000000} /* (10, 15, 14) {real, imag} */,
  {32'h43dffd27, 32'h00000000} /* (10, 15, 13) {real, imag} */,
  {32'h43b209c8, 32'h00000000} /* (10, 15, 12) {real, imag} */,
  {32'h43a75143, 32'h00000000} /* (10, 15, 11) {real, imag} */,
  {32'h438f2d8e, 32'h00000000} /* (10, 15, 10) {real, imag} */,
  {32'hc3582d6c, 32'h00000000} /* (10, 15, 9) {real, imag} */,
  {32'hc3f42bba, 32'h00000000} /* (10, 15, 8) {real, imag} */,
  {32'h440b7acb, 32'h00000000} /* (10, 15, 7) {real, imag} */,
  {32'h4423c04f, 32'h00000000} /* (10, 15, 6) {real, imag} */,
  {32'h44275f7c, 32'h00000000} /* (10, 15, 5) {real, imag} */,
  {32'h434f3e58, 32'h00000000} /* (10, 15, 4) {real, imag} */,
  {32'hc421fbfa, 32'h00000000} /* (10, 15, 3) {real, imag} */,
  {32'h43cc540e, 32'h00000000} /* (10, 15, 2) {real, imag} */,
  {32'h43954940, 32'h00000000} /* (10, 15, 1) {real, imag} */,
  {32'h4356f55b, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'h445931fb, 32'h00000000} /* (10, 14, 15) {real, imag} */,
  {32'h44b19738, 32'h00000000} /* (10, 14, 14) {real, imag} */,
  {32'h44a8cfdb, 32'h00000000} /* (10, 14, 13) {real, imag} */,
  {32'h444c8220, 32'h00000000} /* (10, 14, 12) {real, imag} */,
  {32'h43c8d46f, 32'h00000000} /* (10, 14, 11) {real, imag} */,
  {32'h42cbdcb4, 32'h00000000} /* (10, 14, 10) {real, imag} */,
  {32'hc4516852, 32'h00000000} /* (10, 14, 9) {real, imag} */,
  {32'hc38f907c, 32'h00000000} /* (10, 14, 8) {real, imag} */,
  {32'h443bcb5d, 32'h00000000} /* (10, 14, 7) {real, imag} */,
  {32'h4453a11c, 32'h00000000} /* (10, 14, 6) {real, imag} */,
  {32'h449294af, 32'h00000000} /* (10, 14, 5) {real, imag} */,
  {32'h44155ebc, 32'h00000000} /* (10, 14, 4) {real, imag} */,
  {32'hc42c7040, 32'h00000000} /* (10, 14, 3) {real, imag} */,
  {32'hc4401090, 32'h00000000} /* (10, 14, 2) {real, imag} */,
  {32'h43a21ee1, 32'h00000000} /* (10, 14, 1) {real, imag} */,
  {32'h438f3690, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'h44172e5c, 32'h00000000} /* (10, 13, 15) {real, imag} */,
  {32'h44b616ce, 32'h00000000} /* (10, 13, 14) {real, imag} */,
  {32'h43fd215c, 32'h00000000} /* (10, 13, 13) {real, imag} */,
  {32'h443bfb2d, 32'h00000000} /* (10, 13, 12) {real, imag} */,
  {32'h448cb03d, 32'h00000000} /* (10, 13, 11) {real, imag} */,
  {32'h43e8df9f, 32'h00000000} /* (10, 13, 10) {real, imag} */,
  {32'hc2d595f0, 32'h00000000} /* (10, 13, 9) {real, imag} */,
  {32'h43840433, 32'h00000000} /* (10, 13, 8) {real, imag} */,
  {32'h447156d4, 32'h00000000} /* (10, 13, 7) {real, imag} */,
  {32'h44c85546, 32'h00000000} /* (10, 13, 6) {real, imag} */,
  {32'h4412f792, 32'h00000000} /* (10, 13, 5) {real, imag} */,
  {32'h430cffac, 32'h00000000} /* (10, 13, 4) {real, imag} */,
  {32'h44590fd6, 32'h00000000} /* (10, 13, 3) {real, imag} */,
  {32'hc3239cd6, 32'h00000000} /* (10, 13, 2) {real, imag} */,
  {32'h447a27dc, 32'h00000000} /* (10, 13, 1) {real, imag} */,
  {32'h43fbe65d, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'h43ce7a65, 32'h00000000} /* (10, 12, 15) {real, imag} */,
  {32'hc30ee318, 32'h00000000} /* (10, 12, 14) {real, imag} */,
  {32'hc3b1eacb, 32'h00000000} /* (10, 12, 13) {real, imag} */,
  {32'hc3fbe02c, 32'h00000000} /* (10, 12, 12) {real, imag} */,
  {32'h40fbd3e0, 32'h00000000} /* (10, 12, 11) {real, imag} */,
  {32'hc390259b, 32'h00000000} /* (10, 12, 10) {real, imag} */,
  {32'h4498ab2b, 32'h00000000} /* (10, 12, 9) {real, imag} */,
  {32'h448f930b, 32'h00000000} /* (10, 12, 8) {real, imag} */,
  {32'h44ad7aef, 32'h00000000} /* (10, 12, 7) {real, imag} */,
  {32'h44f2de23, 32'h00000000} /* (10, 12, 6) {real, imag} */,
  {32'h444b3bd6, 32'h00000000} /* (10, 12, 5) {real, imag} */,
  {32'h4427bed6, 32'h00000000} /* (10, 12, 4) {real, imag} */,
  {32'h43380d65, 32'h00000000} /* (10, 12, 3) {real, imag} */,
  {32'h43e53c13, 32'h00000000} /* (10, 12, 2) {real, imag} */,
  {32'h4480b1f9, 32'h00000000} /* (10, 12, 1) {real, imag} */,
  {32'h44242866, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hc3a39dd5, 32'h00000000} /* (10, 11, 15) {real, imag} */,
  {32'h4386399a, 32'h00000000} /* (10, 11, 14) {real, imag} */,
  {32'hc19a8280, 32'h00000000} /* (10, 11, 13) {real, imag} */,
  {32'h4347abb0, 32'h00000000} /* (10, 11, 12) {real, imag} */,
  {32'h434daeb4, 32'h00000000} /* (10, 11, 11) {real, imag} */,
  {32'h43b9af34, 32'h00000000} /* (10, 11, 10) {real, imag} */,
  {32'h450e6310, 32'h00000000} /* (10, 11, 9) {real, imag} */,
  {32'h449d67a3, 32'h00000000} /* (10, 11, 8) {real, imag} */,
  {32'h44911037, 32'h00000000} /* (10, 11, 7) {real, imag} */,
  {32'h44a2304c, 32'h00000000} /* (10, 11, 6) {real, imag} */,
  {32'h44b82dac, 32'h00000000} /* (10, 11, 5) {real, imag} */,
  {32'h44c893d4, 32'h00000000} /* (10, 11, 4) {real, imag} */,
  {32'h445a07e3, 32'h00000000} /* (10, 11, 3) {real, imag} */,
  {32'h43d1700c, 32'h00000000} /* (10, 11, 2) {real, imag} */,
  {32'h43195bb8, 32'h00000000} /* (10, 11, 1) {real, imag} */,
  {32'h4420ab92, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h444970c4, 32'h00000000} /* (10, 10, 15) {real, imag} */,
  {32'h447ebf16, 32'h00000000} /* (10, 10, 14) {real, imag} */,
  {32'hc2635390, 32'h00000000} /* (10, 10, 13) {real, imag} */,
  {32'h441a4ef8, 32'h00000000} /* (10, 10, 12) {real, imag} */,
  {32'hc387a9a2, 32'h00000000} /* (10, 10, 11) {real, imag} */,
  {32'h4199f3a0, 32'h00000000} /* (10, 10, 10) {real, imag} */,
  {32'h442e61d5, 32'h00000000} /* (10, 10, 9) {real, imag} */,
  {32'h449b23b9, 32'h00000000} /* (10, 10, 8) {real, imag} */,
  {32'h44b4a5a6, 32'h00000000} /* (10, 10, 7) {real, imag} */,
  {32'h44678018, 32'h00000000} /* (10, 10, 6) {real, imag} */,
  {32'h449afcce, 32'h00000000} /* (10, 10, 5) {real, imag} */,
  {32'h44b0491d, 32'h00000000} /* (10, 10, 4) {real, imag} */,
  {32'h4440dfad, 32'h00000000} /* (10, 10, 3) {real, imag} */,
  {32'h44c44e6a, 32'h00000000} /* (10, 10, 2) {real, imag} */,
  {32'h449fcb56, 32'h00000000} /* (10, 10, 1) {real, imag} */,
  {32'h44144d1c, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h4433a3c0, 32'h00000000} /* (10, 9, 15) {real, imag} */,
  {32'h448dba7b, 32'h00000000} /* (10, 9, 14) {real, imag} */,
  {32'h43ed1de6, 32'h00000000} /* (10, 9, 13) {real, imag} */,
  {32'hbf575b80, 32'h00000000} /* (10, 9, 12) {real, imag} */,
  {32'h422cc128, 32'h00000000} /* (10, 9, 11) {real, imag} */,
  {32'h440067d8, 32'h00000000} /* (10, 9, 10) {real, imag} */,
  {32'h4437cda4, 32'h00000000} /* (10, 9, 9) {real, imag} */,
  {32'h4422d12c, 32'h00000000} /* (10, 9, 8) {real, imag} */,
  {32'h4479cb66, 32'h00000000} /* (10, 9, 7) {real, imag} */,
  {32'hc3df22b5, 32'h00000000} /* (10, 9, 6) {real, imag} */,
  {32'hc40ba855, 32'h00000000} /* (10, 9, 5) {real, imag} */,
  {32'hc3012964, 32'h00000000} /* (10, 9, 4) {real, imag} */,
  {32'h44297dec, 32'h00000000} /* (10, 9, 3) {real, imag} */,
  {32'h449e53fc, 32'h00000000} /* (10, 9, 2) {real, imag} */,
  {32'h44979101, 32'h00000000} /* (10, 9, 1) {real, imag} */,
  {32'h44b255f0, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'h449381fb, 32'h00000000} /* (10, 8, 15) {real, imag} */,
  {32'h447e6e13, 32'h00000000} /* (10, 8, 14) {real, imag} */,
  {32'h44874d16, 32'h00000000} /* (10, 8, 13) {real, imag} */,
  {32'h42caabd6, 32'h00000000} /* (10, 8, 12) {real, imag} */,
  {32'h440f4807, 32'h00000000} /* (10, 8, 11) {real, imag} */,
  {32'h43856cb0, 32'h00000000} /* (10, 8, 10) {real, imag} */,
  {32'h4481708f, 32'h00000000} /* (10, 8, 9) {real, imag} */,
  {32'h4482405f, 32'h00000000} /* (10, 8, 8) {real, imag} */,
  {32'h44541862, 32'h00000000} /* (10, 8, 7) {real, imag} */,
  {32'hc42df0f3, 32'h00000000} /* (10, 8, 6) {real, imag} */,
  {32'hc402909a, 32'h00000000} /* (10, 8, 5) {real, imag} */,
  {32'h432c2687, 32'h00000000} /* (10, 8, 4) {real, imag} */,
  {32'hc3a0f00e, 32'h00000000} /* (10, 8, 3) {real, imag} */,
  {32'h42ca5f2e, 32'h00000000} /* (10, 8, 2) {real, imag} */,
  {32'h43c97075, 32'h00000000} /* (10, 8, 1) {real, imag} */,
  {32'hc3576688, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h448c46e1, 32'h00000000} /* (10, 7, 15) {real, imag} */,
  {32'h44df3b4e, 32'h00000000} /* (10, 7, 14) {real, imag} */,
  {32'h44725e2b, 32'h00000000} /* (10, 7, 13) {real, imag} */,
  {32'hc338b1d8, 32'h00000000} /* (10, 7, 12) {real, imag} */,
  {32'h435eda94, 32'h00000000} /* (10, 7, 11) {real, imag} */,
  {32'hc28fdde0, 32'h00000000} /* (10, 7, 10) {real, imag} */,
  {32'hc3c2f812, 32'h00000000} /* (10, 7, 9) {real, imag} */,
  {32'h42d7f580, 32'h00000000} /* (10, 7, 8) {real, imag} */,
  {32'h4479a36f, 32'h00000000} /* (10, 7, 7) {real, imag} */,
  {32'hc411a48b, 32'h00000000} /* (10, 7, 6) {real, imag} */,
  {32'h42978598, 32'h00000000} /* (10, 7, 5) {real, imag} */,
  {32'h44360c40, 32'h00000000} /* (10, 7, 4) {real, imag} */,
  {32'h442728d1, 32'h00000000} /* (10, 7, 3) {real, imag} */,
  {32'h4429111a, 32'h00000000} /* (10, 7, 2) {real, imag} */,
  {32'hc40ddbdf, 32'h00000000} /* (10, 7, 1) {real, imag} */,
  {32'h424574e0, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h441edd2a, 32'h00000000} /* (10, 6, 15) {real, imag} */,
  {32'h43cdcf66, 32'h00000000} /* (10, 6, 14) {real, imag} */,
  {32'h43c29d42, 32'h00000000} /* (10, 6, 13) {real, imag} */,
  {32'h44855bce, 32'h00000000} /* (10, 6, 12) {real, imag} */,
  {32'hc3da8589, 32'h00000000} /* (10, 6, 11) {real, imag} */,
  {32'h40898200, 32'h00000000} /* (10, 6, 10) {real, imag} */,
  {32'h43bb15d3, 32'h00000000} /* (10, 6, 9) {real, imag} */,
  {32'h4261a648, 32'h00000000} /* (10, 6, 8) {real, imag} */,
  {32'hc31baaba, 32'h00000000} /* (10, 6, 7) {real, imag} */,
  {32'h443b0989, 32'h00000000} /* (10, 6, 6) {real, imag} */,
  {32'h4412afd0, 32'h00000000} /* (10, 6, 5) {real, imag} */,
  {32'h44893b94, 32'h00000000} /* (10, 6, 4) {real, imag} */,
  {32'h43d51faf, 32'h00000000} /* (10, 6, 3) {real, imag} */,
  {32'hc3cc168a, 32'h00000000} /* (10, 6, 2) {real, imag} */,
  {32'hc41e92a2, 32'h00000000} /* (10, 6, 1) {real, imag} */,
  {32'h440ec088, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'h439389b2, 32'h00000000} /* (10, 5, 15) {real, imag} */,
  {32'h43b5243f, 32'h00000000} /* (10, 5, 14) {real, imag} */,
  {32'hc31119a4, 32'h00000000} /* (10, 5, 13) {real, imag} */,
  {32'hc391bcd1, 32'h00000000} /* (10, 5, 12) {real, imag} */,
  {32'hbe58b800, 32'h00000000} /* (10, 5, 11) {real, imag} */,
  {32'hc486cefa, 32'h00000000} /* (10, 5, 10) {real, imag} */,
  {32'h41475c00, 32'h00000000} /* (10, 5, 9) {real, imag} */,
  {32'h4302d418, 32'h00000000} /* (10, 5, 8) {real, imag} */,
  {32'h43fae41e, 32'h00000000} /* (10, 5, 7) {real, imag} */,
  {32'h441459ce, 32'h00000000} /* (10, 5, 6) {real, imag} */,
  {32'h44d17b1a, 32'h00000000} /* (10, 5, 5) {real, imag} */,
  {32'h445c08b0, 32'h00000000} /* (10, 5, 4) {real, imag} */,
  {32'hc3a061a9, 32'h00000000} /* (10, 5, 3) {real, imag} */,
  {32'hc41dc8c3, 32'h00000000} /* (10, 5, 2) {real, imag} */,
  {32'hc3e146d4, 32'h00000000} /* (10, 5, 1) {real, imag} */,
  {32'h420f7a2a, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h423eaaf0, 32'h00000000} /* (10, 4, 15) {real, imag} */,
  {32'h43062ca8, 32'h00000000} /* (10, 4, 14) {real, imag} */,
  {32'hc2e2c998, 32'h00000000} /* (10, 4, 13) {real, imag} */,
  {32'hc487a9ee, 32'h00000000} /* (10, 4, 12) {real, imag} */,
  {32'hc2a225f4, 32'h00000000} /* (10, 4, 11) {real, imag} */,
  {32'hc43c94f2, 32'h00000000} /* (10, 4, 10) {real, imag} */,
  {32'hc3d15f7a, 32'h00000000} /* (10, 4, 9) {real, imag} */,
  {32'h43291c96, 32'h00000000} /* (10, 4, 8) {real, imag} */,
  {32'hc33ed768, 32'h00000000} /* (10, 4, 7) {real, imag} */,
  {32'h444ac751, 32'h00000000} /* (10, 4, 6) {real, imag} */,
  {32'h443b8aef, 32'h00000000} /* (10, 4, 5) {real, imag} */,
  {32'h43bc0d7e, 32'h00000000} /* (10, 4, 4) {real, imag} */,
  {32'h444ed9dc, 32'h00000000} /* (10, 4, 3) {real, imag} */,
  {32'h4455f10c, 32'h00000000} /* (10, 4, 2) {real, imag} */,
  {32'h43bddeb4, 32'h00000000} /* (10, 4, 1) {real, imag} */,
  {32'h4427bf18, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'hc42cf358, 32'h00000000} /* (10, 3, 15) {real, imag} */,
  {32'hc43c7da6, 32'h00000000} /* (10, 3, 14) {real, imag} */,
  {32'hc2ad1a90, 32'h00000000} /* (10, 3, 13) {real, imag} */,
  {32'hc476c556, 32'h00000000} /* (10, 3, 12) {real, imag} */,
  {32'hc40a9a74, 32'h00000000} /* (10, 3, 11) {real, imag} */,
  {32'h43904ad1, 32'h00000000} /* (10, 3, 10) {real, imag} */,
  {32'hc383ceea, 32'h00000000} /* (10, 3, 9) {real, imag} */,
  {32'h444db63b, 32'h00000000} /* (10, 3, 8) {real, imag} */,
  {32'h42a719b4, 32'h00000000} /* (10, 3, 7) {real, imag} */,
  {32'h444c7bde, 32'h00000000} /* (10, 3, 6) {real, imag} */,
  {32'h43b11866, 32'h00000000} /* (10, 3, 5) {real, imag} */,
  {32'h441b12d0, 32'h00000000} /* (10, 3, 4) {real, imag} */,
  {32'h4439c2c8, 32'h00000000} /* (10, 3, 3) {real, imag} */,
  {32'h435d658d, 32'h00000000} /* (10, 3, 2) {real, imag} */,
  {32'h43ad06c0, 32'h00000000} /* (10, 3, 1) {real, imag} */,
  {32'h43a7b96e, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'hc413b248, 32'h00000000} /* (10, 2, 15) {real, imag} */,
  {32'hc48629ce, 32'h00000000} /* (10, 2, 14) {real, imag} */,
  {32'hc3808fe0, 32'h00000000} /* (10, 2, 13) {real, imag} */,
  {32'hc3a6b4a2, 32'h00000000} /* (10, 2, 12) {real, imag} */,
  {32'h43288cfb, 32'h00000000} /* (10, 2, 11) {real, imag} */,
  {32'h42f1b502, 32'h00000000} /* (10, 2, 10) {real, imag} */,
  {32'hc384e766, 32'h00000000} /* (10, 2, 9) {real, imag} */,
  {32'h44248c1a, 32'h00000000} /* (10, 2, 8) {real, imag} */,
  {32'h44ac15f5, 32'h00000000} /* (10, 2, 7) {real, imag} */,
  {32'h43612d70, 32'h00000000} /* (10, 2, 6) {real, imag} */,
  {32'h44168ee6, 32'h00000000} /* (10, 2, 5) {real, imag} */,
  {32'h43df638e, 32'h00000000} /* (10, 2, 4) {real, imag} */,
  {32'h41c00398, 32'h00000000} /* (10, 2, 3) {real, imag} */,
  {32'h3fb07b80, 32'h00000000} /* (10, 2, 2) {real, imag} */,
  {32'hc45160d9, 32'h00000000} /* (10, 2, 1) {real, imag} */,
  {32'h4329fcc6, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'h424f5fd4, 32'h00000000} /* (10, 1, 15) {real, imag} */,
  {32'hc349aa30, 32'h00000000} /* (10, 1, 14) {real, imag} */,
  {32'hc34e847b, 32'h00000000} /* (10, 1, 13) {real, imag} */,
  {32'hc31624b0, 32'h00000000} /* (10, 1, 12) {real, imag} */,
  {32'h443a973d, 32'h00000000} /* (10, 1, 11) {real, imag} */,
  {32'h440f76ce, 32'h00000000} /* (10, 1, 10) {real, imag} */,
  {32'hc23d6508, 32'h00000000} /* (10, 1, 9) {real, imag} */,
  {32'h4325eb10, 32'h00000000} /* (10, 1, 8) {real, imag} */,
  {32'h43cc5cd6, 32'h00000000} /* (10, 1, 7) {real, imag} */,
  {32'h44358e53, 32'h00000000} /* (10, 1, 6) {real, imag} */,
  {32'hc2a08682, 32'h00000000} /* (10, 1, 5) {real, imag} */,
  {32'h449d17c8, 32'h00000000} /* (10, 1, 4) {real, imag} */,
  {32'h4402537b, 32'h00000000} /* (10, 1, 3) {real, imag} */,
  {32'hc3c5404f, 32'h00000000} /* (10, 1, 2) {real, imag} */,
  {32'h44341740, 32'h00000000} /* (10, 1, 1) {real, imag} */,
  {32'h444ff3bc, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h43e1d3eb, 32'h00000000} /* (10, 0, 15) {real, imag} */,
  {32'h43b731cc, 32'h00000000} /* (10, 0, 14) {real, imag} */,
  {32'h43de52b6, 32'h00000000} /* (10, 0, 13) {real, imag} */,
  {32'h43e6ca86, 32'h00000000} /* (10, 0, 12) {real, imag} */,
  {32'h44595e3c, 32'h00000000} /* (10, 0, 11) {real, imag} */,
  {32'h441d9a03, 32'h00000000} /* (10, 0, 10) {real, imag} */,
  {32'hc3353021, 32'h00000000} /* (10, 0, 9) {real, imag} */,
  {32'hc3b79808, 32'h00000000} /* (10, 0, 8) {real, imag} */,
  {32'h43a270d9, 32'h00000000} /* (10, 0, 7) {real, imag} */,
  {32'h406eac00, 32'h00000000} /* (10, 0, 6) {real, imag} */,
  {32'hc22d0db8, 32'h00000000} /* (10, 0, 5) {real, imag} */,
  {32'h440f2b4d, 32'h00000000} /* (10, 0, 4) {real, imag} */,
  {32'h440f09da, 32'h00000000} /* (10, 0, 3) {real, imag} */,
  {32'hc3e5ed49, 32'h00000000} /* (10, 0, 2) {real, imag} */,
  {32'h43d01902, 32'h00000000} /* (10, 0, 1) {real, imag} */,
  {32'h442ec0dc, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h434ccbc8, 32'h00000000} /* (9, 15, 15) {real, imag} */,
  {32'h43de19f5, 32'h00000000} /* (9, 15, 14) {real, imag} */,
  {32'h431c3430, 32'h00000000} /* (9, 15, 13) {real, imag} */,
  {32'h44392eae, 32'h00000000} /* (9, 15, 12) {real, imag} */,
  {32'h43ca783a, 32'h00000000} /* (9, 15, 11) {real, imag} */,
  {32'h3f8fff00, 32'h00000000} /* (9, 15, 10) {real, imag} */,
  {32'hc3d01258, 32'h00000000} /* (9, 15, 9) {real, imag} */,
  {32'hc3552a63, 32'h00000000} /* (9, 15, 8) {real, imag} */,
  {32'h439c7542, 32'h00000000} /* (9, 15, 7) {real, imag} */,
  {32'h43b80809, 32'h00000000} /* (9, 15, 6) {real, imag} */,
  {32'h43abcdb1, 32'h00000000} /* (9, 15, 5) {real, imag} */,
  {32'h430a3c72, 32'h00000000} /* (9, 15, 4) {real, imag} */,
  {32'h435821b1, 32'h00000000} /* (9, 15, 3) {real, imag} */,
  {32'h441eaa96, 32'h00000000} /* (9, 15, 2) {real, imag} */,
  {32'h4256e8ac, 32'h00000000} /* (9, 15, 1) {real, imag} */,
  {32'h4315ac45, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'h437b7b57, 32'h00000000} /* (9, 14, 15) {real, imag} */,
  {32'h4477aca1, 32'h00000000} /* (9, 14, 14) {real, imag} */,
  {32'h449b9caa, 32'h00000000} /* (9, 14, 13) {real, imag} */,
  {32'h44c6f7ca, 32'h00000000} /* (9, 14, 12) {real, imag} */,
  {32'h42dfdfa0, 32'h00000000} /* (9, 14, 11) {real, imag} */,
  {32'h42aac364, 32'h00000000} /* (9, 14, 10) {real, imag} */,
  {32'h44491895, 32'h00000000} /* (9, 14, 9) {real, imag} */,
  {32'hc3a4e285, 32'h00000000} /* (9, 14, 8) {real, imag} */,
  {32'h43a5f1a2, 32'h00000000} /* (9, 14, 7) {real, imag} */,
  {32'h4466b68d, 32'h00000000} /* (9, 14, 6) {real, imag} */,
  {32'h4506525a, 32'h00000000} /* (9, 14, 5) {real, imag} */,
  {32'hc2dd90c0, 32'h00000000} /* (9, 14, 4) {real, imag} */,
  {32'hc43ceaf7, 32'h00000000} /* (9, 14, 3) {real, imag} */,
  {32'hc40bcb52, 32'h00000000} /* (9, 14, 2) {real, imag} */,
  {32'h4247ebf0, 32'h00000000} /* (9, 14, 1) {real, imag} */,
  {32'h430dc796, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hc4141b58, 32'h00000000} /* (9, 13, 15) {real, imag} */,
  {32'h43fb8e7e, 32'h00000000} /* (9, 13, 14) {real, imag} */,
  {32'h44753e81, 32'h00000000} /* (9, 13, 13) {real, imag} */,
  {32'h43169972, 32'h00000000} /* (9, 13, 12) {real, imag} */,
  {32'hc38b102c, 32'h00000000} /* (9, 13, 11) {real, imag} */,
  {32'hc2011b26, 32'h00000000} /* (9, 13, 10) {real, imag} */,
  {32'h43f83ed2, 32'h00000000} /* (9, 13, 9) {real, imag} */,
  {32'h43e7849c, 32'h00000000} /* (9, 13, 8) {real, imag} */,
  {32'h43d6c927, 32'h00000000} /* (9, 13, 7) {real, imag} */,
  {32'h4450519b, 32'h00000000} /* (9, 13, 6) {real, imag} */,
  {32'h4492fc23, 32'h00000000} /* (9, 13, 5) {real, imag} */,
  {32'h43844626, 32'h00000000} /* (9, 13, 4) {real, imag} */,
  {32'hc45bf42a, 32'h00000000} /* (9, 13, 3) {real, imag} */,
  {32'h42659c06, 32'h00000000} /* (9, 13, 2) {real, imag} */,
  {32'h43bafb3a, 32'h00000000} /* (9, 13, 1) {real, imag} */,
  {32'h4407479e, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'h436bc6b4, 32'h00000000} /* (9, 12, 15) {real, imag} */,
  {32'h43144ae0, 32'h00000000} /* (9, 12, 14) {real, imag} */,
  {32'hc42aafd2, 32'h00000000} /* (9, 12, 13) {real, imag} */,
  {32'h42b8682c, 32'h00000000} /* (9, 12, 12) {real, imag} */,
  {32'h441b8172, 32'h00000000} /* (9, 12, 11) {real, imag} */,
  {32'h4409d4f3, 32'h00000000} /* (9, 12, 10) {real, imag} */,
  {32'h447f76f5, 32'h00000000} /* (9, 12, 9) {real, imag} */,
  {32'h44a1e36a, 32'h00000000} /* (9, 12, 8) {real, imag} */,
  {32'h4450c62f, 32'h00000000} /* (9, 12, 7) {real, imag} */,
  {32'h4398a373, 32'h00000000} /* (9, 12, 6) {real, imag} */,
  {32'h443bb0f2, 32'h00000000} /* (9, 12, 5) {real, imag} */,
  {32'h4482f6cb, 32'h00000000} /* (9, 12, 4) {real, imag} */,
  {32'h4309bfe4, 32'h00000000} /* (9, 12, 3) {real, imag} */,
  {32'hc3fa02d6, 32'h00000000} /* (9, 12, 2) {real, imag} */,
  {32'h44090307, 32'h00000000} /* (9, 12, 1) {real, imag} */,
  {32'h44110330, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'h445777de, 32'h00000000} /* (9, 11, 15) {real, imag} */,
  {32'h440a7827, 32'h00000000} /* (9, 11, 14) {real, imag} */,
  {32'h434f11f0, 32'h00000000} /* (9, 11, 13) {real, imag} */,
  {32'hc455ed14, 32'h00000000} /* (9, 11, 12) {real, imag} */,
  {32'hc3d5fde8, 32'h00000000} /* (9, 11, 11) {real, imag} */,
  {32'h447448ab, 32'h00000000} /* (9, 11, 10) {real, imag} */,
  {32'h447cc866, 32'h00000000} /* (9, 11, 9) {real, imag} */,
  {32'h438082e4, 32'h00000000} /* (9, 11, 8) {real, imag} */,
  {32'h4353bd48, 32'h00000000} /* (9, 11, 7) {real, imag} */,
  {32'h4488a3b6, 32'h00000000} /* (9, 11, 6) {real, imag} */,
  {32'h44c4621e, 32'h00000000} /* (9, 11, 5) {real, imag} */,
  {32'h44b26152, 32'h00000000} /* (9, 11, 4) {real, imag} */,
  {32'h44259484, 32'h00000000} /* (9, 11, 3) {real, imag} */,
  {32'h4486cffc, 32'h00000000} /* (9, 11, 2) {real, imag} */,
  {32'h44b9baed, 32'h00000000} /* (9, 11, 1) {real, imag} */,
  {32'h43e2de3a, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h43b5c1a0, 32'h00000000} /* (9, 10, 15) {real, imag} */,
  {32'h44566e90, 32'h00000000} /* (9, 10, 14) {real, imag} */,
  {32'hc333c62e, 32'h00000000} /* (9, 10, 13) {real, imag} */,
  {32'hc3d7bf79, 32'h00000000} /* (9, 10, 12) {real, imag} */,
  {32'hc35a0750, 32'h00000000} /* (9, 10, 11) {real, imag} */,
  {32'hc425ecb4, 32'h00000000} /* (9, 10, 10) {real, imag} */,
  {32'h44d1e1ea, 32'h00000000} /* (9, 10, 9) {real, imag} */,
  {32'h4449e13a, 32'h00000000} /* (9, 10, 8) {real, imag} */,
  {32'h445e477a, 32'h00000000} /* (9, 10, 7) {real, imag} */,
  {32'h4422382a, 32'h00000000} /* (9, 10, 6) {real, imag} */,
  {32'hc3a2b5ed, 32'h00000000} /* (9, 10, 5) {real, imag} */,
  {32'h4483bda0, 32'h00000000} /* (9, 10, 4) {real, imag} */,
  {32'h44467272, 32'h00000000} /* (9, 10, 3) {real, imag} */,
  {32'h449f50a3, 32'h00000000} /* (9, 10, 2) {real, imag} */,
  {32'h44872772, 32'h00000000} /* (9, 10, 1) {real, imag} */,
  {32'h43b6952d, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'h42e62380, 32'h00000000} /* (9, 9, 15) {real, imag} */,
  {32'h442a419e, 32'h00000000} /* (9, 9, 14) {real, imag} */,
  {32'hc2bad2a0, 32'h00000000} /* (9, 9, 13) {real, imag} */,
  {32'hc4876864, 32'h00000000} /* (9, 9, 12) {real, imag} */,
  {32'h43e001c4, 32'h00000000} /* (9, 9, 11) {real, imag} */,
  {32'hc47998b6, 32'h00000000} /* (9, 9, 10) {real, imag} */,
  {32'h4303bbb4, 32'h00000000} /* (9, 9, 9) {real, imag} */,
  {32'h448a21ca, 32'h00000000} /* (9, 9, 8) {real, imag} */,
  {32'h446be6a4, 32'h00000000} /* (9, 9, 7) {real, imag} */,
  {32'h440a248e, 32'h00000000} /* (9, 9, 6) {real, imag} */,
  {32'h43f96498, 32'h00000000} /* (9, 9, 5) {real, imag} */,
  {32'h44379345, 32'h00000000} /* (9, 9, 4) {real, imag} */,
  {32'h448e566f, 32'h00000000} /* (9, 9, 3) {real, imag} */,
  {32'h4445d6b8, 32'h00000000} /* (9, 9, 2) {real, imag} */,
  {32'h449babf4, 32'h00000000} /* (9, 9, 1) {real, imag} */,
  {32'h4490db02, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h43c5cd07, 32'h00000000} /* (9, 8, 15) {real, imag} */,
  {32'h4451e590, 32'h00000000} /* (9, 8, 14) {real, imag} */,
  {32'h42e40a9c, 32'h00000000} /* (9, 8, 13) {real, imag} */,
  {32'h4300da69, 32'h00000000} /* (9, 8, 12) {real, imag} */,
  {32'hc1d8b6f8, 32'h00000000} /* (9, 8, 11) {real, imag} */,
  {32'hc37e9adc, 32'h00000000} /* (9, 8, 10) {real, imag} */,
  {32'hc3581ac0, 32'h00000000} /* (9, 8, 9) {real, imag} */,
  {32'hc32e3387, 32'h00000000} /* (9, 8, 8) {real, imag} */,
  {32'h445f4f9c, 32'h00000000} /* (9, 8, 7) {real, imag} */,
  {32'h44385d7c, 32'h00000000} /* (9, 8, 6) {real, imag} */,
  {32'h441f230e, 32'h00000000} /* (9, 8, 5) {real, imag} */,
  {32'hc3ea93cc, 32'h00000000} /* (9, 8, 4) {real, imag} */,
  {32'h434d6abb, 32'h00000000} /* (9, 8, 3) {real, imag} */,
  {32'h43a9b976, 32'h00000000} /* (9, 8, 2) {real, imag} */,
  {32'h443678b7, 32'h00000000} /* (9, 8, 1) {real, imag} */,
  {32'h441705a8, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h43b787fa, 32'h00000000} /* (9, 7, 15) {real, imag} */,
  {32'h4439b5ed, 32'h00000000} /* (9, 7, 14) {real, imag} */,
  {32'h44709e1a, 32'h00000000} /* (9, 7, 13) {real, imag} */,
  {32'h44b18d55, 32'h00000000} /* (9, 7, 12) {real, imag} */,
  {32'hc3bcbc31, 32'h00000000} /* (9, 7, 11) {real, imag} */,
  {32'hc4961e24, 32'h00000000} /* (9, 7, 10) {real, imag} */,
  {32'hc2519714, 32'h00000000} /* (9, 7, 9) {real, imag} */,
  {32'h431f07e5, 32'h00000000} /* (9, 7, 8) {real, imag} */,
  {32'h438d1b5e, 32'h00000000} /* (9, 7, 7) {real, imag} */,
  {32'h44291127, 32'h00000000} /* (9, 7, 6) {real, imag} */,
  {32'h43ee4844, 32'h00000000} /* (9, 7, 5) {real, imag} */,
  {32'hc3467bf0, 32'h00000000} /* (9, 7, 4) {real, imag} */,
  {32'h43350086, 32'h00000000} /* (9, 7, 3) {real, imag} */,
  {32'h4347c6f6, 32'h00000000} /* (9, 7, 2) {real, imag} */,
  {32'hc3a7d1ec, 32'h00000000} /* (9, 7, 1) {real, imag} */,
  {32'h430def8b, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h4425873a, 32'h00000000} /* (9, 6, 15) {real, imag} */,
  {32'h44068821, 32'h00000000} /* (9, 6, 14) {real, imag} */,
  {32'h4465a2bf, 32'h00000000} /* (9, 6, 13) {real, imag} */,
  {32'h441e17ab, 32'h00000000} /* (9, 6, 12) {real, imag} */,
  {32'hc327a625, 32'h00000000} /* (9, 6, 11) {real, imag} */,
  {32'hc4428cf9, 32'h00000000} /* (9, 6, 10) {real, imag} */,
  {32'h441207a2, 32'h00000000} /* (9, 6, 9) {real, imag} */,
  {32'hc474a336, 32'h00000000} /* (9, 6, 8) {real, imag} */,
  {32'hc3271a18, 32'h00000000} /* (9, 6, 7) {real, imag} */,
  {32'h44807185, 32'h00000000} /* (9, 6, 6) {real, imag} */,
  {32'h443bf79d, 32'h00000000} /* (9, 6, 5) {real, imag} */,
  {32'h4404be3f, 32'h00000000} /* (9, 6, 4) {real, imag} */,
  {32'hc3ef6906, 32'h00000000} /* (9, 6, 3) {real, imag} */,
  {32'hc45f9d1d, 32'h00000000} /* (9, 6, 2) {real, imag} */,
  {32'h43fbecd3, 32'h00000000} /* (9, 6, 1) {real, imag} */,
  {32'h4216cac0, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'h441838de, 32'h00000000} /* (9, 5, 15) {real, imag} */,
  {32'h440e2bf9, 32'h00000000} /* (9, 5, 14) {real, imag} */,
  {32'hc2f9ca10, 32'h00000000} /* (9, 5, 13) {real, imag} */,
  {32'h440326b2, 32'h00000000} /* (9, 5, 12) {real, imag} */,
  {32'hc3666194, 32'h00000000} /* (9, 5, 11) {real, imag} */,
  {32'h4298f285, 32'h00000000} /* (9, 5, 10) {real, imag} */,
  {32'h4301c48c, 32'h00000000} /* (9, 5, 9) {real, imag} */,
  {32'hc3dd3f59, 32'h00000000} /* (9, 5, 8) {real, imag} */,
  {32'h43493f9f, 32'h00000000} /* (9, 5, 7) {real, imag} */,
  {32'h44d35fda, 32'h00000000} /* (9, 5, 6) {real, imag} */,
  {32'h44d024ab, 32'h00000000} /* (9, 5, 5) {real, imag} */,
  {32'h43da0e98, 32'h00000000} /* (9, 5, 4) {real, imag} */,
  {32'hc32fd5fc, 32'h00000000} /* (9, 5, 3) {real, imag} */,
  {32'hc220378a, 32'h00000000} /* (9, 5, 2) {real, imag} */,
  {32'hc4120abc, 32'h00000000} /* (9, 5, 1) {real, imag} */,
  {32'hc19b9830, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'hc288e2e5, 32'h00000000} /* (9, 4, 15) {real, imag} */,
  {32'hc2c4dfd0, 32'h00000000} /* (9, 4, 14) {real, imag} */,
  {32'h4405fd10, 32'h00000000} /* (9, 4, 13) {real, imag} */,
  {32'h438bb57c, 32'h00000000} /* (9, 4, 12) {real, imag} */,
  {32'hc3687838, 32'h00000000} /* (9, 4, 11) {real, imag} */,
  {32'hc4b3acca, 32'h00000000} /* (9, 4, 10) {real, imag} */,
  {32'hc48bdc1e, 32'h00000000} /* (9, 4, 9) {real, imag} */,
  {32'hc42c3d38, 32'h00000000} /* (9, 4, 8) {real, imag} */,
  {32'hc3300d46, 32'h00000000} /* (9, 4, 7) {real, imag} */,
  {32'h44b5ef5e, 32'h00000000} /* (9, 4, 6) {real, imag} */,
  {32'h44287cc8, 32'h00000000} /* (9, 4, 5) {real, imag} */,
  {32'h448fe5e3, 32'h00000000} /* (9, 4, 4) {real, imag} */,
  {32'h441299ee, 32'h00000000} /* (9, 4, 3) {real, imag} */,
  {32'hc2f7f678, 32'h00000000} /* (9, 4, 2) {real, imag} */,
  {32'hc456c983, 32'h00000000} /* (9, 4, 1) {real, imag} */,
  {32'hc28853c4, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'hc3e766de, 32'h00000000} /* (9, 3, 15) {real, imag} */,
  {32'hc33da3e4, 32'h00000000} /* (9, 3, 14) {real, imag} */,
  {32'hc480681a, 32'h00000000} /* (9, 3, 13) {real, imag} */,
  {32'hc4040a67, 32'h00000000} /* (9, 3, 12) {real, imag} */,
  {32'hc2f63efb, 32'h00000000} /* (9, 3, 11) {real, imag} */,
  {32'hc4da07f2, 32'h00000000} /* (9, 3, 10) {real, imag} */,
  {32'h443800c5, 32'h00000000} /* (9, 3, 9) {real, imag} */,
  {32'hc336ca84, 32'h00000000} /* (9, 3, 8) {real, imag} */,
  {32'h43443694, 32'h00000000} /* (9, 3, 7) {real, imag} */,
  {32'hc2ee8440, 32'h00000000} /* (9, 3, 6) {real, imag} */,
  {32'h4394b00e, 32'h00000000} /* (9, 3, 5) {real, imag} */,
  {32'h42b4b57e, 32'h00000000} /* (9, 3, 4) {real, imag} */,
  {32'hc3a0d9eb, 32'h00000000} /* (9, 3, 3) {real, imag} */,
  {32'hc318ca50, 32'h00000000} /* (9, 3, 2) {real, imag} */,
  {32'h4428e521, 32'h00000000} /* (9, 3, 1) {real, imag} */,
  {32'hc1e35730, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'hc31e2b2f, 32'h00000000} /* (9, 2, 15) {real, imag} */,
  {32'hc37121dc, 32'h00000000} /* (9, 2, 14) {real, imag} */,
  {32'hc49e1238, 32'h00000000} /* (9, 2, 13) {real, imag} */,
  {32'hc45ea23e, 32'h00000000} /* (9, 2, 12) {real, imag} */,
  {32'hc3eeeecc, 32'h00000000} /* (9, 2, 11) {real, imag} */,
  {32'h43f2c7e4, 32'h00000000} /* (9, 2, 10) {real, imag} */,
  {32'hc4836534, 32'h00000000} /* (9, 2, 9) {real, imag} */,
  {32'h43729f18, 32'h00000000} /* (9, 2, 8) {real, imag} */,
  {32'h43c81b84, 32'h00000000} /* (9, 2, 7) {real, imag} */,
  {32'h43abf93e, 32'h00000000} /* (9, 2, 6) {real, imag} */,
  {32'h435647b0, 32'h00000000} /* (9, 2, 5) {real, imag} */,
  {32'h43897f5b, 32'h00000000} /* (9, 2, 4) {real, imag} */,
  {32'hc1926d88, 32'h00000000} /* (9, 2, 3) {real, imag} */,
  {32'h410de3f0, 32'h00000000} /* (9, 2, 2) {real, imag} */,
  {32'h4484cebe, 32'h00000000} /* (9, 2, 1) {real, imag} */,
  {32'hc0e738d0, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'hc3eeab46, 32'h00000000} /* (9, 1, 15) {real, imag} */,
  {32'hc2bed128, 32'h00000000} /* (9, 1, 14) {real, imag} */,
  {32'hc3079354, 32'h00000000} /* (9, 1, 13) {real, imag} */,
  {32'hc348bb88, 32'h00000000} /* (9, 1, 12) {real, imag} */,
  {32'h4469f6d8, 32'h00000000} /* (9, 1, 11) {real, imag} */,
  {32'hc3518b3e, 32'h00000000} /* (9, 1, 10) {real, imag} */,
  {32'hc2307700, 32'h00000000} /* (9, 1, 9) {real, imag} */,
  {32'h443b6a37, 32'h00000000} /* (9, 1, 8) {real, imag} */,
  {32'h4427cafd, 32'h00000000} /* (9, 1, 7) {real, imag} */,
  {32'h43d3e1f0, 32'h00000000} /* (9, 1, 6) {real, imag} */,
  {32'hc400b4cf, 32'h00000000} /* (9, 1, 5) {real, imag} */,
  {32'h44cc0598, 32'h00000000} /* (9, 1, 4) {real, imag} */,
  {32'h44491a0e, 32'h00000000} /* (9, 1, 3) {real, imag} */,
  {32'hc48c78be, 32'h00000000} /* (9, 1, 2) {real, imag} */,
  {32'hc1b72df0, 32'h00000000} /* (9, 1, 1) {real, imag} */,
  {32'h42a18718, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'h43e491f8, 32'h00000000} /* (9, 0, 15) {real, imag} */,
  {32'hc35e7d26, 32'h00000000} /* (9, 0, 14) {real, imag} */,
  {32'hc3569f5c, 32'h00000000} /* (9, 0, 13) {real, imag} */,
  {32'h43896266, 32'h00000000} /* (9, 0, 12) {real, imag} */,
  {32'h431174ba, 32'h00000000} /* (9, 0, 11) {real, imag} */,
  {32'h439eda9e, 32'h00000000} /* (9, 0, 10) {real, imag} */,
  {32'hc255b086, 32'h00000000} /* (9, 0, 9) {real, imag} */,
  {32'hc14a83c0, 32'h00000000} /* (9, 0, 8) {real, imag} */,
  {32'h43d88560, 32'h00000000} /* (9, 0, 7) {real, imag} */,
  {32'h43996d1b, 32'h00000000} /* (9, 0, 6) {real, imag} */,
  {32'h42dfffb8, 32'h00000000} /* (9, 0, 5) {real, imag} */,
  {32'h4353f34f, 32'h00000000} /* (9, 0, 4) {real, imag} */,
  {32'hc25d7490, 32'h00000000} /* (9, 0, 3) {real, imag} */,
  {32'h417c4d10, 32'h00000000} /* (9, 0, 2) {real, imag} */,
  {32'hc31b2c50, 32'h00000000} /* (9, 0, 1) {real, imag} */,
  {32'hc3677cd8, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h432a90df, 32'h00000000} /* (8, 15, 15) {real, imag} */,
  {32'hc2a573f7, 32'h00000000} /* (8, 15, 14) {real, imag} */,
  {32'h4323c5e7, 32'h00000000} /* (8, 15, 13) {real, imag} */,
  {32'hc0fe3660, 32'h00000000} /* (8, 15, 12) {real, imag} */,
  {32'h4412adf3, 32'h00000000} /* (8, 15, 11) {real, imag} */,
  {32'h43c322a6, 32'h00000000} /* (8, 15, 10) {real, imag} */,
  {32'h437505b0, 32'h00000000} /* (8, 15, 9) {real, imag} */,
  {32'hc3f9b385, 32'h00000000} /* (8, 15, 8) {real, imag} */,
  {32'hc3d57e20, 32'h00000000} /* (8, 15, 7) {real, imag} */,
  {32'h431065ee, 32'h00000000} /* (8, 15, 6) {real, imag} */,
  {32'h4285eb00, 32'h00000000} /* (8, 15, 5) {real, imag} */,
  {32'h4275192c, 32'h00000000} /* (8, 15, 4) {real, imag} */,
  {32'hc3e9abea, 32'h00000000} /* (8, 15, 3) {real, imag} */,
  {32'hc40cb35e, 32'h00000000} /* (8, 15, 2) {real, imag} */,
  {32'h437305bc, 32'h00000000} /* (8, 15, 1) {real, imag} */,
  {32'h422626f8, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'h43bbf860, 32'h00000000} /* (8, 14, 15) {real, imag} */,
  {32'h4412b85b, 32'h00000000} /* (8, 14, 14) {real, imag} */,
  {32'hc2d705d0, 32'h00000000} /* (8, 14, 13) {real, imag} */,
  {32'h435b3e28, 32'h00000000} /* (8, 14, 12) {real, imag} */,
  {32'h442a210c, 32'h00000000} /* (8, 14, 11) {real, imag} */,
  {32'hc3c47846, 32'h00000000} /* (8, 14, 10) {real, imag} */,
  {32'hc3838aa8, 32'h00000000} /* (8, 14, 9) {real, imag} */,
  {32'h42213c40, 32'h00000000} /* (8, 14, 8) {real, imag} */,
  {32'hc39fff82, 32'h00000000} /* (8, 14, 7) {real, imag} */,
  {32'h43e01832, 32'h00000000} /* (8, 14, 6) {real, imag} */,
  {32'h43b4c34b, 32'h00000000} /* (8, 14, 5) {real, imag} */,
  {32'hc470bac6, 32'h00000000} /* (8, 14, 4) {real, imag} */,
  {32'h42cb6770, 32'h00000000} /* (8, 14, 3) {real, imag} */,
  {32'hc2ab377a, 32'h00000000} /* (8, 14, 2) {real, imag} */,
  {32'hc415432c, 32'h00000000} /* (8, 14, 1) {real, imag} */,
  {32'hc0f548c0, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'h4310adf3, 32'h00000000} /* (8, 13, 15) {real, imag} */,
  {32'hc43604ee, 32'h00000000} /* (8, 13, 14) {real, imag} */,
  {32'hc3c58860, 32'h00000000} /* (8, 13, 13) {real, imag} */,
  {32'h44067c3b, 32'h00000000} /* (8, 13, 12) {real, imag} */,
  {32'hc2979a0c, 32'h00000000} /* (8, 13, 11) {real, imag} */,
  {32'hc36fa6e8, 32'h00000000} /* (8, 13, 10) {real, imag} */,
  {32'h4470e76c, 32'h00000000} /* (8, 13, 9) {real, imag} */,
  {32'h437c5517, 32'h00000000} /* (8, 13, 8) {real, imag} */,
  {32'hc37eec07, 32'h00000000} /* (8, 13, 7) {real, imag} */,
  {32'h445a48e8, 32'h00000000} /* (8, 13, 6) {real, imag} */,
  {32'h448bafae, 32'h00000000} /* (8, 13, 5) {real, imag} */,
  {32'h440b9491, 32'h00000000} /* (8, 13, 4) {real, imag} */,
  {32'hc4656262, 32'h00000000} /* (8, 13, 3) {real, imag} */,
  {32'h415d2298, 32'h00000000} /* (8, 13, 2) {real, imag} */,
  {32'hc24ac178, 32'h00000000} /* (8, 13, 1) {real, imag} */,
  {32'h43bc50f6, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'h41b9d0c4, 32'h00000000} /* (8, 12, 15) {real, imag} */,
  {32'h4195c268, 32'h00000000} /* (8, 12, 14) {real, imag} */,
  {32'h4388cd20, 32'h00000000} /* (8, 12, 13) {real, imag} */,
  {32'hc1acd2c8, 32'h00000000} /* (8, 12, 12) {real, imag} */,
  {32'hc3b3707e, 32'h00000000} /* (8, 12, 11) {real, imag} */,
  {32'h4412d025, 32'h00000000} /* (8, 12, 10) {real, imag} */,
  {32'h4434eb4b, 32'h00000000} /* (8, 12, 9) {real, imag} */,
  {32'h42ca13d7, 32'h00000000} /* (8, 12, 8) {real, imag} */,
  {32'h43887e54, 32'h00000000} /* (8, 12, 7) {real, imag} */,
  {32'h430deef3, 32'h00000000} /* (8, 12, 6) {real, imag} */,
  {32'hc3949ee4, 32'h00000000} /* (8, 12, 5) {real, imag} */,
  {32'h43922b6e, 32'h00000000} /* (8, 12, 4) {real, imag} */,
  {32'h44155059, 32'h00000000} /* (8, 12, 3) {real, imag} */,
  {32'h440153a5, 32'h00000000} /* (8, 12, 2) {real, imag} */,
  {32'h4393361a, 32'h00000000} /* (8, 12, 1) {real, imag} */,
  {32'h43493298, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'h4401399f, 32'h00000000} /* (8, 11, 15) {real, imag} */,
  {32'h43b95182, 32'h00000000} /* (8, 11, 14) {real, imag} */,
  {32'hc2982be4, 32'h00000000} /* (8, 11, 13) {real, imag} */,
  {32'hc49fa178, 32'h00000000} /* (8, 11, 12) {real, imag} */,
  {32'hc4122b41, 32'h00000000} /* (8, 11, 11) {real, imag} */,
  {32'h438dc63a, 32'h00000000} /* (8, 11, 10) {real, imag} */,
  {32'h448c03c4, 32'h00000000} /* (8, 11, 9) {real, imag} */,
  {32'h431a97c1, 32'h00000000} /* (8, 11, 8) {real, imag} */,
  {32'h43e6568e, 32'h00000000} /* (8, 11, 7) {real, imag} */,
  {32'hc34de438, 32'h00000000} /* (8, 11, 6) {real, imag} */,
  {32'hc34df7be, 32'h00000000} /* (8, 11, 5) {real, imag} */,
  {32'h43f74be3, 32'h00000000} /* (8, 11, 4) {real, imag} */,
  {32'h445abff3, 32'h00000000} /* (8, 11, 3) {real, imag} */,
  {32'h434461ff, 32'h00000000} /* (8, 11, 2) {real, imag} */,
  {32'h43a45857, 32'h00000000} /* (8, 11, 1) {real, imag} */,
  {32'h433724f3, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h439444d3, 32'h00000000} /* (8, 10, 15) {real, imag} */,
  {32'hc3c7c894, 32'h00000000} /* (8, 10, 14) {real, imag} */,
  {32'h4367c6fa, 32'h00000000} /* (8, 10, 13) {real, imag} */,
  {32'hc42138ec, 32'h00000000} /* (8, 10, 12) {real, imag} */,
  {32'hc3c82efc, 32'h00000000} /* (8, 10, 11) {real, imag} */,
  {32'hc2f566e8, 32'h00000000} /* (8, 10, 10) {real, imag} */,
  {32'h44377610, 32'h00000000} /* (8, 10, 9) {real, imag} */,
  {32'h44948f96, 32'h00000000} /* (8, 10, 8) {real, imag} */,
  {32'hc37f9baa, 32'h00000000} /* (8, 10, 7) {real, imag} */,
  {32'h449b6db2, 32'h00000000} /* (8, 10, 6) {real, imag} */,
  {32'h442decd0, 32'h00000000} /* (8, 10, 5) {real, imag} */,
  {32'h43c482dc, 32'h00000000} /* (8, 10, 4) {real, imag} */,
  {32'h4478feb0, 32'h00000000} /* (8, 10, 3) {real, imag} */,
  {32'h44997640, 32'h00000000} /* (8, 10, 2) {real, imag} */,
  {32'h4472f5ca, 32'h00000000} /* (8, 10, 1) {real, imag} */,
  {32'h43c4c919, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'h42358120, 32'h00000000} /* (8, 9, 15) {real, imag} */,
  {32'h4283cf24, 32'h00000000} /* (8, 9, 14) {real, imag} */,
  {32'h4305fdca, 32'h00000000} /* (8, 9, 13) {real, imag} */,
  {32'hc2d540d8, 32'h00000000} /* (8, 9, 12) {real, imag} */,
  {32'hc1818560, 32'h00000000} /* (8, 9, 11) {real, imag} */,
  {32'h4391174a, 32'h00000000} /* (8, 9, 10) {real, imag} */,
  {32'h413e5c60, 32'h00000000} /* (8, 9, 9) {real, imag} */,
  {32'h431697c4, 32'h00000000} /* (8, 9, 8) {real, imag} */,
  {32'h43bde2b0, 32'h00000000} /* (8, 9, 7) {real, imag} */,
  {32'h446d4874, 32'h00000000} /* (8, 9, 6) {real, imag} */,
  {32'h442a9860, 32'h00000000} /* (8, 9, 5) {real, imag} */,
  {32'h44930056, 32'h00000000} /* (8, 9, 4) {real, imag} */,
  {32'h441323d6, 32'h00000000} /* (8, 9, 3) {real, imag} */,
  {32'h438ef324, 32'h00000000} /* (8, 9, 2) {real, imag} */,
  {32'h4457f90c, 32'h00000000} /* (8, 9, 1) {real, imag} */,
  {32'h42d24ad8, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'hc10034c0, 32'h00000000} /* (8, 8, 15) {real, imag} */,
  {32'hc1a79f78, 32'h00000000} /* (8, 8, 14) {real, imag} */,
  {32'h44712622, 32'h00000000} /* (8, 8, 13) {real, imag} */,
  {32'h43e73614, 32'h00000000} /* (8, 8, 12) {real, imag} */,
  {32'h42a0e734, 32'h00000000} /* (8, 8, 11) {real, imag} */,
  {32'hc3d14759, 32'h00000000} /* (8, 8, 10) {real, imag} */,
  {32'hc4a3b3d8, 32'h00000000} /* (8, 8, 9) {real, imag} */,
  {32'h4307b56c, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'h43b7e310, 32'h00000000} /* (8, 8, 7) {real, imag} */,
  {32'h438423a2, 32'h00000000} /* (8, 8, 6) {real, imag} */,
  {32'h4430e470, 32'h00000000} /* (8, 8, 5) {real, imag} */,
  {32'hc3ce89d6, 32'h00000000} /* (8, 8, 4) {real, imag} */,
  {32'hc456edaa, 32'h00000000} /* (8, 8, 3) {real, imag} */,
  {32'hc36f47de, 32'h00000000} /* (8, 8, 2) {real, imag} */,
  {32'h443e9523, 32'h00000000} /* (8, 8, 1) {real, imag} */,
  {32'h43be990c, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h436e75ef, 32'h00000000} /* (8, 7, 15) {real, imag} */,
  {32'h44087502, 32'h00000000} /* (8, 7, 14) {real, imag} */,
  {32'h43476e44, 32'h00000000} /* (8, 7, 13) {real, imag} */,
  {32'h44bf8906, 32'h00000000} /* (8, 7, 12) {real, imag} */,
  {32'h4367212b, 32'h00000000} /* (8, 7, 11) {real, imag} */,
  {32'h43707be0, 32'h00000000} /* (8, 7, 10) {real, imag} */,
  {32'hc17803e0, 32'h00000000} /* (8, 7, 9) {real, imag} */,
  {32'h437a9e41, 32'h00000000} /* (8, 7, 8) {real, imag} */,
  {32'h443b30fe, 32'h00000000} /* (8, 7, 7) {real, imag} */,
  {32'h444f275c, 32'h00000000} /* (8, 7, 6) {real, imag} */,
  {32'hc3624ea6, 32'h00000000} /* (8, 7, 5) {real, imag} */,
  {32'hc361eca0, 32'h00000000} /* (8, 7, 4) {real, imag} */,
  {32'hc3a6ad72, 32'h00000000} /* (8, 7, 3) {real, imag} */,
  {32'hc40c9866, 32'h00000000} /* (8, 7, 2) {real, imag} */,
  {32'hc3ca7f05, 32'h00000000} /* (8, 7, 1) {real, imag} */,
  {32'h437b1d2b, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h432b53db, 32'h00000000} /* (8, 6, 15) {real, imag} */,
  {32'h437d37c1, 32'h00000000} /* (8, 6, 14) {real, imag} */,
  {32'hc307eafc, 32'h00000000} /* (8, 6, 13) {real, imag} */,
  {32'h423e19d0, 32'h00000000} /* (8, 6, 12) {real, imag} */,
  {32'h44291eb5, 32'h00000000} /* (8, 6, 11) {real, imag} */,
  {32'hc456ff7a, 32'h00000000} /* (8, 6, 10) {real, imag} */,
  {32'hc3ff5d3e, 32'h00000000} /* (8, 6, 9) {real, imag} */,
  {32'h436f5418, 32'h00000000} /* (8, 6, 8) {real, imag} */,
  {32'hc40241a9, 32'h00000000} /* (8, 6, 7) {real, imag} */,
  {32'h4431d6e8, 32'h00000000} /* (8, 6, 6) {real, imag} */,
  {32'h44a67a88, 32'h00000000} /* (8, 6, 5) {real, imag} */,
  {32'h43c797be, 32'h00000000} /* (8, 6, 4) {real, imag} */,
  {32'hc4350c57, 32'h00000000} /* (8, 6, 3) {real, imag} */,
  {32'hc3b2eadc, 32'h00000000} /* (8, 6, 2) {real, imag} */,
  {32'h42c940ce, 32'h00000000} /* (8, 6, 1) {real, imag} */,
  {32'hc3eded9c, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'hc2d1f25c, 32'h00000000} /* (8, 5, 15) {real, imag} */,
  {32'h43fa43d2, 32'h00000000} /* (8, 5, 14) {real, imag} */,
  {32'h434e7e7a, 32'h00000000} /* (8, 5, 13) {real, imag} */,
  {32'h43d7ca89, 32'h00000000} /* (8, 5, 12) {real, imag} */,
  {32'hc36167a9, 32'h00000000} /* (8, 5, 11) {real, imag} */,
  {32'hc3e9ff3b, 32'h00000000} /* (8, 5, 10) {real, imag} */,
  {32'hc3b596ab, 32'h00000000} /* (8, 5, 9) {real, imag} */,
  {32'hc4214d9b, 32'h00000000} /* (8, 5, 8) {real, imag} */,
  {32'h42c5a452, 32'h00000000} /* (8, 5, 7) {real, imag} */,
  {32'h4478837d, 32'h00000000} /* (8, 5, 6) {real, imag} */,
  {32'h4491a366, 32'h00000000} /* (8, 5, 5) {real, imag} */,
  {32'h445231d4, 32'h00000000} /* (8, 5, 4) {real, imag} */,
  {32'hc00250c0, 32'h00000000} /* (8, 5, 3) {real, imag} */,
  {32'hc3863809, 32'h00000000} /* (8, 5, 2) {real, imag} */,
  {32'hc3b5d989, 32'h00000000} /* (8, 5, 1) {real, imag} */,
  {32'hc2e92448, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'hc42b6267, 32'h00000000} /* (8, 4, 15) {real, imag} */,
  {32'h44865af0, 32'h00000000} /* (8, 4, 14) {real, imag} */,
  {32'h4451a8e6, 32'h00000000} /* (8, 4, 13) {real, imag} */,
  {32'hc3454c20, 32'h00000000} /* (8, 4, 12) {real, imag} */,
  {32'hc436fa3d, 32'h00000000} /* (8, 4, 11) {real, imag} */,
  {32'hc3b522e4, 32'h00000000} /* (8, 4, 10) {real, imag} */,
  {32'h43493651, 32'h00000000} /* (8, 4, 9) {real, imag} */,
  {32'hc333b78e, 32'h00000000} /* (8, 4, 8) {real, imag} */,
  {32'h446bda9b, 32'h00000000} /* (8, 4, 7) {real, imag} */,
  {32'h445756dd, 32'h00000000} /* (8, 4, 6) {real, imag} */,
  {32'h4391c25c, 32'h00000000} /* (8, 4, 5) {real, imag} */,
  {32'h44717e34, 32'h00000000} /* (8, 4, 4) {real, imag} */,
  {32'h442e7241, 32'h00000000} /* (8, 4, 3) {real, imag} */,
  {32'hc435c878, 32'h00000000} /* (8, 4, 2) {real, imag} */,
  {32'hc3ff4cc2, 32'h00000000} /* (8, 4, 1) {real, imag} */,
  {32'hc34f2ada, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'hc31346ba, 32'h00000000} /* (8, 3, 15) {real, imag} */,
  {32'hc397f57d, 32'h00000000} /* (8, 3, 14) {real, imag} */,
  {32'hc480aef6, 32'h00000000} /* (8, 3, 13) {real, imag} */,
  {32'h43fba9bf, 32'h00000000} /* (8, 3, 12) {real, imag} */,
  {32'hc3521f56, 32'h00000000} /* (8, 3, 11) {real, imag} */,
  {32'hc456b928, 32'h00000000} /* (8, 3, 10) {real, imag} */,
  {32'hc3f4a1de, 32'h00000000} /* (8, 3, 9) {real, imag} */,
  {32'h4316f440, 32'h00000000} /* (8, 3, 8) {real, imag} */,
  {32'h44533cb2, 32'h00000000} /* (8, 3, 7) {real, imag} */,
  {32'h4499460e, 32'h00000000} /* (8, 3, 6) {real, imag} */,
  {32'h445c066d, 32'h00000000} /* (8, 3, 5) {real, imag} */,
  {32'h42e31c9c, 32'h00000000} /* (8, 3, 4) {real, imag} */,
  {32'h41beabac, 32'h00000000} /* (8, 3, 3) {real, imag} */,
  {32'h428750e4, 32'h00000000} /* (8, 3, 2) {real, imag} */,
  {32'hc39bfc2e, 32'h00000000} /* (8, 3, 1) {real, imag} */,
  {32'hc3d41412, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'hc345d993, 32'h00000000} /* (8, 2, 15) {real, imag} */,
  {32'hc416499c, 32'h00000000} /* (8, 2, 14) {real, imag} */,
  {32'hc4c85531, 32'h00000000} /* (8, 2, 13) {real, imag} */,
  {32'hc4710957, 32'h00000000} /* (8, 2, 12) {real, imag} */,
  {32'hc3238ec6, 32'h00000000} /* (8, 2, 11) {real, imag} */,
  {32'hc3c7717c, 32'h00000000} /* (8, 2, 10) {real, imag} */,
  {32'hc312bdf8, 32'h00000000} /* (8, 2, 9) {real, imag} */,
  {32'hc384f499, 32'h00000000} /* (8, 2, 8) {real, imag} */,
  {32'hc38d5622, 32'h00000000} /* (8, 2, 7) {real, imag} */,
  {32'h44b68d4e, 32'h00000000} /* (8, 2, 6) {real, imag} */,
  {32'h4453cc9e, 32'h00000000} /* (8, 2, 5) {real, imag} */,
  {32'h44544c1b, 32'h00000000} /* (8, 2, 4) {real, imag} */,
  {32'h43457800, 32'h00000000} /* (8, 2, 3) {real, imag} */,
  {32'hc2d5ab14, 32'h00000000} /* (8, 2, 2) {real, imag} */,
  {32'hc436c945, 32'h00000000} /* (8, 2, 1) {real, imag} */,
  {32'hc4005062, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'hc3a4cb93, 32'h00000000} /* (8, 1, 15) {real, imag} */,
  {32'hc43eeda6, 32'h00000000} /* (8, 1, 14) {real, imag} */,
  {32'hc4462954, 32'h00000000} /* (8, 1, 13) {real, imag} */,
  {32'h4402d2fa, 32'h00000000} /* (8, 1, 12) {real, imag} */,
  {32'hc4583391, 32'h00000000} /* (8, 1, 11) {real, imag} */,
  {32'hc426d617, 32'h00000000} /* (8, 1, 10) {real, imag} */,
  {32'h44a08f06, 32'h00000000} /* (8, 1, 9) {real, imag} */,
  {32'hc2b1b45c, 32'h00000000} /* (8, 1, 8) {real, imag} */,
  {32'h437f23ba, 32'h00000000} /* (8, 1, 7) {real, imag} */,
  {32'h44750af8, 32'h00000000} /* (8, 1, 6) {real, imag} */,
  {32'h444bb082, 32'h00000000} /* (8, 1, 5) {real, imag} */,
  {32'h42dfc754, 32'h00000000} /* (8, 1, 4) {real, imag} */,
  {32'hc3a4d976, 32'h00000000} /* (8, 1, 3) {real, imag} */,
  {32'hc347d2bb, 32'h00000000} /* (8, 1, 2) {real, imag} */,
  {32'hc413d5ec, 32'h00000000} /* (8, 1, 1) {real, imag} */,
  {32'hc4381a84, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'hc3ff39c5, 32'h00000000} /* (8, 0, 15) {real, imag} */,
  {32'hc35e5a62, 32'h00000000} /* (8, 0, 14) {real, imag} */,
  {32'h43bef58f, 32'h00000000} /* (8, 0, 13) {real, imag} */,
  {32'h434ddb8f, 32'h00000000} /* (8, 0, 12) {real, imag} */,
  {32'hc3ae6536, 32'h00000000} /* (8, 0, 11) {real, imag} */,
  {32'hc3311a8d, 32'h00000000} /* (8, 0, 10) {real, imag} */,
  {32'h4360df98, 32'h00000000} /* (8, 0, 9) {real, imag} */,
  {32'h44240074, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'h44302bda, 32'h00000000} /* (8, 0, 7) {real, imag} */,
  {32'h44135470, 32'h00000000} /* (8, 0, 6) {real, imag} */,
  {32'h4433ae00, 32'h00000000} /* (8, 0, 5) {real, imag} */,
  {32'h42ff67ba, 32'h00000000} /* (8, 0, 4) {real, imag} */,
  {32'hc27a7dfc, 32'h00000000} /* (8, 0, 3) {real, imag} */,
  {32'hc2011490, 32'h00000000} /* (8, 0, 2) {real, imag} */,
  {32'hc427ab5b, 32'h00000000} /* (8, 0, 1) {real, imag} */,
  {32'hc3c02e89, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h420f8560, 32'h00000000} /* (7, 15, 15) {real, imag} */,
  {32'hc140d7a0, 32'h00000000} /* (7, 15, 14) {real, imag} */,
  {32'hc35bc94c, 32'h00000000} /* (7, 15, 13) {real, imag} */,
  {32'hc419ff78, 32'h00000000} /* (7, 15, 12) {real, imag} */,
  {32'hc2b61888, 32'h00000000} /* (7, 15, 11) {real, imag} */,
  {32'hc3a44bea, 32'h00000000} /* (7, 15, 10) {real, imag} */,
  {32'hc3ae4839, 32'h00000000} /* (7, 15, 9) {real, imag} */,
  {32'hc3b0ed7e, 32'h00000000} /* (7, 15, 8) {real, imag} */,
  {32'h4403dd34, 32'h00000000} /* (7, 15, 7) {real, imag} */,
  {32'h4451cd58, 32'h00000000} /* (7, 15, 6) {real, imag} */,
  {32'h438536c0, 32'h00000000} /* (7, 15, 5) {real, imag} */,
  {32'hc451a09e, 32'h00000000} /* (7, 15, 4) {real, imag} */,
  {32'hc42bf6cd, 32'h00000000} /* (7, 15, 3) {real, imag} */,
  {32'hc40bddb9, 32'h00000000} /* (7, 15, 2) {real, imag} */,
  {32'hc2cacc14, 32'h00000000} /* (7, 15, 1) {real, imag} */,
  {32'hc3bd491e, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'h43910316, 32'h00000000} /* (7, 14, 15) {real, imag} */,
  {32'h41f7a368, 32'h00000000} /* (7, 14, 14) {real, imag} */,
  {32'hc44f56b4, 32'h00000000} /* (7, 14, 13) {real, imag} */,
  {32'hc4838754, 32'h00000000} /* (7, 14, 12) {real, imag} */,
  {32'hc307442a, 32'h00000000} /* (7, 14, 11) {real, imag} */,
  {32'hc478e76a, 32'h00000000} /* (7, 14, 10) {real, imag} */,
  {32'hc45712bc, 32'h00000000} /* (7, 14, 9) {real, imag} */,
  {32'h430f5b44, 32'h00000000} /* (7, 14, 8) {real, imag} */,
  {32'h43436a0e, 32'h00000000} /* (7, 14, 7) {real, imag} */,
  {32'h43c736bc, 32'h00000000} /* (7, 14, 6) {real, imag} */,
  {32'h4444d490, 32'h00000000} /* (7, 14, 5) {real, imag} */,
  {32'hc46deda4, 32'h00000000} /* (7, 14, 4) {real, imag} */,
  {32'hc3ab9010, 32'h00000000} /* (7, 14, 3) {real, imag} */,
  {32'hc2b083d0, 32'h00000000} /* (7, 14, 2) {real, imag} */,
  {32'h41216200, 32'h00000000} /* (7, 14, 1) {real, imag} */,
  {32'h428ff0d1, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hc38e2a36, 32'h00000000} /* (7, 13, 15) {real, imag} */,
  {32'hc2cfd5b0, 32'h00000000} /* (7, 13, 14) {real, imag} */,
  {32'hc3f8d18a, 32'h00000000} /* (7, 13, 13) {real, imag} */,
  {32'h43f009f5, 32'h00000000} /* (7, 13, 12) {real, imag} */,
  {32'h42162bb2, 32'h00000000} /* (7, 13, 11) {real, imag} */,
  {32'hc3e98f5f, 32'h00000000} /* (7, 13, 10) {real, imag} */,
  {32'h44711131, 32'h00000000} /* (7, 13, 9) {real, imag} */,
  {32'h4443b494, 32'h00000000} /* (7, 13, 8) {real, imag} */,
  {32'hc3d87892, 32'h00000000} /* (7, 13, 7) {real, imag} */,
  {32'h44f4882f, 32'h00000000} /* (7, 13, 6) {real, imag} */,
  {32'h438cf1d2, 32'h00000000} /* (7, 13, 5) {real, imag} */,
  {32'h431cee8a, 32'h00000000} /* (7, 13, 4) {real, imag} */,
  {32'h42d828f3, 32'h00000000} /* (7, 13, 3) {real, imag} */,
  {32'h4280823c, 32'h00000000} /* (7, 13, 2) {real, imag} */,
  {32'h43e5c8d2, 32'h00000000} /* (7, 13, 1) {real, imag} */,
  {32'hc2b997cc, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'h41ac23f0, 32'h00000000} /* (7, 12, 15) {real, imag} */,
  {32'hc1efd124, 32'h00000000} /* (7, 12, 14) {real, imag} */,
  {32'h432e0efe, 32'h00000000} /* (7, 12, 13) {real, imag} */,
  {32'hc3cb4fa1, 32'h00000000} /* (7, 12, 12) {real, imag} */,
  {32'hc44b96c0, 32'h00000000} /* (7, 12, 11) {real, imag} */,
  {32'hc41f3418, 32'h00000000} /* (7, 12, 10) {real, imag} */,
  {32'h4467c7d6, 32'h00000000} /* (7, 12, 9) {real, imag} */,
  {32'hc31a7510, 32'h00000000} /* (7, 12, 8) {real, imag} */,
  {32'h42c62088, 32'h00000000} /* (7, 12, 7) {real, imag} */,
  {32'hc2ce8f6f, 32'h00000000} /* (7, 12, 6) {real, imag} */,
  {32'h42841684, 32'h00000000} /* (7, 12, 5) {real, imag} */,
  {32'h4302d636, 32'h00000000} /* (7, 12, 4) {real, imag} */,
  {32'h43813c3c, 32'h00000000} /* (7, 12, 3) {real, imag} */,
  {32'h43fba891, 32'h00000000} /* (7, 12, 2) {real, imag} */,
  {32'hc35716fa, 32'h00000000} /* (7, 12, 1) {real, imag} */,
  {32'h43cd8628, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'h427eca28, 32'h00000000} /* (7, 11, 15) {real, imag} */,
  {32'h43bbd890, 32'h00000000} /* (7, 11, 14) {real, imag} */,
  {32'hc2b94294, 32'h00000000} /* (7, 11, 13) {real, imag} */,
  {32'hc42a0375, 32'h00000000} /* (7, 11, 12) {real, imag} */,
  {32'hc41cf7e9, 32'h00000000} /* (7, 11, 11) {real, imag} */,
  {32'hc320e1b8, 32'h00000000} /* (7, 11, 10) {real, imag} */,
  {32'hc2de849e, 32'h00000000} /* (7, 11, 9) {real, imag} */,
  {32'h431a1bcd, 32'h00000000} /* (7, 11, 8) {real, imag} */,
  {32'h43ef0217, 32'h00000000} /* (7, 11, 7) {real, imag} */,
  {32'hc2e1bd22, 32'h00000000} /* (7, 11, 6) {real, imag} */,
  {32'h442ea070, 32'h00000000} /* (7, 11, 5) {real, imag} */,
  {32'h4466978f, 32'h00000000} /* (7, 11, 4) {real, imag} */,
  {32'h445834e3, 32'h00000000} /* (7, 11, 3) {real, imag} */,
  {32'h4392186d, 32'h00000000} /* (7, 11, 2) {real, imag} */,
  {32'hc2ecb09a, 32'h00000000} /* (7, 11, 1) {real, imag} */,
  {32'h4343d9bd, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'hc26755f0, 32'h00000000} /* (7, 10, 15) {real, imag} */,
  {32'hc2e4d116, 32'h00000000} /* (7, 10, 14) {real, imag} */,
  {32'h44230416, 32'h00000000} /* (7, 10, 13) {real, imag} */,
  {32'hc3a63b92, 32'h00000000} /* (7, 10, 12) {real, imag} */,
  {32'hc3d632b4, 32'h00000000} /* (7, 10, 11) {real, imag} */,
  {32'h4459eab0, 32'h00000000} /* (7, 10, 10) {real, imag} */,
  {32'h44349961, 32'h00000000} /* (7, 10, 9) {real, imag} */,
  {32'h43ba1fd9, 32'h00000000} /* (7, 10, 8) {real, imag} */,
  {32'h44497ec9, 32'h00000000} /* (7, 10, 7) {real, imag} */,
  {32'h4376c22b, 32'h00000000} /* (7, 10, 6) {real, imag} */,
  {32'h44982923, 32'h00000000} /* (7, 10, 5) {real, imag} */,
  {32'h44d5fc18, 32'h00000000} /* (7, 10, 4) {real, imag} */,
  {32'h449851a8, 32'h00000000} /* (7, 10, 3) {real, imag} */,
  {32'h449132d8, 32'h00000000} /* (7, 10, 2) {real, imag} */,
  {32'hc225eea0, 32'h00000000} /* (7, 10, 1) {real, imag} */,
  {32'h3ff91a00, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'h41f1f2e0, 32'h00000000} /* (7, 9, 15) {real, imag} */,
  {32'hc322dce1, 32'h00000000} /* (7, 9, 14) {real, imag} */,
  {32'hc393bb98, 32'h00000000} /* (7, 9, 13) {real, imag} */,
  {32'h420a67cc, 32'h00000000} /* (7, 9, 12) {real, imag} */,
  {32'h4404df32, 32'h00000000} /* (7, 9, 11) {real, imag} */,
  {32'hc3873bd2, 32'h00000000} /* (7, 9, 10) {real, imag} */,
  {32'h437174f4, 32'h00000000} /* (7, 9, 9) {real, imag} */,
  {32'h433ff0de, 32'h00000000} /* (7, 9, 8) {real, imag} */,
  {32'hc41d073a, 32'h00000000} /* (7, 9, 7) {real, imag} */,
  {32'h43cfa3a0, 32'h00000000} /* (7, 9, 6) {real, imag} */,
  {32'h44ade4aa, 32'h00000000} /* (7, 9, 5) {real, imag} */,
  {32'h43e02b1e, 32'h00000000} /* (7, 9, 4) {real, imag} */,
  {32'h43cafb73, 32'h00000000} /* (7, 9, 3) {real, imag} */,
  {32'h43c865a0, 32'h00000000} /* (7, 9, 2) {real, imag} */,
  {32'h447dead3, 32'h00000000} /* (7, 9, 1) {real, imag} */,
  {32'h430d3e72, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'hc2ed0368, 32'h00000000} /* (7, 8, 15) {real, imag} */,
  {32'hc2e10fbc, 32'h00000000} /* (7, 8, 14) {real, imag} */,
  {32'hc269d020, 32'h00000000} /* (7, 8, 13) {real, imag} */,
  {32'h42b5cd99, 32'h00000000} /* (7, 8, 12) {real, imag} */,
  {32'hc321d9fa, 32'h00000000} /* (7, 8, 11) {real, imag} */,
  {32'hc12361f7, 32'h00000000} /* (7, 8, 10) {real, imag} */,
  {32'h43d315be, 32'h00000000} /* (7, 8, 9) {real, imag} */,
  {32'h43b04ab3, 32'h00000000} /* (7, 8, 8) {real, imag} */,
  {32'h44003ab1, 32'h00000000} /* (7, 8, 7) {real, imag} */,
  {32'h44187f52, 32'h00000000} /* (7, 8, 6) {real, imag} */,
  {32'h441fccf5, 32'h00000000} /* (7, 8, 5) {real, imag} */,
  {32'h4348795a, 32'h00000000} /* (7, 8, 4) {real, imag} */,
  {32'h4454033c, 32'h00000000} /* (7, 8, 3) {real, imag} */,
  {32'h3ea14ce0, 32'h00000000} /* (7, 8, 2) {real, imag} */,
  {32'h440851a4, 32'h00000000} /* (7, 8, 1) {real, imag} */,
  {32'h4356588a, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'h425d3ede, 32'h00000000} /* (7, 7, 15) {real, imag} */,
  {32'hc464e0a8, 32'h00000000} /* (7, 7, 14) {real, imag} */,
  {32'hc30491fd, 32'h00000000} /* (7, 7, 13) {real, imag} */,
  {32'hc3699d51, 32'h00000000} /* (7, 7, 12) {real, imag} */,
  {32'h4334ba7c, 32'h00000000} /* (7, 7, 11) {real, imag} */,
  {32'h4400d9ba, 32'h00000000} /* (7, 7, 10) {real, imag} */,
  {32'hc2d2dbe0, 32'h00000000} /* (7, 7, 9) {real, imag} */,
  {32'hc3de7eb4, 32'h00000000} /* (7, 7, 8) {real, imag} */,
  {32'h4332799c, 32'h00000000} /* (7, 7, 7) {real, imag} */,
  {32'h43cc546c, 32'h00000000} /* (7, 7, 6) {real, imag} */,
  {32'h42df2ada, 32'h00000000} /* (7, 7, 5) {real, imag} */,
  {32'hc3c1ac18, 32'h00000000} /* (7, 7, 4) {real, imag} */,
  {32'hc24b446e, 32'h00000000} /* (7, 7, 3) {real, imag} */,
  {32'h438d59f8, 32'h00000000} /* (7, 7, 2) {real, imag} */,
  {32'hc4a8dedc, 32'h00000000} /* (7, 7, 1) {real, imag} */,
  {32'hc41a63d0, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'hc45c91d2, 32'h00000000} /* (7, 6, 15) {real, imag} */,
  {32'hc447d7d2, 32'h00000000} /* (7, 6, 14) {real, imag} */,
  {32'hc42cb083, 32'h00000000} /* (7, 6, 13) {real, imag} */,
  {32'hc44e57c5, 32'h00000000} /* (7, 6, 12) {real, imag} */,
  {32'hc297cc40, 32'h00000000} /* (7, 6, 11) {real, imag} */,
  {32'hc3899a47, 32'h00000000} /* (7, 6, 10) {real, imag} */,
  {32'h43eff5f0, 32'h00000000} /* (7, 6, 9) {real, imag} */,
  {32'h443f3f67, 32'h00000000} /* (7, 6, 8) {real, imag} */,
  {32'hc3f0efd4, 32'h00000000} /* (7, 6, 7) {real, imag} */,
  {32'h43ceba5c, 32'h00000000} /* (7, 6, 6) {real, imag} */,
  {32'h4286dea8, 32'h00000000} /* (7, 6, 5) {real, imag} */,
  {32'h438dfcee, 32'h00000000} /* (7, 6, 4) {real, imag} */,
  {32'hc4309aa4, 32'h00000000} /* (7, 6, 3) {real, imag} */,
  {32'hc4833a08, 32'h00000000} /* (7, 6, 2) {real, imag} */,
  {32'h430645c0, 32'h00000000} /* (7, 6, 1) {real, imag} */,
  {32'h420b8710, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'hc3b27d86, 32'h00000000} /* (7, 5, 15) {real, imag} */,
  {32'hc406caa1, 32'h00000000} /* (7, 5, 14) {real, imag} */,
  {32'hc3c76ba5, 32'h00000000} /* (7, 5, 13) {real, imag} */,
  {32'hc428f1d1, 32'h00000000} /* (7, 5, 12) {real, imag} */,
  {32'hc373e92e, 32'h00000000} /* (7, 5, 11) {real, imag} */,
  {32'hc4202576, 32'h00000000} /* (7, 5, 10) {real, imag} */,
  {32'h440ca592, 32'h00000000} /* (7, 5, 9) {real, imag} */,
  {32'h42734fb8, 32'h00000000} /* (7, 5, 8) {real, imag} */,
  {32'h44109e58, 32'h00000000} /* (7, 5, 7) {real, imag} */,
  {32'h443595e1, 32'h00000000} /* (7, 5, 6) {real, imag} */,
  {32'h445cd01e, 32'h00000000} /* (7, 5, 5) {real, imag} */,
  {32'h448093b6, 32'h00000000} /* (7, 5, 4) {real, imag} */,
  {32'hc422d1f0, 32'h00000000} /* (7, 5, 3) {real, imag} */,
  {32'hc4486f96, 32'h00000000} /* (7, 5, 2) {real, imag} */,
  {32'hc39f060f, 32'h00000000} /* (7, 5, 1) {real, imag} */,
  {32'hc3ebb5fd, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'hc441b37a, 32'h00000000} /* (7, 4, 15) {real, imag} */,
  {32'hc2f20010, 32'h00000000} /* (7, 4, 14) {real, imag} */,
  {32'h430f3618, 32'h00000000} /* (7, 4, 13) {real, imag} */,
  {32'h43183194, 32'h00000000} /* (7, 4, 12) {real, imag} */,
  {32'h43fafe2d, 32'h00000000} /* (7, 4, 11) {real, imag} */,
  {32'hc46908b0, 32'h00000000} /* (7, 4, 10) {real, imag} */,
  {32'h44a605be, 32'h00000000} /* (7, 4, 9) {real, imag} */,
  {32'h40863500, 32'h00000000} /* (7, 4, 8) {real, imag} */,
  {32'hc34d5e3c, 32'h00000000} /* (7, 4, 7) {real, imag} */,
  {32'h44ab6c26, 32'h00000000} /* (7, 4, 6) {real, imag} */,
  {32'h448fa0cf, 32'h00000000} /* (7, 4, 5) {real, imag} */,
  {32'h447c34d1, 32'h00000000} /* (7, 4, 4) {real, imag} */,
  {32'hc336d0d6, 32'h00000000} /* (7, 4, 3) {real, imag} */,
  {32'hc4b9eef0, 32'h00000000} /* (7, 4, 2) {real, imag} */,
  {32'hc42689e3, 32'h00000000} /* (7, 4, 1) {real, imag} */,
  {32'hc38eac30, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'hc45ce1f2, 32'h00000000} /* (7, 3, 15) {real, imag} */,
  {32'h4450177c, 32'h00000000} /* (7, 3, 14) {real, imag} */,
  {32'h44825748, 32'h00000000} /* (7, 3, 13) {real, imag} */,
  {32'hc3d21871, 32'h00000000} /* (7, 3, 12) {real, imag} */,
  {32'h4405fb58, 32'h00000000} /* (7, 3, 11) {real, imag} */,
  {32'hc19088c0, 32'h00000000} /* (7, 3, 10) {real, imag} */,
  {32'hc3fc8f28, 32'h00000000} /* (7, 3, 9) {real, imag} */,
  {32'h430e8a8a, 32'h00000000} /* (7, 3, 8) {real, imag} */,
  {32'h43d7f880, 32'h00000000} /* (7, 3, 7) {real, imag} */,
  {32'h44354854, 32'h00000000} /* (7, 3, 6) {real, imag} */,
  {32'h44ac283a, 32'h00000000} /* (7, 3, 5) {real, imag} */,
  {32'hc0ccfdc0, 32'h00000000} /* (7, 3, 4) {real, imag} */,
  {32'hc3c2a708, 32'h00000000} /* (7, 3, 3) {real, imag} */,
  {32'hc43a6e33, 32'h00000000} /* (7, 3, 2) {real, imag} */,
  {32'hc490e4e0, 32'h00000000} /* (7, 3, 1) {real, imag} */,
  {32'hc3fe6f99, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'hc27bd48d, 32'h00000000} /* (7, 2, 15) {real, imag} */,
  {32'hc3f602c3, 32'h00000000} /* (7, 2, 14) {real, imag} */,
  {32'h43286324, 32'h00000000} /* (7, 2, 13) {real, imag} */,
  {32'h441cea0e, 32'h00000000} /* (7, 2, 12) {real, imag} */,
  {32'hc431207a, 32'h00000000} /* (7, 2, 11) {real, imag} */,
  {32'hc4361ed2, 32'h00000000} /* (7, 2, 10) {real, imag} */,
  {32'hc40c75b3, 32'h00000000} /* (7, 2, 9) {real, imag} */,
  {32'hc3f8eafc, 32'h00000000} /* (7, 2, 8) {real, imag} */,
  {32'hc1d72f46, 32'h00000000} /* (7, 2, 7) {real, imag} */,
  {32'h442727a4, 32'h00000000} /* (7, 2, 6) {real, imag} */,
  {32'h447b6427, 32'h00000000} /* (7, 2, 5) {real, imag} */,
  {32'h42f7a43c, 32'h00000000} /* (7, 2, 4) {real, imag} */,
  {32'hc3d47425, 32'h00000000} /* (7, 2, 3) {real, imag} */,
  {32'hc46777ae, 32'h00000000} /* (7, 2, 2) {real, imag} */,
  {32'hc4cb6186, 32'h00000000} /* (7, 2, 1) {real, imag} */,
  {32'hc4806ccd, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'h428ec78c, 32'h00000000} /* (7, 1, 15) {real, imag} */,
  {32'hc3dced89, 32'h00000000} /* (7, 1, 14) {real, imag} */,
  {32'hc42e1502, 32'h00000000} /* (7, 1, 13) {real, imag} */,
  {32'h43646462, 32'h00000000} /* (7, 1, 12) {real, imag} */,
  {32'hc44fedea, 32'h00000000} /* (7, 1, 11) {real, imag} */,
  {32'hc3866f81, 32'h00000000} /* (7, 1, 10) {real, imag} */,
  {32'hc3ecff40, 32'h00000000} /* (7, 1, 9) {real, imag} */,
  {32'hc465a732, 32'h00000000} /* (7, 1, 8) {real, imag} */,
  {32'h4447297a, 32'h00000000} /* (7, 1, 7) {real, imag} */,
  {32'h4437d19e, 32'h00000000} /* (7, 1, 6) {real, imag} */,
  {32'h43d1042f, 32'h00000000} /* (7, 1, 5) {real, imag} */,
  {32'h446a8ae0, 32'h00000000} /* (7, 1, 4) {real, imag} */,
  {32'h43964994, 32'h00000000} /* (7, 1, 3) {real, imag} */,
  {32'hc46114f8, 32'h00000000} /* (7, 1, 2) {real, imag} */,
  {32'hc4b2e980, 32'h00000000} /* (7, 1, 1) {real, imag} */,
  {32'hc3d371d4, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'hc41bbf35, 32'h00000000} /* (7, 0, 15) {real, imag} */,
  {32'hc3f92636, 32'h00000000} /* (7, 0, 14) {real, imag} */,
  {32'hc3f67c23, 32'h00000000} /* (7, 0, 13) {real, imag} */,
  {32'hc32e27ce, 32'h00000000} /* (7, 0, 12) {real, imag} */,
  {32'h41a56f30, 32'h00000000} /* (7, 0, 11) {real, imag} */,
  {32'hc3578989, 32'h00000000} /* (7, 0, 10) {real, imag} */,
  {32'h43e35b44, 32'h00000000} /* (7, 0, 9) {real, imag} */,
  {32'h43942cbc, 32'h00000000} /* (7, 0, 8) {real, imag} */,
  {32'hc2e7206e, 32'h00000000} /* (7, 0, 7) {real, imag} */,
  {32'h43f7e240, 32'h00000000} /* (7, 0, 6) {real, imag} */,
  {32'h4409da52, 32'h00000000} /* (7, 0, 5) {real, imag} */,
  {32'h43b1a413, 32'h00000000} /* (7, 0, 4) {real, imag} */,
  {32'hc2b36074, 32'h00000000} /* (7, 0, 3) {real, imag} */,
  {32'hc365d627, 32'h00000000} /* (7, 0, 2) {real, imag} */,
  {32'hc3683989, 32'h00000000} /* (7, 0, 1) {real, imag} */,
  {32'h4351d301, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'hc3b3ef2a, 32'h00000000} /* (6, 15, 15) {real, imag} */,
  {32'hc3305a2a, 32'h00000000} /* (6, 15, 14) {real, imag} */,
  {32'hc43e5aea, 32'h00000000} /* (6, 15, 13) {real, imag} */,
  {32'hc41fc380, 32'h00000000} /* (6, 15, 12) {real, imag} */,
  {32'hc3c8e31c, 32'h00000000} /* (6, 15, 11) {real, imag} */,
  {32'hc3bb048e, 32'h00000000} /* (6, 15, 10) {real, imag} */,
  {32'hc34f8b3c, 32'h00000000} /* (6, 15, 9) {real, imag} */,
  {32'h43bbdb02, 32'h00000000} /* (6, 15, 8) {real, imag} */,
  {32'h422d0394, 32'h00000000} /* (6, 15, 7) {real, imag} */,
  {32'h42db2434, 32'h00000000} /* (6, 15, 6) {real, imag} */,
  {32'hc388e2e0, 32'h00000000} /* (6, 15, 5) {real, imag} */,
  {32'hc454a0f0, 32'h00000000} /* (6, 15, 4) {real, imag} */,
  {32'hc30fe8ef, 32'h00000000} /* (6, 15, 3) {real, imag} */,
  {32'hc40da53f, 32'h00000000} /* (6, 15, 2) {real, imag} */,
  {32'hc3bd5bea, 32'h00000000} /* (6, 15, 1) {real, imag} */,
  {32'hc2bf0518, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'hc324d256, 32'h00000000} /* (6, 14, 15) {real, imag} */,
  {32'hc468436c, 32'h00000000} /* (6, 14, 14) {real, imag} */,
  {32'hc4491caa, 32'h00000000} /* (6, 14, 13) {real, imag} */,
  {32'hc3cf0732, 32'h00000000} /* (6, 14, 12) {real, imag} */,
  {32'hc3af62f1, 32'h00000000} /* (6, 14, 11) {real, imag} */,
  {32'hc40a445b, 32'h00000000} /* (6, 14, 10) {real, imag} */,
  {32'hc2dd0021, 32'h00000000} /* (6, 14, 9) {real, imag} */,
  {32'h4379254c, 32'h00000000} /* (6, 14, 8) {real, imag} */,
  {32'hc32be030, 32'h00000000} /* (6, 14, 7) {real, imag} */,
  {32'h43a0f764, 32'h00000000} /* (6, 14, 6) {real, imag} */,
  {32'hc3abd62c, 32'h00000000} /* (6, 14, 5) {real, imag} */,
  {32'hc356ba0c, 32'h00000000} /* (6, 14, 4) {real, imag} */,
  {32'hc38bd32b, 32'h00000000} /* (6, 14, 3) {real, imag} */,
  {32'hc41451d7, 32'h00000000} /* (6, 14, 2) {real, imag} */,
  {32'hc30250b2, 32'h00000000} /* (6, 14, 1) {real, imag} */,
  {32'h4230d148, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hc3e7160c, 32'h00000000} /* (6, 13, 15) {real, imag} */,
  {32'hc3ca408d, 32'h00000000} /* (6, 13, 14) {real, imag} */,
  {32'hc4389a48, 32'h00000000} /* (6, 13, 13) {real, imag} */,
  {32'hc465ea39, 32'h00000000} /* (6, 13, 12) {real, imag} */,
  {32'hc4218617, 32'h00000000} /* (6, 13, 11) {real, imag} */,
  {32'h43fbd5d1, 32'h00000000} /* (6, 13, 10) {real, imag} */,
  {32'hc356bca8, 32'h00000000} /* (6, 13, 9) {real, imag} */,
  {32'hc43be73e, 32'h00000000} /* (6, 13, 8) {real, imag} */,
  {32'h43d74988, 32'h00000000} /* (6, 13, 7) {real, imag} */,
  {32'h42a8470c, 32'h00000000} /* (6, 13, 6) {real, imag} */,
  {32'hc2f0d154, 32'h00000000} /* (6, 13, 5) {real, imag} */,
  {32'hc4147c91, 32'h00000000} /* (6, 13, 4) {real, imag} */,
  {32'hc40ac777, 32'h00000000} /* (6, 13, 3) {real, imag} */,
  {32'hc1505ee0, 32'h00000000} /* (6, 13, 2) {real, imag} */,
  {32'hc303ea80, 32'h00000000} /* (6, 13, 1) {real, imag} */,
  {32'hc40155f4, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'hc2e4e8fd, 32'h00000000} /* (6, 12, 15) {real, imag} */,
  {32'hc43377ee, 32'h00000000} /* (6, 12, 14) {real, imag} */,
  {32'hc2efdbc0, 32'h00000000} /* (6, 12, 13) {real, imag} */,
  {32'hc473e0ad, 32'h00000000} /* (6, 12, 12) {real, imag} */,
  {32'h427e2bd8, 32'h00000000} /* (6, 12, 11) {real, imag} */,
  {32'hc3c446f2, 32'h00000000} /* (6, 12, 10) {real, imag} */,
  {32'hc4066192, 32'h00000000} /* (6, 12, 9) {real, imag} */,
  {32'h441477aa, 32'h00000000} /* (6, 12, 8) {real, imag} */,
  {32'hc3870740, 32'h00000000} /* (6, 12, 7) {real, imag} */,
  {32'h440c385a, 32'h00000000} /* (6, 12, 6) {real, imag} */,
  {32'hc1c382c2, 32'h00000000} /* (6, 12, 5) {real, imag} */,
  {32'h43e09c4e, 32'h00000000} /* (6, 12, 4) {real, imag} */,
  {32'h440e8d9c, 32'h00000000} /* (6, 12, 3) {real, imag} */,
  {32'hc2fb1846, 32'h00000000} /* (6, 12, 2) {real, imag} */,
  {32'hc3ba6d18, 32'h00000000} /* (6, 12, 1) {real, imag} */,
  {32'hc2d4e492, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'h446493fa, 32'h00000000} /* (6, 11, 15) {real, imag} */,
  {32'h4484d001, 32'h00000000} /* (6, 11, 14) {real, imag} */,
  {32'hc42c8a4b, 32'h00000000} /* (6, 11, 13) {real, imag} */,
  {32'hc338ba5a, 32'h00000000} /* (6, 11, 12) {real, imag} */,
  {32'hc4852294, 32'h00000000} /* (6, 11, 11) {real, imag} */,
  {32'hc470a482, 32'h00000000} /* (6, 11, 10) {real, imag} */,
  {32'hc41aa6f1, 32'h00000000} /* (6, 11, 9) {real, imag} */,
  {32'h427bb29c, 32'h00000000} /* (6, 11, 8) {real, imag} */,
  {32'hc3b3bc45, 32'h00000000} /* (6, 11, 7) {real, imag} */,
  {32'h43af6d3c, 32'h00000000} /* (6, 11, 6) {real, imag} */,
  {32'h443a0de5, 32'h00000000} /* (6, 11, 5) {real, imag} */,
  {32'h4434b6d8, 32'h00000000} /* (6, 11, 4) {real, imag} */,
  {32'h44911e00, 32'h00000000} /* (6, 11, 3) {real, imag} */,
  {32'h41d28130, 32'h00000000} /* (6, 11, 2) {real, imag} */,
  {32'h442ad0f9, 32'h00000000} /* (6, 11, 1) {real, imag} */,
  {32'hc272f684, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h44034227, 32'h00000000} /* (6, 10, 15) {real, imag} */,
  {32'h4215f43c, 32'h00000000} /* (6, 10, 14) {real, imag} */,
  {32'hc48ce70f, 32'h00000000} /* (6, 10, 13) {real, imag} */,
  {32'hc3de385c, 32'h00000000} /* (6, 10, 12) {real, imag} */,
  {32'hc3eedc9c, 32'h00000000} /* (6, 10, 11) {real, imag} */,
  {32'hc400d930, 32'h00000000} /* (6, 10, 10) {real, imag} */,
  {32'h4322b700, 32'h00000000} /* (6, 10, 9) {real, imag} */,
  {32'hc242fc84, 32'h00000000} /* (6, 10, 8) {real, imag} */,
  {32'hbfcfde00, 32'h00000000} /* (6, 10, 7) {real, imag} */,
  {32'h43a04ffa, 32'h00000000} /* (6, 10, 6) {real, imag} */,
  {32'h441a0f92, 32'h00000000} /* (6, 10, 5) {real, imag} */,
  {32'h44c88f2d, 32'h00000000} /* (6, 10, 4) {real, imag} */,
  {32'h4509f474, 32'h00000000} /* (6, 10, 3) {real, imag} */,
  {32'h440eb46c, 32'h00000000} /* (6, 10, 2) {real, imag} */,
  {32'h444eab56, 32'h00000000} /* (6, 10, 1) {real, imag} */,
  {32'h43c16b90, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'h4482701a, 32'h00000000} /* (6, 9, 15) {real, imag} */,
  {32'hc40d2d13, 32'h00000000} /* (6, 9, 14) {real, imag} */,
  {32'hc4a2b611, 32'h00000000} /* (6, 9, 13) {real, imag} */,
  {32'hc37828e4, 32'h00000000} /* (6, 9, 12) {real, imag} */,
  {32'h4415731d, 32'h00000000} /* (6, 9, 11) {real, imag} */,
  {32'hc23eeff8, 32'h00000000} /* (6, 9, 10) {real, imag} */,
  {32'h445acb20, 32'h00000000} /* (6, 9, 9) {real, imag} */,
  {32'h449be41c, 32'h00000000} /* (6, 9, 8) {real, imag} */,
  {32'h44424177, 32'h00000000} /* (6, 9, 7) {real, imag} */,
  {32'h442e8a33, 32'h00000000} /* (6, 9, 6) {real, imag} */,
  {32'h4441c142, 32'h00000000} /* (6, 9, 5) {real, imag} */,
  {32'h44916bec, 32'h00000000} /* (6, 9, 4) {real, imag} */,
  {32'h43cd9609, 32'h00000000} /* (6, 9, 3) {real, imag} */,
  {32'h444df32a, 32'h00000000} /* (6, 9, 2) {real, imag} */,
  {32'h443a155c, 32'h00000000} /* (6, 9, 1) {real, imag} */,
  {32'hc3844f34, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'h444c49fe, 32'h00000000} /* (6, 8, 15) {real, imag} */,
  {32'hc3882306, 32'h00000000} /* (6, 8, 14) {real, imag} */,
  {32'hc49e6857, 32'h00000000} /* (6, 8, 13) {real, imag} */,
  {32'hc3cb5472, 32'h00000000} /* (6, 8, 12) {real, imag} */,
  {32'hc3eea7e0, 32'h00000000} /* (6, 8, 11) {real, imag} */,
  {32'hc2cd638d, 32'h00000000} /* (6, 8, 10) {real, imag} */,
  {32'h43a25943, 32'h00000000} /* (6, 8, 9) {real, imag} */,
  {32'h4284bc31, 32'h00000000} /* (6, 8, 8) {real, imag} */,
  {32'h44361c8a, 32'h00000000} /* (6, 8, 7) {real, imag} */,
  {32'h44061637, 32'h00000000} /* (6, 8, 6) {real, imag} */,
  {32'h4442a7c2, 32'h00000000} /* (6, 8, 5) {real, imag} */,
  {32'hc2ecf3e0, 32'h00000000} /* (6, 8, 4) {real, imag} */,
  {32'h43a25082, 32'h00000000} /* (6, 8, 3) {real, imag} */,
  {32'h42835a23, 32'h00000000} /* (6, 8, 2) {real, imag} */,
  {32'hc4014b0d, 32'h00000000} /* (6, 8, 1) {real, imag} */,
  {32'hc3208e9c, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'hc39df17f, 32'h00000000} /* (6, 7, 15) {real, imag} */,
  {32'hc44b3385, 32'h00000000} /* (6, 7, 14) {real, imag} */,
  {32'hc497216f, 32'h00000000} /* (6, 7, 13) {real, imag} */,
  {32'hc4cc66cb, 32'h00000000} /* (6, 7, 12) {real, imag} */,
  {32'hc469bf7c, 32'h00000000} /* (6, 7, 11) {real, imag} */,
  {32'hc3be07dd, 32'h00000000} /* (6, 7, 10) {real, imag} */,
  {32'hc3b37751, 32'h00000000} /* (6, 7, 9) {real, imag} */,
  {32'hc4395732, 32'h00000000} /* (6, 7, 8) {real, imag} */,
  {32'h42d9e420, 32'h00000000} /* (6, 7, 7) {real, imag} */,
  {32'h43ce5a36, 32'h00000000} /* (6, 7, 6) {real, imag} */,
  {32'hc40c6372, 32'h00000000} /* (6, 7, 5) {real, imag} */,
  {32'hc39ec7cc, 32'h00000000} /* (6, 7, 4) {real, imag} */,
  {32'h44338f92, 32'h00000000} /* (6, 7, 3) {real, imag} */,
  {32'h42d8cb94, 32'h00000000} /* (6, 7, 2) {real, imag} */,
  {32'h43e6ad75, 32'h00000000} /* (6, 7, 1) {real, imag} */,
  {32'h43d5e22c, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'hc37e4a3c, 32'h00000000} /* (6, 6, 15) {real, imag} */,
  {32'hc41a7547, 32'h00000000} /* (6, 6, 14) {real, imag} */,
  {32'hc468ea20, 32'h00000000} /* (6, 6, 13) {real, imag} */,
  {32'hc4b91e65, 32'h00000000} /* (6, 6, 12) {real, imag} */,
  {32'h42870424, 32'h00000000} /* (6, 6, 11) {real, imag} */,
  {32'h4359f2f1, 32'h00000000} /* (6, 6, 10) {real, imag} */,
  {32'hc417ea4e, 32'h00000000} /* (6, 6, 9) {real, imag} */,
  {32'hc37113a6, 32'h00000000} /* (6, 6, 8) {real, imag} */,
  {32'h4270f968, 32'h00000000} /* (6, 6, 7) {real, imag} */,
  {32'h4414d001, 32'h00000000} /* (6, 6, 6) {real, imag} */,
  {32'hc358882e, 32'h00000000} /* (6, 6, 5) {real, imag} */,
  {32'hc3da6e20, 32'h00000000} /* (6, 6, 4) {real, imag} */,
  {32'hc3bf3f4e, 32'h00000000} /* (6, 6, 3) {real, imag} */,
  {32'h42db6a76, 32'h00000000} /* (6, 6, 2) {real, imag} */,
  {32'hc325aada, 32'h00000000} /* (6, 6, 1) {real, imag} */,
  {32'hc2d58da4, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'hc45243cb, 32'h00000000} /* (6, 5, 15) {real, imag} */,
  {32'hc45968a1, 32'h00000000} /* (6, 5, 14) {real, imag} */,
  {32'hc38c5042, 32'h00000000} /* (6, 5, 13) {real, imag} */,
  {32'hc48bf76d, 32'h00000000} /* (6, 5, 12) {real, imag} */,
  {32'hc40bf3b4, 32'h00000000} /* (6, 5, 11) {real, imag} */,
  {32'hc41df48f, 32'h00000000} /* (6, 5, 10) {real, imag} */,
  {32'h41d9a520, 32'h00000000} /* (6, 5, 9) {real, imag} */,
  {32'h42d237e6, 32'h00000000} /* (6, 5, 8) {real, imag} */,
  {32'h44115657, 32'h00000000} /* (6, 5, 7) {real, imag} */,
  {32'h442ecc45, 32'h00000000} /* (6, 5, 6) {real, imag} */,
  {32'h43102aa4, 32'h00000000} /* (6, 5, 5) {real, imag} */,
  {32'hc324fc88, 32'h00000000} /* (6, 5, 4) {real, imag} */,
  {32'hc48b14d6, 32'h00000000} /* (6, 5, 3) {real, imag} */,
  {32'hc48cd363, 32'h00000000} /* (6, 5, 2) {real, imag} */,
  {32'hc49c4606, 32'h00000000} /* (6, 5, 1) {real, imag} */,
  {32'hc3bc9342, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'hc4036a79, 32'h00000000} /* (6, 4, 15) {real, imag} */,
  {32'h437466f1, 32'h00000000} /* (6, 4, 14) {real, imag} */,
  {32'hc32837ae, 32'h00000000} /* (6, 4, 13) {real, imag} */,
  {32'h43319910, 32'h00000000} /* (6, 4, 12) {real, imag} */,
  {32'hc42c60c8, 32'h00000000} /* (6, 4, 11) {real, imag} */,
  {32'hc3224ee8, 32'h00000000} /* (6, 4, 10) {real, imag} */,
  {32'h43d2d9a1, 32'h00000000} /* (6, 4, 9) {real, imag} */,
  {32'hc20c1650, 32'h00000000} /* (6, 4, 8) {real, imag} */,
  {32'hc346600c, 32'h00000000} /* (6, 4, 7) {real, imag} */,
  {32'h43e0a7b0, 32'h00000000} /* (6, 4, 6) {real, imag} */,
  {32'h43ef36d3, 32'h00000000} /* (6, 4, 5) {real, imag} */,
  {32'h433d97b6, 32'h00000000} /* (6, 4, 4) {real, imag} */,
  {32'hc4da2b0c, 32'h00000000} /* (6, 4, 3) {real, imag} */,
  {32'hc4905db3, 32'h00000000} /* (6, 4, 2) {real, imag} */,
  {32'hc40cb863, 32'h00000000} /* (6, 4, 1) {real, imag} */,
  {32'hc4263855, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'hc436f175, 32'h00000000} /* (6, 3, 15) {real, imag} */,
  {32'h422fb770, 32'h00000000} /* (6, 3, 14) {real, imag} */,
  {32'h4458e84b, 32'h00000000} /* (6, 3, 13) {real, imag} */,
  {32'hc42225ca, 32'h00000000} /* (6, 3, 12) {real, imag} */,
  {32'h443be95c, 32'h00000000} /* (6, 3, 11) {real, imag} */,
  {32'hc341caab, 32'h00000000} /* (6, 3, 10) {real, imag} */,
  {32'hc3e7e6a2, 32'h00000000} /* (6, 3, 9) {real, imag} */,
  {32'hc1f5e950, 32'h00000000} /* (6, 3, 8) {real, imag} */,
  {32'hc42ae76f, 32'h00000000} /* (6, 3, 7) {real, imag} */,
  {32'hc3847654, 32'h00000000} /* (6, 3, 6) {real, imag} */,
  {32'h44175b51, 32'h00000000} /* (6, 3, 5) {real, imag} */,
  {32'hc43ce9ce, 32'h00000000} /* (6, 3, 4) {real, imag} */,
  {32'hc4aa459a, 32'h00000000} /* (6, 3, 3) {real, imag} */,
  {32'hc33cb631, 32'h00000000} /* (6, 3, 2) {real, imag} */,
  {32'hc41f873f, 32'h00000000} /* (6, 3, 1) {real, imag} */,
  {32'hc439bac6, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'hc4881d96, 32'h00000000} /* (6, 2, 15) {real, imag} */,
  {32'hc41b4dd8, 32'h00000000} /* (6, 2, 14) {real, imag} */,
  {32'h42c88e78, 32'h00000000} /* (6, 2, 13) {real, imag} */,
  {32'hc4147772, 32'h00000000} /* (6, 2, 12) {real, imag} */,
  {32'hc3600000, 32'h00000000} /* (6, 2, 11) {real, imag} */,
  {32'hc471ed53, 32'h00000000} /* (6, 2, 10) {real, imag} */,
  {32'hc3fe397c, 32'h00000000} /* (6, 2, 9) {real, imag} */,
  {32'hc46e4e6b, 32'h00000000} /* (6, 2, 8) {real, imag} */,
  {32'h43ca18e6, 32'h00000000} /* (6, 2, 7) {real, imag} */,
  {32'h4445c62e, 32'h00000000} /* (6, 2, 6) {real, imag} */,
  {32'hc45f658a, 32'h00000000} /* (6, 2, 5) {real, imag} */,
  {32'hc311d2e5, 32'h00000000} /* (6, 2, 4) {real, imag} */,
  {32'h42cb5e64, 32'h00000000} /* (6, 2, 3) {real, imag} */,
  {32'hc43defaf, 32'h00000000} /* (6, 2, 2) {real, imag} */,
  {32'hc4a0f82b, 32'h00000000} /* (6, 2, 1) {real, imag} */,
  {32'hc4590b3d, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'hc46907a5, 32'h00000000} /* (6, 1, 15) {real, imag} */,
  {32'hc254669a, 32'h00000000} /* (6, 1, 14) {real, imag} */,
  {32'h4316882c, 32'h00000000} /* (6, 1, 13) {real, imag} */,
  {32'hc3de67e2, 32'h00000000} /* (6, 1, 12) {real, imag} */,
  {32'hc4c0e163, 32'h00000000} /* (6, 1, 11) {real, imag} */,
  {32'hc4739044, 32'h00000000} /* (6, 1, 10) {real, imag} */,
  {32'h43875a91, 32'h00000000} /* (6, 1, 9) {real, imag} */,
  {32'h42029a30, 32'h00000000} /* (6, 1, 8) {real, imag} */,
  {32'hc449fe3f, 32'h00000000} /* (6, 1, 7) {real, imag} */,
  {32'hc3472f82, 32'h00000000} /* (6, 1, 6) {real, imag} */,
  {32'h4403a55a, 32'h00000000} /* (6, 1, 5) {real, imag} */,
  {32'h44cf4e78, 32'h00000000} /* (6, 1, 4) {real, imag} */,
  {32'h43be5c64, 32'h00000000} /* (6, 1, 3) {real, imag} */,
  {32'hc4436bc2, 32'h00000000} /* (6, 1, 2) {real, imag} */,
  {32'hc499232c, 32'h00000000} /* (6, 1, 1) {real, imag} */,
  {32'hc48840de, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'hc3d51c3d, 32'h00000000} /* (6, 0, 15) {real, imag} */,
  {32'hc3a72a99, 32'h00000000} /* (6, 0, 14) {real, imag} */,
  {32'hc3481cdc, 32'h00000000} /* (6, 0, 13) {real, imag} */,
  {32'hc39dd9e1, 32'h00000000} /* (6, 0, 12) {real, imag} */,
  {32'hc40dddaf, 32'h00000000} /* (6, 0, 11) {real, imag} */,
  {32'hc3881f09, 32'h00000000} /* (6, 0, 10) {real, imag} */,
  {32'hc2584de4, 32'h00000000} /* (6, 0, 9) {real, imag} */,
  {32'hc31d7336, 32'h00000000} /* (6, 0, 8) {real, imag} */,
  {32'hc32f7c86, 32'h00000000} /* (6, 0, 7) {real, imag} */,
  {32'hc3aed517, 32'h00000000} /* (6, 0, 6) {real, imag} */,
  {32'h44820cec, 32'h00000000} /* (6, 0, 5) {real, imag} */,
  {32'h43a6c8ab, 32'h00000000} /* (6, 0, 4) {real, imag} */,
  {32'hc4084ae5, 32'h00000000} /* (6, 0, 3) {real, imag} */,
  {32'hc3dc7f4f, 32'h00000000} /* (6, 0, 2) {real, imag} */,
  {32'hc3f07924, 32'h00000000} /* (6, 0, 1) {real, imag} */,
  {32'hc3d285c9, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'hc4b3aba0, 32'h00000000} /* (5, 15, 15) {real, imag} */,
  {32'hc47131dc, 32'h00000000} /* (5, 15, 14) {real, imag} */,
  {32'hc3b5f87c, 32'h00000000} /* (5, 15, 13) {real, imag} */,
  {32'hc39a2df5, 32'h00000000} /* (5, 15, 12) {real, imag} */,
  {32'hc46dc77f, 32'h00000000} /* (5, 15, 11) {real, imag} */,
  {32'hc4029109, 32'h00000000} /* (5, 15, 10) {real, imag} */,
  {32'hc34e1b98, 32'h00000000} /* (5, 15, 9) {real, imag} */,
  {32'hc3b57bf0, 32'h00000000} /* (5, 15, 8) {real, imag} */,
  {32'hc384439e, 32'h00000000} /* (5, 15, 7) {real, imag} */,
  {32'hc314c88e, 32'h00000000} /* (5, 15, 6) {real, imag} */,
  {32'h42a04770, 32'h00000000} /* (5, 15, 5) {real, imag} */,
  {32'h444c38f6, 32'h00000000} /* (5, 15, 4) {real, imag} */,
  {32'hc3abfe92, 32'h00000000} /* (5, 15, 3) {real, imag} */,
  {32'hc45fa947, 32'h00000000} /* (5, 15, 2) {real, imag} */,
  {32'hc3dcfa98, 32'h00000000} /* (5, 15, 1) {real, imag} */,
  {32'hc260c6b0, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'hc48c1221, 32'h00000000} /* (5, 14, 15) {real, imag} */,
  {32'hc3ac660e, 32'h00000000} /* (5, 14, 14) {real, imag} */,
  {32'hc48a114e, 32'h00000000} /* (5, 14, 13) {real, imag} */,
  {32'hc46b5f32, 32'h00000000} /* (5, 14, 12) {real, imag} */,
  {32'hc3f3edf5, 32'h00000000} /* (5, 14, 11) {real, imag} */,
  {32'hc4338bcc, 32'h00000000} /* (5, 14, 10) {real, imag} */,
  {32'hc23ad268, 32'h00000000} /* (5, 14, 9) {real, imag} */,
  {32'hc4189eb5, 32'h00000000} /* (5, 14, 8) {real, imag} */,
  {32'h42de82d4, 32'h00000000} /* (5, 14, 7) {real, imag} */,
  {32'h43102265, 32'h00000000} /* (5, 14, 6) {real, imag} */,
  {32'hc2a94380, 32'h00000000} /* (5, 14, 5) {real, imag} */,
  {32'hc302c8fa, 32'h00000000} /* (5, 14, 4) {real, imag} */,
  {32'hc42dc192, 32'h00000000} /* (5, 14, 3) {real, imag} */,
  {32'hc4c13bc6, 32'h00000000} /* (5, 14, 2) {real, imag} */,
  {32'h42189a18, 32'h00000000} /* (5, 14, 1) {real, imag} */,
  {32'h4441908d, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hc39f066e, 32'h00000000} /* (5, 13, 15) {real, imag} */,
  {32'hc41b88fc, 32'h00000000} /* (5, 13, 14) {real, imag} */,
  {32'hc433816c, 32'h00000000} /* (5, 13, 13) {real, imag} */,
  {32'hc4ba83c7, 32'h00000000} /* (5, 13, 12) {real, imag} */,
  {32'hc4369bd1, 32'h00000000} /* (5, 13, 11) {real, imag} */,
  {32'hc3a0ed23, 32'h00000000} /* (5, 13, 10) {real, imag} */,
  {32'hc473a73c, 32'h00000000} /* (5, 13, 9) {real, imag} */,
  {32'hc3bf1706, 32'h00000000} /* (5, 13, 8) {real, imag} */,
  {32'h421f3ba4, 32'h00000000} /* (5, 13, 7) {real, imag} */,
  {32'h41b40360, 32'h00000000} /* (5, 13, 6) {real, imag} */,
  {32'hc40516dc, 32'h00000000} /* (5, 13, 5) {real, imag} */,
  {32'hc4954089, 32'h00000000} /* (5, 13, 4) {real, imag} */,
  {32'hc212f720, 32'h00000000} /* (5, 13, 3) {real, imag} */,
  {32'hc3a7e3ab, 32'h00000000} /* (5, 13, 2) {real, imag} */,
  {32'hc46e2864, 32'h00000000} /* (5, 13, 1) {real, imag} */,
  {32'hc410dfbc, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'hc4107e47, 32'h00000000} /* (5, 12, 15) {real, imag} */,
  {32'h43c9a8c4, 32'h00000000} /* (5, 12, 14) {real, imag} */,
  {32'h43a5b66e, 32'h00000000} /* (5, 12, 13) {real, imag} */,
  {32'hc4b5d78e, 32'h00000000} /* (5, 12, 12) {real, imag} */,
  {32'hc47ced44, 32'h00000000} /* (5, 12, 11) {real, imag} */,
  {32'hc484426c, 32'h00000000} /* (5, 12, 10) {real, imag} */,
  {32'hc4b70221, 32'h00000000} /* (5, 12, 9) {real, imag} */,
  {32'hc41f8c3c, 32'h00000000} /* (5, 12, 8) {real, imag} */,
  {32'h43d52002, 32'h00000000} /* (5, 12, 7) {real, imag} */,
  {32'hc410f42d, 32'h00000000} /* (5, 12, 6) {real, imag} */,
  {32'hc350e21c, 32'h00000000} /* (5, 12, 5) {real, imag} */,
  {32'h428aeec0, 32'h00000000} /* (5, 12, 4) {real, imag} */,
  {32'hc359adc2, 32'h00000000} /* (5, 12, 3) {real, imag} */,
  {32'h42d4d014, 32'h00000000} /* (5, 12, 2) {real, imag} */,
  {32'hc431560e, 32'h00000000} /* (5, 12, 1) {real, imag} */,
  {32'hc4075830, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h43d1606f, 32'h00000000} /* (5, 11, 15) {real, imag} */,
  {32'hc4240946, 32'h00000000} /* (5, 11, 14) {real, imag} */,
  {32'hc4e22dea, 32'h00000000} /* (5, 11, 13) {real, imag} */,
  {32'hc3b210b4, 32'h00000000} /* (5, 11, 12) {real, imag} */,
  {32'hc1d6cc80, 32'h00000000} /* (5, 11, 11) {real, imag} */,
  {32'hc4a9e958, 32'h00000000} /* (5, 11, 10) {real, imag} */,
  {32'hc48fbbfd, 32'h00000000} /* (5, 11, 9) {real, imag} */,
  {32'hc470ece6, 32'h00000000} /* (5, 11, 8) {real, imag} */,
  {32'hc30feb2a, 32'h00000000} /* (5, 11, 7) {real, imag} */,
  {32'h44353d8e, 32'h00000000} /* (5, 11, 6) {real, imag} */,
  {32'h438a6350, 32'h00000000} /* (5, 11, 5) {real, imag} */,
  {32'h42998258, 32'h00000000} /* (5, 11, 4) {real, imag} */,
  {32'h4402525b, 32'h00000000} /* (5, 11, 3) {real, imag} */,
  {32'hc2e11028, 32'h00000000} /* (5, 11, 2) {real, imag} */,
  {32'hc35c9e46, 32'h00000000} /* (5, 11, 1) {real, imag} */,
  {32'hc3b5a6d5, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'hc3212de1, 32'h00000000} /* (5, 10, 15) {real, imag} */,
  {32'hc456ffce, 32'h00000000} /* (5, 10, 14) {real, imag} */,
  {32'hc487a484, 32'h00000000} /* (5, 10, 13) {real, imag} */,
  {32'hc45243f4, 32'h00000000} /* (5, 10, 12) {real, imag} */,
  {32'hc3c0546c, 32'h00000000} /* (5, 10, 11) {real, imag} */,
  {32'hc402501f, 32'h00000000} /* (5, 10, 10) {real, imag} */,
  {32'hc38d7bcb, 32'h00000000} /* (5, 10, 9) {real, imag} */,
  {32'hc390cbb1, 32'h00000000} /* (5, 10, 8) {real, imag} */,
  {32'hc3b824e0, 32'h00000000} /* (5, 10, 7) {real, imag} */,
  {32'h44495d1e, 32'h00000000} /* (5, 10, 6) {real, imag} */,
  {32'h4444241e, 32'h00000000} /* (5, 10, 5) {real, imag} */,
  {32'h4449e956, 32'h00000000} /* (5, 10, 4) {real, imag} */,
  {32'h43409928, 32'h00000000} /* (5, 10, 3) {real, imag} */,
  {32'h440ce327, 32'h00000000} /* (5, 10, 2) {real, imag} */,
  {32'h43ecde8d, 32'h00000000} /* (5, 10, 1) {real, imag} */,
  {32'h42bb2aa3, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'h42a9d394, 32'h00000000} /* (5, 9, 15) {real, imag} */,
  {32'h4236cbf8, 32'h00000000} /* (5, 9, 14) {real, imag} */,
  {32'h440ac6c9, 32'h00000000} /* (5, 9, 13) {real, imag} */,
  {32'hc4af41f4, 32'h00000000} /* (5, 9, 12) {real, imag} */,
  {32'hc3dac899, 32'h00000000} /* (5, 9, 11) {real, imag} */,
  {32'h4412ebea, 32'h00000000} /* (5, 9, 10) {real, imag} */,
  {32'h43674ddf, 32'h00000000} /* (5, 9, 9) {real, imag} */,
  {32'hc344742a, 32'h00000000} /* (5, 9, 8) {real, imag} */,
  {32'h43dbb7f7, 32'h00000000} /* (5, 9, 7) {real, imag} */,
  {32'hc3dc9fc6, 32'h00000000} /* (5, 9, 6) {real, imag} */,
  {32'h43a7c526, 32'h00000000} /* (5, 9, 5) {real, imag} */,
  {32'h4389ae1a, 32'h00000000} /* (5, 9, 4) {real, imag} */,
  {32'hc31db22e, 32'h00000000} /* (5, 9, 3) {real, imag} */,
  {32'h42d3b01e, 32'h00000000} /* (5, 9, 2) {real, imag} */,
  {32'h43267483, 32'h00000000} /* (5, 9, 1) {real, imag} */,
  {32'hc1e9a090, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'h4408cde2, 32'h00000000} /* (5, 8, 15) {real, imag} */,
  {32'h41aebabc, 32'h00000000} /* (5, 8, 14) {real, imag} */,
  {32'hc4920c79, 32'h00000000} /* (5, 8, 13) {real, imag} */,
  {32'hc4c1ec1f, 32'h00000000} /* (5, 8, 12) {real, imag} */,
  {32'hc3fd702a, 32'h00000000} /* (5, 8, 11) {real, imag} */,
  {32'h4395b78a, 32'h00000000} /* (5, 8, 10) {real, imag} */,
  {32'h42b02514, 32'h00000000} /* (5, 8, 9) {real, imag} */,
  {32'h43317169, 32'h00000000} /* (5, 8, 8) {real, imag} */,
  {32'h446dde22, 32'h00000000} /* (5, 8, 7) {real, imag} */,
  {32'hc2ed9617, 32'h00000000} /* (5, 8, 6) {real, imag} */,
  {32'h43572306, 32'h00000000} /* (5, 8, 5) {real, imag} */,
  {32'h44350182, 32'h00000000} /* (5, 8, 4) {real, imag} */,
  {32'hc3b1f916, 32'h00000000} /* (5, 8, 3) {real, imag} */,
  {32'h43058600, 32'h00000000} /* (5, 8, 2) {real, imag} */,
  {32'h431c03da, 32'h00000000} /* (5, 8, 1) {real, imag} */,
  {32'h440db4c6, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'h43a3dce0, 32'h00000000} /* (5, 7, 15) {real, imag} */,
  {32'hc1915c10, 32'h00000000} /* (5, 7, 14) {real, imag} */,
  {32'hc476365c, 32'h00000000} /* (5, 7, 13) {real, imag} */,
  {32'hc4c678bf, 32'h00000000} /* (5, 7, 12) {real, imag} */,
  {32'hc4fadbfb, 32'h00000000} /* (5, 7, 11) {real, imag} */,
  {32'h42e03d7a, 32'h00000000} /* (5, 7, 10) {real, imag} */,
  {32'hc1c9a760, 32'h00000000} /* (5, 7, 9) {real, imag} */,
  {32'h43ef5764, 32'h00000000} /* (5, 7, 8) {real, imag} */,
  {32'h41b325c0, 32'h00000000} /* (5, 7, 7) {real, imag} */,
  {32'h442bca76, 32'h00000000} /* (5, 7, 6) {real, imag} */,
  {32'h443e95ca, 32'h00000000} /* (5, 7, 5) {real, imag} */,
  {32'hc28cb630, 32'h00000000} /* (5, 7, 4) {real, imag} */,
  {32'hc3a43324, 32'h00000000} /* (5, 7, 3) {real, imag} */,
  {32'hc40e10db, 32'h00000000} /* (5, 7, 2) {real, imag} */,
  {32'h440de70c, 32'h00000000} /* (5, 7, 1) {real, imag} */,
  {32'hc3e40ba6, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'hc38b3bf5, 32'h00000000} /* (5, 6, 15) {real, imag} */,
  {32'h41923328, 32'h00000000} /* (5, 6, 14) {real, imag} */,
  {32'hc48106c1, 32'h00000000} /* (5, 6, 13) {real, imag} */,
  {32'hc48b5b4f, 32'h00000000} /* (5, 6, 12) {real, imag} */,
  {32'hc470c5b8, 32'h00000000} /* (5, 6, 11) {real, imag} */,
  {32'h42bc1ab8, 32'h00000000} /* (5, 6, 10) {real, imag} */,
  {32'hc3ef174e, 32'h00000000} /* (5, 6, 9) {real, imag} */,
  {32'hc1356a50, 32'h00000000} /* (5, 6, 8) {real, imag} */,
  {32'h431560de, 32'h00000000} /* (5, 6, 7) {real, imag} */,
  {32'hc3933f00, 32'h00000000} /* (5, 6, 6) {real, imag} */,
  {32'h44104551, 32'h00000000} /* (5, 6, 5) {real, imag} */,
  {32'hc3f3aa5d, 32'h00000000} /* (5, 6, 4) {real, imag} */,
  {32'hc47802e4, 32'h00000000} /* (5, 6, 3) {real, imag} */,
  {32'hc4f2f244, 32'h00000000} /* (5, 6, 2) {real, imag} */,
  {32'hc46c5e63, 32'h00000000} /* (5, 6, 1) {real, imag} */,
  {32'hc380e840, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'hc46ac376, 32'h00000000} /* (5, 5, 15) {real, imag} */,
  {32'hc242f64a, 32'h00000000} /* (5, 5, 14) {real, imag} */,
  {32'hc41c724e, 32'h00000000} /* (5, 5, 13) {real, imag} */,
  {32'hc4341388, 32'h00000000} /* (5, 5, 12) {real, imag} */,
  {32'hc389cb72, 32'h00000000} /* (5, 5, 11) {real, imag} */,
  {32'hc3e9cfd9, 32'h00000000} /* (5, 5, 10) {real, imag} */,
  {32'hc3b07298, 32'h00000000} /* (5, 5, 9) {real, imag} */,
  {32'h421365e0, 32'h00000000} /* (5, 5, 8) {real, imag} */,
  {32'h428c7a5c, 32'h00000000} /* (5, 5, 7) {real, imag} */,
  {32'h429edd55, 32'h00000000} /* (5, 5, 6) {real, imag} */,
  {32'hc390478f, 32'h00000000} /* (5, 5, 5) {real, imag} */,
  {32'hc437925c, 32'h00000000} /* (5, 5, 4) {real, imag} */,
  {32'hc459d48f, 32'h00000000} /* (5, 5, 3) {real, imag} */,
  {32'hc48c6c75, 32'h00000000} /* (5, 5, 2) {real, imag} */,
  {32'hc5066883, 32'h00000000} /* (5, 5, 1) {real, imag} */,
  {32'hc3811216, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'h439dcbd6, 32'h00000000} /* (5, 4, 15) {real, imag} */,
  {32'h434c8d04, 32'h00000000} /* (5, 4, 14) {real, imag} */,
  {32'hc444711f, 32'h00000000} /* (5, 4, 13) {real, imag} */,
  {32'hc424e6ff, 32'h00000000} /* (5, 4, 12) {real, imag} */,
  {32'hc3d54974, 32'h00000000} /* (5, 4, 11) {real, imag} */,
  {32'h43b690cf, 32'h00000000} /* (5, 4, 10) {real, imag} */,
  {32'h43f0e92c, 32'h00000000} /* (5, 4, 9) {real, imag} */,
  {32'hc3ac5b8b, 32'h00000000} /* (5, 4, 8) {real, imag} */,
  {32'hc30364ab, 32'h00000000} /* (5, 4, 7) {real, imag} */,
  {32'h42cc713f, 32'h00000000} /* (5, 4, 6) {real, imag} */,
  {32'h444f8fcd, 32'h00000000} /* (5, 4, 5) {real, imag} */,
  {32'hc3c379f6, 32'h00000000} /* (5, 4, 4) {real, imag} */,
  {32'hc4e125d9, 32'h00000000} /* (5, 4, 3) {real, imag} */,
  {32'hc46c8a1c, 32'h00000000} /* (5, 4, 2) {real, imag} */,
  {32'hc4576710, 32'h00000000} /* (5, 4, 1) {real, imag} */,
  {32'hc49c7fc2, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'hc43b225e, 32'h00000000} /* (5, 3, 15) {real, imag} */,
  {32'h43611d60, 32'h00000000} /* (5, 3, 14) {real, imag} */,
  {32'h4332e130, 32'h00000000} /* (5, 3, 13) {real, imag} */,
  {32'hc3cf0b08, 32'h00000000} /* (5, 3, 12) {real, imag} */,
  {32'h4436a62e, 32'h00000000} /* (5, 3, 11) {real, imag} */,
  {32'h441cc20b, 32'h00000000} /* (5, 3, 10) {real, imag} */,
  {32'hc40428e5, 32'h00000000} /* (5, 3, 9) {real, imag} */,
  {32'hc424072f, 32'h00000000} /* (5, 3, 8) {real, imag} */,
  {32'hc38eb64d, 32'h00000000} /* (5, 3, 7) {real, imag} */,
  {32'hc3c23d68, 32'h00000000} /* (5, 3, 6) {real, imag} */,
  {32'hc303c5fa, 32'h00000000} /* (5, 3, 5) {real, imag} */,
  {32'hc50d1271, 32'h00000000} /* (5, 3, 4) {real, imag} */,
  {32'hc48782c5, 32'h00000000} /* (5, 3, 3) {real, imag} */,
  {32'hc4ab8292, 32'h00000000} /* (5, 3, 2) {real, imag} */,
  {32'hc3af0ef1, 32'h00000000} /* (5, 3, 1) {real, imag} */,
  {32'hc3f1916a, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'hc4966b79, 32'h00000000} /* (5, 2, 15) {real, imag} */,
  {32'hc480a5a7, 32'h00000000} /* (5, 2, 14) {real, imag} */,
  {32'h438f0791, 32'h00000000} /* (5, 2, 13) {real, imag} */,
  {32'hc401d406, 32'h00000000} /* (5, 2, 12) {real, imag} */,
  {32'h4339d8a0, 32'h00000000} /* (5, 2, 11) {real, imag} */,
  {32'hc4d96a58, 32'h00000000} /* (5, 2, 10) {real, imag} */,
  {32'hc27755c0, 32'h00000000} /* (5, 2, 9) {real, imag} */,
  {32'h43966f5a, 32'h00000000} /* (5, 2, 8) {real, imag} */,
  {32'h42c592f0, 32'h00000000} /* (5, 2, 7) {real, imag} */,
  {32'hc3906a41, 32'h00000000} /* (5, 2, 6) {real, imag} */,
  {32'h4410e006, 32'h00000000} /* (5, 2, 5) {real, imag} */,
  {32'h43c702a0, 32'h00000000} /* (5, 2, 4) {real, imag} */,
  {32'hc3aa67e4, 32'h00000000} /* (5, 2, 3) {real, imag} */,
  {32'hc467b0b1, 32'h00000000} /* (5, 2, 2) {real, imag} */,
  {32'hc49fb19b, 32'h00000000} /* (5, 2, 1) {real, imag} */,
  {32'hc48325cc, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'hc491c6cf, 32'h00000000} /* (5, 1, 15) {real, imag} */,
  {32'hc34e19d7, 32'h00000000} /* (5, 1, 14) {real, imag} */,
  {32'h431a8c99, 32'h00000000} /* (5, 1, 13) {real, imag} */,
  {32'h4337e0f4, 32'h00000000} /* (5, 1, 12) {real, imag} */,
  {32'hc415369a, 32'h00000000} /* (5, 1, 11) {real, imag} */,
  {32'h43cfd3f3, 32'h00000000} /* (5, 1, 10) {real, imag} */,
  {32'h43eb18b0, 32'h00000000} /* (5, 1, 9) {real, imag} */,
  {32'hc3961cf5, 32'h00000000} /* (5, 1, 8) {real, imag} */,
  {32'hc4405066, 32'h00000000} /* (5, 1, 7) {real, imag} */,
  {32'h41db6418, 32'h00000000} /* (5, 1, 6) {real, imag} */,
  {32'h439164f0, 32'h00000000} /* (5, 1, 5) {real, imag} */,
  {32'hc24616e0, 32'h00000000} /* (5, 1, 4) {real, imag} */,
  {32'hc4a44391, 32'h00000000} /* (5, 1, 3) {real, imag} */,
  {32'hc48b7699, 32'h00000000} /* (5, 1, 2) {real, imag} */,
  {32'hc43260c2, 32'h00000000} /* (5, 1, 1) {real, imag} */,
  {32'hc4967d1d, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'hc4005e3d, 32'h00000000} /* (5, 0, 15) {real, imag} */,
  {32'hc3a163f8, 32'h00000000} /* (5, 0, 14) {real, imag} */,
  {32'hc3889429, 32'h00000000} /* (5, 0, 13) {real, imag} */,
  {32'hc4511fac, 32'h00000000} /* (5, 0, 12) {real, imag} */,
  {32'hc3845a4f, 32'h00000000} /* (5, 0, 11) {real, imag} */,
  {32'hc41da47f, 32'h00000000} /* (5, 0, 10) {real, imag} */,
  {32'hc40c7308, 32'h00000000} /* (5, 0, 9) {real, imag} */,
  {32'h440aea66, 32'h00000000} /* (5, 0, 8) {real, imag} */,
  {32'hc2503ea4, 32'h00000000} /* (5, 0, 7) {real, imag} */,
  {32'hc1f38c20, 32'h00000000} /* (5, 0, 6) {real, imag} */,
  {32'h43296162, 32'h00000000} /* (5, 0, 5) {real, imag} */,
  {32'hc3ef3a91, 32'h00000000} /* (5, 0, 4) {real, imag} */,
  {32'h424a58aa, 32'h00000000} /* (5, 0, 3) {real, imag} */,
  {32'hc3bcf315, 32'h00000000} /* (5, 0, 2) {real, imag} */,
  {32'hc4587a30, 32'h00000000} /* (5, 0, 1) {real, imag} */,
  {32'hc4220d4a, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hc3f18e20, 32'h00000000} /* (4, 15, 15) {real, imag} */,
  {32'hc40bc682, 32'h00000000} /* (4, 15, 14) {real, imag} */,
  {32'h431456f0, 32'h00000000} /* (4, 15, 13) {real, imag} */,
  {32'h43880006, 32'h00000000} /* (4, 15, 12) {real, imag} */,
  {32'hc29f3edc, 32'h00000000} /* (4, 15, 11) {real, imag} */,
  {32'hc323da75, 32'h00000000} /* (4, 15, 10) {real, imag} */,
  {32'hc3988fb9, 32'h00000000} /* (4, 15, 9) {real, imag} */,
  {32'hc3ba41fa, 32'h00000000} /* (4, 15, 8) {real, imag} */,
  {32'hc3951640, 32'h00000000} /* (4, 15, 7) {real, imag} */,
  {32'h433208dc, 32'h00000000} /* (4, 15, 6) {real, imag} */,
  {32'h43f9c60a, 32'h00000000} /* (4, 15, 5) {real, imag} */,
  {32'h42a91636, 32'h00000000} /* (4, 15, 4) {real, imag} */,
  {32'hc3119f94, 32'h00000000} /* (4, 15, 3) {real, imag} */,
  {32'hc3d4ca74, 32'h00000000} /* (4, 15, 2) {real, imag} */,
  {32'hc3db2f2d, 32'h00000000} /* (4, 15, 1) {real, imag} */,
  {32'hc3e3bca2, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'hc43ef347, 32'h00000000} /* (4, 14, 15) {real, imag} */,
  {32'hc4b2a55d, 32'h00000000} /* (4, 14, 14) {real, imag} */,
  {32'hc3f9a29b, 32'h00000000} /* (4, 14, 13) {real, imag} */,
  {32'hc42701f4, 32'h00000000} /* (4, 14, 12) {real, imag} */,
  {32'hc32ac263, 32'h00000000} /* (4, 14, 11) {real, imag} */,
  {32'hc4924e40, 32'h00000000} /* (4, 14, 10) {real, imag} */,
  {32'hc4ad2995, 32'h00000000} /* (4, 14, 9) {real, imag} */,
  {32'hc42cf725, 32'h00000000} /* (4, 14, 8) {real, imag} */,
  {32'hc30559bc, 32'h00000000} /* (4, 14, 7) {real, imag} */,
  {32'h43ccaffd, 32'h00000000} /* (4, 14, 6) {real, imag} */,
  {32'hc2b2677c, 32'h00000000} /* (4, 14, 5) {real, imag} */,
  {32'h420a8880, 32'h00000000} /* (4, 14, 4) {real, imag} */,
  {32'hc2ea641a, 32'h00000000} /* (4, 14, 3) {real, imag} */,
  {32'hc3e52e6e, 32'h00000000} /* (4, 14, 2) {real, imag} */,
  {32'h43bd1233, 32'h00000000} /* (4, 14, 1) {real, imag} */,
  {32'h43806a2a, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'hc3ad8af1, 32'h00000000} /* (4, 13, 15) {real, imag} */,
  {32'hc486362b, 32'h00000000} /* (4, 13, 14) {real, imag} */,
  {32'hc4745fe9, 32'h00000000} /* (4, 13, 13) {real, imag} */,
  {32'h4401fb02, 32'h00000000} /* (4, 13, 12) {real, imag} */,
  {32'hc48cb09c, 32'h00000000} /* (4, 13, 11) {real, imag} */,
  {32'hc468f06c, 32'h00000000} /* (4, 13, 10) {real, imag} */,
  {32'hc4a10ea9, 32'h00000000} /* (4, 13, 9) {real, imag} */,
  {32'h41b29048, 32'h00000000} /* (4, 13, 8) {real, imag} */,
  {32'h44632150, 32'h00000000} /* (4, 13, 7) {real, imag} */,
  {32'h43fe0490, 32'h00000000} /* (4, 13, 6) {real, imag} */,
  {32'h42033430, 32'h00000000} /* (4, 13, 5) {real, imag} */,
  {32'h438a8beb, 32'h00000000} /* (4, 13, 4) {real, imag} */,
  {32'h44134216, 32'h00000000} /* (4, 13, 3) {real, imag} */,
  {32'hc3919cf4, 32'h00000000} /* (4, 13, 2) {real, imag} */,
  {32'hc3e71b80, 32'h00000000} /* (4, 13, 1) {real, imag} */,
  {32'hc28a58ea, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'hc43cac4f, 32'h00000000} /* (4, 12, 15) {real, imag} */,
  {32'hc410b585, 32'h00000000} /* (4, 12, 14) {real, imag} */,
  {32'h44090f56, 32'h00000000} /* (4, 12, 13) {real, imag} */,
  {32'h420ca07c, 32'h00000000} /* (4, 12, 12) {real, imag} */,
  {32'hc451734c, 32'h00000000} /* (4, 12, 11) {real, imag} */,
  {32'hc431f061, 32'h00000000} /* (4, 12, 10) {real, imag} */,
  {32'hc3c4cdc2, 32'h00000000} /* (4, 12, 9) {real, imag} */,
  {32'hc251961e, 32'h00000000} /* (4, 12, 8) {real, imag} */,
  {32'hc4121e45, 32'h00000000} /* (4, 12, 7) {real, imag} */,
  {32'h43b46a32, 32'h00000000} /* (4, 12, 6) {real, imag} */,
  {32'h44c7d58d, 32'h00000000} /* (4, 12, 5) {real, imag} */,
  {32'hc39a4eaa, 32'h00000000} /* (4, 12, 4) {real, imag} */,
  {32'hc2802d64, 32'h00000000} /* (4, 12, 3) {real, imag} */,
  {32'hc4004e3b, 32'h00000000} /* (4, 12, 2) {real, imag} */,
  {32'h43c8f546, 32'h00000000} /* (4, 12, 1) {real, imag} */,
  {32'hc387d43d, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'hc3ddbc0a, 32'h00000000} /* (4, 11, 15) {real, imag} */,
  {32'hc3e0876b, 32'h00000000} /* (4, 11, 14) {real, imag} */,
  {32'h430dc7c0, 32'h00000000} /* (4, 11, 13) {real, imag} */,
  {32'hc39f820e, 32'h00000000} /* (4, 11, 12) {real, imag} */,
  {32'hc49cab2a, 32'h00000000} /* (4, 11, 11) {real, imag} */,
  {32'hc43d7410, 32'h00000000} /* (4, 11, 10) {real, imag} */,
  {32'hc3d45e70, 32'h00000000} /* (4, 11, 9) {real, imag} */,
  {32'hc48a071a, 32'h00000000} /* (4, 11, 8) {real, imag} */,
  {32'h4457c8d3, 32'h00000000} /* (4, 11, 7) {real, imag} */,
  {32'h4490056c, 32'h00000000} /* (4, 11, 6) {real, imag} */,
  {32'h44c88018, 32'h00000000} /* (4, 11, 5) {real, imag} */,
  {32'h44077c6f, 32'h00000000} /* (4, 11, 4) {real, imag} */,
  {32'hc3109d5c, 32'h00000000} /* (4, 11, 3) {real, imag} */,
  {32'h433de814, 32'h00000000} /* (4, 11, 2) {real, imag} */,
  {32'h41000d00, 32'h00000000} /* (4, 11, 1) {real, imag} */,
  {32'h437b7a24, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'hc2a46d4d, 32'h00000000} /* (4, 10, 15) {real, imag} */,
  {32'hc33a130b, 32'h00000000} /* (4, 10, 14) {real, imag} */,
  {32'h4352c478, 32'h00000000} /* (4, 10, 13) {real, imag} */,
  {32'h42c2c39a, 32'h00000000} /* (4, 10, 12) {real, imag} */,
  {32'hc3d3305d, 32'h00000000} /* (4, 10, 11) {real, imag} */,
  {32'hc19d7228, 32'h00000000} /* (4, 10, 10) {real, imag} */,
  {32'hc4564c88, 32'h00000000} /* (4, 10, 9) {real, imag} */,
  {32'h43451d38, 32'h00000000} /* (4, 10, 8) {real, imag} */,
  {32'hc137a328, 32'h00000000} /* (4, 10, 7) {real, imag} */,
  {32'h43315d5b, 32'h00000000} /* (4, 10, 6) {real, imag} */,
  {32'h443d15fd, 32'h00000000} /* (4, 10, 5) {real, imag} */,
  {32'h440fdf09, 32'h00000000} /* (4, 10, 4) {real, imag} */,
  {32'h41c7d210, 32'h00000000} /* (4, 10, 3) {real, imag} */,
  {32'hc3f6d414, 32'h00000000} /* (4, 10, 2) {real, imag} */,
  {32'hc3904778, 32'h00000000} /* (4, 10, 1) {real, imag} */,
  {32'h439d9b94, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'hc3bdb0c6, 32'h00000000} /* (4, 9, 15) {real, imag} */,
  {32'hc3e1cbe9, 32'h00000000} /* (4, 9, 14) {real, imag} */,
  {32'h42dc01f3, 32'h00000000} /* (4, 9, 13) {real, imag} */,
  {32'hc455b2ca, 32'h00000000} /* (4, 9, 12) {real, imag} */,
  {32'hc453c909, 32'h00000000} /* (4, 9, 11) {real, imag} */,
  {32'hc2f4c928, 32'h00000000} /* (4, 9, 10) {real, imag} */,
  {32'hc412bffc, 32'h00000000} /* (4, 9, 9) {real, imag} */,
  {32'h4396e098, 32'h00000000} /* (4, 9, 8) {real, imag} */,
  {32'h441595cd, 32'h00000000} /* (4, 9, 7) {real, imag} */,
  {32'hc427b06f, 32'h00000000} /* (4, 9, 6) {real, imag} */,
  {32'h404add20, 32'h00000000} /* (4, 9, 5) {real, imag} */,
  {32'hc41811da, 32'h00000000} /* (4, 9, 4) {real, imag} */,
  {32'hc34caddc, 32'h00000000} /* (4, 9, 3) {real, imag} */,
  {32'hc3a09c29, 32'h00000000} /* (4, 9, 2) {real, imag} */,
  {32'h420f21a8, 32'h00000000} /* (4, 9, 1) {real, imag} */,
  {32'h4413b1df, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'h4481bc25, 32'h00000000} /* (4, 8, 15) {real, imag} */,
  {32'h423df408, 32'h00000000} /* (4, 8, 14) {real, imag} */,
  {32'hc3f75168, 32'h00000000} /* (4, 8, 13) {real, imag} */,
  {32'hc450097a, 32'h00000000} /* (4, 8, 12) {real, imag} */,
  {32'hc4672510, 32'h00000000} /* (4, 8, 11) {real, imag} */,
  {32'hc2bbc7e0, 32'h00000000} /* (4, 8, 10) {real, imag} */,
  {32'hc2cfe162, 32'h00000000} /* (4, 8, 9) {real, imag} */,
  {32'hc483624c, 32'h00000000} /* (4, 8, 8) {real, imag} */,
  {32'h4292e9fc, 32'h00000000} /* (4, 8, 7) {real, imag} */,
  {32'h4428b134, 32'h00000000} /* (4, 8, 6) {real, imag} */,
  {32'h4410bc84, 32'h00000000} /* (4, 8, 5) {real, imag} */,
  {32'hc3b22234, 32'h00000000} /* (4, 8, 4) {real, imag} */,
  {32'hc487ff4b, 32'h00000000} /* (4, 8, 3) {real, imag} */,
  {32'hc4180757, 32'h00000000} /* (4, 8, 2) {real, imag} */,
  {32'h43c93708, 32'h00000000} /* (4, 8, 1) {real, imag} */,
  {32'h43bb946e, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'hc0d9a8d0, 32'h00000000} /* (4, 7, 15) {real, imag} */,
  {32'h43939b3e, 32'h00000000} /* (4, 7, 14) {real, imag} */,
  {32'hc414bb66, 32'h00000000} /* (4, 7, 13) {real, imag} */,
  {32'hc40ebfee, 32'h00000000} /* (4, 7, 12) {real, imag} */,
  {32'hc46a83b6, 32'h00000000} /* (4, 7, 11) {real, imag} */,
  {32'hc41fdf30, 32'h00000000} /* (4, 7, 10) {real, imag} */,
  {32'h447e6685, 32'h00000000} /* (4, 7, 9) {real, imag} */,
  {32'hc338133c, 32'h00000000} /* (4, 7, 8) {real, imag} */,
  {32'h432c82d2, 32'h00000000} /* (4, 7, 7) {real, imag} */,
  {32'hc38e94d2, 32'h00000000} /* (4, 7, 6) {real, imag} */,
  {32'h43229bf0, 32'h00000000} /* (4, 7, 5) {real, imag} */,
  {32'hc43f612a, 32'h00000000} /* (4, 7, 4) {real, imag} */,
  {32'hc425f946, 32'h00000000} /* (4, 7, 3) {real, imag} */,
  {32'hc39de3f5, 32'h00000000} /* (4, 7, 2) {real, imag} */,
  {32'hc47053f7, 32'h00000000} /* (4, 7, 1) {real, imag} */,
  {32'hc139ec80, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'hc36b688f, 32'h00000000} /* (4, 6, 15) {real, imag} */,
  {32'hc43df9dc, 32'h00000000} /* (4, 6, 14) {real, imag} */,
  {32'hc4942dc9, 32'h00000000} /* (4, 6, 13) {real, imag} */,
  {32'hc4d93f5c, 32'h00000000} /* (4, 6, 12) {real, imag} */,
  {32'hc4841e8e, 32'h00000000} /* (4, 6, 11) {real, imag} */,
  {32'hc4527a23, 32'h00000000} /* (4, 6, 10) {real, imag} */,
  {32'h44040754, 32'h00000000} /* (4, 6, 9) {real, imag} */,
  {32'h42f09ba8, 32'h00000000} /* (4, 6, 8) {real, imag} */,
  {32'h41ecad58, 32'h00000000} /* (4, 6, 7) {real, imag} */,
  {32'h4412bcd2, 32'h00000000} /* (4, 6, 6) {real, imag} */,
  {32'hc44bb8bb, 32'h00000000} /* (4, 6, 5) {real, imag} */,
  {32'hc3a6205a, 32'h00000000} /* (4, 6, 4) {real, imag} */,
  {32'hc4646041, 32'h00000000} /* (4, 6, 3) {real, imag} */,
  {32'hc49f19e6, 32'h00000000} /* (4, 6, 2) {real, imag} */,
  {32'hc4a44151, 32'h00000000} /* (4, 6, 1) {real, imag} */,
  {32'hc426b0d5, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'hc3fa3c6d, 32'h00000000} /* (4, 5, 15) {real, imag} */,
  {32'hc44179ae, 32'h00000000} /* (4, 5, 14) {real, imag} */,
  {32'hc486ccdd, 32'h00000000} /* (4, 5, 13) {real, imag} */,
  {32'hc386dd18, 32'h00000000} /* (4, 5, 12) {real, imag} */,
  {32'hc323673b, 32'h00000000} /* (4, 5, 11) {real, imag} */,
  {32'hc30077bc, 32'h00000000} /* (4, 5, 10) {real, imag} */,
  {32'hc1c5eb28, 32'h00000000} /* (4, 5, 9) {real, imag} */,
  {32'h43e8023c, 32'h00000000} /* (4, 5, 8) {real, imag} */,
  {32'h43804a95, 32'h00000000} /* (4, 5, 7) {real, imag} */,
  {32'h44943733, 32'h00000000} /* (4, 5, 6) {real, imag} */,
  {32'hc1094380, 32'h00000000} /* (4, 5, 5) {real, imag} */,
  {32'hc3b5f9b0, 32'h00000000} /* (4, 5, 4) {real, imag} */,
  {32'hc39b9f02, 32'h00000000} /* (4, 5, 3) {real, imag} */,
  {32'hc48adee4, 32'h00000000} /* (4, 5, 2) {real, imag} */,
  {32'hc3ac4338, 32'h00000000} /* (4, 5, 1) {real, imag} */,
  {32'hc4658c5e, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'hc4624a32, 32'h00000000} /* (4, 4, 15) {real, imag} */,
  {32'hc45dd248, 32'h00000000} /* (4, 4, 14) {real, imag} */,
  {32'hc4284444, 32'h00000000} /* (4, 4, 13) {real, imag} */,
  {32'h4308fcac, 32'h00000000} /* (4, 4, 12) {real, imag} */,
  {32'h4410d3ea, 32'h00000000} /* (4, 4, 11) {real, imag} */,
  {32'h43af54b7, 32'h00000000} /* (4, 4, 10) {real, imag} */,
  {32'h43eb982e, 32'h00000000} /* (4, 4, 9) {real, imag} */,
  {32'hc40b4458, 32'h00000000} /* (4, 4, 8) {real, imag} */,
  {32'hc48f3b47, 32'h00000000} /* (4, 4, 7) {real, imag} */,
  {32'hc36f4bd0, 32'h00000000} /* (4, 4, 6) {real, imag} */,
  {32'hc1ca5e30, 32'h00000000} /* (4, 4, 5) {real, imag} */,
  {32'hc45fccb1, 32'h00000000} /* (4, 4, 4) {real, imag} */,
  {32'hc48e265e, 32'h00000000} /* (4, 4, 3) {real, imag} */,
  {32'hc480db69, 32'h00000000} /* (4, 4, 2) {real, imag} */,
  {32'hc458a74b, 32'h00000000} /* (4, 4, 1) {real, imag} */,
  {32'hc3a2c6af, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'hc47728f7, 32'h00000000} /* (4, 3, 15) {real, imag} */,
  {32'hc443902a, 32'h00000000} /* (4, 3, 14) {real, imag} */,
  {32'hc450e53c, 32'h00000000} /* (4, 3, 13) {real, imag} */,
  {32'h43d35730, 32'h00000000} /* (4, 3, 12) {real, imag} */,
  {32'h43ec9d8f, 32'h00000000} /* (4, 3, 11) {real, imag} */,
  {32'hc3b0ca84, 32'h00000000} /* (4, 3, 10) {real, imag} */,
  {32'h441bc47c, 32'h00000000} /* (4, 3, 9) {real, imag} */,
  {32'hc3fbfea0, 32'h00000000} /* (4, 3, 8) {real, imag} */,
  {32'hc2fc2c28, 32'h00000000} /* (4, 3, 7) {real, imag} */,
  {32'hc3b46d80, 32'h00000000} /* (4, 3, 6) {real, imag} */,
  {32'hc4870d30, 32'h00000000} /* (4, 3, 5) {real, imag} */,
  {32'hc4a4dbc2, 32'h00000000} /* (4, 3, 4) {real, imag} */,
  {32'hc4b14206, 32'h00000000} /* (4, 3, 3) {real, imag} */,
  {32'hc4aaf94a, 32'h00000000} /* (4, 3, 2) {real, imag} */,
  {32'hc4f4b920, 32'h00000000} /* (4, 3, 1) {real, imag} */,
  {32'hc314e090, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'hc48d733f, 32'h00000000} /* (4, 2, 15) {real, imag} */,
  {32'hc4625a5a, 32'h00000000} /* (4, 2, 14) {real, imag} */,
  {32'hc2e70920, 32'h00000000} /* (4, 2, 13) {real, imag} */,
  {32'h44800f64, 32'h00000000} /* (4, 2, 12) {real, imag} */,
  {32'h420c8960, 32'h00000000} /* (4, 2, 11) {real, imag} */,
  {32'hc3c76a05, 32'h00000000} /* (4, 2, 10) {real, imag} */,
  {32'hc3f93b26, 32'h00000000} /* (4, 2, 9) {real, imag} */,
  {32'hc3634e26, 32'h00000000} /* (4, 2, 8) {real, imag} */,
  {32'hc310ffe8, 32'h00000000} /* (4, 2, 7) {real, imag} */,
  {32'hc415921a, 32'h00000000} /* (4, 2, 6) {real, imag} */,
  {32'hc42abd6d, 32'h00000000} /* (4, 2, 5) {real, imag} */,
  {32'hc4a587f4, 32'h00000000} /* (4, 2, 4) {real, imag} */,
  {32'hc4b8d0a3, 32'h00000000} /* (4, 2, 3) {real, imag} */,
  {32'hc4a074ef, 32'h00000000} /* (4, 2, 2) {real, imag} */,
  {32'hc433527d, 32'h00000000} /* (4, 2, 1) {real, imag} */,
  {32'hc432d7aa, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'hc42cb271, 32'h00000000} /* (4, 1, 15) {real, imag} */,
  {32'hc39423f1, 32'h00000000} /* (4, 1, 14) {real, imag} */,
  {32'h4408c9ae, 32'h00000000} /* (4, 1, 13) {real, imag} */,
  {32'hc2825f80, 32'h00000000} /* (4, 1, 12) {real, imag} */,
  {32'hc3bbcbec, 32'h00000000} /* (4, 1, 11) {real, imag} */,
  {32'h43345398, 32'h00000000} /* (4, 1, 10) {real, imag} */,
  {32'hc309cdb0, 32'h00000000} /* (4, 1, 9) {real, imag} */,
  {32'hc2761d08, 32'h00000000} /* (4, 1, 8) {real, imag} */,
  {32'hc37365c3, 32'h00000000} /* (4, 1, 7) {real, imag} */,
  {32'hc3b12cdb, 32'h00000000} /* (4, 1, 6) {real, imag} */,
  {32'h43ae910c, 32'h00000000} /* (4, 1, 5) {real, imag} */,
  {32'hc42c95e4, 32'h00000000} /* (4, 1, 4) {real, imag} */,
  {32'hc428cca4, 32'h00000000} /* (4, 1, 3) {real, imag} */,
  {32'hc4868e74, 32'h00000000} /* (4, 1, 2) {real, imag} */,
  {32'hc498b9ea, 32'h00000000} /* (4, 1, 1) {real, imag} */,
  {32'hc42f7154, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'hc425643d, 32'h00000000} /* (4, 0, 15) {real, imag} */,
  {32'hc38cd322, 32'h00000000} /* (4, 0, 14) {real, imag} */,
  {32'hc3721b8c, 32'h00000000} /* (4, 0, 13) {real, imag} */,
  {32'hc463d857, 32'h00000000} /* (4, 0, 12) {real, imag} */,
  {32'hc478dc45, 32'h00000000} /* (4, 0, 11) {real, imag} */,
  {32'hc35f5560, 32'h00000000} /* (4, 0, 10) {real, imag} */,
  {32'hc2f5b738, 32'h00000000} /* (4, 0, 9) {real, imag} */,
  {32'h43a307ac, 32'h00000000} /* (4, 0, 8) {real, imag} */,
  {32'hc2a6ead8, 32'h00000000} /* (4, 0, 7) {real, imag} */,
  {32'h4335968c, 32'h00000000} /* (4, 0, 6) {real, imag} */,
  {32'h4392cef8, 32'h00000000} /* (4, 0, 5) {real, imag} */,
  {32'hc2ccbfc8, 32'h00000000} /* (4, 0, 4) {real, imag} */,
  {32'hc3bd5f96, 32'h00000000} /* (4, 0, 3) {real, imag} */,
  {32'hc4762b66, 32'h00000000} /* (4, 0, 2) {real, imag} */,
  {32'hc4676c55, 32'h00000000} /* (4, 0, 1) {real, imag} */,
  {32'hc4130857, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hc3c4e45e, 32'h00000000} /* (3, 15, 15) {real, imag} */,
  {32'hc451f914, 32'h00000000} /* (3, 15, 14) {real, imag} */,
  {32'hc3a3186e, 32'h00000000} /* (3, 15, 13) {real, imag} */,
  {32'hc2bb4c68, 32'h00000000} /* (3, 15, 12) {real, imag} */,
  {32'h438f4123, 32'h00000000} /* (3, 15, 11) {real, imag} */,
  {32'h4204379e, 32'h00000000} /* (3, 15, 10) {real, imag} */,
  {32'hc1b299a0, 32'h00000000} /* (3, 15, 9) {real, imag} */,
  {32'h43187738, 32'h00000000} /* (3, 15, 8) {real, imag} */,
  {32'h43a63894, 32'h00000000} /* (3, 15, 7) {real, imag} */,
  {32'h42461f38, 32'h00000000} /* (3, 15, 6) {real, imag} */,
  {32'h43419c5c, 32'h00000000} /* (3, 15, 5) {real, imag} */,
  {32'hc48f07fc, 32'h00000000} /* (3, 15, 4) {real, imag} */,
  {32'hc3688bca, 32'h00000000} /* (3, 15, 3) {real, imag} */,
  {32'hc31a8cda, 32'h00000000} /* (3, 15, 2) {real, imag} */,
  {32'hc433c6a1, 32'h00000000} /* (3, 15, 1) {real, imag} */,
  {32'hc436ebac, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'hc2f7aaee, 32'h00000000} /* (3, 14, 15) {real, imag} */,
  {32'hc44172ca, 32'h00000000} /* (3, 14, 14) {real, imag} */,
  {32'hc457c8f2, 32'h00000000} /* (3, 14, 13) {real, imag} */,
  {32'h434af2bd, 32'h00000000} /* (3, 14, 12) {real, imag} */,
  {32'h445cd467, 32'h00000000} /* (3, 14, 11) {real, imag} */,
  {32'hc405c89b, 32'h00000000} /* (3, 14, 10) {real, imag} */,
  {32'hc43de808, 32'h00000000} /* (3, 14, 9) {real, imag} */,
  {32'h44634908, 32'h00000000} /* (3, 14, 8) {real, imag} */,
  {32'hc300e40d, 32'h00000000} /* (3, 14, 7) {real, imag} */,
  {32'hc4052fec, 32'h00000000} /* (3, 14, 6) {real, imag} */,
  {32'h43cc6791, 32'h00000000} /* (3, 14, 5) {real, imag} */,
  {32'h439a519e, 32'h00000000} /* (3, 14, 4) {real, imag} */,
  {32'hc3f4070e, 32'h00000000} /* (3, 14, 3) {real, imag} */,
  {32'hc38f0e86, 32'h00000000} /* (3, 14, 2) {real, imag} */,
  {32'hc4694ed8, 32'h00000000} /* (3, 14, 1) {real, imag} */,
  {32'h42059c60, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'hc341a5ee, 32'h00000000} /* (3, 13, 15) {real, imag} */,
  {32'hc45f44de, 32'h00000000} /* (3, 13, 14) {real, imag} */,
  {32'hc38f19df, 32'h00000000} /* (3, 13, 13) {real, imag} */,
  {32'h442b478c, 32'h00000000} /* (3, 13, 12) {real, imag} */,
  {32'hc0ead040, 32'h00000000} /* (3, 13, 11) {real, imag} */,
  {32'hc41a6621, 32'h00000000} /* (3, 13, 10) {real, imag} */,
  {32'hc3f1a500, 32'h00000000} /* (3, 13, 9) {real, imag} */,
  {32'h436b4004, 32'h00000000} /* (3, 13, 8) {real, imag} */,
  {32'hc37ce4ce, 32'h00000000} /* (3, 13, 7) {real, imag} */,
  {32'h43a8784c, 32'h00000000} /* (3, 13, 6) {real, imag} */,
  {32'h43f9d9bd, 32'h00000000} /* (3, 13, 5) {real, imag} */,
  {32'h42b89e54, 32'h00000000} /* (3, 13, 4) {real, imag} */,
  {32'h4423a546, 32'h00000000} /* (3, 13, 3) {real, imag} */,
  {32'hc324c353, 32'h00000000} /* (3, 13, 2) {real, imag} */,
  {32'h4381862e, 32'h00000000} /* (3, 13, 1) {real, imag} */,
  {32'h432b6928, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'hc1e1a830, 32'h00000000} /* (3, 12, 15) {real, imag} */,
  {32'hc38d254a, 32'h00000000} /* (3, 12, 14) {real, imag} */,
  {32'h44359ab8, 32'h00000000} /* (3, 12, 13) {real, imag} */,
  {32'h445468d1, 32'h00000000} /* (3, 12, 12) {real, imag} */,
  {32'hc41e8e93, 32'h00000000} /* (3, 12, 11) {real, imag} */,
  {32'hc3f179c4, 32'h00000000} /* (3, 12, 10) {real, imag} */,
  {32'hc417daf8, 32'h00000000} /* (3, 12, 9) {real, imag} */,
  {32'hc3e1fd95, 32'h00000000} /* (3, 12, 8) {real, imag} */,
  {32'h43326398, 32'h00000000} /* (3, 12, 7) {real, imag} */,
  {32'h44665faf, 32'h00000000} /* (3, 12, 6) {real, imag} */,
  {32'h4468529a, 32'h00000000} /* (3, 12, 5) {real, imag} */,
  {32'hc3979ae2, 32'h00000000} /* (3, 12, 4) {real, imag} */,
  {32'hc38ba926, 32'h00000000} /* (3, 12, 3) {real, imag} */,
  {32'hc1f3ac40, 32'h00000000} /* (3, 12, 2) {real, imag} */,
  {32'hc34906ea, 32'h00000000} /* (3, 12, 1) {real, imag} */,
  {32'hc2ac268c, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'hc305958e, 32'h00000000} /* (3, 11, 15) {real, imag} */,
  {32'hc38c2930, 32'h00000000} /* (3, 11, 14) {real, imag} */,
  {32'h43fb87f4, 32'h00000000} /* (3, 11, 13) {real, imag} */,
  {32'hc30fc59c, 32'h00000000} /* (3, 11, 12) {real, imag} */,
  {32'h44278c1e, 32'h00000000} /* (3, 11, 11) {real, imag} */,
  {32'hc3a53e90, 32'h00000000} /* (3, 11, 10) {real, imag} */,
  {32'hc282d232, 32'h00000000} /* (3, 11, 9) {real, imag} */,
  {32'h43fa4248, 32'h00000000} /* (3, 11, 8) {real, imag} */,
  {32'hc43d6ba2, 32'h00000000} /* (3, 11, 7) {real, imag} */,
  {32'hc21f01ac, 32'h00000000} /* (3, 11, 6) {real, imag} */,
  {32'h44503f82, 32'h00000000} /* (3, 11, 5) {real, imag} */,
  {32'h4475fb61, 32'h00000000} /* (3, 11, 4) {real, imag} */,
  {32'h43d43760, 32'h00000000} /* (3, 11, 3) {real, imag} */,
  {32'hc325af80, 32'h00000000} /* (3, 11, 2) {real, imag} */,
  {32'hc3f84c1c, 32'h00000000} /* (3, 11, 1) {real, imag} */,
  {32'h43c26b0c, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'h43d32790, 32'h00000000} /* (3, 10, 15) {real, imag} */,
  {32'hc4817c8b, 32'h00000000} /* (3, 10, 14) {real, imag} */,
  {32'hc404e639, 32'h00000000} /* (3, 10, 13) {real, imag} */,
  {32'h44096b86, 32'h00000000} /* (3, 10, 12) {real, imag} */,
  {32'h4345a700, 32'h00000000} /* (3, 10, 11) {real, imag} */,
  {32'h43c22df8, 32'h00000000} /* (3, 10, 10) {real, imag} */,
  {32'h434cde06, 32'h00000000} /* (3, 10, 9) {real, imag} */,
  {32'hc42c3ee8, 32'h00000000} /* (3, 10, 8) {real, imag} */,
  {32'hc2292b6c, 32'h00000000} /* (3, 10, 7) {real, imag} */,
  {32'hc41d26d6, 32'h00000000} /* (3, 10, 6) {real, imag} */,
  {32'hc2ad7ef8, 32'h00000000} /* (3, 10, 5) {real, imag} */,
  {32'h445094ce, 32'h00000000} /* (3, 10, 4) {real, imag} */,
  {32'h422c0cba, 32'h00000000} /* (3, 10, 3) {real, imag} */,
  {32'hc34d3914, 32'h00000000} /* (3, 10, 2) {real, imag} */,
  {32'h431b9dba, 32'h00000000} /* (3, 10, 1) {real, imag} */,
  {32'h4380389e, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'h440e4ea1, 32'h00000000} /* (3, 9, 15) {real, imag} */,
  {32'h43c51c43, 32'h00000000} /* (3, 9, 14) {real, imag} */,
  {32'hc38b789a, 32'h00000000} /* (3, 9, 13) {real, imag} */,
  {32'hc317fced, 32'h00000000} /* (3, 9, 12) {real, imag} */,
  {32'hc3ec1209, 32'h00000000} /* (3, 9, 11) {real, imag} */,
  {32'hc35542be, 32'h00000000} /* (3, 9, 10) {real, imag} */,
  {32'hc2a67bd8, 32'h00000000} /* (3, 9, 9) {real, imag} */,
  {32'hc3a509e0, 32'h00000000} /* (3, 9, 8) {real, imag} */,
  {32'h43916076, 32'h00000000} /* (3, 9, 7) {real, imag} */,
  {32'h43740d36, 32'h00000000} /* (3, 9, 6) {real, imag} */,
  {32'hc31b07ca, 32'h00000000} /* (3, 9, 5) {real, imag} */,
  {32'h43fff368, 32'h00000000} /* (3, 9, 4) {real, imag} */,
  {32'hc3706156, 32'h00000000} /* (3, 9, 3) {real, imag} */,
  {32'hc42adf1a, 32'h00000000} /* (3, 9, 2) {real, imag} */,
  {32'h43c62bc1, 32'h00000000} /* (3, 9, 1) {real, imag} */,
  {32'h43be2dfa, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'h43b01464, 32'h00000000} /* (3, 8, 15) {real, imag} */,
  {32'h44375424, 32'h00000000} /* (3, 8, 14) {real, imag} */,
  {32'hc1fa63f8, 32'h00000000} /* (3, 8, 13) {real, imag} */,
  {32'hc3bfc208, 32'h00000000} /* (3, 8, 12) {real, imag} */,
  {32'hc28d3dd4, 32'h00000000} /* (3, 8, 11) {real, imag} */,
  {32'hc38d06de, 32'h00000000} /* (3, 8, 10) {real, imag} */,
  {32'h439c4c66, 32'h00000000} /* (3, 8, 9) {real, imag} */,
  {32'h441a4dec, 32'h00000000} /* (3, 8, 8) {real, imag} */,
  {32'hc3a2cf00, 32'h00000000} /* (3, 8, 7) {real, imag} */,
  {32'h44a9e284, 32'h00000000} /* (3, 8, 6) {real, imag} */,
  {32'h43e2ca94, 32'h00000000} /* (3, 8, 5) {real, imag} */,
  {32'hc2bd5c90, 32'h00000000} /* (3, 8, 4) {real, imag} */,
  {32'hc3ea27cb, 32'h00000000} /* (3, 8, 3) {real, imag} */,
  {32'hc4c9c62a, 32'h00000000} /* (3, 8, 2) {real, imag} */,
  {32'hc3dea4ea, 32'h00000000} /* (3, 8, 1) {real, imag} */,
  {32'h434124ea, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'h43055690, 32'h00000000} /* (3, 7, 15) {real, imag} */,
  {32'hc1ac5590, 32'h00000000} /* (3, 7, 14) {real, imag} */,
  {32'h42b5cc48, 32'h00000000} /* (3, 7, 13) {real, imag} */,
  {32'hc42f336e, 32'h00000000} /* (3, 7, 12) {real, imag} */,
  {32'hc43210fa, 32'h00000000} /* (3, 7, 11) {real, imag} */,
  {32'h43a5b057, 32'h00000000} /* (3, 7, 10) {real, imag} */,
  {32'h44651d6c, 32'h00000000} /* (3, 7, 9) {real, imag} */,
  {32'h42b0bf90, 32'h00000000} /* (3, 7, 8) {real, imag} */,
  {32'hc3effce4, 32'h00000000} /* (3, 7, 7) {real, imag} */,
  {32'hc385f455, 32'h00000000} /* (3, 7, 6) {real, imag} */,
  {32'hc41e6b7f, 32'h00000000} /* (3, 7, 5) {real, imag} */,
  {32'hc449f8ee, 32'h00000000} /* (3, 7, 4) {real, imag} */,
  {32'hc4356d1e, 32'h00000000} /* (3, 7, 3) {real, imag} */,
  {32'hc4778a78, 32'h00000000} /* (3, 7, 2) {real, imag} */,
  {32'hc4759c14, 32'h00000000} /* (3, 7, 1) {real, imag} */,
  {32'hc409b4ae, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'h417bd670, 32'h00000000} /* (3, 6, 15) {real, imag} */,
  {32'hc4a6d528, 32'h00000000} /* (3, 6, 14) {real, imag} */,
  {32'hc4613be4, 32'h00000000} /* (3, 6, 13) {real, imag} */,
  {32'hc30596a8, 32'h00000000} /* (3, 6, 12) {real, imag} */,
  {32'hc3d8932e, 32'h00000000} /* (3, 6, 11) {real, imag} */,
  {32'h429ab5c8, 32'h00000000} /* (3, 6, 10) {real, imag} */,
  {32'hc394ac63, 32'h00000000} /* (3, 6, 9) {real, imag} */,
  {32'hc3d5dfbb, 32'h00000000} /* (3, 6, 8) {real, imag} */,
  {32'hc37bd7f1, 32'h00000000} /* (3, 6, 7) {real, imag} */,
  {32'hc2a76ac8, 32'h00000000} /* (3, 6, 6) {real, imag} */,
  {32'hc4074ab4, 32'h00000000} /* (3, 6, 5) {real, imag} */,
  {32'hc4a759d1, 32'h00000000} /* (3, 6, 4) {real, imag} */,
  {32'hc3bf203e, 32'h00000000} /* (3, 6, 3) {real, imag} */,
  {32'hc4b127ea, 32'h00000000} /* (3, 6, 2) {real, imag} */,
  {32'hc3eb6387, 32'h00000000} /* (3, 6, 1) {real, imag} */,
  {32'hc4133a6c, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hc437a206, 32'h00000000} /* (3, 5, 15) {real, imag} */,
  {32'hc448965a, 32'h00000000} /* (3, 5, 14) {real, imag} */,
  {32'hc407c083, 32'h00000000} /* (3, 5, 13) {real, imag} */,
  {32'hc3e2256a, 32'h00000000} /* (3, 5, 12) {real, imag} */,
  {32'hc4407f8c, 32'h00000000} /* (3, 5, 11) {real, imag} */,
  {32'hc1c8fcc0, 32'h00000000} /* (3, 5, 10) {real, imag} */,
  {32'h442cd414, 32'h00000000} /* (3, 5, 9) {real, imag} */,
  {32'hc39577ae, 32'h00000000} /* (3, 5, 8) {real, imag} */,
  {32'h43bdc1c4, 32'h00000000} /* (3, 5, 7) {real, imag} */,
  {32'h439395f8, 32'h00000000} /* (3, 5, 6) {real, imag} */,
  {32'hc492a094, 32'h00000000} /* (3, 5, 5) {real, imag} */,
  {32'hc42fbd4f, 32'h00000000} /* (3, 5, 4) {real, imag} */,
  {32'hc4779bb0, 32'h00000000} /* (3, 5, 3) {real, imag} */,
  {32'hc4a74335, 32'h00000000} /* (3, 5, 2) {real, imag} */,
  {32'h4223b480, 32'h00000000} /* (3, 5, 1) {real, imag} */,
  {32'hc3184399, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hc489c451, 32'h00000000} /* (3, 4, 15) {real, imag} */,
  {32'hc45f6225, 32'h00000000} /* (3, 4, 14) {real, imag} */,
  {32'hc3e66ec4, 32'h00000000} /* (3, 4, 13) {real, imag} */,
  {32'hc329827c, 32'h00000000} /* (3, 4, 12) {real, imag} */,
  {32'h4383bdf8, 32'h00000000} /* (3, 4, 11) {real, imag} */,
  {32'h442d1c86, 32'h00000000} /* (3, 4, 10) {real, imag} */,
  {32'hc4762838, 32'h00000000} /* (3, 4, 9) {real, imag} */,
  {32'h43d751d4, 32'h00000000} /* (3, 4, 8) {real, imag} */,
  {32'hc3e81bf0, 32'h00000000} /* (3, 4, 7) {real, imag} */,
  {32'hc4aba862, 32'h00000000} /* (3, 4, 6) {real, imag} */,
  {32'hc40b4a8c, 32'h00000000} /* (3, 4, 5) {real, imag} */,
  {32'hc478317d, 32'h00000000} /* (3, 4, 4) {real, imag} */,
  {32'hc465f53a, 32'h00000000} /* (3, 4, 3) {real, imag} */,
  {32'hc493ff54, 32'h00000000} /* (3, 4, 2) {real, imag} */,
  {32'hc4a8a458, 32'h00000000} /* (3, 4, 1) {real, imag} */,
  {32'hc415effa, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hc40d1a2a, 32'h00000000} /* (3, 3, 15) {real, imag} */,
  {32'hc48b728f, 32'h00000000} /* (3, 3, 14) {real, imag} */,
  {32'hc48e4ec0, 32'h00000000} /* (3, 3, 13) {real, imag} */,
  {32'hc2a59940, 32'h00000000} /* (3, 3, 12) {real, imag} */,
  {32'h4409e52e, 32'h00000000} /* (3, 3, 11) {real, imag} */,
  {32'hc419416d, 32'h00000000} /* (3, 3, 10) {real, imag} */,
  {32'hc363a849, 32'h00000000} /* (3, 3, 9) {real, imag} */,
  {32'hc23c4c00, 32'h00000000} /* (3, 3, 8) {real, imag} */,
  {32'hc3939335, 32'h00000000} /* (3, 3, 7) {real, imag} */,
  {32'hc496e08b, 32'h00000000} /* (3, 3, 6) {real, imag} */,
  {32'hc3bf864f, 32'h00000000} /* (3, 3, 5) {real, imag} */,
  {32'hc4593d78, 32'h00000000} /* (3, 3, 4) {real, imag} */,
  {32'hc4885aa3, 32'h00000000} /* (3, 3, 3) {real, imag} */,
  {32'hc422cf3b, 32'h00000000} /* (3, 3, 2) {real, imag} */,
  {32'hc35135cb, 32'h00000000} /* (3, 3, 1) {real, imag} */,
  {32'hc47f0e6c, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hc4898b10, 32'h00000000} /* (3, 2, 15) {real, imag} */,
  {32'hc43cb98c, 32'h00000000} /* (3, 2, 14) {real, imag} */,
  {32'hc280e7c0, 32'h00000000} /* (3, 2, 13) {real, imag} */,
  {32'h4288c7c8, 32'h00000000} /* (3, 2, 12) {real, imag} */,
  {32'h42e5a2a0, 32'h00000000} /* (3, 2, 11) {real, imag} */,
  {32'h42f97688, 32'h00000000} /* (3, 2, 10) {real, imag} */,
  {32'h4272f930, 32'h00000000} /* (3, 2, 9) {real, imag} */,
  {32'hc3baecd8, 32'h00000000} /* (3, 2, 8) {real, imag} */,
  {32'hc3c93722, 32'h00000000} /* (3, 2, 7) {real, imag} */,
  {32'hc28e5ebc, 32'h00000000} /* (3, 2, 6) {real, imag} */,
  {32'hc47e3d32, 32'h00000000} /* (3, 2, 5) {real, imag} */,
  {32'hc4c2efc2, 32'h00000000} /* (3, 2, 4) {real, imag} */,
  {32'hc4c305aa, 32'h00000000} /* (3, 2, 3) {real, imag} */,
  {32'hc48573dc, 32'h00000000} /* (3, 2, 2) {real, imag} */,
  {32'hc48724c0, 32'h00000000} /* (3, 2, 1) {real, imag} */,
  {32'hc3fd482c, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hc433129d, 32'h00000000} /* (3, 1, 15) {real, imag} */,
  {32'hc43f568a, 32'h00000000} /* (3, 1, 14) {real, imag} */,
  {32'h440b7e86, 32'h00000000} /* (3, 1, 13) {real, imag} */,
  {32'h443c7f95, 32'h00000000} /* (3, 1, 12) {real, imag} */,
  {32'h43bd4287, 32'h00000000} /* (3, 1, 11) {real, imag} */,
  {32'hc3ace80d, 32'h00000000} /* (3, 1, 10) {real, imag} */,
  {32'hc44ccd13, 32'h00000000} /* (3, 1, 9) {real, imag} */,
  {32'hc2e3692c, 32'h00000000} /* (3, 1, 8) {real, imag} */,
  {32'hc41002fb, 32'h00000000} /* (3, 1, 7) {real, imag} */,
  {32'h428a77a4, 32'h00000000} /* (3, 1, 6) {real, imag} */,
  {32'hc3ca70e8, 32'h00000000} /* (3, 1, 5) {real, imag} */,
  {32'hc4b48c68, 32'h00000000} /* (3, 1, 4) {real, imag} */,
  {32'hc344d812, 32'h00000000} /* (3, 1, 3) {real, imag} */,
  {32'h43c39797, 32'h00000000} /* (3, 1, 2) {real, imag} */,
  {32'hc4a5870e, 32'h00000000} /* (3, 1, 1) {real, imag} */,
  {32'hc4029304, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'hc47e1e34, 32'h00000000} /* (3, 0, 15) {real, imag} */,
  {32'h411a1b40, 32'h00000000} /* (3, 0, 14) {real, imag} */,
  {32'h449bb1f8, 32'h00000000} /* (3, 0, 13) {real, imag} */,
  {32'h43c6d8e8, 32'h00000000} /* (3, 0, 12) {real, imag} */,
  {32'hc2d7b458, 32'h00000000} /* (3, 0, 11) {real, imag} */,
  {32'hc23415cc, 32'h00000000} /* (3, 0, 10) {real, imag} */,
  {32'hc3d6466b, 32'h00000000} /* (3, 0, 9) {real, imag} */,
  {32'hc2f2880d, 32'h00000000} /* (3, 0, 8) {real, imag} */,
  {32'hc469e4a4, 32'h00000000} /* (3, 0, 7) {real, imag} */,
  {32'hc3c4814e, 32'h00000000} /* (3, 0, 6) {real, imag} */,
  {32'h43063ee4, 32'h00000000} /* (3, 0, 5) {real, imag} */,
  {32'h441f5a24, 32'h00000000} /* (3, 0, 4) {real, imag} */,
  {32'hc457bead, 32'h00000000} /* (3, 0, 3) {real, imag} */,
  {32'hc34cc055, 32'h00000000} /* (3, 0, 2) {real, imag} */,
  {32'h43730852, 32'h00000000} /* (3, 0, 1) {real, imag} */,
  {32'hc3ba3815, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc405ac32, 32'h00000000} /* (2, 15, 15) {real, imag} */,
  {32'hc35490f2, 32'h00000000} /* (2, 15, 14) {real, imag} */,
  {32'h4205e000, 32'h00000000} /* (2, 15, 13) {real, imag} */,
  {32'hc32395f8, 32'h00000000} /* (2, 15, 12) {real, imag} */,
  {32'h43828c31, 32'h00000000} /* (2, 15, 11) {real, imag} */,
  {32'h43926a43, 32'h00000000} /* (2, 15, 10) {real, imag} */,
  {32'h4351c5d9, 32'h00000000} /* (2, 15, 9) {real, imag} */,
  {32'h432a104a, 32'h00000000} /* (2, 15, 8) {real, imag} */,
  {32'h44438d4e, 32'h00000000} /* (2, 15, 7) {real, imag} */,
  {32'hc319189a, 32'h00000000} /* (2, 15, 6) {real, imag} */,
  {32'hc40e05b6, 32'h00000000} /* (2, 15, 5) {real, imag} */,
  {32'hc3a9946e, 32'h00000000} /* (2, 15, 4) {real, imag} */,
  {32'hc49fd2ae, 32'h00000000} /* (2, 15, 3) {real, imag} */,
  {32'hc4602e10, 32'h00000000} /* (2, 15, 2) {real, imag} */,
  {32'hc3bf6c34, 32'h00000000} /* (2, 15, 1) {real, imag} */,
  {32'hc4570200, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'h4307e639, 32'h00000000} /* (2, 14, 15) {real, imag} */,
  {32'h437d088b, 32'h00000000} /* (2, 14, 14) {real, imag} */,
  {32'hc404d696, 32'h00000000} /* (2, 14, 13) {real, imag} */,
  {32'hc35d944b, 32'h00000000} /* (2, 14, 12) {real, imag} */,
  {32'hc389066a, 32'h00000000} /* (2, 14, 11) {real, imag} */,
  {32'hc22d9bb8, 32'h00000000} /* (2, 14, 10) {real, imag} */,
  {32'hc3d5b9a5, 32'h00000000} /* (2, 14, 9) {real, imag} */,
  {32'h43c5b0a8, 32'h00000000} /* (2, 14, 8) {real, imag} */,
  {32'h43848248, 32'h00000000} /* (2, 14, 7) {real, imag} */,
  {32'hc2f8868a, 32'h00000000} /* (2, 14, 6) {real, imag} */,
  {32'hc27cbde4, 32'h00000000} /* (2, 14, 5) {real, imag} */,
  {32'hc43463cb, 32'h00000000} /* (2, 14, 4) {real, imag} */,
  {32'hc3aa4eb2, 32'h00000000} /* (2, 14, 3) {real, imag} */,
  {32'hc42a676a, 32'h00000000} /* (2, 14, 2) {real, imag} */,
  {32'hc41cf4ce, 32'h00000000} /* (2, 14, 1) {real, imag} */,
  {32'hc1f9fd38, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h4401b0bb, 32'h00000000} /* (2, 13, 15) {real, imag} */,
  {32'hc44be8da, 32'h00000000} /* (2, 13, 14) {real, imag} */,
  {32'hc3d5720f, 32'h00000000} /* (2, 13, 13) {real, imag} */,
  {32'h41a35b40, 32'h00000000} /* (2, 13, 12) {real, imag} */,
  {32'hc2aee6b4, 32'h00000000} /* (2, 13, 11) {real, imag} */,
  {32'hc418e3b8, 32'h00000000} /* (2, 13, 10) {real, imag} */,
  {32'hc4ac3570, 32'h00000000} /* (2, 13, 9) {real, imag} */,
  {32'h42fa5760, 32'h00000000} /* (2, 13, 8) {real, imag} */,
  {32'h43cad089, 32'h00000000} /* (2, 13, 7) {real, imag} */,
  {32'hc1eebb20, 32'h00000000} /* (2, 13, 6) {real, imag} */,
  {32'h42f44fa4, 32'h00000000} /* (2, 13, 5) {real, imag} */,
  {32'hc2011320, 32'h00000000} /* (2, 13, 4) {real, imag} */,
  {32'hc3de3f43, 32'h00000000} /* (2, 13, 3) {real, imag} */,
  {32'hc4808496, 32'h00000000} /* (2, 13, 2) {real, imag} */,
  {32'hc324c75c, 32'h00000000} /* (2, 13, 1) {real, imag} */,
  {32'h4432a422, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'h434ae802, 32'h00000000} /* (2, 12, 15) {real, imag} */,
  {32'hc34542a4, 32'h00000000} /* (2, 12, 14) {real, imag} */,
  {32'h4394a3be, 32'h00000000} /* (2, 12, 13) {real, imag} */,
  {32'h43a55c4e, 32'h00000000} /* (2, 12, 12) {real, imag} */,
  {32'hc40905ab, 32'h00000000} /* (2, 12, 11) {real, imag} */,
  {32'hc3744936, 32'h00000000} /* (2, 12, 10) {real, imag} */,
  {32'h4254971c, 32'h00000000} /* (2, 12, 9) {real, imag} */,
  {32'h42abd224, 32'h00000000} /* (2, 12, 8) {real, imag} */,
  {32'h4400a176, 32'h00000000} /* (2, 12, 7) {real, imag} */,
  {32'h43dc23b8, 32'h00000000} /* (2, 12, 6) {real, imag} */,
  {32'h4489fc5c, 32'h00000000} /* (2, 12, 5) {real, imag} */,
  {32'h43da4a64, 32'h00000000} /* (2, 12, 4) {real, imag} */,
  {32'hc41d8725, 32'h00000000} /* (2, 12, 3) {real, imag} */,
  {32'hc426cb7c, 32'h00000000} /* (2, 12, 2) {real, imag} */,
  {32'h437f3c61, 32'h00000000} /* (2, 12, 1) {real, imag} */,
  {32'hbfaf6700, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h4369c2b6, 32'h00000000} /* (2, 11, 15) {real, imag} */,
  {32'h44138f5c, 32'h00000000} /* (2, 11, 14) {real, imag} */,
  {32'h44b7e7ac, 32'h00000000} /* (2, 11, 13) {real, imag} */,
  {32'h43fb2529, 32'h00000000} /* (2, 11, 12) {real, imag} */,
  {32'h439db5e1, 32'h00000000} /* (2, 11, 11) {real, imag} */,
  {32'hc41591f4, 32'h00000000} /* (2, 11, 10) {real, imag} */,
  {32'hc3456c48, 32'h00000000} /* (2, 11, 9) {real, imag} */,
  {32'h43df6f7c, 32'h00000000} /* (2, 11, 8) {real, imag} */,
  {32'hc409f6d4, 32'h00000000} /* (2, 11, 7) {real, imag} */,
  {32'hc45e970c, 32'h00000000} /* (2, 11, 6) {real, imag} */,
  {32'h43bab76a, 32'h00000000} /* (2, 11, 5) {real, imag} */,
  {32'h4253cf88, 32'h00000000} /* (2, 11, 4) {real, imag} */,
  {32'hc27f2318, 32'h00000000} /* (2, 11, 3) {real, imag} */,
  {32'h42189830, 32'h00000000} /* (2, 11, 2) {real, imag} */,
  {32'hc2f5fc90, 32'h00000000} /* (2, 11, 1) {real, imag} */,
  {32'h43d3f60a, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'h44573a1f, 32'h00000000} /* (2, 10, 15) {real, imag} */,
  {32'h44351d59, 32'h00000000} /* (2, 10, 14) {real, imag} */,
  {32'hc361dce0, 32'h00000000} /* (2, 10, 13) {real, imag} */,
  {32'h439b13b0, 32'h00000000} /* (2, 10, 12) {real, imag} */,
  {32'h4427b892, 32'h00000000} /* (2, 10, 11) {real, imag} */,
  {32'h433af184, 32'h00000000} /* (2, 10, 10) {real, imag} */,
  {32'hc42ac354, 32'h00000000} /* (2, 10, 9) {real, imag} */,
  {32'hc4799aa2, 32'h00000000} /* (2, 10, 8) {real, imag} */,
  {32'hc44bbc29, 32'h00000000} /* (2, 10, 7) {real, imag} */,
  {32'h44414793, 32'h00000000} /* (2, 10, 6) {real, imag} */,
  {32'h41c382fc, 32'h00000000} /* (2, 10, 5) {real, imag} */,
  {32'h41d67fe0, 32'h00000000} /* (2, 10, 4) {real, imag} */,
  {32'hc48273fa, 32'h00000000} /* (2, 10, 3) {real, imag} */,
  {32'h41f23a84, 32'h00000000} /* (2, 10, 2) {real, imag} */,
  {32'h430ccc36, 32'h00000000} /* (2, 10, 1) {real, imag} */,
  {32'h441198be, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'h441c2ba5, 32'h00000000} /* (2, 9, 15) {real, imag} */,
  {32'h448250c2, 32'h00000000} /* (2, 9, 14) {real, imag} */,
  {32'h4482e584, 32'h00000000} /* (2, 9, 13) {real, imag} */,
  {32'h439ace55, 32'h00000000} /* (2, 9, 12) {real, imag} */,
  {32'h43cf3498, 32'h00000000} /* (2, 9, 11) {real, imag} */,
  {32'h443f6be2, 32'h00000000} /* (2, 9, 10) {real, imag} */,
  {32'h43d616c2, 32'h00000000} /* (2, 9, 9) {real, imag} */,
  {32'hc26756e0, 32'h00000000} /* (2, 9, 8) {real, imag} */,
  {32'h4422d4ef, 32'h00000000} /* (2, 9, 7) {real, imag} */,
  {32'h42cb691c, 32'h00000000} /* (2, 9, 6) {real, imag} */,
  {32'h446f1bcf, 32'h00000000} /* (2, 9, 5) {real, imag} */,
  {32'h4409346c, 32'h00000000} /* (2, 9, 4) {real, imag} */,
  {32'h446850e4, 32'h00000000} /* (2, 9, 3) {real, imag} */,
  {32'hc31c05ca, 32'h00000000} /* (2, 9, 2) {real, imag} */,
  {32'h4422fccd, 32'h00000000} /* (2, 9, 1) {real, imag} */,
  {32'h43b1812e, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'h447fb5ed, 32'h00000000} /* (2, 8, 15) {real, imag} */,
  {32'h4507c4d4, 32'h00000000} /* (2, 8, 14) {real, imag} */,
  {32'h442a927e, 32'h00000000} /* (2, 8, 13) {real, imag} */,
  {32'h422c0408, 32'h00000000} /* (2, 8, 12) {real, imag} */,
  {32'h4406136b, 32'h00000000} /* (2, 8, 11) {real, imag} */,
  {32'h4392cf08, 32'h00000000} /* (2, 8, 10) {real, imag} */,
  {32'h441cbebf, 32'h00000000} /* (2, 8, 9) {real, imag} */,
  {32'h423230d4, 32'h00000000} /* (2, 8, 8) {real, imag} */,
  {32'h44666953, 32'h00000000} /* (2, 8, 7) {real, imag} */,
  {32'hc135a180, 32'h00000000} /* (2, 8, 6) {real, imag} */,
  {32'hc34ee206, 32'h00000000} /* (2, 8, 5) {real, imag} */,
  {32'h440826d2, 32'h00000000} /* (2, 8, 4) {real, imag} */,
  {32'h43f13c2b, 32'h00000000} /* (2, 8, 3) {real, imag} */,
  {32'hc3ac12b8, 32'h00000000} /* (2, 8, 2) {real, imag} */,
  {32'hc419ab1d, 32'h00000000} /* (2, 8, 1) {real, imag} */,
  {32'h436fdd7f, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'h43cec92c, 32'h00000000} /* (2, 7, 15) {real, imag} */,
  {32'h43ee1f6e, 32'h00000000} /* (2, 7, 14) {real, imag} */,
  {32'h449b3e55, 32'h00000000} /* (2, 7, 13) {real, imag} */,
  {32'hc2e9cd6a, 32'h00000000} /* (2, 7, 12) {real, imag} */,
  {32'h446a9612, 32'h00000000} /* (2, 7, 11) {real, imag} */,
  {32'hc429441b, 32'h00000000} /* (2, 7, 10) {real, imag} */,
  {32'hc3471dce, 32'h00000000} /* (2, 7, 9) {real, imag} */,
  {32'h4435339e, 32'h00000000} /* (2, 7, 8) {real, imag} */,
  {32'h4299c4e6, 32'h00000000} /* (2, 7, 7) {real, imag} */,
  {32'hc44633a3, 32'h00000000} /* (2, 7, 6) {real, imag} */,
  {32'hc46050e2, 32'h00000000} /* (2, 7, 5) {real, imag} */,
  {32'hc31feea3, 32'h00000000} /* (2, 7, 4) {real, imag} */,
  {32'hc3cc4610, 32'h00000000} /* (2, 7, 3) {real, imag} */,
  {32'hc458440d, 32'h00000000} /* (2, 7, 2) {real, imag} */,
  {32'hc3cc2241, 32'h00000000} /* (2, 7, 1) {real, imag} */,
  {32'h447477e4, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'h43c8facc, 32'h00000000} /* (2, 6, 15) {real, imag} */,
  {32'hc3e2dada, 32'h00000000} /* (2, 6, 14) {real, imag} */,
  {32'h4320d64e, 32'h00000000} /* (2, 6, 13) {real, imag} */,
  {32'h44af15fc, 32'h00000000} /* (2, 6, 12) {real, imag} */,
  {32'hc3a6c078, 32'h00000000} /* (2, 6, 11) {real, imag} */,
  {32'hc3d0ee71, 32'h00000000} /* (2, 6, 10) {real, imag} */,
  {32'hc20e9066, 32'h00000000} /* (2, 6, 9) {real, imag} */,
  {32'hc34f9eb8, 32'h00000000} /* (2, 6, 8) {real, imag} */,
  {32'hc3c0e078, 32'h00000000} /* (2, 6, 7) {real, imag} */,
  {32'hc354a15c, 32'h00000000} /* (2, 6, 6) {real, imag} */,
  {32'hc4346ecc, 32'h00000000} /* (2, 6, 5) {real, imag} */,
  {32'hc436d249, 32'h00000000} /* (2, 6, 4) {real, imag} */,
  {32'hc4174860, 32'h00000000} /* (2, 6, 3) {real, imag} */,
  {32'hc4891352, 32'h00000000} /* (2, 6, 2) {real, imag} */,
  {32'hc2f259b7, 32'h00000000} /* (2, 6, 1) {real, imag} */,
  {32'h434eb0c0, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hc4070373, 32'h00000000} /* (2, 5, 15) {real, imag} */,
  {32'hc4516282, 32'h00000000} /* (2, 5, 14) {real, imag} */,
  {32'hc3682cd8, 32'h00000000} /* (2, 5, 13) {real, imag} */,
  {32'h432098e8, 32'h00000000} /* (2, 5, 12) {real, imag} */,
  {32'hc2d379d8, 32'h00000000} /* (2, 5, 11) {real, imag} */,
  {32'h43235a32, 32'h00000000} /* (2, 5, 10) {real, imag} */,
  {32'hc29324c4, 32'h00000000} /* (2, 5, 9) {real, imag} */,
  {32'h42a7173c, 32'h00000000} /* (2, 5, 8) {real, imag} */,
  {32'hc374a98d, 32'h00000000} /* (2, 5, 7) {real, imag} */,
  {32'hc498bd1f, 32'h00000000} /* (2, 5, 6) {real, imag} */,
  {32'hc4b34817, 32'h00000000} /* (2, 5, 5) {real, imag} */,
  {32'hc402f830, 32'h00000000} /* (2, 5, 4) {real, imag} */,
  {32'hc4b79a8c, 32'h00000000} /* (2, 5, 3) {real, imag} */,
  {32'hc43ff3da, 32'h00000000} /* (2, 5, 2) {real, imag} */,
  {32'h444cb162, 32'h00000000} /* (2, 5, 1) {real, imag} */,
  {32'hc34a193e, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hc400c1d6, 32'h00000000} /* (2, 4, 15) {real, imag} */,
  {32'hc426f938, 32'h00000000} /* (2, 4, 14) {real, imag} */,
  {32'hc00f7200, 32'h00000000} /* (2, 4, 13) {real, imag} */,
  {32'hc3cc0116, 32'h00000000} /* (2, 4, 12) {real, imag} */,
  {32'h43b8099b, 32'h00000000} /* (2, 4, 11) {real, imag} */,
  {32'h4406879e, 32'h00000000} /* (2, 4, 10) {real, imag} */,
  {32'h42e42058, 32'h00000000} /* (2, 4, 9) {real, imag} */,
  {32'h43e7907c, 32'h00000000} /* (2, 4, 8) {real, imag} */,
  {32'hc3d1778a, 32'h00000000} /* (2, 4, 7) {real, imag} */,
  {32'hc455058c, 32'h00000000} /* (2, 4, 6) {real, imag} */,
  {32'hc46a21dc, 32'h00000000} /* (2, 4, 5) {real, imag} */,
  {32'hc4b54f42, 32'h00000000} /* (2, 4, 4) {real, imag} */,
  {32'hc3d4fd0b, 32'h00000000} /* (2, 4, 3) {real, imag} */,
  {32'hc455a010, 32'h00000000} /* (2, 4, 2) {real, imag} */,
  {32'h43b35719, 32'h00000000} /* (2, 4, 1) {real, imag} */,
  {32'hc3e7bba0, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hc481f844, 32'h00000000} /* (2, 3, 15) {real, imag} */,
  {32'hc4827de8, 32'h00000000} /* (2, 3, 14) {real, imag} */,
  {32'h442ae45d, 32'h00000000} /* (2, 3, 13) {real, imag} */,
  {32'h42c683ac, 32'h00000000} /* (2, 3, 12) {real, imag} */,
  {32'h439229ef, 32'h00000000} /* (2, 3, 11) {real, imag} */,
  {32'h446643b5, 32'h00000000} /* (2, 3, 10) {real, imag} */,
  {32'hc35a0697, 32'h00000000} /* (2, 3, 9) {real, imag} */,
  {32'hc2ba77e0, 32'h00000000} /* (2, 3, 8) {real, imag} */,
  {32'hc4637e60, 32'h00000000} /* (2, 3, 7) {real, imag} */,
  {32'hc460caa6, 32'h00000000} /* (2, 3, 6) {real, imag} */,
  {32'hc4599fdf, 32'h00000000} /* (2, 3, 5) {real, imag} */,
  {32'hc3fbb155, 32'h00000000} /* (2, 3, 4) {real, imag} */,
  {32'hc3eaec91, 32'h00000000} /* (2, 3, 3) {real, imag} */,
  {32'hbfc77600, 32'h00000000} /* (2, 3, 2) {real, imag} */,
  {32'hc3874e1c, 32'h00000000} /* (2, 3, 1) {real, imag} */,
  {32'hc24cfe70, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hc3e3d816, 32'h00000000} /* (2, 2, 15) {real, imag} */,
  {32'h42f5d0f2, 32'h00000000} /* (2, 2, 14) {real, imag} */,
  {32'hc30f0d86, 32'h00000000} /* (2, 2, 13) {real, imag} */,
  {32'h442da4be, 32'h00000000} /* (2, 2, 12) {real, imag} */,
  {32'h441d66af, 32'h00000000} /* (2, 2, 11) {real, imag} */,
  {32'hc2f5bb58, 32'h00000000} /* (2, 2, 10) {real, imag} */,
  {32'hc42527bb, 32'h00000000} /* (2, 2, 9) {real, imag} */,
  {32'h4175e2d0, 32'h00000000} /* (2, 2, 8) {real, imag} */,
  {32'h437a175c, 32'h00000000} /* (2, 2, 7) {real, imag} */,
  {32'hc35122b5, 32'h00000000} /* (2, 2, 6) {real, imag} */,
  {32'hc447d29a, 32'h00000000} /* (2, 2, 5) {real, imag} */,
  {32'hc4806f83, 32'h00000000} /* (2, 2, 4) {real, imag} */,
  {32'hc3d2068a, 32'h00000000} /* (2, 2, 3) {real, imag} */,
  {32'hc49eac6a, 32'h00000000} /* (2, 2, 2) {real, imag} */,
  {32'hc3f9e4f3, 32'h00000000} /* (2, 2, 1) {real, imag} */,
  {32'hc3ab3420, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hc45fcd2f, 32'h00000000} /* (2, 1, 15) {real, imag} */,
  {32'hc42ef71a, 32'h00000000} /* (2, 1, 14) {real, imag} */,
  {32'h41888c00, 32'h00000000} /* (2, 1, 13) {real, imag} */,
  {32'h430f1508, 32'h00000000} /* (2, 1, 12) {real, imag} */,
  {32'h4451cbe7, 32'h00000000} /* (2, 1, 11) {real, imag} */,
  {32'h431cf118, 32'h00000000} /* (2, 1, 10) {real, imag} */,
  {32'h43c290fe, 32'h00000000} /* (2, 1, 9) {real, imag} */,
  {32'hc4a2c45c, 32'h00000000} /* (2, 1, 8) {real, imag} */,
  {32'h439711aa, 32'h00000000} /* (2, 1, 7) {real, imag} */,
  {32'h44071542, 32'h00000000} /* (2, 1, 6) {real, imag} */,
  {32'hc43a48ce, 32'h00000000} /* (2, 1, 5) {real, imag} */,
  {32'hc4253d92, 32'h00000000} /* (2, 1, 4) {real, imag} */,
  {32'hc47b21e1, 32'h00000000} /* (2, 1, 3) {real, imag} */,
  {32'hc47eed7c, 32'h00000000} /* (2, 1, 2) {real, imag} */,
  {32'hc4279f35, 32'h00000000} /* (2, 1, 1) {real, imag} */,
  {32'hc3cc1162, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hc3e08c90, 32'h00000000} /* (2, 0, 15) {real, imag} */,
  {32'hc44a7581, 32'h00000000} /* (2, 0, 14) {real, imag} */,
  {32'hc2e0fdc0, 32'h00000000} /* (2, 0, 13) {real, imag} */,
  {32'h44886839, 32'h00000000} /* (2, 0, 12) {real, imag} */,
  {32'h43e12662, 32'h00000000} /* (2, 0, 11) {real, imag} */,
  {32'h420f0128, 32'h00000000} /* (2, 0, 10) {real, imag} */,
  {32'h4389ade2, 32'h00000000} /* (2, 0, 9) {real, imag} */,
  {32'hc3c5ce54, 32'h00000000} /* (2, 0, 8) {real, imag} */,
  {32'h4295b720, 32'h00000000} /* (2, 0, 7) {real, imag} */,
  {32'h438fa9fe, 32'h00000000} /* (2, 0, 6) {real, imag} */,
  {32'hc403cb9c, 32'h00000000} /* (2, 0, 5) {real, imag} */,
  {32'hc4078642, 32'h00000000} /* (2, 0, 4) {real, imag} */,
  {32'hc2647950, 32'h00000000} /* (2, 0, 3) {real, imag} */,
  {32'h4304857d, 32'h00000000} /* (2, 0, 2) {real, imag} */,
  {32'hc3a5f2d6, 32'h00000000} /* (2, 0, 1) {real, imag} */,
  {32'hc3dc2bda, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc2b2f811, 32'h00000000} /* (1, 15, 15) {real, imag} */,
  {32'hc383895a, 32'h00000000} /* (1, 15, 14) {real, imag} */,
  {32'h4137a0c0, 32'h00000000} /* (1, 15, 13) {real, imag} */,
  {32'hc28d84b0, 32'h00000000} /* (1, 15, 12) {real, imag} */,
  {32'h43adccbd, 32'h00000000} /* (1, 15, 11) {real, imag} */,
  {32'h4416ba97, 32'h00000000} /* (1, 15, 10) {real, imag} */,
  {32'hc3a20a02, 32'h00000000} /* (1, 15, 9) {real, imag} */,
  {32'h43363493, 32'h00000000} /* (1, 15, 8) {real, imag} */,
  {32'h430babe2, 32'h00000000} /* (1, 15, 7) {real, imag} */,
  {32'hc2e89a1b, 32'h00000000} /* (1, 15, 6) {real, imag} */,
  {32'hc42bf559, 32'h00000000} /* (1, 15, 5) {real, imag} */,
  {32'hc43d9eac, 32'h00000000} /* (1, 15, 4) {real, imag} */,
  {32'hc43a6516, 32'h00000000} /* (1, 15, 3) {real, imag} */,
  {32'hc422ce6d, 32'h00000000} /* (1, 15, 2) {real, imag} */,
  {32'hc407c5ad, 32'h00000000} /* (1, 15, 1) {real, imag} */,
  {32'hc3bdb81c, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'hc2879574, 32'h00000000} /* (1, 14, 15) {real, imag} */,
  {32'hc2e78048, 32'h00000000} /* (1, 14, 14) {real, imag} */,
  {32'h4258e6c0, 32'h00000000} /* (1, 14, 13) {real, imag} */,
  {32'hc24598d4, 32'h00000000} /* (1, 14, 12) {real, imag} */,
  {32'h44119060, 32'h00000000} /* (1, 14, 11) {real, imag} */,
  {32'h43607220, 32'h00000000} /* (1, 14, 10) {real, imag} */,
  {32'h430afe9c, 32'h00000000} /* (1, 14, 9) {real, imag} */,
  {32'hc28aa5f4, 32'h00000000} /* (1, 14, 8) {real, imag} */,
  {32'h436a8876, 32'h00000000} /* (1, 14, 7) {real, imag} */,
  {32'h44669123, 32'h00000000} /* (1, 14, 6) {real, imag} */,
  {32'hc3ec3398, 32'h00000000} /* (1, 14, 5) {real, imag} */,
  {32'h425ce2e8, 32'h00000000} /* (1, 14, 4) {real, imag} */,
  {32'hc489ec46, 32'h00000000} /* (1, 14, 3) {real, imag} */,
  {32'hc49190df, 32'h00000000} /* (1, 14, 2) {real, imag} */,
  {32'h4328bcb4, 32'h00000000} /* (1, 14, 1) {real, imag} */,
  {32'hc3a6cedd, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'h422c4ffa, 32'h00000000} /* (1, 13, 15) {real, imag} */,
  {32'h4286b8ee, 32'h00000000} /* (1, 13, 14) {real, imag} */,
  {32'hc40b2798, 32'h00000000} /* (1, 13, 13) {real, imag} */,
  {32'h43b58c00, 32'h00000000} /* (1, 13, 12) {real, imag} */,
  {32'h4402870a, 32'h00000000} /* (1, 13, 11) {real, imag} */,
  {32'hc30053c9, 32'h00000000} /* (1, 13, 10) {real, imag} */,
  {32'hc33a881b, 32'h00000000} /* (1, 13, 9) {real, imag} */,
  {32'h437ad91c, 32'h00000000} /* (1, 13, 8) {real, imag} */,
  {32'hc2d16fcb, 32'h00000000} /* (1, 13, 7) {real, imag} */,
  {32'h435d3351, 32'h00000000} /* (1, 13, 6) {real, imag} */,
  {32'h4342525a, 32'h00000000} /* (1, 13, 5) {real, imag} */,
  {32'hc3912390, 32'h00000000} /* (1, 13, 4) {real, imag} */,
  {32'h40fc8e40, 32'h00000000} /* (1, 13, 3) {real, imag} */,
  {32'hc40585b1, 32'h00000000} /* (1, 13, 2) {real, imag} */,
  {32'hc337fccd, 32'h00000000} /* (1, 13, 1) {real, imag} */,
  {32'h4454611f, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'hc1035c00, 32'h00000000} /* (1, 12, 15) {real, imag} */,
  {32'hc3a61f1d, 32'h00000000} /* (1, 12, 14) {real, imag} */,
  {32'h4414a488, 32'h00000000} /* (1, 12, 13) {real, imag} */,
  {32'h4417daeb, 32'h00000000} /* (1, 12, 12) {real, imag} */,
  {32'hc32c5aea, 32'h00000000} /* (1, 12, 11) {real, imag} */,
  {32'hc3432520, 32'h00000000} /* (1, 12, 10) {real, imag} */,
  {32'hc3f045f3, 32'h00000000} /* (1, 12, 9) {real, imag} */,
  {32'hc434fafc, 32'h00000000} /* (1, 12, 8) {real, imag} */,
  {32'hc4956d62, 32'h00000000} /* (1, 12, 7) {real, imag} */,
  {32'hc482c811, 32'h00000000} /* (1, 12, 6) {real, imag} */,
  {32'hc3ed7850, 32'h00000000} /* (1, 12, 5) {real, imag} */,
  {32'hc3894f52, 32'h00000000} /* (1, 12, 4) {real, imag} */,
  {32'h441f647e, 32'h00000000} /* (1, 12, 3) {real, imag} */,
  {32'h441170f1, 32'h00000000} /* (1, 12, 2) {real, imag} */,
  {32'h4408e8d1, 32'h00000000} /* (1, 12, 1) {real, imag} */,
  {32'h43dbf848, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'h4370f3b0, 32'h00000000} /* (1, 11, 15) {real, imag} */,
  {32'h442aef2e, 32'h00000000} /* (1, 11, 14) {real, imag} */,
  {32'h44ee0ada, 32'h00000000} /* (1, 11, 13) {real, imag} */,
  {32'h44b74e46, 32'h00000000} /* (1, 11, 12) {real, imag} */,
  {32'h425c08c8, 32'h00000000} /* (1, 11, 11) {real, imag} */,
  {32'h43dce173, 32'h00000000} /* (1, 11, 10) {real, imag} */,
  {32'h43b69c95, 32'h00000000} /* (1, 11, 9) {real, imag} */,
  {32'h408214a0, 32'h00000000} /* (1, 11, 8) {real, imag} */,
  {32'hc3c89384, 32'h00000000} /* (1, 11, 7) {real, imag} */,
  {32'h42f409ec, 32'h00000000} /* (1, 11, 6) {real, imag} */,
  {32'h43b01460, 32'h00000000} /* (1, 11, 5) {real, imag} */,
  {32'h43b08c44, 32'h00000000} /* (1, 11, 4) {real, imag} */,
  {32'hc401e464, 32'h00000000} /* (1, 11, 3) {real, imag} */,
  {32'hc44bc774, 32'h00000000} /* (1, 11, 2) {real, imag} */,
  {32'h441969aa, 32'h00000000} /* (1, 11, 1) {real, imag} */,
  {32'h43b4b7ea, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'h446216ce, 32'h00000000} /* (1, 10, 15) {real, imag} */,
  {32'h44c272ba, 32'h00000000} /* (1, 10, 14) {real, imag} */,
  {32'h44236818, 32'h00000000} /* (1, 10, 13) {real, imag} */,
  {32'h448d57cd, 32'h00000000} /* (1, 10, 12) {real, imag} */,
  {32'h44446ee7, 32'h00000000} /* (1, 10, 11) {real, imag} */,
  {32'h440e17e7, 32'h00000000} /* (1, 10, 10) {real, imag} */,
  {32'h4476a18e, 32'h00000000} /* (1, 10, 9) {real, imag} */,
  {32'h448b2f8e, 32'h00000000} /* (1, 10, 8) {real, imag} */,
  {32'hc35b4918, 32'h00000000} /* (1, 10, 7) {real, imag} */,
  {32'h43608874, 32'h00000000} /* (1, 10, 6) {real, imag} */,
  {32'hc3acf9f9, 32'h00000000} /* (1, 10, 5) {real, imag} */,
  {32'hc41fc546, 32'h00000000} /* (1, 10, 4) {real, imag} */,
  {32'h4360affc, 32'h00000000} /* (1, 10, 3) {real, imag} */,
  {32'hc37be8e4, 32'h00000000} /* (1, 10, 2) {real, imag} */,
  {32'hc363f13e, 32'h00000000} /* (1, 10, 1) {real, imag} */,
  {32'hc3008dce, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'h44845fa6, 32'h00000000} /* (1, 9, 15) {real, imag} */,
  {32'h43ce7308, 32'h00000000} /* (1, 9, 14) {real, imag} */,
  {32'h43711dcf, 32'h00000000} /* (1, 9, 13) {real, imag} */,
  {32'h4469ca46, 32'h00000000} /* (1, 9, 12) {real, imag} */,
  {32'h43de37e8, 32'h00000000} /* (1, 9, 11) {real, imag} */,
  {32'h448c1d9e, 32'h00000000} /* (1, 9, 10) {real, imag} */,
  {32'h43e2675f, 32'h00000000} /* (1, 9, 9) {real, imag} */,
  {32'hc348f3a4, 32'h00000000} /* (1, 9, 8) {real, imag} */,
  {32'h44205311, 32'h00000000} /* (1, 9, 7) {real, imag} */,
  {32'h3fa3c300, 32'h00000000} /* (1, 9, 6) {real, imag} */,
  {32'h43d45246, 32'h00000000} /* (1, 9, 5) {real, imag} */,
  {32'h43dc6915, 32'h00000000} /* (1, 9, 4) {real, imag} */,
  {32'h438ff3ac, 32'h00000000} /* (1, 9, 3) {real, imag} */,
  {32'h42bd8ab0, 32'h00000000} /* (1, 9, 2) {real, imag} */,
  {32'h44315bfa, 32'h00000000} /* (1, 9, 1) {real, imag} */,
  {32'h447be219, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'h44468fa2, 32'h00000000} /* (1, 8, 15) {real, imag} */,
  {32'h440e709c, 32'h00000000} /* (1, 8, 14) {real, imag} */,
  {32'h43463ba6, 32'h00000000} /* (1, 8, 13) {real, imag} */,
  {32'h440e6481, 32'h00000000} /* (1, 8, 12) {real, imag} */,
  {32'hc0fa5800, 32'h00000000} /* (1, 8, 11) {real, imag} */,
  {32'h4431757b, 32'h00000000} /* (1, 8, 10) {real, imag} */,
  {32'h438a0fda, 32'h00000000} /* (1, 8, 9) {real, imag} */,
  {32'hc3e5b932, 32'h00000000} /* (1, 8, 8) {real, imag} */,
  {32'h43590e6a, 32'h00000000} /* (1, 8, 7) {real, imag} */,
  {32'hc433f134, 32'h00000000} /* (1, 8, 6) {real, imag} */,
  {32'h439c5cf4, 32'h00000000} /* (1, 8, 5) {real, imag} */,
  {32'h445087c1, 32'h00000000} /* (1, 8, 4) {real, imag} */,
  {32'h440352b4, 32'h00000000} /* (1, 8, 3) {real, imag} */,
  {32'h43fe74da, 32'h00000000} /* (1, 8, 2) {real, imag} */,
  {32'h43511cc2, 32'h00000000} /* (1, 8, 1) {real, imag} */,
  {32'h44359147, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'hc2e1a646, 32'h00000000} /* (1, 7, 15) {real, imag} */,
  {32'h433752d8, 32'h00000000} /* (1, 7, 14) {real, imag} */,
  {32'h4379d0cc, 32'h00000000} /* (1, 7, 13) {real, imag} */,
  {32'h43d9865e, 32'h00000000} /* (1, 7, 12) {real, imag} */,
  {32'hc304fb73, 32'h00000000} /* (1, 7, 11) {real, imag} */,
  {32'hc1ef52b8, 32'h00000000} /* (1, 7, 10) {real, imag} */,
  {32'hc43f3a4d, 32'h00000000} /* (1, 7, 9) {real, imag} */,
  {32'hc333571c, 32'h00000000} /* (1, 7, 8) {real, imag} */,
  {32'h43ad7c1a, 32'h00000000} /* (1, 7, 7) {real, imag} */,
  {32'hc4cf21c3, 32'h00000000} /* (1, 7, 6) {real, imag} */,
  {32'hc4128ca5, 32'h00000000} /* (1, 7, 5) {real, imag} */,
  {32'hc367d888, 32'h00000000} /* (1, 7, 4) {real, imag} */,
  {32'h41946586, 32'h00000000} /* (1, 7, 3) {real, imag} */,
  {32'h4397895c, 32'h00000000} /* (1, 7, 2) {real, imag} */,
  {32'h4433ceed, 32'h00000000} /* (1, 7, 1) {real, imag} */,
  {32'h44db557a, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'hc33c64ba, 32'h00000000} /* (1, 6, 15) {real, imag} */,
  {32'hc1f9ec70, 32'h00000000} /* (1, 6, 14) {real, imag} */,
  {32'h43a14c2c, 32'h00000000} /* (1, 6, 13) {real, imag} */,
  {32'h43d6a809, 32'h00000000} /* (1, 6, 12) {real, imag} */,
  {32'h43d213c2, 32'h00000000} /* (1, 6, 11) {real, imag} */,
  {32'h43a06832, 32'h00000000} /* (1, 6, 10) {real, imag} */,
  {32'h425152a0, 32'h00000000} /* (1, 6, 9) {real, imag} */,
  {32'hc37f9098, 32'h00000000} /* (1, 6, 8) {real, imag} */,
  {32'h43c87553, 32'h00000000} /* (1, 6, 7) {real, imag} */,
  {32'hc46330b6, 32'h00000000} /* (1, 6, 6) {real, imag} */,
  {32'hc4b44c02, 32'h00000000} /* (1, 6, 5) {real, imag} */,
  {32'h42668b78, 32'h00000000} /* (1, 6, 4) {real, imag} */,
  {32'hc4576e31, 32'h00000000} /* (1, 6, 3) {real, imag} */,
  {32'hc4bca570, 32'h00000000} /* (1, 6, 2) {real, imag} */,
  {32'h43cce530, 32'h00000000} /* (1, 6, 1) {real, imag} */,
  {32'h44b49e74, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'hc3726d03, 32'h00000000} /* (1, 5, 15) {real, imag} */,
  {32'hc4177efb, 32'h00000000} /* (1, 5, 14) {real, imag} */,
  {32'h42df7c2c, 32'h00000000} /* (1, 5, 13) {real, imag} */,
  {32'h441ed469, 32'h00000000} /* (1, 5, 12) {real, imag} */,
  {32'h4456f641, 32'h00000000} /* (1, 5, 11) {real, imag} */,
  {32'h4225fbfd, 32'h00000000} /* (1, 5, 10) {real, imag} */,
  {32'hc439dff6, 32'h00000000} /* (1, 5, 9) {real, imag} */,
  {32'h43ab1690, 32'h00000000} /* (1, 5, 8) {real, imag} */,
  {32'hc35dfb47, 32'h00000000} /* (1, 5, 7) {real, imag} */,
  {32'hc3aa3592, 32'h00000000} /* (1, 5, 6) {real, imag} */,
  {32'hc46e5896, 32'h00000000} /* (1, 5, 5) {real, imag} */,
  {32'hc3f4d546, 32'h00000000} /* (1, 5, 4) {real, imag} */,
  {32'h41d2a8a0, 32'h00000000} /* (1, 5, 3) {real, imag} */,
  {32'h42d73ade, 32'h00000000} /* (1, 5, 2) {real, imag} */,
  {32'h4434b542, 32'h00000000} /* (1, 5, 1) {real, imag} */,
  {32'h4450e086, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'hc4a65917, 32'h00000000} /* (1, 4, 15) {real, imag} */,
  {32'hc45ed7eb, 32'h00000000} /* (1, 4, 14) {real, imag} */,
  {32'h44401b3a, 32'h00000000} /* (1, 4, 13) {real, imag} */,
  {32'h42649e80, 32'h00000000} /* (1, 4, 12) {real, imag} */,
  {32'h4317002d, 32'h00000000} /* (1, 4, 11) {real, imag} */,
  {32'h4436dc32, 32'h00000000} /* (1, 4, 10) {real, imag} */,
  {32'hc432c5f0, 32'h00000000} /* (1, 4, 9) {real, imag} */,
  {32'hc3f00a54, 32'h00000000} /* (1, 4, 8) {real, imag} */,
  {32'h43ecbde4, 32'h00000000} /* (1, 4, 7) {real, imag} */,
  {32'hc46c3905, 32'h00000000} /* (1, 4, 6) {real, imag} */,
  {32'hc4871b7b, 32'h00000000} /* (1, 4, 5) {real, imag} */,
  {32'hc403421b, 32'h00000000} /* (1, 4, 4) {real, imag} */,
  {32'hc3c6956e, 32'h00000000} /* (1, 4, 3) {real, imag} */,
  {32'h43f2b7ac, 32'h00000000} /* (1, 4, 2) {real, imag} */,
  {32'h43d88dd7, 32'h00000000} /* (1, 4, 1) {real, imag} */,
  {32'h43cbb15c, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hc3e0e8d0, 32'h00000000} /* (1, 3, 15) {real, imag} */,
  {32'h4421610e, 32'h00000000} /* (1, 3, 14) {real, imag} */,
  {32'h43d060dc, 32'h00000000} /* (1, 3, 13) {real, imag} */,
  {32'h438fe7aa, 32'h00000000} /* (1, 3, 12) {real, imag} */,
  {32'h4481b86b, 32'h00000000} /* (1, 3, 11) {real, imag} */,
  {32'h439494e2, 32'h00000000} /* (1, 3, 10) {real, imag} */,
  {32'h445b3bee, 32'h00000000} /* (1, 3, 9) {real, imag} */,
  {32'hc2f4d5ae, 32'h00000000} /* (1, 3, 8) {real, imag} */,
  {32'hc2cf69e0, 32'h00000000} /* (1, 3, 7) {real, imag} */,
  {32'hc493cacb, 32'h00000000} /* (1, 3, 6) {real, imag} */,
  {32'hc522b138, 32'h00000000} /* (1, 3, 5) {real, imag} */,
  {32'hc48eec2e, 32'h00000000} /* (1, 3, 4) {real, imag} */,
  {32'hc4587b64, 32'h00000000} /* (1, 3, 3) {real, imag} */,
  {32'hc3e412ae, 32'h00000000} /* (1, 3, 2) {real, imag} */,
  {32'hc4235f7e, 32'h00000000} /* (1, 3, 1) {real, imag} */,
  {32'hc30f1899, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hc4615a5c, 32'h00000000} /* (1, 2, 15) {real, imag} */,
  {32'hc3903ce9, 32'h00000000} /* (1, 2, 14) {real, imag} */,
  {32'hc20e9288, 32'h00000000} /* (1, 2, 13) {real, imag} */,
  {32'h43957060, 32'h00000000} /* (1, 2, 12) {real, imag} */,
  {32'h448e9536, 32'h00000000} /* (1, 2, 11) {real, imag} */,
  {32'h43d4cc98, 32'h00000000} /* (1, 2, 10) {real, imag} */,
  {32'h4319b0c0, 32'h00000000} /* (1, 2, 9) {real, imag} */,
  {32'h42677038, 32'h00000000} /* (1, 2, 8) {real, imag} */,
  {32'h4419074a, 32'h00000000} /* (1, 2, 7) {real, imag} */,
  {32'hc39ef9af, 32'h00000000} /* (1, 2, 6) {real, imag} */,
  {32'hc4317430, 32'h00000000} /* (1, 2, 5) {real, imag} */,
  {32'hc4089f10, 32'h00000000} /* (1, 2, 4) {real, imag} */,
  {32'hc419f768, 32'h00000000} /* (1, 2, 3) {real, imag} */,
  {32'hc481c440, 32'h00000000} /* (1, 2, 2) {real, imag} */,
  {32'hc4c61dd8, 32'h00000000} /* (1, 2, 1) {real, imag} */,
  {32'h423bb888, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hc4320b06, 32'h00000000} /* (1, 1, 15) {real, imag} */,
  {32'hc4add5c1, 32'h00000000} /* (1, 1, 14) {real, imag} */,
  {32'h4296e7d8, 32'h00000000} /* (1, 1, 13) {real, imag} */,
  {32'h44838700, 32'h00000000} /* (1, 1, 12) {real, imag} */,
  {32'h43bf803a, 32'h00000000} /* (1, 1, 11) {real, imag} */,
  {32'h42b4f490, 32'h00000000} /* (1, 1, 10) {real, imag} */,
  {32'hc3f317f7, 32'h00000000} /* (1, 1, 9) {real, imag} */,
  {32'h4420eeb9, 32'h00000000} /* (1, 1, 8) {real, imag} */,
  {32'h42dea070, 32'h00000000} /* (1, 1, 7) {real, imag} */,
  {32'hc1f74a40, 32'h00000000} /* (1, 1, 6) {real, imag} */,
  {32'h444395ef, 32'h00000000} /* (1, 1, 5) {real, imag} */,
  {32'hc420d9d4, 32'h00000000} /* (1, 1, 4) {real, imag} */,
  {32'hc4318ff9, 32'h00000000} /* (1, 1, 3) {real, imag} */,
  {32'hc488c48f, 32'h00000000} /* (1, 1, 2) {real, imag} */,
  {32'h434418ae, 32'h00000000} /* (1, 1, 1) {real, imag} */,
  {32'hc3b52b06, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hc384b831, 32'h00000000} /* (1, 0, 15) {real, imag} */,
  {32'h429b76ba, 32'h00000000} /* (1, 0, 14) {real, imag} */,
  {32'hc2cfb810, 32'h00000000} /* (1, 0, 13) {real, imag} */,
  {32'h43e9f94a, 32'h00000000} /* (1, 0, 12) {real, imag} */,
  {32'h43a9c6cc, 32'h00000000} /* (1, 0, 11) {real, imag} */,
  {32'hc3ca6d6b, 32'h00000000} /* (1, 0, 10) {real, imag} */,
  {32'hc3918106, 32'h00000000} /* (1, 0, 9) {real, imag} */,
  {32'hc396f8eb, 32'h00000000} /* (1, 0, 8) {real, imag} */,
  {32'hc25ea598, 32'h00000000} /* (1, 0, 7) {real, imag} */,
  {32'h432b0c05, 32'h00000000} /* (1, 0, 6) {real, imag} */,
  {32'hc3a84328, 32'h00000000} /* (1, 0, 5) {real, imag} */,
  {32'hc41d19c5, 32'h00000000} /* (1, 0, 4) {real, imag} */,
  {32'hc48322d4, 32'h00000000} /* (1, 0, 3) {real, imag} */,
  {32'hc428e32e, 32'h00000000} /* (1, 0, 2) {real, imag} */,
  {32'hc3aaff1e, 32'h00000000} /* (1, 0, 1) {real, imag} */,
  {32'hc41b208e, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'h4343009c, 32'h00000000} /* (0, 15, 15) {real, imag} */,
  {32'h42455df0, 32'h00000000} /* (0, 15, 14) {real, imag} */,
  {32'hc363ba88, 32'h00000000} /* (0, 15, 13) {real, imag} */,
  {32'h4382fa78, 32'h00000000} /* (0, 15, 12) {real, imag} */,
  {32'h43251c54, 32'h00000000} /* (0, 15, 11) {real, imag} */,
  {32'hc3f75197, 32'h00000000} /* (0, 15, 10) {real, imag} */,
  {32'hc41ca6e4, 32'h00000000} /* (0, 15, 9) {real, imag} */,
  {32'hc2b884fc, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'hc12e3ac8, 32'h00000000} /* (0, 15, 7) {real, imag} */,
  {32'hc331efa4, 32'h00000000} /* (0, 15, 6) {real, imag} */,
  {32'hc3a0a564, 32'h00000000} /* (0, 15, 5) {real, imag} */,
  {32'hc4097cd8, 32'h00000000} /* (0, 15, 4) {real, imag} */,
  {32'hc4053d1b, 32'h00000000} /* (0, 15, 3) {real, imag} */,
  {32'hc3c76e61, 32'h00000000} /* (0, 15, 2) {real, imag} */,
  {32'hc350b6c0, 32'h00000000} /* (0, 15, 1) {real, imag} */,
  {32'hc3cfd3e1, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h4412951e, 32'h00000000} /* (0, 14, 15) {real, imag} */,
  {32'h431dae14, 32'h00000000} /* (0, 14, 14) {real, imag} */,
  {32'hc3c87762, 32'h00000000} /* (0, 14, 13) {real, imag} */,
  {32'hc28ec6ce, 32'h00000000} /* (0, 14, 12) {real, imag} */,
  {32'h44928926, 32'h00000000} /* (0, 14, 11) {real, imag} */,
  {32'hc3413bc8, 32'h00000000} /* (0, 14, 10) {real, imag} */,
  {32'hc435ba52, 32'h00000000} /* (0, 14, 9) {real, imag} */,
  {32'hc25354d8, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'hc3c5f2f9, 32'h00000000} /* (0, 14, 7) {real, imag} */,
  {32'h43238564, 32'h00000000} /* (0, 14, 6) {real, imag} */,
  {32'h3fa38b00, 32'h00000000} /* (0, 14, 5) {real, imag} */,
  {32'hc40718a9, 32'h00000000} /* (0, 14, 4) {real, imag} */,
  {32'hc3df7508, 32'h00000000} /* (0, 14, 3) {real, imag} */,
  {32'hc3b3d638, 32'h00000000} /* (0, 14, 2) {real, imag} */,
  {32'h43a169fc, 32'h00000000} /* (0, 14, 1) {real, imag} */,
  {32'h439db2f5, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h42458828, 32'h00000000} /* (0, 13, 15) {real, imag} */,
  {32'h43d4bed4, 32'h00000000} /* (0, 13, 14) {real, imag} */,
  {32'h431894f5, 32'h00000000} /* (0, 13, 13) {real, imag} */,
  {32'h4419cefa, 32'h00000000} /* (0, 13, 12) {real, imag} */,
  {32'h43aa6ffb, 32'h00000000} /* (0, 13, 11) {real, imag} */,
  {32'h3e326000, 32'h00000000} /* (0, 13, 10) {real, imag} */,
  {32'h42e85f64, 32'h00000000} /* (0, 13, 9) {real, imag} */,
  {32'hc3489824, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'hc398dd0b, 32'h00000000} /* (0, 13, 7) {real, imag} */,
  {32'hc3e7e190, 32'h00000000} /* (0, 13, 6) {real, imag} */,
  {32'hc327319f, 32'h00000000} /* (0, 13, 5) {real, imag} */,
  {32'hc38ef108, 32'h00000000} /* (0, 13, 4) {real, imag} */,
  {32'hc3ad5da1, 32'h00000000} /* (0, 13, 3) {real, imag} */,
  {32'h43858268, 32'h00000000} /* (0, 13, 2) {real, imag} */,
  {32'h43e19ec3, 32'h00000000} /* (0, 13, 1) {real, imag} */,
  {32'h433b13ba, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'h4251b4c8, 32'h00000000} /* (0, 12, 15) {real, imag} */,
  {32'h43c898a3, 32'h00000000} /* (0, 12, 14) {real, imag} */,
  {32'h4435edb0, 32'h00000000} /* (0, 12, 13) {real, imag} */,
  {32'h43ced6d9, 32'h00000000} /* (0, 12, 12) {real, imag} */,
  {32'h43c9d139, 32'h00000000} /* (0, 12, 11) {real, imag} */,
  {32'hc3fa86a8, 32'h00000000} /* (0, 12, 10) {real, imag} */,
  {32'hc429475a, 32'h00000000} /* (0, 12, 9) {real, imag} */,
  {32'hc4a8bac8, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'hc403a104, 32'h00000000} /* (0, 12, 7) {real, imag} */,
  {32'hc3badd25, 32'h00000000} /* (0, 12, 6) {real, imag} */,
  {32'hc3a3ee7c, 32'h00000000} /* (0, 12, 5) {real, imag} */,
  {32'hc3e702d9, 32'h00000000} /* (0, 12, 4) {real, imag} */,
  {32'h441abc14, 32'h00000000} /* (0, 12, 3) {real, imag} */,
  {32'h44284dce, 32'h00000000} /* (0, 12, 2) {real, imag} */,
  {32'h443aa20e, 32'h00000000} /* (0, 12, 1) {real, imag} */,
  {32'h443ebb15, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h437c130e, 32'h00000000} /* (0, 11, 15) {real, imag} */,
  {32'h43e63432, 32'h00000000} /* (0, 11, 14) {real, imag} */,
  {32'h438e5aca, 32'h00000000} /* (0, 11, 13) {real, imag} */,
  {32'hc262e7c8, 32'h00000000} /* (0, 11, 12) {real, imag} */,
  {32'h43a42dec, 32'h00000000} /* (0, 11, 11) {real, imag} */,
  {32'h43915467, 32'h00000000} /* (0, 11, 10) {real, imag} */,
  {32'h4229d024, 32'h00000000} /* (0, 11, 9) {real, imag} */,
  {32'hc03dc240, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'h41039018, 32'h00000000} /* (0, 11, 7) {real, imag} */,
  {32'hc382e89e, 32'h00000000} /* (0, 11, 6) {real, imag} */,
  {32'hc310e78a, 32'h00000000} /* (0, 11, 5) {real, imag} */,
  {32'h425a3238, 32'h00000000} /* (0, 11, 4) {real, imag} */,
  {32'hc38e0686, 32'h00000000} /* (0, 11, 3) {real, imag} */,
  {32'hc34b01ae, 32'h00000000} /* (0, 11, 2) {real, imag} */,
  {32'h4404d536, 32'h00000000} /* (0, 11, 1) {real, imag} */,
  {32'h43d05cec, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h4362cd81, 32'h00000000} /* (0, 10, 15) {real, imag} */,
  {32'h43d9326c, 32'h00000000} /* (0, 10, 14) {real, imag} */,
  {32'h4408c415, 32'h00000000} /* (0, 10, 13) {real, imag} */,
  {32'h43d5ed99, 32'h00000000} /* (0, 10, 12) {real, imag} */,
  {32'h44160d9a, 32'h00000000} /* (0, 10, 11) {real, imag} */,
  {32'h435a126f, 32'h00000000} /* (0, 10, 10) {real, imag} */,
  {32'h442c6424, 32'h00000000} /* (0, 10, 9) {real, imag} */,
  {32'h425163c4, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'hc250022c, 32'h00000000} /* (0, 10, 7) {real, imag} */,
  {32'hc3419b43, 32'h00000000} /* (0, 10, 6) {real, imag} */,
  {32'hc42a0a61, 32'h00000000} /* (0, 10, 5) {real, imag} */,
  {32'h42e4aa44, 32'h00000000} /* (0, 10, 4) {real, imag} */,
  {32'h431d91d7, 32'h00000000} /* (0, 10, 3) {real, imag} */,
  {32'hc38e212c, 32'h00000000} /* (0, 10, 2) {real, imag} */,
  {32'hc22b0508, 32'h00000000} /* (0, 10, 1) {real, imag} */,
  {32'h43ada99c, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'h43ea9a28, 32'h00000000} /* (0, 9, 15) {real, imag} */,
  {32'h42d99d6c, 32'h00000000} /* (0, 9, 14) {real, imag} */,
  {32'hc31c6cdb, 32'h00000000} /* (0, 9, 13) {real, imag} */,
  {32'h43ea0aea, 32'h00000000} /* (0, 9, 12) {real, imag} */,
  {32'h442673da, 32'h00000000} /* (0, 9, 11) {real, imag} */,
  {32'h44384b65, 32'h00000000} /* (0, 9, 10) {real, imag} */,
  {32'h439e0420, 32'h00000000} /* (0, 9, 9) {real, imag} */,
  {32'hc41a8c9e, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'hc3c1801a, 32'h00000000} /* (0, 9, 7) {real, imag} */,
  {32'h448a8ffe, 32'h00000000} /* (0, 9, 6) {real, imag} */,
  {32'hc0e01160, 32'h00000000} /* (0, 9, 5) {real, imag} */,
  {32'h4392bb2a, 32'h00000000} /* (0, 9, 4) {real, imag} */,
  {32'h43a86f33, 32'h00000000} /* (0, 9, 3) {real, imag} */,
  {32'h43aa8fc2, 32'h00000000} /* (0, 9, 2) {real, imag} */,
  {32'h4431b440, 32'h00000000} /* (0, 9, 1) {real, imag} */,
  {32'h442e3db2, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'h439781e6, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'h43d20445, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'hc3bc420c, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'h43a2998e, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'h43246328, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'h43aaf1d4, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hc3a4d749, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'hc3e783fb, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hc39f04ce, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hc4138496, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'h425ffa80, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'hc33f0e48, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'h43647d28, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'h444d03aa, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'h43d91683, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'h442228fa, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h437bd97e, 32'h00000000} /* (0, 7, 15) {real, imag} */,
  {32'h42919d10, 32'h00000000} /* (0, 7, 14) {real, imag} */,
  {32'hc2928574, 32'h00000000} /* (0, 7, 13) {real, imag} */,
  {32'h42508628, 32'h00000000} /* (0, 7, 12) {real, imag} */,
  {32'h4331f5e4, 32'h00000000} /* (0, 7, 11) {real, imag} */,
  {32'h44077231, 32'h00000000} /* (0, 7, 10) {real, imag} */,
  {32'h43d9e126, 32'h00000000} /* (0, 7, 9) {real, imag} */,
  {32'hc2a0a046, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'hc3cd3d39, 32'h00000000} /* (0, 7, 7) {real, imag} */,
  {32'hc3fbe0e4, 32'h00000000} /* (0, 7, 6) {real, imag} */,
  {32'hc4272154, 32'h00000000} /* (0, 7, 5) {real, imag} */,
  {32'hc2064158, 32'h00000000} /* (0, 7, 4) {real, imag} */,
  {32'h4395331a, 32'h00000000} /* (0, 7, 3) {real, imag} */,
  {32'h4391ff71, 32'h00000000} /* (0, 7, 2) {real, imag} */,
  {32'h43d57626, 32'h00000000} /* (0, 7, 1) {real, imag} */,
  {32'h43ff1c10, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'h4376c79d, 32'h00000000} /* (0, 6, 15) {real, imag} */,
  {32'hc3a074a8, 32'h00000000} /* (0, 6, 14) {real, imag} */,
  {32'hc32fc29a, 32'h00000000} /* (0, 6, 13) {real, imag} */,
  {32'h4388d9fc, 32'h00000000} /* (0, 6, 12) {real, imag} */,
  {32'h42181018, 32'h00000000} /* (0, 6, 11) {real, imag} */,
  {32'h43c27de2, 32'h00000000} /* (0, 6, 10) {real, imag} */,
  {32'h437621c7, 32'h00000000} /* (0, 6, 9) {real, imag} */,
  {32'hc3b1adf2, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'hc38af74a, 32'h00000000} /* (0, 6, 7) {real, imag} */,
  {32'hc3ed667c, 32'h00000000} /* (0, 6, 6) {real, imag} */,
  {32'hc40f9e7a, 32'h00000000} /* (0, 6, 5) {real, imag} */,
  {32'hc4096f16, 32'h00000000} /* (0, 6, 4) {real, imag} */,
  {32'hc43f4382, 32'h00000000} /* (0, 6, 3) {real, imag} */,
  {32'hc45849ef, 32'h00000000} /* (0, 6, 2) {real, imag} */,
  {32'h43fbb1ba, 32'h00000000} /* (0, 6, 1) {real, imag} */,
  {32'h44050101, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'h41d94a00, 32'h00000000} /* (0, 5, 15) {real, imag} */,
  {32'hc3c2c309, 32'h00000000} /* (0, 5, 14) {real, imag} */,
  {32'h41a486c8, 32'h00000000} /* (0, 5, 13) {real, imag} */,
  {32'h43304f6c, 32'h00000000} /* (0, 5, 12) {real, imag} */,
  {32'h44225eca, 32'h00000000} /* (0, 5, 11) {real, imag} */,
  {32'h4404d2da, 32'h00000000} /* (0, 5, 10) {real, imag} */,
  {32'h42606fb2, 32'h00000000} /* (0, 5, 9) {real, imag} */,
  {32'h43cf58b6, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'hc30c0544, 32'h00000000} /* (0, 5, 7) {real, imag} */,
  {32'h438c0519, 32'h00000000} /* (0, 5, 6) {real, imag} */,
  {32'hc3fe298c, 32'h00000000} /* (0, 5, 5) {real, imag} */,
  {32'hc3856091, 32'h00000000} /* (0, 5, 4) {real, imag} */,
  {32'hc3beddf7, 32'h00000000} /* (0, 5, 3) {real, imag} */,
  {32'h430e5918, 32'h00000000} /* (0, 5, 2) {real, imag} */,
  {32'h4357f162, 32'h00000000} /* (0, 5, 1) {real, imag} */,
  {32'h42da73b0, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'h433c720e, 32'h00000000} /* (0, 4, 15) {real, imag} */,
  {32'h4395db55, 32'h00000000} /* (0, 4, 14) {real, imag} */,
  {32'h4360d80a, 32'h00000000} /* (0, 4, 13) {real, imag} */,
  {32'h43f000b1, 32'h00000000} /* (0, 4, 12) {real, imag} */,
  {32'hc1a9a6b0, 32'h00000000} /* (0, 4, 11) {real, imag} */,
  {32'h43fd5506, 32'h00000000} /* (0, 4, 10) {real, imag} */,
  {32'h439c0f64, 32'h00000000} /* (0, 4, 9) {real, imag} */,
  {32'h433c874a, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'hc3478fce, 32'h00000000} /* (0, 4, 7) {real, imag} */,
  {32'hc415b054, 32'h00000000} /* (0, 4, 6) {real, imag} */,
  {32'hc413220c, 32'h00000000} /* (0, 4, 5) {real, imag} */,
  {32'hc47fd2d4, 32'h00000000} /* (0, 4, 4) {real, imag} */,
  {32'hc3a8aaff, 32'h00000000} /* (0, 4, 3) {real, imag} */,
  {32'hc2881fe0, 32'h00000000} /* (0, 4, 2) {real, imag} */,
  {32'h42110730, 32'h00000000} /* (0, 4, 1) {real, imag} */,
  {32'hc36b2eae, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hc16f0c20, 32'h00000000} /* (0, 3, 15) {real, imag} */,
  {32'h43a229d2, 32'h00000000} /* (0, 3, 14) {real, imag} */,
  {32'h44596666, 32'h00000000} /* (0, 3, 13) {real, imag} */,
  {32'h4339147e, 32'h00000000} /* (0, 3, 12) {real, imag} */,
  {32'h441816a6, 32'h00000000} /* (0, 3, 11) {real, imag} */,
  {32'hc2a83d9a, 32'h00000000} /* (0, 3, 10) {real, imag} */,
  {32'h43ba1b67, 32'h00000000} /* (0, 3, 9) {real, imag} */,
  {32'h438024c4, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h441e951e, 32'h00000000} /* (0, 3, 7) {real, imag} */,
  {32'hc429e1a1, 32'h00000000} /* (0, 3, 6) {real, imag} */,
  {32'hc48285b8, 32'h00000000} /* (0, 3, 5) {real, imag} */,
  {32'hc3e579af, 32'h00000000} /* (0, 3, 4) {real, imag} */,
  {32'hc4197f1e, 32'h00000000} /* (0, 3, 3) {real, imag} */,
  {32'hc40cafa5, 32'h00000000} /* (0, 3, 2) {real, imag} */,
  {32'hc46ffebc, 32'h00000000} /* (0, 3, 1) {real, imag} */,
  {32'hc43090f6, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hc3bb210f, 32'h00000000} /* (0, 2, 15) {real, imag} */,
  {32'hc2a8ba20, 32'h00000000} /* (0, 2, 14) {real, imag} */,
  {32'h441a7fcf, 32'h00000000} /* (0, 2, 13) {real, imag} */,
  {32'hc2689c08, 32'h00000000} /* (0, 2, 12) {real, imag} */,
  {32'h446bfaf9, 32'h00000000} /* (0, 2, 11) {real, imag} */,
  {32'h4446e610, 32'h00000000} /* (0, 2, 10) {real, imag} */,
  {32'h43fc01e8, 32'h00000000} /* (0, 2, 9) {real, imag} */,
  {32'h43b28861, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'h43e8ffe9, 32'h00000000} /* (0, 2, 7) {real, imag} */,
  {32'hc49990f5, 32'h00000000} /* (0, 2, 6) {real, imag} */,
  {32'hc2faf62a, 32'h00000000} /* (0, 2, 5) {real, imag} */,
  {32'h43ceecb3, 32'h00000000} /* (0, 2, 4) {real, imag} */,
  {32'hc43704cb, 32'h00000000} /* (0, 2, 3) {real, imag} */,
  {32'hc44390dc, 32'h00000000} /* (0, 2, 2) {real, imag} */,
  {32'hc44c718c, 32'h00000000} /* (0, 2, 1) {real, imag} */,
  {32'hc3d48a0f, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hc428b152, 32'h00000000} /* (0, 1, 15) {real, imag} */,
  {32'hc3d663c2, 32'h00000000} /* (0, 1, 14) {real, imag} */,
  {32'h435744bb, 32'h00000000} /* (0, 1, 13) {real, imag} */,
  {32'h4439bb42, 32'h00000000} /* (0, 1, 12) {real, imag} */,
  {32'h429e8740, 32'h00000000} /* (0, 1, 11) {real, imag} */,
  {32'hc3a1cb6c, 32'h00000000} /* (0, 1, 10) {real, imag} */,
  {32'h44248650, 32'h00000000} /* (0, 1, 9) {real, imag} */,
  {32'hc2e99f7e, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'hc34cf008, 32'h00000000} /* (0, 1, 7) {real, imag} */,
  {32'h424206a4, 32'h00000000} /* (0, 1, 6) {real, imag} */,
  {32'hc20099b4, 32'h00000000} /* (0, 1, 5) {real, imag} */,
  {32'hc3c62c44, 32'h00000000} /* (0, 1, 4) {real, imag} */,
  {32'hc41c4d74, 32'h00000000} /* (0, 1, 3) {real, imag} */,
  {32'hc484ea47, 32'h00000000} /* (0, 1, 2) {real, imag} */,
  {32'hc385d634, 32'h00000000} /* (0, 1, 1) {real, imag} */,
  {32'hc2854a0e, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hc42c02a0, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'hc383c1c5, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'h43372925, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h441ce2bc, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'h43721458, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'hc25819fa, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'hc42bd97c, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'hc302e5da, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'hc30560fc, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'hc3dd66c3, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'hc3d58904, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'hc40ade14, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'hc3d1d6f4, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'hc393c1b8, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'hc3f57b20, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'hc326d50e, 32'h00000000} /* (0, 0, 0) {real, imag} */};
