-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MKstdB+VmobPDQl/eIW0TO8BM6xq3Xy6yuiKLzr/WipbboOMy0fjGDLDsNp5h5Sx4ZxDeoxbIibE
q037INCNdXjqIQpo9WUYJaioo72bdbLQrwt2RJXslbnifntIRnZfvlCLjBfqM0g5ynjemVjd43/O
DtmaOZQICLab++D5RjaAunMo9uII5Dhwtvad/Cqhb41O9+OTpmUjUS8uGuV6KJHs2A89jrIccyTm
AGPHT3zff8pNO/i9NtH+DvoZZJYJDXSSW34F4bL8J5Wi/vi0rLT0NX2YJ11sw6RwkPWA/SczefsF
9H6RrJvumDb8vCn+CUEImG51/M01+n4GBB+DwQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 42976)
`protect data_block
4CYFqW5Jvf5lCZUByOXhSoQIqH8w6Rlv1gs8UcoYx7p9ofSa/uB/cjqS8zl+2zPYTIF2Jv6HPzF3
WsubGuYvJ3BdSsxzUbQqZ1JCI8D0E8ucwBZnRNVSGeIrS0wUsFsiNfLvFna6FV7pepObMMU9n2T4
pdi1+O35yh00QNMGQ4bAtX8DynZHZJLHoH3TpKnmbtM2/fqxCEmyKc3JHMIlGfaiPt/VrCCHnzX4
/MV7IxtbCColkqu9aX+wm5Ugfr+bR7u2xQvQt1LkE+KVePN/STVqAVQxuCHZbgKnHTcX2IKXUoLO
0587zZhMTyE43Z0v/NRIMRAl/rFNnOaxQGhQucSZgfmfOwjhnWdBH7fh5PZ2ZNxPv81aMaNOR9jx
LFScecnTK+ZXkD1j93aGWHkvirEqocGTiU728nMF4MRBA0TjpIHqOxguQP8kGQeefWC8dCULRqRE
XErnxUnxgLN4sdo9W9h8ZaUJrN6nOGeKgvUBGT3wbAp1vvqzAyiG6z/o625AjzIip+3oMYnnRj8h
Uv3iv3RMXeMsZNBUw9DY6ygkXB0qXQLs/AU+8KeDxSSeUQd9i9/mReSjRsQbmumGYMCOnJliQk4m
1DFDWQ9NROtezj5OBhmtfCibaFrywicHTLgP6/umTb+iXJ00kyuMem1Aj+/h8eOYfTADKk/wTfhz
0MSjH2YhDIRi7GimQfCZGa7VtmmykL+18kvaIWrCjNXYFHK70xQA1ioijtQ6UtW8LpY6fj8WusLQ
ZlH867gVqVCGjpFGrLJxJqvEMV+6Dlk6HVjZw9WtwcIPOnuXJ5gvA7i9PUyQ8z1pPhJMF5E2uqyB
j01DSOSJBuo+lGtohRMUjKUdV6gxrH54RtoTBfEEefN7q4dAkX4tV3Ep1D19PxqIg+eTRXgrlovZ
ISi6JKrPaoKfCH4nECa0oQfnV+mFnKN7UkgOw1mfmkTUOAfqIIMsUz4SpkBiKUkqqU2I3Hq2otfK
amV3r2+TxxBB1Pq4ntKclWZ/DiFVXlLsu9vFrfDVVs6tQhVNHnU5gl2s8IexBYP0B3LY627slSZ2
JzU9ipMrWoM9mKF+67oH4JiOUxI3RcwEyQIzMy1J3Q7ezJcIiTzTOddUEyvZLZh5x/bYHAYnjIwZ
zxBoWyE6FiO69fpXUPMp9bzLGFbb3QwLdgB6BvlnuHFFpDnSi6i162fIU3cXc+NjhL6w/aSuLyTS
BWdGSaS0r/MnGa/bUWk/x3MRqZqhdt/LjvLoARKdBQscG0cJ6oVhzv+vz5L8WeHefrziZgS4eWcZ
LnAND3pyG+fT4GzndhPs25RFdZ4qNBOK4/yi42DbXoM2WYSizfaqmOcPmnVqfUHEb2s9Y46bxWPh
+9Wu9VXa7UtxU7uGIiIFpRL7JeNQjHOvcZEXfKAFuTX+m2qbH7oCr5GIk3hbLcPhnoB6o92bdbQT
qxQAqMYGVacCl9dgiXA4Qhr4Ko82wfjTzabCDhPxhHOd799bl/Ddm+AG9n+i/y890BqQSSW5GDE0
Ftl+vo0Jy2hoC3QQ6zknfEVeObQ6x+qM9vNsm2+g7s0xbmCOh9EASxBC1nJ/rCTOAwV/yFhc3ilr
ffAmrEKzSMp8Ny/iVOeEClBNKmK9obqGnuGLL+g43AgrijtYvHMeinlCGk9gkYVzBcVuyMLKeLxP
NlOveAM7LTsLq8tZPkQz0dE9Mpv4nZwjCe5InubzoLWfwIBdbnyc9mC6y37S939t2u9WDGuD7Q5A
1XsZXKFAEris7yr519sdx/XM67dLCyGwlv3J4Xs5P/zcj1hQ2mWgIRgSpwJnkYXmKR5lfHiXLP6n
WDQB0VMsER2OXxW3D+hM3Yr4FatDtPNzrXcpGAm08+4p0xRbu37TmV4n4OQhCOcYpph9RWqKJr7D
3KCkUiBN7VFaQnVvrQsdUhF9fc5AvaLwQU+Bm7G4pW9hKyCkxfdPEPA9BYwD+fRxvGCb/MzGqRa7
k9fP7r71JnDrjBAYSOau5Y1PYHMGrskgdVgI9jnTOTv9TuOKQHthY5Em9bTS1D70+DrgoCjOH9pT
b2bgrm84/qRb7/+wrgyp63y3F77hB34XuMljXXQujy7GeJuPz8sn4rBANHn04NGg7gmcU+z5sxfC
xr7Nw26W94DbPZu+1zhv/CVM/NA8/h2UFUtV1Ahw1B4Kzpc89OMJZNKfQbnW8ELfasCnLj7GcuPt
SI/z4mJbd523w2N3jhS6PmODh7T5uLkv7wDCv2DIAhZ783Zp6G3YjfDKXpE/7GNJ9o6n3zRVL7aC
WkA9TgchFj/nOERezyi8xBrN6E1O++AOlvh/9RX9xKIWVaA5wuE1t6upG+sKHb5i3pvYkULpLUhe
csPbZwZHvAgfD7imyOFfO9k4ahsuIsh58ixovAkxd8Gi0LIdcVGxDq0trhVHcF2xC6MCRx3RSuwi
wzjf6Cmd4NEVJfZvPERGXXGgRPUNW8EETHSumTz7yn5LTE16EyfOIp+stTB/hAW2dfauz/+XLzTd
pW4QAh3TFMsLBkqHkxxYqvCwosb8ullZqL1/BOHNv8HcRam2VwkQZkCYw/FTNiq9oKOxt8lW9aaP
CufIzPTGFTwf97aa6+1rqhv8ILUvYeagYjLFfnoWXT2s21gHWH9GRAlP4gGIN5yYMUQCuIMBlzHM
uPEqskkDmAAnrZi+2d3DDYxf6Hbn+nMlyRepj3HbVB3FGDkhYsMuu/gHKwxbR50fhl9fs7SYeX39
Rshfo/zv3LOfiuffgR3cN2eVCL181Y1z203rkmT06dEKOU9lqps4p/m9aq9TyFGiDxIm10Kbts5X
B1Xh8YkhYQ/CAjCwxHfuyk0sNJ3Eam+wZMcVDGv6ys2nxlbtIzXLfI+wvhgWNqBsGp5R6EtWRq8c
Q1oM3ohysnws0IgOdBAoitqXoUfTqxoPOosiG6XIBx3ZNplCdS8z4b0ZqrVnYe48oIgiK92vA8xz
ut5Fyp61T6ZsY5rxMlLVt3FEovaiOl1drdAhTTNOi78vvCsvSzeZsG7Kov6NEfK+mMJDam+8tc/x
uwBY5dsmsg7vhNSFfWs+m0Fcf8uIrWjdXyz1BP3m0DyGXbE8rEADmYo9t2y5wwkZK0/ayU4CJw4E
A6SGxiNiwqrckmKjETJKprgOkx/VYR1YGfd59jhcyHdycdTDqfs/05dfJH19tN3uIBXZpsVPSep7
UHHNl00ZWSPflOAFm4LQzYtJAN5+vjiXXrXs73n+mCUfhiPo/SbLGCK1TLxOB5Xm9LHRGeqZ8h7r
kkzTkOrls7pq/DrqylvW4VLKTvaGJMqODmLDacTKIU8dLludFcQBN/aGXr6UtK1wx0EO4OSDfQrw
Ig3uY15nRFAp3N/Q+BIIRCFWg4TKSRhG9v15/V5LpchtyLMg03USqkwybcGbBRqGHlVylH7LN3q1
cxYEtUBRcHqYyw1SFg+ucxSUqdxxj9dFPQHPmpq1/NcRNVtmBk5WLq3pNrOwrg2rA7AafsJOqeKZ
PJZYEOlmYAeRKiEoNkT+g4fuwI+vFZmY1I9Cq72cP11q39sxpmEv9ie9DeNwgTb2s1qXFwckuB28
VnDvtLNc97VR6uscmI5VZFjN31zLfli4AYD1Q1zxV0Yy3q4Xxn8jspQQfy2HwCDMleWS0XMrNJYj
O9H/4M+iQa5BhWJjHeG0xKeKHhmPq3iyCNqYssbenc98hccTvCj6On4Tw/63XWiUlakTtl8LVPFM
Kypf9QSo9Y3abb2kydxIRXY0SAzHJuzsQJKkqvf6cQierb3kvsTfpzrCBgK49SX/JiOJ2vvbCS4D
W56+9VYl3/XD4dceGWtcBHX6AGI3o8TNK6NTFilnSgJWzKW8XP8qJ63ivExTn0trNQQKroacUpN+
0ON6v3Kw91Ss+56Ud1qHaFirnlngRwMei9M078Zs2Or2OHPHrkH+A/Ork8hXVtzIkj7KFAwn0pJG
l0qIFsO19z0d1YgVeWSIJyyjsY06xFhjesRjBXhfsEfshm9wtx9VeSGQ4nJg4182oGonDwwYK02Y
g2pN6Cl/EoBAyo6ZPzNQ+gl8CfTgOulMpP17beB7lUTb5vecBRTqW+Coa1B8RSgoQHRG3PELeFzv
Eyb+ba6kDgq4OzGT1teJcZh2uykFLfG+q2vYXEMSAEqzomE6E/u4Zx1jBEsZUOg/JHg+bjt+Oa7v
Qk1eCMm4PxLLCyuavzcEnlfJbp5B90DKH5nvF+O0uJBqdhT0WAQYV0+xBdQxYx91Fgva976c4l4+
XB6lGOOuHyb+SUFHPGYd6Ho0cHKA80MjqsAK87xPlHQkVjY5nPgT+ZRZ3y8gqZGqxZoyiCR1X7RY
pp6qxUYzU5BU0oXNoc2wU2H0zxJf9KOhLzAC/PMY//wbwu7Wjgafia9TN8su/N2LG1ho0uxGzHAt
K2rbC4hH2/nTp6nxaFQr6oB5ouOuqVYcNVOBKy0HZpa3ddA3YrzQgC1Sx75KlajwwNbRQgyghX2N
Hfp7DCRWamY2y/y0Ve5nOOwfS9RpS6kszIA23iTJd3XQWqNf8HNP3Q5LoIu51bOWHu/rnva3NCcL
PNB+9RUnvi7URm6ktTTX/wr0EVABEAooK4KeQT7J+LtVdKP5RQKfObO+0c83CJ6L6/uH43sHnW6W
wlvFz/PUErZ0r2kjAKJu5BBl6xbo7frmiHx5uojSM+PCmtYhhwew12Z413J79c8wRjIpZGueovbH
Z/CJwXXNEl0aNd78BSCJLpMLg6QfudxAgK/0YtDZEE8fUu3ZI/HsUZMy2Pz+YDrLj+qb04cykvWa
KU5oEpGtKHcS+OMjusVRyWKAErFPWMR86XcPdDtvjojZdQ4I+KxSQit3aCubK8P7a8Vw9eZDBnSX
TcbHskJxX+wB61KCUDFt4h1OFHFwwxpfNsCVG1oo47YHZUA4dvN9vwEl1VxBf1mEAk08Dg1DMoJP
sOvdb2A3VndY7KtpI9alYbjwyKDYfFBP6FP6f9fTfSHa/zwthLtXErbCPhM3I/TsZKAbOdsU/7Sj
wwglG58lN5eRWYP4GmKq7fURB7wWWq2dOu9JDAZ7TizxTTdy7Ilm+C4aXAsuR0hD9gaOyYkmh8Bi
OJ1OTDOT9fiZuI4y4cdRr4g0Xq9H/Kuyzrsc8NSxph4oFxAmvfknA7vpGhlLOWZZUqEbrSI5/+Ei
fqypiuMmqWKbAtu5TJSyCH5iCH36FvKkVBQbaz7pZlXdIgiaqIkbhNwJp7+zG2DvdNEv/0UMaMQn
TIrqggWdE/1wz6Z2FC+cGXKqDE5em0sqxHy/lr+DEabtRDtfn6U0mx/ePT2VF/qr5+V2jGgC5xbC
NWkrkkujMZUFYZjQhwrtwpytQLXsl4joqjQ/pPAKvmBah+t+7U/TjeffrwRJ4kNvJe2Kz64toYNb
bl/YvA1i3XHx/5Y2/k2rB2HN4TW0gWo+WuiVJYufd4pJpH1Tbp6KfWgPc4LKUjm11qC/ysG57Tdq
5+CcZ0PRzsG20tIm0iicQgq8eKWsT1iD8J47AwMhw1Xoun7IQNqZ40limqUQviZkgIynohuheTcl
oZ6LZXhaFEmqIBnotURPw4yGE79OFgogLTjuA98IcT+xSzCi+GIgW1jjCJLPevXCKe0pVvTaqXpy
BC6ScSlvYLLG4AllHG1pwXyxkt/8xsEoZZba6MyEwEA6MCj/zJjn0TGHcEryHmuKX53zezj9m5mp
w1n/z7lTh5so76Z++UWGmXPs4bI61d2pvSTe7eTyXKqmBubl1/yTWzpBHpFLXmaWkHjdLdXlyVUg
WXPDKqs+LDpjk30oZQ8gldBik7R3MbEocAatZgkEmXAyFiWYORI0rGhZ4sMNj/I7MdsXZKhzNIPO
B7qL4Ws436ENB1QZXQI62vGt0qGszxFnQ7YoyVpegTkSNMdyQfoi8B3+dlrtBBAnfmQb1RyH9KFs
GsQwk3OcFICZd/TUJLRsI9u8HsBRrmMY97lxxnKy/kUFmnxG73sxppBq1LhmZDIsZexPKPfdLxTM
8cNJhaJnGOLdMZsrifkq+i4Kk/whhNhMG+JJvc7AVzCHSYc2m9kRUEzq8WQpHJEhsUf/vuNsgWfB
0fWDtsiXYgGmjRQJE5NjuceWaD9iTwN1y/EkkNTJxMe/BpNp8IUUOQiq3G+bYZgRXKXUrkPlxiIq
n7IQNWb+PMjNERoGBhyZ+MTK+IW8xXZua3uwqMA/MI5uypc+BJ3PpboZIN4xdTyit5bOSYBDlYND
2261VfTmp/zGD3DcYVxHayWwZ3eQSiSRl0+kYk02yfqEoycEvVDYm97cTEZRaRiRHtTq5LD2ny0f
bnx0MXZikga2rlnRazq6iCEegd+umYQXmP5mxw1uON3OmE+oyE9zo5YEQVwbCqgRFQuq9bEfLN13
mID6NIeSNkpymc50V89bA1umOth92cOThgZNkWt+RM7ghSmb/S3kEJvVEYv+h+f+dB85sQ9iVQlL
lmzqFXnQJelZ+5/NmCZCt6Z+aJxj1/c5beXIn0X1ovUZFq/YT+MAOcdnoLyOU0uR42XcSQHvn86m
0E1SzEYMz8CWVSjv6odENo7j40wufoFg/7C7kdUHMvc1+hXy589MNp6ZaNfMK7eB9m1l5l6+8MRK
G/jOLHZAHjncWQHguLJs0c4fB8k+WEwSQ3pJpKkerlaOsyb0uIvezlcQW0PA4qjKPO7ZqNRHprkC
p6EfdmCe7ht1WYnl0+PbleQ82tdNe3N8dGm5tyfjXcAhQeNPYymKXlIdaCoM1W8/u3yKnHsaKRKs
lSNr0Rx9hX6Z7hjgkwI882iQSUu9G3NnNG8ANJDOk/a8uh5t2nHO6JWrJ/eZ1juBV9SdIT+IzLyf
G+Fhq+HDQ4SiZdFz945drNySMd04eekIwhBJ63GQi3EwzUDIo0DlP4PNkhinKp2PZN9OCzPBGwvC
p+yy5JuUn/MpNd0j8lcDo4Zw10JFrSevVklpN+FRU/8NmSMc1WbCjYkX6PWShLuP6t3L83h41tWz
V59VoVIUTZ8JJXPp57A1td1pQZwP1weGFKBk/2AqJYyQ3tzDEB7DzXD2XW+fy6hD4chvq5iWpBhf
OT78LEVImiNMD77RJMlD4pvQETw72aYNocVQ3Zyamn9DQxIckYNRZ/J+fOknKn8OXgcRV6GgLLFf
RtAM9aPk6Ygl086X6N9JPtpDos0xRULsFXeT4AVSMIWv683lMmEgZlckzIwuJqCpmiQXGfnhLJ/B
ATmX3BH5HchmYB7P8ZwSdhjfUG0C7jO5KxcAiE9y+/UEuOsYb1ji6eKTkoa/qIBz6aX0j2FVyyHb
HWuVCGTEs8UZWyo81x8psvtMo81GsKaXTyRJa2Iyjk4rs1Y3ktLMKAP+piL13X1UpriBHQg/c9ab
ZLlmHkoiw7OkEFrWkdTdp67mbnvwplSwVFGnWBLKXvcXrDxzG4Eym6RXtW8GcIEQqZ3cE7cL5bQ2
riAdRMGCZrMZxMz9w/2purupffqsgEwypFdY/Hl6ofpcNJY4ioA86yR0lq/i3nZjNdc2ZXKLuGPS
FhO7iGfrSRD5o1eioSYw1g1bch2y0W2Yu4IoEWW1xCJQDVoohJqKipc00vmzGkM9ulMcbrsXxIWl
GJHv697Ssg9vYCUwchakVYkTISOmF6f2bk5JgeIoUMEzIKTvkEwKUeoIRwFSG0Kmg9h0Z0rYS5v6
p2qf5yzLf2whrNh9JlscY2N9lpAcoJeLiacniFodSYqUYLFXImNhFCR/21rTCFOyCHrWUN9+NE16
iYKZWRETMw54h/RLKEJlaJE6HLjzkyTbodMToHMmvCa3+C9qzHrrx4VZNH5FPnG+DqU73h5T/+1A
PpQzYgcKrsLf0GfBJY2ZlOy9AweFaUznma6midIVuCnFe0tjTE/2fIaI2uDxt0sPGWcyDfLEpyMu
HNUbUQ7epf3HN81rOLkoOPSsc6QxSXuuqLzp2vqxbGKqxvRykpafWOHkqlhXOYKBQbn2MbFktDw5
yVb+hvtT+bGAP8cmWorm+0ktDQecViZJLaEB4Fok7r7xEEvbTCOfEf6kKS9yANnw7IY2H2Hxa/ql
+pxpAUaiZW4NlPXiF/v6kEprb/d9GJDgqbM5X34yLt5DG9M5yBpGO0AR/lx4Z6aGnnBFdTTgZGoz
jya0iVnzq3gHjIUzz2LiL9+pWU7GdPz4Omj5DTuavV8cLJUPiQqnNMDLCyZO9mwbjOVnCFLYGrmN
81oKiTnmOI2NY5C38PLSSsa88WizCE2K0Rx/zb4qvnHuto9qpVjP50n/OEXUNC0JyluTKtrsWKb3
ieRcx0VDjsH1dBdrJR7hqCECwN4TaUW8HYI+WlhRUI1fsdp2l/qv44QQhaSbWLShYMgcYRX6Uzb1
UDhFF8KJs1Cf5Efnre4G5erwByMJcrcKQi0QW/3Cq6RzgMcW8rRrowkPhffuCMC8ScVWdz/wsuUM
eW8jYrAQnJyAEEp/Z9cdBHM/10I0mLL4UX0t19heC1yMhDY9PItUAf1HWx09bFQKVCGdnCIRLp3W
dzeXMN9ZQXJAmTpNZZBKvTGhEtgbTV/SjWIMHtUk3mqUxwU1GrlV7m0Tpt51hq5WU3IV4gQi3/hG
kL85P+VkNm5D8C09wuEdv/f9GBvBuHeIcwdRNDg44/0kMbqUpJq2bcQMPD0lYn0cbfhGR9BgYoeB
0AuFiCqhLdm94gPGepwQAY6WctyHCAoY3ku2y0c7X2OfdTWeykXTZhrewIVmEb7ASwE232U7nsC4
9TzBGs1xaWWsE0oZ3JiQvIYF/jnJDtHmzxSCUau9POh0zoOGJXHRo/fjghB5hxXR2qhkGjyVfviu
PSUqpudtTuDmTSbV1bb0QCJAPlbunXe+jImCXUf8z3L/qI0VBywycYCzneTp9KPCsYodVAOemC1W
PyIPj8DW6E0EdG1rb6icNZOsa5iTdGT2UjPcwmV+brYQLOamWOTkUFw7dBuX11094nd7sK/IQfaZ
34tPdxW6dNLbs61yf2BY6+y0lNAsmI0LO66z98b53cz/rjodz4tsxiMebwcUxS36stYeHcXhgMcS
aoxSdkCG5Mqh7bjpAQ2VbgI4+w/jG/S9NfqxIlTZliAKl4cKErNOj+GaOG2T3VPuBOZ24hxKjDyS
ljtoubtfB8saqOMUSNaR4DjkHaMtaGqScGCnP31mTFGfDGzZH3XcpZqg8jiRIXRZyvsnvvhH6sNH
qd1tlZ4Gxk7QcDJ4JJ2+cz1oRwW2XiL1/pa2dfRQIO4gmUcsqgP5Uh/yhTMr6NmDS88syKV3bLA0
OBB8XjA4bAaieTzprfsIASPkcXlItgEvm4IYfTjn7SLfCRDlSuHbe/ivTE8NlemVc4FtprHND9x0
JCxnGo8+TeJuzGUfMh4WWBI12uhirhIttCx+j714uW8vLbZKY1vJzJ8O9/+tK0IErc5QfXl0ZLAb
kjFkiztB0w+l2FCRA4+h7SdBCglANhMfMQeDMUN957d9B+H6wpZQemKwaNpatb+dfq0D0jvIY9/i
vDJQRnLMLL2nlASqhIRD14Qi2iQlnvug0EqKDVz/qVX+8rNZHguvwjb+AgMt3Avi+1gSHCdFjUSB
S4zUEXAm25oef2schjYeMISjnMChrwSbjug7zk60BBl3JEjQes/eKwD8vh9r2dz0vmkfSvGxF027
d1hOnbG7HmdfOCdIly9IPJHft4d3UaB63ciiJ2Vrn/Giwkaep58A5rpbNIurSwViuOKMvgOuGXNK
SaOE/zZc1AaekBiKHOxQfEw0eWusod+I46KGbXG75umpOqHYdEGBhJvLXLC2N0QJU9pp3asy+S32
SY5ptdS/Uf3z9Nhg2Bo7t4WeAxSpQFRhCrKcexcYyVPqtHtFcnDNqKcSr6X0Cp9cd0uunt1YQdVO
s1sqP2qV9o3Rq9ReX1L8tALRulbXpSADa3kLUFAQxPJfylpJEqztHUbkBHcAxhVPiQ0ehOOnXfcI
kQ+MGEPdsy3jHmqBQZX5jPX0xV3v+BtuFMz4fWw9MzM74d1wv1mX0NY1jc9bs1QIhqMiBtnb6ooE
JES4oKw0SNEy+/yvv4ej2j40rFZZprtn1zehR2rembzDY6yBga3RIQEk1L3PkkySrhRObeiQj/Mc
hIvHp53AVIX3HCcmesP8GsB9XWzR6dlJsCe+xZnzDOuUIqPE6Az8+dTNj5RbIo2kvlBUNCXWVQf6
Jfj+apJ9R/HOGgeleE3dxvFc+KMdkTl+QmNIBDt3GjUwOx7gYxIfkMedpcHUbdPS7QhX4wwHjRWr
5Mn8vBcwS+Nz7NS6u/biKg+Nb1vVmEY8aTIIhy/zEVhjp0M0twMkMvxXQTkgtC0Qic9+T2akoR7Q
qIOmBi/fPYBLq6tE4DXi5iAjxkDgKMrHaA//dmZryCi+kFLj8nSUWiNAPdAFDZI0KOayYW1HgEjN
KQ/vhhL4nAChhCdIGg+XY8kC2CwY9W8mLWIx0NoV9ZjSPKbE2N9bAjeEi9S6H7aAl2/sKyKFK+bP
rb8/6HT1P7qloPf6nyLHjYsSNx8qD+/clTN5ylVzalmQNl+1hIbZT4GRZWtIEYg/wsVu7GLFc2cZ
TEKpEUrsXc4mc7f3xX79ZZfi4CXIfMUbksNoTYLyWBKi25Ooh0GLNcXUGZi5KAMyv+I4pPZee6EH
bGKAVA1UoKCT1VaVZLrOLP492S4wIgxG1D1KHcTWz5dl3bCWeY+IuSMcS9pmWSIm+NTyX0UeD3LO
ZSF71SqVgawGh7EkEUNgILUeU2m7rbSchxBYcdrhqiWto61Jm8WTK2Ay9c9deaZzed8NltZmu6+H
nM4OMlFMiElP6827myrhWEDlHcp5rb1oV98dAwqnB5EtiKoEm36KqcBXk9Qkd3aU9UXR+ssqYm7Z
bN5bmOdCSEXtvsJhDX1I9xN2AIjWxynRa5xvF0YQdvvt0rf60q23o0tnJjzYFgaJPXX28L8Bo7wt
htBo1fRJjQ/U1XaY20w741jmAcIXS9of+nEsg6sUOdckFQOfDNW3+R7uKwQzbG6jzDAQfzq0lXKM
z8FjWtCG+/GHA+fbCUZ32m09OCdB0OEz5X1sM1MyUhVOxKEQlFNohIQ6YpiOyC+xqwRxa33Y77Um
fiN/3pJaiGdGhN69GrMVd+aHMVMidsgDEN/w+ZzizlCx5J14LiaurN5f4p1apWVGA70+aQAvPQnL
i1zYnBA54Arl2eF0LQrEgQnjQHN4oLTUse2eheisCtP2SSbMkPUSCT35iPQ+0zb7JQQoCYSnlq5P
6d5OYWzNpcOzHxYzG9upjOKLLbAGdgK1/B22pYmFCS9M/yUo4w3Lr5H6bf78crN0Qv38b58Eqm+P
7ZK+3oiU0db/QxZ5w1chU6cxdK7IrvNMXKxUkC7YsYeh8N186a4C0bbANQyKhWw8MFnHkSTqxJM2
TUuBgAqJJ0A+1ldeTF5CZFFRSceNhZQA/Q/I96s7yWE6246fxrhtCa1IteBn7Xpuw2Ie1l6luQ0y
9Ok2iBYD+8NttV/8KhnMh34P1ZOVn4uVTNCwKkEXrFHo1/pcyJBtKJGGSxZ3LUgZSinU/1OE9V9a
NQ8cmVqcUwshX+yQytfpd+wcOg8UegnTmbfflbTCF3SnXb3TAU34dZ5N5ga+1B/56F9ggokR6I8B
yvzJMYqnWqNO6+VFdr1yQjR2u9OGZUV6NbyuIhTc/A0U/AqhlgatjP/c3XqDJ5pnJ51yJeeVxY3x
wp+l0wjkZSriL8IgICl3tLBJAfMp61gyjT5M1XISCliYrg8+vZSYH1+qm27M/XH2XsnMYJDXD2AB
Z/LH0e7LsAt0Q5yRsVfoQVrUXnajrVPe6mm1DgQMSKSb6QEsMyKG6wNpWXjItG6WeC/SHsNpaDcu
jowSdOof8iqhLVOsFTu5NaC62cLYRuwROCrpmtVoUGkcpEccZn97XKfMiVWpq4/EXAyz92nlBwmK
VTMiwa+MGAXqbyM7EuHkJ6/EsmExGo1eKbd28mEbFaOH2rm6cRJqxAiJdTxwGssomzVhZNfeH8m9
4h4db+AKS/Rcvaxs+VDoG1vyOJTdS4gucwpDNFM+R44NLugy/HKpCwld/GJjY4XvWQxGyJGBW7hl
PvMnqb8FzcYscWbzW4IIUbQ1S1nBIhv/mbgwX4goSTe/XuDEiwTXWHTRLX4phxqZNUa0b4PSvDoG
d4K/j7sabheCdNwJzSpL6ApNfvSJ39+zuPlrGbFDvEZ8aQ6EduImpJsYHUgjEnV0mprQKMUVc0a6
7Cc1oC9zMI4UnhWbu5Kt4cisjdOYsv0QJXttQAk5gN9Tyk7WGTU3SUcHAwh4cph7NE5uOabgRB3x
LuWinFK59WzUVwv4X04TXNoY36NDdi+jTIvbN4VJYRDAvEL54nYd/uv4mjZVUsfI4MkD+ztb1Frl
RbdQn5nlsLrAH9zjmy922kpRUQHlYdouvC/w8HKOgyV1bzjhDljLtKetijBcx96r64uXl2i67K6O
vDhpwjuMYPPzaIaaVWQ1x/NlPhWE3xnifJmG9dDLOo/XwUJi2Dd+wXyyI3qEJ9LCD1dX0pi5sdxa
+DDHrGzIhs5kaVMB8HOUOocohQFc3TvtD/96ifzsFpOQRjOytMuf4kfO5XUEz70hiNbZ1BmrHHxm
b2ilmvmu2Hac9rZYva3e4R4wmdRrxoY6NCpGxPhBEP7sKF5B0FS2dcdxgrqOSST2Ry/rBxS0yn49
z6XsNxIA7ouOkpXl5IxsfKNfGj2KGRl17Hv5kI3wFmAtJdZiouxbfZhNOPmPncxEaS+7YsyvdYDc
sb/LWn3nX5CHuOQk3ERj0b48YqIRdJQ1dMi5bO4vuVWse0WSE3hJD/l9kcdMvJgDtuhIBpbBl4uE
FtvYTyuvIypQIsfh9mtJ8VTU6svow3/xo4Th3oSsUka+rZROnG1a3HVmE26xaYJ/5gebLgplVsGz
Qa+8N5MWdVgEewm8064MhbXTwu/dQpBCpDF4obJwgx3NdpWOnvuU9JIyidTFmfR2Y5yG4zujKgQn
rImcPMxfbq13bqKw3/aMSnwJ3YT8Ixdv3vO1X1+p1hC+BUXf0ZfbiOrUtYsHtDKF9sWYKcJpgqNQ
5ijNNnunGtzm13KxbRGzcKdJSJV4ozaryrB6KixH0z6zITiQxVk7cEmCmI893WmMhIoWOGLbvlEH
Y55WdHWPmDqxUWmEXZRKoLhAxuAPQQVzn6EVJAG6daAv6jmUcYWcIsS9UoArpexIEy1f9QgwDV4M
tKjgCuvLlg27l68cp0lduLIz3tPbBi1WUeqAMWPU4xu0ynF+8jC3wQFuqnWAWzU7exHXHEOSieTC
zo3LeOMgIdPUxmPwUi7ly23fyvELupggNxb/sWrGTbJ7zmXO8JIE132si0ksQzoNMTyR1muhVVH9
laSw3F92aJ5jKxMMqwJnF9Lnki0+BJ4GL1lYGGvfVaXyMTcKNLvJ1JUghRVtHl7eU2+RmFtzV7aJ
EG9QI12ECpK4tDx5FN7b88GC2buNez1ZEP5e0kNdrXT8Fhje2l2VjBXJ4gc0usMLME9oU2a5z9Rx
BIUDDEMq7/3B7r3kIuHgWGvKtxjJ6RisdoBF2bEDbyB2q+feGocVjD8aZqaYYJAIJuwiW2JPCx/g
KrnkwkjGDDDO5KZC5H3ti2GZt3UnbeResNDODpzDtKt4rZYYKYvKakW1zmg5hrxkP5fjGDQoSdZb
ftCmdQRS7e7vbrOi+X6bn0pr4M/k1DLKC5Mchzwh0Iqu7fhNDZg9UHVP7pfgj/jxNfovQ6gm0ncS
LtrwYOoObjSHbf8/aEhhEFJtvdVUHo7GroZ8yzgurWlGZLpdJc1QdDWf1j71b37eRsaYEORKvYPV
JsQO2R9pizwy+BvMHpFFCm47rGl7lQw+ag2Meip4VcNjMn3RLfCDHTpDzgVizGp6SVD6GNcd4qZs
AeIJDFoUr/vTk0Mh8cTSmvAMKHv5TDnnQZKLNrYKnwX+htDwrATlhF6uXPVuWx90L20tDVFbL4rX
I/sfmqQMQuH3/JaAgZW+l4DMW2BJuWT82dCj6YytwyPt9oMJxiwRMzlzVAR4lNvWYO3qQk/x+cs0
WhDZ9fFhE/EaEN9nyVlQmTOwMTfjeCMfusAN8zciqC96a0hP3QBMMxIczCkilSYRO9VzWqr936Po
psZJ0JCjHbBBnHHtBWYzA1XEYzODvBoovqUKoRXlUVJnyVn38F7igBCp8TE8Fsm/7zmOdcmXLUXH
PwzbsgE/9g8gNfP5EW6Vouzj4QBqAwRdX7nJp5WvvW6BK9B9jDe2+xjxuc4Fr+IMiiFfVgBrvE6l
QLtc+LcZx1nsKKe7Ax1opEOlS7Hmdzi+glBFT+fiWciOe36qpehEXD9K2rrrv5lInughM73p980M
aLkUY5A7EeYzs1GexVmt8sucKQPkLLZDd6DHEfn26vCwhEFJjogzxqTbSZfa1PJe9Ica7Vx5oa3+
7ZV23Y8ZjiFfCKMrY67AmWvT53DbHQsmJuXWNV6c2TfR+3ZxU6cDDbKr16KdQ88MZdVQYLzJgbLg
6OlppUsAhSQo9c55VRmfi+8TKCAkk0akY8kIlaoPw8+q2fLgn6oxol1vnVdU4eTVzhwiCZmj8ekJ
bwHk0vfRorkgiofm+LbdzlXXm2QRPkbCB12N+jv6zpN1XXtqm/Ztp+W/kKq05A66YtbQHsQD/zkf
gf37BirFkGvCrF8hiyijqGztgRQQ+dDxL0rwygBOJlNvqOs38H/3F7H5tqwnJntkoyMVpCkvYo+a
jBUyMpQs9UPTnY8GErMqVjmJzNxFrzJJTEbByBYWBabDkJTOPFln01M4PmRM8hZbm5NPORMEXeb5
uZGRAW8bqt1FC6fvItY93kEzG60BUXqgTUO9tr+cobAR0HTuVt677To9lZcfGuHSweMDb+RGlYAF
ndcLugAL5u36WchdgE/HE+z7YPEVOxROqgI0vXJ2XKVgAXblczk+393I2UCTgm5AWHbHO8lRO/9w
PAeNxq7GykLQjYCUniQ4CYSbnpNSPuepO3zvRCI/K+znd2MoH6sY9RdEi8PUEY9KgqbtBtvz4ZBY
/4UDLih3KOkSOp3U1DpNAXvX+ivbiVy0/QrHqjd1K6n9avdfrhvfuVgr46EOQemnxz4my3ryHQTh
UTP/bKW/QZ9mTskIVMZvPE7cNjUuPQOtk2wyltzVZ/WrkEhLrSFvcpW7t+s8tgTsqy2sv85Pr3cW
/pWDcltRhdPoKkFOIU6xf+piSW1Ov6wurdu8xCZKw/D/bZiHfoi7IL+AkCVksT1kTNzSwj+VdQ6v
APtUt2pRlsv705cJ8kTBZsTD3Z1RNptoZdcbsjkN20CpT1nI90hkR7JPt7Y7qg1WDz1gpdVCyIjH
gj2x1QE9QYdRF3k7bW5HZnd7tBpI+Gr+Uzds/wiY/jTb/xtyp+9GPFeis7OQuKUIum9f2REJJg1C
mtWFPXHikemn5GVgfEdOfoX3ZUbjAZB4mSIq4pRjUeGAWzADc9Q0on0cDivYZmlPY3FpxXWmo9x/
sPLp1N6Ht23NCPGO4kFw+CK6ZKoiM365BIfzQLHXFc/vFnrh4Xtssm//vWDA/FEiIJTf+S9b4ylR
pTjH4RGOO7j0NrvXe5m3r26GJRESbCymyJGKctdUdyHsVjwhAu6EkNMBx5GpqIFFBiIpSmkMFEwJ
R/EFCsCXynG2szt5FJpDFfIHcbAIh/K5WuRUbwBi/p0JIm6hPcOtOtISTA6N8TZzaNo/UtH0hJFt
mRHz2M5AcOakIGLVx3TucSpsWAsQ9ea/aC9UDZ3nFdTV8ATSOboGr+bpxJ1nuYWe2ve4EEJ2GHZw
+prl2OX0TZ1tvA7yg0JvWorGwkwcIDlKzONwa/6aOLqj5wkh2Lmn/i/16r+ODWklyV3wUedKf8EV
7mvjkXXwm1+EKVx2n3LElesN1mtbteDhdei9V3XYSuiDJdWM3vGEmj022zfWA90BMt1loAoFvyFI
NLJY53OXqXHmK2tZJ1f3NfgbsEzK00Mnzg12b/srWNTo3pPe3scxgHzs0dL0P92USAONRZN8i/4G
b5ZUToNxIELPJ+6DxFu8/oEFJdTiScQzC99DzdIYoIrwOuJnEKuMZ8Kq4UaQaqOk0ojhTm3c4y0A
dh/AtpgfB5gdDHULNHyV29Ut6JzVq8y2/f9EAIA3UcVCIso4isyhFCO0prCtn1W9cao0Quk8J8RY
KM9wwg3UeywUQmIdg49eP4h2qtDIFxQqQHdCWlLyjN8ciz6jdvaNycLLSuth5cW4xMdmnmjvb9/v
4jza0N6/1iBITAQ7b4tuw96x7nmu0ZuB2boVQ6eOU3lRWPzvYoUpl9XHXQK7dpdTUVgBRvFBmWZE
lCKhWS20JiSeB9fs3mr5lebnpmx5OrTlzyEzrQSeTssyGkhMugk5NwyDrM/VbcIPCoRTJd1p3+ZA
UiH+rHkNvBSmpRHujE4qrH3FfpmSOh6wbiGpB7cYmHiXYyXx1YBpHpjhN74q0clL+1T39hHLH58g
nsnotK+nlp3oiLjmpUh4fobFz4IMtiazwiUK/R+btkdtXM1E/lstfRZI48buTTK9d4r8v9L3wyb+
u5eoNKDow/cXExzynq/owJhIc++u9KgPL/tiGDWT8K3ceVc92XELd5/ALIvBt1MKANtOtnLMtAQI
Ij6AIYVoq4raU4CZKfq0ZNtrqExh9hL1pqU3Ybr+YDWLUC7lzdSy+xfp2QyQTo/UoMi+Bid4SEx3
GCDmi5nVMQbQglTrBbMIaAEeA4UzLFOuTdUQ3HQF3U7BG3rG8qeEbYHSr8njMa9uTx0Ukw9sIFoH
6KxXmqmIITtkp7Ry9BeULI2uGaYSw6IZTaKDJg5YLeihhLKgFJD/PXg7EyYOUTfvpsDNbDUR82ki
MNLuMVvkN/0ANEpMa9PLFdk3po9euiay/LBJuhFCDu6efL+sluSgiEn9l2/Tge1ZBSHCMxcZHbhF
nkxvi3SYBfoTvU8qr1QL73TOcvnrJ8LL7EBSZtx4PfzbTN0m/vSCUA/LghiYzoHGTN6CaMuwjtGg
RI1Dj72Lar8IvMoeNFry6qYw8RsWcYFqFqqFjnWPNDJLH9SmPp96jP6tbbTtJeTXeWIZX9zPquK+
MutZ5ACsQmGpd4GJfizVs2z3RcK/9HqGtD6QC65QaIwAQ+LozqEJAMj0lkPfh4gqeZYjEpMEC0dZ
zEcvDww+H1Lb0dQZANs/0sd0LnKahOw4ppyZ0LS3gFsNnhv3hv5yUDNAe7O9iLyhthyMaOwYiUI4
i8j30GiL1txFMHAUxyvJ0H+sTDBA/bnitIp4irGSTFExRKMPFFEQJLyxmEhoIOdtQhTGIj0Pg9oi
PSpyFzgQHtxnu9PkgAiSbB5lLXmBnetkm2q0jxj6DgOAXN0xcy2X3/YxewPTEyX+6oxAAHXGwIcT
c6n3KYiCJQHPI7u2uyEdY8g2N07CM/RsYiaYijRmSQSRDNpNr1ncR5HckhCHgRZUR33J9BbebqRH
wfReB00tf6euLBI/8cG3Oee3CUP9EQ2WZf8VmOOUOC1auAAU2lGgGKeHxLyYpzvE0vaCQRAAKiSk
XxvTlMYA29CdWX9V4yDF/FuM/T/yVfoTjEYyB1Hf41Xr3sVxVUoZD0ILJSeb90X4tiOtvAkZtVgh
uspat9IDFY42pDfI4w4mAEs79kmXD40G7eUqQsnFx+zejy4e+ITz/wo9OmpHGCq3tBYebAwiNIPf
1tK4PQUSCFhezB0SKchDn0q0rK4+oKn85fS7s1Nf4ev025Dia+y7u/DSNpYXGdbWjx1IxjEdq3fZ
WPh4yw+ph2d3BaVDOp079M003862rDWiWCpb/isc9jPqjWehGDaSfjFRNpf3SBheokOfbcQ7AxE/
ZY1VoLzZjrmHrsd7c4U2RtkcaeL94cfAYSQwHWIt52hbaWiN7k8P7tD/CYwJ+RZfMOin7fE/X+95
P81qQg4Lb6IfK7CMIfgEkfsaA3myUclQXZR+H0btG7M4zZwYmmjzoXq5474hvQKDMK+IhLUYH8FJ
VF6pH05SRM3HtK4JSCtCenl5Z9tx6JYWuAvVYVtnenDfRkxZr5g12K0Wy8AdA5cGvyRodC9AO+qT
aCUHouRODXCxg79I3fkVSClymMNS508e6dJDYC4/9v2eRvGqfZ2JM3W9ALRsKkJu4Xsetoph9WXe
uilVkxR4G9Ejz7BxRynA4ByUxCWVdpJa+OsH/8oay0qGtZunKPTu3t67eWQ0+siqjHadsCFtpLnN
4m191W4LEBXXasZTfsIPmUjFxAIEF8xEVQmC2uS15cOWW4XuViVtL+3hKE5qJbejNmq9wn2sbYLu
RA7HcdjNNpyCjeuG0jtcHRwuBdSi79KVLKCvVZZ186TYq/lGLCde8Yj6I6ph8BDRenSmvzxkuekN
NHf0zWM9iNyxqbwukPQ+3qYKeKpVbjKciQNPtJr729ExSCI92KKyXT0+5KJAENi9pRCOlN+BMJNH
Z5C0TyLRimfC51RTgqKgvb0Gh5o0ENn3O23K1496nPTfW6cp3UwjvtJwfcr2eB+fkVbAf8y2y9zm
VVfdJgCds2O7VKDildBN+b7sJZzzhkYUpeAUNM4UT0MnrYEb7SFcxBngxiS3juYJht8oDq+hbT2z
XoLLcWjIBus1QgHd3zLtfxPPDaFrYVSd1ZlNoEdo0z0TMvBAfdsaPmkeQBeytXElTPNzkbohOkUV
PGgcWBpYQDzAuwVfUhNagVBqa9DN20tSPxZxMrrqX+nXLx6Kid/cY+uG5Ar/GIAlUvTEO5+Bl7CC
jwcTfmLy4CSIbR0AW2YruF6RNjHjDjHneIEaWS9IRpDr+/FScw+fbdrO6Dzp9kA7e5GBtepd4oHH
UHNzI1SBvlREaGRn19Rjp02WZ+62EB1e87XtTPN7oZ1Mvy9lCSodtLSN9nQIL53r3KxcvDNP53eN
/V3aHEYSTtWByOvzgdX3XN0nYWqWK2oxesT4FSrqHBzgQ7wJAhAm3hIl+vYJ/SXwyxyNdTW6gPUq
UkPhNgTzhWGN8P6Y3bOnvYU8+4joAgaCzT7ap0FBEtgwQGepqS/zfoMdohcuvkAMTLIfqMzdKgro
9F/s0Rvgui266IxbeNMF3ipoTq2xRJliwnbPO7KP+6eeb8H1FRggmk1ulbjqlFqUqPOoR/iMSRLd
bvqfVbgX9O+MqfS7Q4l3inZbr61+samQNBFrJ2I3Ha8g/4Lgj+7qQjXZLuc/jvvUcTYiaKi0CuSg
fByBQv3H9i0DIsYFlQNgnASaGD8n52H1y929spwVC6kLHb0PEFUgeTLW+rru2Q+8b3Fl7l/R4+1c
eshJRCGgojtCuiYT/qh7pyiOSj+uy5tDLoe9awH/mQN2TcKpu+ck0FalrV+vgYDPAjM1l7DTH86Y
nOpZchEAD5h3h1yldQiCR5AzNaLf5O3x7memajc3qY2H4/tUCaK1vcaUlgpu5Bzxi4kxKdUq+3Ra
zgVEZ7sNQD7Pryfxwm/OSRVaLvxfy24DZOq4NwbDRw9/rHjyE5hZEQl/+mQABCJD4QPGuBaKM3bk
xADxinkPWpzuLCmv43kggIiU84GCmpNDRSbLc82Dn+mGjGPVluvX3HIDspNKTcpAyUyRgp7ecSr6
K+uHcA3vF3KDye7yVVH6qwp6LggJ2hYoMNvmPt8cTp+leqMBsgAoYTte5AV6Oov8by1q2yh2kbTD
5uovLZ/Vn3KK8oS6V0oGPt1NtfpI0mTHjmvxDz0lhHeRItAm5OozvAd5OU5Evsxp9YJcGHOeSv3A
yEhENcGwGPlB+pqAFsbjGssvG166pkPvhM3VFPEuu+3jS2BhwEQMeTTveC4sQ44uYZqqtqk5+aQI
e9xyHoOeAT9ZCLhR4wWdGmUKFP2GVxiHR45u6JVyo29jSTy3tSrczvFtDs1aVy8beQhCunTtdoz1
kKSfB+osyN0mnvHqHIpejDFuxmCY7raT/QgdNQliNvv6I38roB9PX/xwxsxSj722VnhShXuushL6
ZUJOEM0frgTwaswH6z578PhImWSFwx8ffDVErjXiLWHxXxzQmVg2+yaqmYlL83+vDBOniS93v1lh
AlZlG4bCvscJwqFXP9E37PdsCbOA+9rX5DVtTzWn3hyAxcofIp4UCVfW+csrGlk1qvxMtxCgtfOZ
MAW8ki0E9wjekgmlAAEvyQwqGps7DDMuFtNiDJukULr2rFilSc1KNK4ROvBPAPALGsH00g3rycI+
QX+Cl03AQv2vK6REaSU9aUIs5QbndWhe9mC0MPgr0ZwFRDYwV9gK8hX86MiaCaNSNXOPO+1xs4EK
edFp2zYT6bIecuocDruV0bZjKj/WpbW7GOl91rWPeU7d4SEHf/NFDONE627aHBIf2NUTx2AaGFzK
+DLmsxgwL/2x92GzcmVKrUMPupaS01skVKFjE6DO+qrMNEHlsjEvekiJZUCdGntlH5S1nOus3wlM
eceHqxXUoJfM9d74KshGWG6/rwJ5zarqPt2lqRDUrG8cZFzoScurWbaELKhSCnqqcSgcKJo4OjZ9
1qlemh5S99LiIhbn8Jb40YXBAudm/BlmRyaUAhrCm5+Pjqw6/ekr2EP2cBW0Zn4KLAvWnTjFuwog
pmmFSFjYJgGvh9xjla0J96wjwM3blWIpYE2ryMz3axYSkpFHnCYQ3vxb6+I14Rt7cnGfouEzufJf
nRF4qnmHvtMXDGqpMaCWgX9aRt0jY3St/00UwZ93E9cFdN1WnacFkk0FV0XOH2ze12D94Uoqb1QX
44XEjGfMjkDaCk4JgFQxuHJ1cszaOKkRv/krlgaGkGHr0lCc9Fke7fltUnXJaShFJwmRwXYHcm09
YeHjI3oPNOjTlprYTwsJJSGHCZidlY+y9f7xylfEKNeHQ1oqQ0iJ8xyU9uySyog7ISpUZHFRQ0zd
BeOsELBPku+7stYs7GK7HAC7anNH7xiieHVE1VanBXf//76zwT7bGwvSGcqyByLJzRh9Ln1n+AfP
X1Ik7NV7NugtjP6o6Z+zqXC5H8KB6hR/YPFPxBBHIa/mnJCbNx2m2eH5un9Eg7IvAwbJoBbvP8Sa
z9YwA/yM+0yzUFw+aac6059HhU5EtQPP6sXusPabhDTZnPTFdBmUT4ov8zSVke5L27b5/Vh+orSs
6jQk3rQcj/olT+eAibLDiEvGvYN98hukLRKJbdcc1z5RKaTMs2O63Y2yFGAL/0+VIFjbBAhGy+mY
qOLk5YJx94IETXgneOT19ZXdHwG10pUTVQ3il35aiA65T3pknui6xcQzXWcwY+LKMhl6zyfAHGb7
DGQ+1GGbo3EU+TdJv8NOk+5nmqyJzPvErm/gzWZWLWipGfC0bEZBd3zUUQ7SQO2J6/A4xpMs0lWT
mcjV8CvqEoWKuD78uYx6J7idSx/WAa73AYAEZPspBqatVFiavXSKf0ToL40Ryl84EQeQPIiKf+D4
jhes1CJAynhtNDCAcy7X+bKn5PtEiN86twOf6UgVq0DqUMUEXdvY1ONwVlhxC+duKuo4juGy4cFN
MgmvfAKUcnYEohbOcab+sDM2RQTTg3coqlbboRnQXV1I4tKVj/3sWl3/fPLX5Mw6N7qqRr6MGFWY
g3Ahwp5Do62jsEZCEEOjQ6HfQDuhejeoVYjMFM7Vj+/GQcJFePZr27WHtASYx7oXb7/HJlJpo4Zw
rM/sfA2UBBadnDBcfK6RUI4pO3VnZf2xjgLRQLUK5zK0uD7gc2V2lh5DYTToGgzLTvJhTrhUMkfd
mqhP8RPf3gG4X1sY+1YhwHKZUyf4tcik2LW+FBRAY4Iaf/ZA7WIssAItpYttMxqn3Wmc+FwHi0oV
95y65L4amGiKuyz4M6FOh4mEXtNwbioTLQt0wDfEXd7Muw1pP2KbGz9vKWEVEQ8mixIsmkz5ESAh
a6GaLpgtmDGx0YSFpb6Z6stvStUTTzjWiO3H36xqX28jOX+MRyB5VrK6/atXwr0FYGaroqbKHgtO
L6Im1CXIH2N45b/Zc8J3xXu214cVyu/+TfDwoOfKvU2UAEu/CIRrYmfUYfBqiqmoig68MmMJlS6J
B9pAYQhFangB11j/nhSf/EYPZPJeGqNKV+Db82oS2UA2uVzO/vOg1M5VGDVfCh7K9RoarZWquj8h
5wk9VxoFf4EX9wm6FqDpTKODuEmKUIZb9e21krW9k5hhOn3/OSpKU5eoucNNAmWk3RI2387bYILh
/QZWV5s5GEwyrvAjLdwA3dlF8lDazXYwbepOgh/Qk0s+4JPpc5zXQRQl0xXlkEplPrVSgdr6xgUs
Izz3Fixg4Agl2QOIBjeGy8Ln0Ux73fZIpspB5ojGNGzB89qxtmgUi3s/vh06pNlUxLCGp0KZsQ+A
tajuoXOmGopNUmPyzzzN9JFRny6IGmVj1KEStnTT8AEvHvcLvsTJbgnUq4CUbsrkyrK+ikea4u9P
8eXertIX+pVWBatZuDPU6iiv5B8ZZojm0QlN7Uy1+fA041FzA31lhp8YPufuOxtKgCtnHJpc52TP
me90J4+/s+X7YlOrrq0t1RWdUlLMGTr+XU1hFTVxBU2IzPdFCZ+7MFwnTwjo3P5MfmNcnM938QWF
us3CoDh5qRtDtNf5t077J3etYY3AvAigoD77dgYItS5sBcNJqQV8a7tqIYqdLlWeMd2JiIrxGa+7
D/GYOC6luHeqECe4b9HaDXbZGT0TMdXPt042UU+Ty1iYYP8lu/rBUcoGfAPCdmFvFNoKojtwIn+M
HfAOE9LJgoqTpvpvD0Rj0JsjypXXjOQ1csL08FqayvnhmFhzr/oFfBUvrGoibGmaYYRZIVX81nsf
7EOuX99RiIi5jiIH+xDcUxc4FrQTgP/pwlfDYbRaqs3lwlnjdSzy6pOlvcL6LjcXmSJfPn3zaKor
VL9G7twVntsWO5VxisoWEULR7321umm+7yuy4DbQoX288ai6ERV+7uoAzjxiYBRwSOqr8XYyObPR
AXLo2rDBotspk42iQMBBzgFbE9VBF57bfk88ZS3ztvE/JfNF5+aPqtKqdxrCK/CjgRx4BjvgyQw/
/NCAKlNYy7FKhgr/CSEkvky31BQCSMUg+4ND7hL1ZqT34KybZmlSzn+ud7z7OIaEeCzquUEQRuEa
k32jtS1FCVG00dLp6OxdCEK+y7PLWQ6Pv5a/lq80V1Wzzs8a9xz0KJ2Ytg7vrhvg/sklQs0utKou
3lkUfXkKVpQRWkhN3/y4DJP8eJA2Wr13RT6RYhbAJU+uIO4/N+cp7STxR+qsuZ2u8cP1YcLwzPaq
ABwi1hNJ3VhPxP4SRes4ZatCuD18HUkrLjcVcu+HGl3M/EcVLLbLEIMxptwUcByhH7n679X6aI6+
3bCU+rzzr/jc8Yt84590dNXuq3KJuOvtpWh43XEOSLJHRfC+NWWjEaXqAhdG84eCO/4jaX7m7xRV
ZvNtrLueB9YtFNgDguHv9Y8pcwD4Gl7c6vCWMpuUR19vhxsLaZKKDacPCspofiPEJyVLeWMk+VX7
+WwUamzVBMbNbuQkU57Cmy6RSJ1SAsr0sNSZgWfwD5xqm/nZ4EvVv+ytKPnibz2jl/Kj4tlsg5qe
BTzHYDdn0LRoxQbo6WlEHMpN0l7Ss1ojM9pJecy8xFdh15mp+F3fqJdDXkSaqgueJbPJ7baCd9bL
08jC+J+wtIbXmlJLwxwuRAtl01440WkvAMoDFrPMjUxQXQChOWuiwMj4eyNbtEc07FzxoC4nzw98
2tEPvaepiJyqCs6wJCdqeDoP0bSu6tlryVbMYbL/dJ7zgTp+0ze2PNHnxCRu88IJaf3riCYr83ZP
1AZhjItCCMb5lPx0y2bTk53wfvmfNyn9pQ1LxudmqcFFl7GmLzGaO9IQqN35gl7PpzWyLcugCn1N
LeBtM/by8Lj7kmY/fsIwuWS7EB8L+05fcm4GjJEQnQsJwE3iyS74x55Sm4NKcoVFg4u8xdAtXR91
m+7N51vt8Xz8E3VTq2UpcaiyDDY0Q3DSEcjL4u1dQe/f5QBmBHmuRx0LlWU9OHqIZm0HQhthLXPZ
h1JE3bZlf9a4fKm/vhpL0o5LaIHSfz47SYqw04DFHj2UtGdkKvpLd4HX6UUl4BjCOAFHD9CJ20//
jxmSErsxK0EW/UvEqbPic/MN+3XVT2YaS1qpsqJxQA8XPW97KQaaCy1MX0FitH52khDsloCyj6rs
YSeljKWAJlU6fwgRjiEAKoXFYggxBdVKoMoQszA2Sf/R6znA/IVO/YUg3ojAaHazwqpzgm5s/U/3
fQSTq1xwE7S97C6KQ1sQp9tIzaUyW9UdMWIbZZR6sIgJFq9c2A31pynq4TwMyM6bvcpkJTqHrHj3
KW2gmcNDbZfyWjgv0gudFwJT+cmVyMnXoHXGaHw/nPyp2VSnUcM+sItzWNOOTxSihO9g4yqeEQbh
RR9qx/FIUj7xbSYhHLRN4OlVksSxEqIo4gBwT65WKoisFXSB1lbNp4rARvYzJ4m61LGiUt4NNQxe
zlMlnNRj27+WUn4sGc9vKENiQ5tt+sVb9bDeLlBS293uze6vksIkKuQyN7LShBmCgz1o4GCuSger
YFMceI+BivJSmZXFPwfL8iyxDaui1C+G2YGEMwW1tTOVt/Aom3u4s1Df9Dc06Gs1hKEM+z1KCBRr
M1LZc5RXRbYC4hraMTYJ+ngdv8ng7e0f1YqBUGg9GMCjg35PNcifnkvdqnMyHwEBCYqskbrr3YZ2
qmVZOSe7VUTm1YgPiUcBg4UhjC4ZCz104ByLDbobCa3dbXlE3vsClwSZzJ+flqbfm9dHqrC1xO+9
e1z8t9YxQ8zs/T/7rsOneTd8yIhJYdvCLKyI29Kr5xeb3zjd1Wjr57ZOUoZvOmgVyg5affdLSkZr
7jA1O5d44hYMEtP6odyfqf5vFhVYQpf4KgaVSZzpX9CRP1TIq3DyZKQo7Kw8jaLMSTuAOVai5Ob7
ju9LcrB/ud6VDs8vZAGQky1qPrSYQs3+gamJspfmYa1MWWE4HJJqSGunZKnMzFitloJuHOS19L21
t5HDnXFqXHFYhJl4zFxv4WKatKy1K9+HnC8dwC8sLI+0ACYOPlgMWtSJ78EruvsZErGrwSCnT1/O
USTLRclBAoDoVc7TfBJDXvUcWKRF1StlTBlTroU+QRkDpUvkndyv84krdAh8fsCNaA/f+8x8gDaB
jJk8ZtOBePhZs+LH4z1scWuz1uf2jcGahpCDAb1D35w6KgHC373uaaYMwKFb8d6Vyhmi5ul/AqxU
9sWc/oH86BaATOOlpKKc4fK3ZRxSlj/xADi3XyA4WT7SrTcXgWj1XzxgVHEt1sVfBcDDKyLl6Xl1
AURqQO8YpPsqdD4FcR+o9nlStxj0t9rGZjLuOxOSUkh0SK5wIlWuXKgAnT+cthKbaGmTOLZExx2E
3LXRpKwSgjC5TWxyJPS9+kBlY9/NF/YB0Ut5e4CueC5T+T+tcYW5J7gMErBH5r3td6bwLPJyziop
8IHfpSM8OyfRNAABzn29284o4Ux/+WG21Uh4NlxinQYgfnMePqrmnoSpNa2kQYJ3JZjYXxMfkmbV
XRXXt1N3/gc8CtXIE/WAIjIdFscb9mum/tRnMWSx3AfxIBDLMvePc9d0WKtL6tNCPPO4Os9b6el/
+9vJOxhKtFJgHtBdmb4hKme0bmgdLN9WHDPDdhgMJqdAjJH+mtXAU0wgQKhsjRAL9LHRSjuIE1Ar
Vdmw8Ej2HmbbRKyCZDYlJxTDUqnSyhEcgCrwCfmU0L8NE5aTIZdwbS9j8c+8IMMdgV7l2i9GKn5Z
TfSJHoQKCEzw1OFEFH7j0hCjNc+1LOn4JPhXIM8lar0pn+IF3fnp96EMBe2I3kJLrhQOte/1U0Yh
z1Xt4drMAlFdMtb+tN5hZ3L7gNhY7Z65CGr56302gx63rZPHQyuerpoB0RQY4tpztUf9EqHtsQaH
qSjdAsf4cM0LZHJ6AkX4T8nFof/DpPvidWw2ZckK5f5lvh/bp7oyS19wHwGv1oAkfBJuOwMQe3xn
YGhUafO8YAk2p8SmnUxGBF7M8hBbwS6N1IsVy5sKARK3QV0LSqyAEc+XqzDfjL4J4NlOWbvcZG/u
31r2ZnvjV0KguwT9atA/7cJ51a5A6SuoaHo8AaIYc6e1oA4eeaTC1BCQlX2ECN6vampiHBHMHUmT
kpz18+YG2nR4s6jjeI4SqJn8gGkD6dfNm+YmKM8fTODkUEtvNSy/OFt6MS9BPbgPHTcaZmCuQ1sr
flHWYZ8l1sUvxbl8tSs/NIqHzaEfqUyqR8gEAaMA/DQDSfLbZ+LFC4H+tqs1It+txGCzXCo702XW
JgPWnHJ2zWCDnMwmaDhI4zzpEZF7U11KjeJZRShjzBdBJ3pvRUzpD61iYNi689EDqGIDii82WhEW
0O1r9ejFdIejKwR1UW9Jigr6N9Qe4SYNhKeVM1goQyiKOiwNgFYgpx0la6UVqttB1XZaKeQa3k4b
9+3NNA2IgXD7+zq8oQXU/JRXezbOkbp6FFj76+fpJGR3vVgSCKNTk1BUTeufOGtEcq7g0gT5e25H
oP25ERYzR80cIKc1pBU2sOO4RuCfhhwqBn+qR/5uc9U7RLQNuluvHxa3P7mBbFIfT3QLiMm6eKqn
9ff70CwTYb07TWe7HdcAC2NmtRRjd/XmplKL2UAm13c6ZFGXpmNMhCBlFndRKpkg399IOdNJJYaq
xPrjEOmbTvfg0QJgjJ+Z1BjnZ5wDynK+hvIjXLaMNAHtzhohKBHnnjh+w9KEy/N5qyY7pldaIgDC
JvAhBeg31KI9VqB1m2+XOEj5+dsjkmCmGTRzEBIbft9LftOAnY36T8IxQrEeevC95RFQzGdtyaSz
eG6Wqg9TPNYrL8OFmls7TfoWJ85d3OwZmJzqhBoOG6ZUnUnxJ+oz/J+OOcFHJPtnLU46nS9yevN9
1h3bUXDNOMeLTiTknr8QmjN1p78n9iNNOVe339OB6mAreps1oxPmAWJwV1TGTzcq+FPiWoArH2dq
WUjXHwQBrMH8WsbInMucvl/QQzQP/rVa2eUkFudub9QcALns3qT8YCBVXbvSCeYIJD3HpLD94xnD
VWF0mSXz/amQXibbAjNfGLa78XDBXoUkjRiqWk2/MPukWt156HR9bUqWyO9g0QVpE4N2PYV9/WOv
nNC+lD7Vbe/Clm/mHWkkYS6SLWTl11mbFGGL2CCYZOsll6AnaYwArwiX9u9QQiMAeQggZD18C7mk
fObaWDITNawX2grdR/dTXTVbv5PC7et0mPIVqZNb9msA22tgGj54VBYMiENRR5wVfJhFK4k0b7gN
4wUkSQSXj+uNk6MrK7R4UjI68WQxQN+wF/yz0vIPDi8gfar2V0Znla6i80fXJF2QdEtLv2Ns83ko
yhTSYW8URtr20DY//Xfi/ExlW+xU2e/AeQng+yXHlUf1/62OzTVGHoTmX3lv2BPcxldyUt1nDE2u
mlFekFmLX/6UFU7MvMsBu4T036jhaCDLXkNQzzM0j3iCoMEFjrq1SZTJDlExSxBw1ctrWrP2h+Mv
qXIkdhCsMcVhU3Uvdon9X3SakJ/VGPrvtNw4hXgKu9Kput+7jB1jW7jBDTDL2K1LGSyhg+xLnODW
zq6YeBb6MekZUQv9azgA4G31Ji5EIEzef2xY5gZZkdnBbd/UpIchHiDOQdDynBdf0mi9cykDeIo2
M0Ahx95JDjzf7tEynNJdGuTyFMvMQ4h4OAWHmIKUmrQq9ifObQ1u8StI3M7tXqGoqBgI8jxkGK7o
DhdTLCBPAYZDOlA2+zvG7zytdrqYcl94pU1+s8uZ2aJ7WmrQsVN9qHHV/KfcAz+UjjBePG0rPPf9
ObwEG5JV+e8TMXJVsuUJcusRi5NIGJq/ez7kLMa0ZYOB3qCeatQRbwmsgExe5FQ0YjfQfVVs68mr
5jeaNSh7YFs5tVNbWAtKEukHiDwkTayTb/BeOrBHvvGfmL1b5YTQPEXSA87WMN1FMUeNuaXdB2Ys
/JMN6EV5yhDjTTWnHoVru2d0CoZUR9sxpThWHQmHW9w3jEtufgGgWfLeXpH59qzh7/8VnPt3f+M+
qpRWTQCukVzE6DTjkLin9UDi9dRKjjMWCR4WYZPXH8prqH6yGPV3q9kKisI9H1TG4dJpg2aFKSg7
nLABnIBej6JVuvCacWuok8MCWaIFel+ozdwWqq7krjSATJApODxquY0tEbpPV2r0sM+W1zMpaPli
SeR1r/SEIUoJJrEDzrrlhOYMzAJkD3jiSJ249SUj0XgWj9u4verOLgSuOb/ZKi0FX+uvcSCA3KqE
PGhlkoL8GdXbIC5X+jiO5hmG/nB86ii7dYTCttm14YDaBGOmR2QxRHjvV2aAWaXm4j6hSmwJ57xP
9eN3powzu2YgzDcxdkgQp096KR3nODf23iymHSWIwqn4jnjQrg89Z6+UDPmwhwDTKw9omEUsYnfK
Nqg2tZBbKrNxfzyp2sO7q+Hr3Qzt1TxwlWxJStBS1nQuIOxrdJNYneRugn+iWSv8yqtzF61iyqSS
kfa2CjKSyQQrkHYOa9YwzQMgLDysmgkPE0nNH+si60VcVcHTh+bcyFPN8XNh0deoWY4FQJqv+VuC
WsV6n7y4C/7GfMMq+cek8eT0dv2NIvKzBQPK3zpEmEMwhYXqAN/qolqqlLQ7uPIMf8pO1mWSLVBr
Agxu0IW8s5pstMVi4OWv6hXMgohzQSL/+66IWanKcD5wAp+DxGo9bidQbn6AuxebF4zOLhfkY99a
A7FPXH9M096wRk3o1a3Eqah4R76wQQ76Pe4WrAe9mziHGlOdRoZL0X9MEIIdTDbvDUUJhC1ELpsc
TyuDU/b3AnYOpMW6gHiw58a6kz+jpMXEYcSPRtWacJvJU2aVw7dFclQpf6ByFZsM+mof/ukyk8V3
+7X6WBNheG/715nToOON/bfKwCvBYhf6LQ3wInPZbi63XgxuiXGp6iJIkALyvcofSOkW9vmB2gOQ
lY2o9JY9+uJvOzv1zbKGzJCW4WbX2ZNAWD8o1CAL0VTsHlvJfxNZEiZkTAfobgbBXz8snyXp0ozl
RstVYje0Hf5Y6RzVpdHGVe1iqhc/FU+Fsf8l4vaZPl/3NB/JgDONMHIa9Z8I2lzdyxXuiIYVZPeG
R964WqqRw1HN0GEEAMinmHPk6JDXEROVoRP3puM2X003z32acteCW3J1g6bgKVtJ/Nykt1xgLQZF
wcOkUC/dslOKPWtnwgyGUgrTztMKoTHh/eSHoeRPeoMW8XxY/oitamv65+IySCmLaa1kofX5NJ6V
kju8OkAW9vP8ACX9jsAraA8wTFDNYHtkgFR4uoqLbP24l+s/dZbuqbHMZssEnIdmn7p/naYkESRz
K3jaICdFZN18etN3OpmW+elQyJBksIH1Ap2hgeIaAXeVm1+bCkOtGDqgy2w9sVmPdoDE+hmV+ZGs
EXT4zS6Cj8T+aH+rctvLuDuRMWJfxkg3eZ2IoXx8iSLR4icVDpaOp9YX8YQGmPlVezycpoBanTFd
zu61tzo+gClcZKYc6h7RvFiu44BV2nIj0jeZpOwsq8HwkTGF3yfHPVas5RO0xRBHERUi2mIRgWWO
lSRt9DGU4mfWc5zFrxkfoyIdVQXF8LQbQKzwq7YqX6W3YRdRYqTo3mtqRmIc/nT9Hd3Xh1mxUvar
6OUBmZ/DBIZlQtNCCQ+wTfxNHOwRTf98/T7wtSa0XyKx6GTjEMN7VKp1GGheabk7cvqRxAuzDbA6
9Jk/vjGWvxYy3T+wLfn4fum6bYH/G7WgQR/G3494220oeYdQG1ldHNf5ww4Ef3fkpl+VpAYc1qaP
UJqg9YtNvuIzBfB5y3QmfCnnO0Bl9QTJ8MU3S7VUCE9aXkRz9BsQm7/h8kRsa6fj057fBZkNwR+Z
j20JKDRqQ70LqJn8CIzotYG4ZusLSo/cmRWtUB1sqCnXaZvKG62nGyuosTYlIOVSuLBBRImvWqVw
KoXb+cuA5TYBUx8Ov3z4WKfI0BlVlRGLTs0V+dXNsu7qJuNNR0wE6xY0kkHJ6wG0fHSslwcPvuQC
XfcHt3kVMSI5Ibn3yNQ+eOr0lGpUuta+jh+WxK4VqbKW7LUQC01nVe8Ve+I/5zzYlNsJkspfSNq9
qKd57RGi0nKTarShIMijLZao6QyTpcMcFDc2kgXFJo1d6ZF38mnXlOLoUbnTfRokEae3lFnTuh12
M8sz+C1Fa2DSKhH4wf9KNkJKMewQ5EF1Q2CaAd8nBlo9XC4Howj0zAk73VhC/c1WP/tkeq8bsrbz
EOxUTKbxlekQFjJaGJp7CZADO/A/jk6kWhDqjCziFJro/jmjt5MjBfjlgEe+LtlfKIEropi3KAsJ
qRjuDDaTlr9yYIMqQNcd4gk66KOxIxceDdzMHlls5IIHev6FKe1b1wHr2tOn13OIn6zcJfQciv7t
5ud1ynG97/m4UZToPg7W7kiS5xL/qck9pdhpV4HQsCSTmiSyPEdgESclEJHt1IlVb/f0aWtl7ai4
KyYPww7MwYvRlDcsfAz8h0kKHFVPdNJVI8XUjHrDUJYKL9n/EYtSUt489iJGL7KcSDUUxuirNggy
pQ8dmJn0gTy6jzotPMqitK8gKXKiC/Xq4yYDjbj0KmNTmFdkS8IdvQdzSEmFc4psDMokIlroAgLU
PMBojJf7r/QfYGo2CMFhwcw6Rb/3n74U2nDGBvGN4z69TvL3ipdLRKffHt/ubN0JF5xDl2FQU2c+
B+vxnjLJrAi34YORZgvc9aZWlJf0U7VE2XchItBuDdnBMkqXAY8udwE5VM3wRr9DnDhjogQTbEqu
yyZZxo/+PWkJtGaiXQRE5QL3ShO64p9BClM94uvIFsgPUgqv+Lu/EzkSE3+aeb27MTyynHYDMr4n
yfiCsd3oy/vq/tbJJbBvInK3CeOH8/4jdxJGD3J3nNT2iMSNxwN1/uraywnu2U3Q8w2Odadl/HvN
sUTPGHTu7rRxWt9nEpHD0wkR6oKtVVCVl38FigMdg74KhFRNIqIsL/aFlUT6v9GTaiCc2ukRHe9H
s3tG5lKmhqVla6i6Lir9yCzFsKKfOsOQ26kD/hLGIpVxUm/DuIQN2ktJbYe77UGasN0lmvOGPGcw
oFEl3P80JssBaEo8ynXR1FQxV2bBdS/ILt7uVFM6Wr95X44KgeGLvNzw99u7z2VMP9aLOvjj2mY0
D5wcRH8wOeaKxV84/H5VUC7e/XtGayyyPn5phsguCRQH6BxCxkHqFd7GKz8MTjMOjUIo+lB3W82r
v/3Ql0N/PJuNDXga9GwGqUq/VTlUpedKkK1yFID4quRrkIw/tMz65Qg566yJOzo19hLvOXkfA6+t
9OhgXe7y48kb6EY6ZxIQLZokzj+PJKVfbTTS/Psk2BGJJfB3L+JJgNBF1y9g4NCXTYhRirwBdaJW
SnG8bF50Oz+HSrilIrz9WwP8gg4ad+4HNmBb25k78DO1ZftJToJorBIQ0AMbLykpZo/KyYOrXdRK
Rmz5dd20pH2xxBIIXLm5vf2DbLb4Kzou7/G2pWhuKPDkFZETVTOE2g1JPE6P+t2AUW5Fvi9La2kB
qXGs683fLocGI41etfjdFBViawE729TonKhHWH8fsFH9NAGosZ49/dgZ5tdMsTkGUc8iHgxHh/Je
edXkDns+LaVA9HxP8HvFr/aYYBMWrm1FCEmLKIc/y6Ju4aaZWaws41FN11bwqO78ftmR00tnC9h5
HCG1aOVZvPa1R79VCamIJhD1RBrtJon137LkTg/GLcoBc7utM3jMzEMZVqyNU4VgiLMoMC4+GUzj
4WAwqs6Sm8+vo9090u/Vif6zpZTRuSEhtpY8CYSpgJ4Jk5tTA9N37CwCi57fktkqsyBbL3ZyQU9L
bI+FgiAvmpcbgcyeWm4+uKCLDxx51e9bNyDLSjWhP0Wz0RyK5ZAhznJgXlOTVDe1u7xZKdzu7LPA
zCJtwnYLM8jzSG0svyWduohA/b042RKoWuDvlStK7AVb6MQ7L37NxUXCM444XkDd+FNiB82idkg1
R7v0KHfMQDIBZ55imXZDjq8ruNZ/7dAvhXLghiLf+3l4YCivgB1M5is9tQ84WtdR1KFR+G5vxIbF
blJJAWg0z4E3t1IN+vINhQ3pFGAXwY0/mRebRZFE2Otur8VS345gr4zDOeVGOXCLA+mUJkCkzRBg
XaflkWweQZvJ22LN95yFJTZDi/gS9uiXFqiZoRaUuqofBp2UjpNM0D0/r2h/B/pK8M/DHu7LOFDp
Hb19wp4O+4g1jRXJODeqM8iuTlbUKEr0nxST2uurpb0AQtCuOmz589T7NJGPSvseG9kzz1qJFfV5
1WYbXeQBgTCQxUDfMD9gtmRSpIGYdKdXG+FvPB+nfEmT89iA5zNsIRJ04EtTymgIAMdzn0HQoEhh
mfj+yD4nfRfaIuwcKH/emfCIMRaSsZdPbKghfehJN2ZFeBqgsXCK4z9WohA+A06Jy1pktTUYqFqu
IwiXQbDx2kez7NBMqAb3FxL3wgYvudd7k/SJsG2z6tl2UVMF7AstmSxw2lx029HM7OuH6jia1cOR
nfcsPF7XXW06aHjrB7DMmzcM+ssJ6jxD/Al3rWPYdweMDkGWjD0mEi2XFCIVpN/0scB/ka0aFg2l
EvoeJg3snZnob+N9BOua6QyuQAwcseyHn+9ALyDq53NW4RPl8CYRhz3ERvsBjf62+XqP336VEMbe
9LzuPn8xunAFMN6Nt1s56Wm7Lw/OrOs2QQy4WAwy8u2Z28YZfyNuaBMX+dMVdKmMVlRJX3WcT0b5
ndKxHRVEPvzi8+FP8te9G/cA4hneUdAMrQArMUpsBKopXll/sU3BA/8EEAs7vhr4fAvUk+gFGDoh
eubVgeyFHMPOJclou8Nv7fQygaSgdUfgbQOEtWklm5sxX21IDMTc97T60AnUvhe4rjGAE4xYYJon
DmoZCP3LdI/JoCa9yJulEaS6YZ6Sn7lMZzDfNI8Cb3ZfefDYb/9mF6vjmKrM4/BcjhzgEE+jvzZG
eSXvnTh0yYNTJlVR0z2SLgIQuU0G9EmzL0Hfp6h40Exr8W4CXcPN7yLVuCl3jC8rlmMeyQF3mPSD
GdM60kQYWCldKdNmEKg3LX61foOmFMieQQkTX40n2uJdaUBBKx4OrqJZDeVZsP8l3zflbsAnGnXz
+fyQlHweEz/nfvA9OirWNZgeYIAtopVoOwe+KZbQXLzzTc0Ih/RVFAYOtENmb4uoqJ50y57JgJ2d
YSOiGMO71/6p7gnisqHEAkdRo+CrqZ+dwc4GzDqOrGFge7F7yFFa2lDQa1ni//mRNGzvd9asogt0
h1wKyyIYtQWOjzTib7HJw+bF5RdSD7LiX6rPwZP20ohdxKWKjQ6F8hwUdSepH4yaYzX0vueny8HQ
+Je/RSLaNdTYoHLrHFRIXQ54j+ceeJJeEQfaKQ54I3dYT9HGMEreoq/c4gDWwXmaJ2hbwHay9n48
smHuLPTbgtXfyeIkB0k8/S7j9wbVrIJ1/fUNY7O4UfrV095Y4IpNaSdZsAV/lJMSfOTufn7S9KOt
YGfiuywbclaEocyrN7PVKCJl/+s8gmJvU37mkj2yHnoqxCYHCuO15IAg59+cW69J7nP9D1FgRkGg
yf5vCTpZH7p/c+j23ePgPceezJSXEp30o5UyaR2G7gNa6k8XdswOrVjMJNJ6kMirX7eMbo2wfNbC
Pbz+6rw9sMkSJTJlQt2OvJ2LsMn3j8B43B3LHYiyOtW7tTPq6nsbu9tIvSbiErEgA6SVngryLoMV
iahYoQDdjMZLlVNGVA3KmpcR9FqR1QCOa2sOhYAMhA0TWO7oWpfHwZJd1jKkQnbk5ZCAhAA4Az2l
PAM7bXZy/U4R7uXJbgMza68a9d/ClbXkrUMgD5jsC/WW5PxDicRFbHnXtmFxmydDytdsphh45jcv
Ndw2EAcKoKIWx3Le5injTdiURla+7F71dgyikAEyz69lNmxOIDlbiSB3+e/upF7pkx6UmztBqhyh
3HKdh55iOqrKKeAV7lbJVNF7DV82ABYmBsUEaDEeinTTCjTZZZFcEa0txCLFyyxka8Tg/z+Dumep
jY8/BZ3ciQgmWBSSilA8iQXlQb2v4rE2Mih/qAuxreGwDktlSQe6yZYbmiYVGCLZM2pV8IvAyHvd
w6KhoJJhCyrjw8Mgod4n8irPlDcs2cN8MeTHtbkLR7jRbhwCoP/R+OWWI6uuzg4COMCLXnjB7I4H
hJJLcp279yieaAuRTZBn07Y0tBapggMve8ZRNLq5jH7YRf/gdGx+AUt7ufJVEDJPFxSJrFVre9GK
KBX75tgJ6NAVCLAaGrLiRk/Oas2gLH0UM1LOifDRDYUBcQZa13ONGeFH/9o8QxzfFnlCLFMqg47X
Luul/jffJllvZlzZy2htx0ce03F8IrtO+cbbLjrSUSk6piDgL+MOYczdLdEKtZlbBB9Y5HohHEMi
6TeNJKDOv08tEQBvAlhKrZyHLcYjHDlzG5s3vX0G0CoXG2AmL+wYB+sMxDYFScJfVB25uKntZi65
hcubO7DTXNBnMovBUWK7+aK5OhPyW4CXCRU9f7HtLZzFrhR1uC8jCARbNR66nmILOBErXBmxOWN0
H+pLtJEVemXT/0TR6dkKH5l2JNU5gcbr4Hy05CKz/YsoW3qaEVCk462IBggDkCArv0HNCy35A2zW
7Y7oS2Z40/D2Yp5PJ2R2G6g2uk4zjdcgXsJGD+8zuHvhd3XkRzqFgok0P1m8dkH0XfDX9RARHr+b
NhKXEIstx07obgxVFYCuHpPzaZdzc5BVHEPAa39opTmHq/ZLQ9BLuf28dyZ22GIo2jFCmaj7AkDJ
7U2Ucg69vnueVNpu6JrjSOcqa2MsNp/PYXMQuw/deCILxcDJqjMl2lKFg407NTOmD9HDvJUR02mQ
rMK7YHZM1CPSZ2slcUqzwdo+R/VtEeMtOum/XSLFYvnxVpyAlkGmWX7MSHRVfLxXhMUze5+3cYlc
WW/pzopO1226V94zZcRrXmq9siBui0xwWm4W9HsBwaRXJi7JbCPQwm6EUKUrtnFMBAVCYn56fjBZ
4LjMoLiM/vjfWTaVB+OkF6V2br2M6Ws7xOHaU/Z7hF8qJzLG6FThCo0OP6jqee0JA4vnWX3/dcVL
7w2hc46WnYAaqy3H5exYlQr6MdFU5Pwe97uAxnUNRR2y9tGshAvhpkBq1CYcqbRuOVJgRqr0YG3p
DwYXlzb0tq3rA47GQLRtiCJkQG4VHES7S4HR8ULZTkqD+Jjuy4T/3hXm6WllOYHPUXHpaJpl5DcO
x9t4ix3dgWKI9we9gezndsvCPlVmjyUZYg0qw5ED4iDyrcTvmydl2zTYQXVppC9XDGKTI6ZXlyZf
yzwYwmDTNPor1ELj0vxQfc2AlmNbkDKFcjq+j8E+bSxH6k7TB43O9/Q3rBxA0bHR3R5tfBg+bTVj
/7rbiJRKNDZ9awT7c3EndW61enXAdZL+TtXHjVD72KI8Bj1eNJ/Cq9IaUuRhV48N9szQbr6URH43
6p7ruC+AADwjszm3LhDuXtI/spRnPNqQI69XC7rYHYZgJQC5OP1QoU/B7QuAQdv+vCInu/GQdlxb
zCDJNf6nrS27LCNhPnsNmE2ijJhjogZNdqY5t0mabdQNW3zh3EL8rOhOUvCdwmQvX5KU6u1lkWbe
XdeUx5zyHH4UczqP6Nk8vkCF4OvP+Z36hcIPvplEKY8wYWDwXCx2CYPW4GbpHn+8nwBYM2M3gFEz
wFeZ8MnolVQdQgaBXYJSlAp6gy3WfQXsw5/fqDGPfYpMQPV17qKBiNf4lBPxwWorXMiSgtawdqOY
vUsrjxsDZscZS5yPecZBZmW8eQc/uLr6ZwjIdKefOzhhz8usmT56Wmo/Gc2gODclecpRFgVZQw91
WOgwx8mvrIeX7bICMXRxtYnkKQTePMt3TBXvPaBPbpMjZTw92ydYZXWXdVbs8eyAjq5HLOxsZZSp
K0QIO+HCpEgAj0SD7JEIRxPxXJRFMXhfcX9jBruS0ZCyjRqGxCsT85dkiMZOG8x0zIBijxZb+ZSD
uchCdZE898C8xCNsf+QtLpUOA62OX96Oa/Gv7wEiO0XaN11LoSjnWp/Jhi6xokiKkIabfYTutXFI
x7+ZBbw0xNcbv8Hp5s+cEik6n1IExQlvql62/D1X9PlohZXTpIAcyx8oEc4vABzIvkUInfnzGJET
rDj8lfJnoGe5EAe4E1qZ2WGZClGJ2cbgMHHDRqLNtHtoqyQH7UH610aEX3Ksrz4yZFDavEx+Fz4J
Se3xVeUbPAVhsK2+yrbDguSK4wrByeWHBCGPlHQMm2oYmQbXC2l+1M8ZUw/h/YnV3AZ/uhXWUpmo
yhtZlm7X6LVhTd4f/IUMTAaTZ2RV07h7TCuXFE7nHYMHAmgXX5M2FiRPqlnmrU30ruIqCVbJ7Ax4
7ahnrqxuB4SUaeNksROSWf8d/GKozp9VJV9craJfX9NPKKKeGX3ZOdI9KnYwrGNZhaIEpENwWz26
+Kib4QEpevjz3cZLdHWssxRTEJyM4MRiV0I/6qzu4Ki7YhDw0cnV2FYQniQm+nAZezrLJE2d3Iqp
Itkl9SIAUHvUcICcYGLzAvEAufJ9XK/QOHIBMiN3DRWoc+uLY13/sEVw2WeR44HCYuTNSAZNA+bH
jkmeKP/HHDntW/BfccBmpDBh/wnRwd8oUpKrPRU1otlVTTXNoAN+9ZEL2YiGaebF+1SibdT/5zUO
LAcxh+1ofavTc9V2WcMMFloIy8V1Rs0xi7PlFQWRRa0dxL4NO4YImPBKif3yVM45dYasV7YXYGEk
B/8qMGyURqljf4pEz/26i+qe/YOhuTetdcL1vtPbY3ShBJGtiNwp4invbbydymtY+JUZXb/lDI8r
uDfoS+FUWHwngt0hs2msmO6XQl3CY/rtD6QNqWxRG9XhYbmXGOpBkm+zchv2Lf0i6JMEtqsoA2Gu
qePj1k2rIZsGgQ8EnfdBqcrTkwpw1g4fipJs13EO3RwfDzhfx8Fn3AheBrdgF1plDNs6XSBEbdRS
11/pROjnLItjQA0qvQsIcrqSNEEq8rqQQSJAdCTLvSPMCW/ndDpjHzwGgDTggPAcwaUQC5R6MsMO
m2hz257USQCyJgXZlGkitJDRIq+np3QVFOOEQkgj0LeakUcOM1ZZ2wJ6k16IcHEqARN5qsHSN++F
Kz+X6lK3fkIJAvhqvuHgBdYqjnS1sJYtHWBQdl8lwv0i/HuhzJGoeB972+IwDNUaa8d0FZz4wVwg
O8QMfOOJqr4WhKXMcisrzr/jHXOcHYwErS7tdDDSrYTtmzULf1K0E/pURwBW7r+wWPENFDND3PQc
X30PboFfEfZpnIugFTw2I+pOmKncOPACGpBUUtFTrzLimYZX7L/ud0R9IEypNKiRPzuUnLwNC8O+
tcmv1jbzzRFjCSInyh1vZqgOwVinZsTh34ym4vMBa94zk0AE3CpncOoQWnLtQE/z9ZkRKFJQtVJY
FnM3hi9zGfeKiEbEH0Jh9nFAa5aJ9UqXk06s4CoJ+iNbSzHQFaE9O/lByqJb2kMBRCj3k8LmlowO
6OHFotPWbpJykTUn6Q3ts5tT69ufSmC5cvE2U/8MFcoN+kfemz4OpYRf32pfA2hMJItXtHWvgYha
GcGKsiBd9EHAdZRj2TPd2rQATFeyQa9jHF04zDjgeZ09JC3WqlrHaPJKj8U1BJ4fSd4q+f6kHbxW
kT+VISujBbOAkx5/SCPPoXd6sqYcLf7IiJ/35p58yrJC/coVlzPKV0VGRrkyiGQ7KkuFWphse0O0
GE5YuIgu+ivENJTD8JQnd8NR3YaLGbpw3DMiBfsOFJEZ5CKWSQq9G1XPDAtdCs5N7nlct8dZh0yA
W9VeFYoeinlXsUhxyYEKm4qAoGdMXnS0sLyWgV9ey9jx9hrnM++HSbn8ozhHfNvJWzYAaBjm8tXC
bzLLJsLDkPAoi7j6XxU+3MTGhpYCST+b7wm8j7vq7RcqRC9mSQm1LFdv9J88SkWQ2x617Fe0aOyS
cFQJ0O/qOEUVsBNnw/FpSIl4e/7L9XFDIOU87A9+qDiczSM6aEtCEt1O06A9YRDJ/okBPilJZsNd
eVlCQ9CC+iB+QrnvO7HpCxWSvisvq714OtvCwlwLQ8N+xWNGIp8Ni5M7mj3qowLcSzF/PzgsBrLU
rCktsaUSlfeNSY9FA6gmMPgh8kDSRWbCvmL2Ks8o3CLAHeuCxWbaobA1oeELSdWkNWBHsVZQQb/s
XfjkbFWknUucyK6fr5eHEP+Inhzlqt2LXLimBCnSuWS+oPdsRG89/lCq9QkFnAZFpzUYaB9AuPQg
JnTUbHSFHXGnVrmvW5YVM3U9OoLt5H2/NP8+RVoYNR6KzRSb29LZzf9Ctr+i4tPjw4XOhqEZhlaB
8biTyalHY33+ihaoW83B7Uay2JVQRSdbR4ss2CjusgoW+Arz2hGd79I6IM0O8QjJ+NqThyayBOZQ
FmZIb7kP7p7f48Gp5w0bItimy+Xk5KO9uOCPVG5ode7R+XZwB6ya90FvWty5vFOKMe6hNz0k3PFt
Fx+5kqDEU08aGUoWaxUFBTpGNVpkA3wz1vB7l3bpzc1xnwbgou62al9gs6i9D0CBS0Jz2UAO/gnz
Zn+svwvasrsKpGqYrxUTebndTElaXgpT/YQfcEMxJzIBOS1M3XXCkhS0JP1OFm6yBrBESEmsolUY
ZUgDa5BQTJgyZg3TRpgt+y3Sq8c/3x9scaHr1IW23P9k0g0bcmoq88m4VD2wyw1DM2aYIADYkb9j
P+tev7M4pgLhbaIt5TVRU3kColZm7EmBU81DJ/ydALyeEG2n/snBxlq04xXzsinmPyp3A6+MJF2A
kezAVQDg2kKFFVm5eblgWqbuVcffNoklRWW4hBj5kenKqjxRbx8Urbq8+xKAg5BvLxiXvT3CzWyo
zgZk2iE7dX7HCCYgNvY2NM/eKTCAuf1+2XmZl2o0u8ndXgoZQ51mGcw21GPYL7vkvZbw45cXiRbE
P/Nhjv4l8z9R5el6/pd7zndVhNriQYbP6lQBLAydkDqNClxxlKVeC8Q6TUCLZoglGowPxw/dOB7O
pfA7dmm8EZHdbmziomh2QH71hO+OYYzBuZhwO5XnpC/PHQ6VPxs/2/CDrvcJrzhFWiWvx5GZuA0p
1DVIuyp79eeGqlS0xEMLU8OBij1wSVT+7F9MfBt5KDw7O7qcjH+HyNWP0h3+NjARrfCIE0FqWZrO
sh4Vu2642wO7DF4nF2fO/Q5q3+1uwEfbnoj43yq4jdSzsv94zJiA/gJ0CSBC4aIcYSWr+3llbBvX
FTo/kieQs9BQmOdzehl6E4tSLJcy2u4GSsSNnHXz28qovO9XOOVPKQz4K0X0MtbrcfNYuGo7BKV2
xArmqqRI55QBfDuxuVPvSK94T4HhxxsILgIETf8AH2l3+nkvAH9NDf859y9fk+7HKLwipmAOJKVf
aNeJ+Zxnr0OeUmVJW0aCLFeodJMoYvOF9I5G50Sa0sXM4+ywg4rSShLmqCGA7NbIgMX9iJvScC0L
SHJaez0MHFQKP5Y/vvzoZAcZXQrX/IF9//oz0zaUDC3Gx4Gk0WI9iQQA52fS6sxW5qQ+ykNTWDKU
aBfL3M+I4/vqHEfX5aH543z0NLEQdJTOZhX2MJr4sx1OxGLw4cvNRv7XjoGOkCwqSlGeAOYF+7Z1
lXzJW0RKrSFE5jSBXhSZH/MvrH8hyvcnJdEX+v3HVvArOd7NvBJwe4oHk0ay+mpvTwsG43FCIVpp
9HDhrLbO6oEFOAw/bMNb/8O+TAFQCJjCAd6J0ZjWsmSdAAU+qZTdMOBEoKAs0IBjOiZ4Gx/JNF4A
X4BcO+Pvq3ZsOmFs638dgFm3sAJRHibJlgb7Xt99PQk2cHiq5xkChQU61/uQ9nfJq/wdPG2Nqsl8
w8ZEzncWcqg8VhlEEZ/kETYuEWXXpGGa0zf1B0bFpYa1afls1NnKyVTo9nbuuk0GUswG0xBMjLyb
2qkyzywblwD6Dc3ov7fk8p9Pxo86byW+yj6AA3dczqv24VoCkI+5p1mb8fUnIjyRhlDjkkSlSvTW
ZlK5OEfdVVRDaQPUeN9WuNLr5Sy8YP5qpZclO6mXC41mUiweL+IYm1+z6H3P1uKeL2O8NKLtmwLY
uUWHTimQSyisWxXHAofoH/vxsnMJUcd7jLlkeWF1eOxmR6aKKQ2C3KBm15E2NODqRVYP7yxoqr+E
3RUvGI2igXRxSfu4yBId2rT9qDEnjja2zjVP0BymMpQwFgv/F9FHLu5dtijDes6WboTy+4n0VgDK
fV/Toul6JNoU/8iskR4HR24fiyqeYVWC/cgPYgnbAk2xOnAJc85053JQAzpMi6Og8tAJf/EkEoXe
WyhMhyNN3++p25njAHcFDIMmgxeS69RlBzMn8VSNZ62PPn5JsgSScEbiC5JDQyFiCUWHeXI+e8X7
oaJuPI5zEhrjMsQ0zmIS/JkF+kTzt8s7x3/JgREw1aW+8SikegiW0ph7TtT9VKkoXzfXPbRJaA5X
pLoO9xkcbf+5VuCUng+HTjts0i/6BZ1LUUIMK/Of9xMMRU3wtBo8bR30oHb0Y3qScD1TG0uEvpau
fJBN+o+NeSnvn/rAOI7ChCA/VjV9Agx9b23/9S58nHA//GF/IdNAVbwE5Q43Ad8oD8OCAmapNqbA
Ywqer8rZkt4AvlJdYN2xro8xM6S65UtJBa7h3nNHRIHqTeyFlOr4WHcgeeu3BTzDGX4k31bnHeIh
GizBlSH900dtlPceKRCO4Q7Qv89VBNBJXY5p6THQB+Ezo8Vx5tBYtKTTHGc+ztL0164+hy58pHxl
MDZYRx8gTKwOUDtSYH/dWIGY9zROqGBLeIyaz0Yx7MF9jqre3K+7ymEGu6lV8RaFA0YW62IGS5T0
ttQ7NGDhzzMeQ9jgxDFUKCcZOMC9Uvin3YQcdXSVGXNymEDO1GPeh64+r3SmjD3QS7/PrIjMu3CG
uVlqufbQiBPe85NgM1WtACIoP7lquDzZMWWarNGbMnqqFhC4xkfgkPFXzIcNUevO9YQppsa8Pg2M
R2Q2iGANoTod+hId2nWxB1ZOFJVRKWNv1QRaTEvxIR+kB96BHsQyvXp0PbFxPGwLaMajyVYycWvA
l5pxq95jdamzz6ec4ag1Q1mJQH0R7D7TshUpjDgbkR9r76yb1T+LWsss7AOp2pj35K0Dup3ALRFZ
QJJtQ4BkGBcKGIT6ZI+yGmXyms3NRneuqCbX0RY/2mO+gh4o7+90qZnEUse7nitrSoCl/Zx3zqiv
AB8u0eK+QOLEqOeZM5J3cxwE5DcJ0DQKkkbogK4yFpDWzZOIA1xIOBOB1nqJMTJ6tQw8UMW20JSh
ABuywSCE6CpzQIn4KYDRGrrCdtKGBpfanmM3t8DNrnG3p556rTgiKEdhq9Rxo9R9NoyBzQUnYBKb
PLzfhOz0QI8LGibeG1DdlFzbocSDgwFQ3l+Mc7xw3Lk88AHWVwwNCQWuRiVtr41GeX+hwjkxrYYn
biKVwiykvqgkQE6GRBGtVSbIGnrgTFSSZEnPmX1TWJ0M5RLco4YR6771jWU7VySGtnUKPjeTtbAb
b292JwYGIfQlx8yWZtdGD72dbfvDFnw6y2feIRTmNTe5IB14v6unNoTEiqNGwlmiPFZh5xObLbiB
2FDA4jaWgZD8wx2pd76WRqH49KO9I14KGXLbgo+xLOvvQdQirIjWS+ozNw9mLejXnYyTErqr/I+J
Mk9Uuz2FrVaPlZ3O+9HEuiKKO2hzc1tHBqoOAaIfVKTYuhjGKAoYnBgAMb5AM8ICWiPu2H4wWIci
HEEBr6iagaQMNTXZdOH5C2kLuSaB0EzM4sMTZDkZ4T/wMccC3/k8mkj//+onekFB29IBq+pwG6Xt
IJQo5hu80bmOD3o4jbM2mtdZCiF13d2OZ8iJmPIeab7We6FuoIWzLs72ofhjTdYKkAXxM4IJRpjW
V7QwABSGSE3rhdhZWQ2QR4SRB+aFc05JOAtpRFe/PsCoK8je8nX819cIWPYx6xu3ulMNmFay1jte
nrq6xeeMGbDYYkGu/5bq10ue3HMSkByWRxa0ehxRi1X7S5N0Dgruguu1vaXpRzOnp/G0Os4pbFn1
UdGO/O7s1a3hpnZy28GfD6g50XBq/b0IDCr4oPlERpwtAbw+zhaLGPxHz2nZhQ0KouAmrYPbnkCK
U89AZoDMn2cwUnmQH7/O42mjY5lQgcMlgNcgUdcS1+dMtG8g64+nFFmxaayzzbk88q1nxdE2GDk2
B6mQDuVL+e6yVvGaITarleW/ANAgPiPwvShRRYh/gMtx8Hri9qKLJh/D25JCEySkYDlnUHy9shCW
4vsMGm32NnVgBtS8Hsof1DvrAKd8jJoqP3kdvd5YPT3A7vZkSUqKVilogRxJVX82IJKWfa4sG8v3
fS2aNC7G52a2kXjz39AidqV4vXY8O64qjxJrJ+bek2yJ44Q9CxthVghdqw7xLqXkAFfPJxiP2b19
HDgQYrFBJua02GAO0zAoQ5zBpQ4RC5YemcrtHTN9crBc+bVw8orL7une1CZruXf5BW8PYSdqdRWx
BnipKELMo5brB+ZEOXBHUYqx8SfMsKVlVs9Adw2DnpXRwrFiwGPyLmxj1qVcXQS7JjPQhANunvd0
GKD14vnUmlSj5fYY5obGlwRlKFK3APmtwyypRSX3E3ccGPM+O5rXRD0jgozF7iyhEafUhxMLD8qN
Mh7ectOVTYOAZKKVu6njzC1RXV+f/KFqWuEXtSNKlIi12sUMFUzgfwYUk/ARQhXn1MubfVaOEZj0
UQMNHNsDa4CXx9C+Ks6mUyyxFnJN50qIBYcTugjaXHpjlBpnwHl0S1IjuRfGMOUoImySxRMDRw0k
KUhIsT0O6J5A2x6Pg0SwZfhmp3vGupJcWvQ3u+lklwzJnvjZgYZqjkweuD0DpUuHaecPiCzOLpfW
bkTwvcRctmJWLND+30K4kUR1022TgCDO1KvT9eJCpjsTUf/rt45YSJL7Xa4Ny39EdAp0CmNQFf9s
jogO2nWqgD6FF96wKrQ/b3q1q3TqKYf+GLljt6//UWO806/y5sN2iJ2msVEQVu6K/bbzO4LdaU8L
M8vXK9JVOAYZNFGvdbl4qsfQVde4gBrmEUThfLTlOcfkHbTdJHCnhefc+u/6Efnf3edxJdzAKF87
OJJpdalSvR8wQzTaNMX1b/Bk8hybLsOvRB7bJ07eSJ9S9Ct5A5jonfqAbLfXZVx7fBcOfpBHaWhX
XTe4RY93tOxqRqIl4U+IkkjWOWE3PpLljfZSXfoGwJkiWaNMHFrIVhPCIbjMxTgWZZaSGn8XgYZ4
crkRiyBYQFENsgtHmGIjmKcBKZVB+Tj40d3P2QAH4o5oKvCloeHQB97kaNvGMN+frBVk525r4FgW
eGshFCbOyVx4fmely4LFj4YwaXMyeoZbn5ot1EloWU7JxB/RKXdNBvi6MLaexdNb4fuaEFAuo5oe
pDN2awFWl1DDOENuIBOhIEcO7zEwi2BL0wI5xP/S+/tylivXvLlviK7E6GRm5V+I2/PfNRJ2paqb
DhHeIrsGqNF4+89Bi35v0iiAN0P5L4IfDwttviqfVprxzaD8Fh1z/qSk10gUCE4cDcoJ3Ss5MlMM
iwq9/xAzTifpgbSBo51+ipr1O8BGfvIm8x4RBc1KTdD82Vwmjmv25Mvg3pTuath+gEark83cnfpW
43oxWzvjd1VHQtD9mnW7VM89qUZ3G9FlmpBGV/DocojffXafOqrc8F2Dle/LELOC2665Sr7k8oMy
CEC38Dkp+KFSm16VQtsg8Jkv+ilzXmh8Ky0vYC7ZwBloEO83ki4+Vu/U9fwx56lxtXxU+NXlhHSh
wiilpEg1SEdVFd0RRmwoQk/BbYDNuCIkuAzd9QN2NVmd0PcDStjqzBVEJRT63BVUHfM5JvKsp1P9
9ZqezJCnU1BsToWJ6E1pELK4k/XrtL4B5GgFGGEFXwc0oFHQF1aD/y2PwF+mJy8cuX/AEOQsMTx9
gznTSjRkBX69rwqkgm4mMps+HJ48fluWo43KHfnjzxT82hQ4yW6+hhsKftrK2XuRCUEnuHzoAtn6
kYLq+QBVhMMgctvnSGwyWQtPcjEVEg6ML1JDgE+MJdAAmvSmVorKgjrxzpk/5kJgwRAsZgo4aeeU
9zGY6v9yBpeI8Ch1DQNtfbzUfA3sZesLQ95XgzUVA15doIMzpQeCRuo6XLnpEKfpGR9JrKG/4w+q
gwSdC19dkrekDOAMyRhhLXEr3N6d3BENkha3lSkDcXOHWAbd1doWLRdX3G9ked3Cprz0/9nzQ0LV
V5yzwKOTZo72vOlggh2vAA6nMk1PaZ8hGs3ytaWfsktSeaVpukwD/2/K4jnr4c2BKb334xdqVapT
ihcChnNpsYVThGti2W4UYejhZBmYC6WjkoQEgXesZB4MlCEEtk2N1aYz4EIkAHWsEy9u/zNPwB/b
0oMdFLAKMGGUb9BRAM8sTU+Pe/eKRvU2UOjavTdaHbzN2nj8QvYqoWA5mrfxUls5Tz1b41xcOMw0
K52zBtWbB5hUvrLNVB0Vm3Sz7s3HCj4Dx3sCqQkGXyGWmDH0uWGWL7VAPE7e7Q4LnnKcwC1qrX1G
hGnCeGDjf1d/gbPl3FV7lQ1CY5EjTg+13lE5yxh3Yo8neaNMeCzP8rt8Av18vjkFvaD1lrDTab5D
IUByeW6SPe3ArQxCeUQMIeztTzgKBAimlLKH5k6zlTPwZKhrzRtNXgkWf53jlem2FsVwA1rWcmhT
qdMbrb2qAQUwGk+VMXAvyXDb9zsv5Kn29QgEIPKqtVTREoiQ11IyLkG3rXc/EZuIEnvje8e4w0pQ
5t3P4kLMeROqzV/DWT11mVrpiE4pRxnj1jOuPNO7nkv7QmM+012JHxKRLHX2HDc53QI4SCkZ2ZO+
kRPnuMRuF00gC+AAxpW8/Al6igVh22/ium5remB6EZEsqKj0wLDj+0lqjkLrnf0mYD0b/UK2MeIb
8ZwKn50F+jD9qE4ntRBIunvPBUbv2l59+//ce1gYE6/pehXiiFpT0zTVe6dZnhQnCFAyXgEuuc4/
8IiRx1eoaw7dlN2CWLIURpKVbQtG7PY1DfVVhfxxJ56mvxSh6mPvugeXPi+Z6M5g/UVwTBeJvJlz
Ktu9HN5y6IZsxXvOCOBxCHPXyP7Noe+NFCVtuOGr3oc8SFNhX4cxMuSTPPdmwcBUteKDSIp+uRkW
VR/OJXLZSLnVX1yFhLDJJRS6Qt1p6SUPtvhx1qy/1nsF+3feff6rAn8GHcyVilDX2p9YIoU81xjf
JerP/gXCPnuXcIYwcPl5EHNsuXnoKMDSGdO01alhoysIwM+gchjv5TcEyiY+P1DgQg/c4erHWMbx
mwuffDsebTA1g8QpctQmCGSrwPivSkYVVP2glHXEQCayooVIfY8RCSTLjINQKlFfJ6+it9Bt9HyX
XyzyeFQxxIxPjrde4Jo1TJSjvovzX7p+s5cza/2Sc+LA07jvwlwEzC6tXVv1Q1wrP1ug/O2ug4MK
iugysVaTfoGLItXJVWy4wB54NV0VvjWZzdxSX2+88+2wPwhl6Vm6iVYLty97vm0SUvAoJiW+60hx
4PxZ1boR+l5AkIEmEwJXUU6bvi0i0S0Trike0iTTrd1X5+0XBe7xE91QooY23Qsx1+I5W9TUIaVw
JmMQ0gpVTqN6/0xEeMil0PGeLnKRMq7YLkbRJsDU7PmJCnDOinWa3Sswhf0GH66BPYXSj5mNkQsp
KHeB1KbuWebgeG1cK2mNq8EDAUHx99rqB1dBeQ6P1s17nbkeBpsmXm7JSYP1pzizDZ1ll+HNSw4q
uhQcPY50E+P3+pvlpg5m40dQ0FBFPx+bjk/8QrAV1oLCNbBRqvLvKSlXs+URjWJUQj73ch7dUF2k
qOm0MR9k9T1QlNP39UB6bSsBvSB7SSS4xugfRMop1RXrSo+1kfc6tzCzwT2bFwSNkxAD0yghFIQ3
bXSDf3ZIPsruqkOXA8f2hhVtmXcs4JrHlc5sqNwRmfy7AjnMYBxiJoqs6UDzW2+eK8dLDoqJRHzD
o16PBpFWo4PK0QbTfnsuexJQvdNvABzp8FOC5QX94GC2NdF/2s+RO9LSxxIcLLkC6/vE6e5DDClQ
Tg6/kZktswGGLlPH63cGBLR5f3mQNbLOZnB12my6jtgRZSJTWpb8L3E3RM/Lm1nchYUU8JsIV4eA
F+gx7iZ5u/XteR1M/vDF3APw3xokkjvkPx9VbWnQAsCNyD2E4YIlE2ZCNlyShgFgBYr1xep8jCHW
iXmgi/SfphrXF6XFn5I42m8076ulx0ZUlgbtrWMWKLRhwKhXL0QjgfsBY1pVp5kXzREskRF7uvJQ
Nz1XcstEEyJdgEjZcnYj8uU7F5Mi5hTj+fv3WCSbtt1cq5/ok6uQDxBjuEQOZISshW+y7BfjGlPE
AQ+bZozOdy9YpgOAGJ7AGJg/iJ+LyEbmDHG8Zimw7DmZ8BpBMJYucGVU9YFxnT79O7ykDlCa00bV
/b+sLCH/GjHuEzRMTUv+0BKb5hQNxT9nWZEBqh2THwoPKN+BHy928XLckJ5ROe/TpCpWiWsjuAJv
JoGGNsJ7W5WbG1lOoyqw5cmwK5bvfmcXzXnY1Pz1A6IwVTO9PJPsNcxbAZ7w1VIPFJfBaD1KSREo
udSMsV/esT2t8WiT80UdHa5mc350LolUyjQlpEtHlwqYWGNz6u6qlpBYyoNdGg8ty6ZGzBUaeZU9
t57KfMrmpP1PlKtqNMZT5Cut0rBrQTpebjxUKx9VHOutiA6gqwJOxoyodcm5KHKdtnLNLoroMZu/
YuOLq0KHJQcSkxQVLh5PVpuTnaWWkk17DYosOGIo0qsDyLDPFZog+ZPIbfljeHHySMAEGxZ+pmVt
HMp4T2r67wFYfjmOVLqrSD9tmACf6KwS0Nm5frzR+XuaLOPKSCpBYDZUw7yn347mui5zVeDZzI3u
pG9pmSAjvAtjY8Jt/aLEFYQRSoE2FkxJQHft+tQm+MhYwYMwoaLMbh1Z5VoCI0TA7Pg/DSgFvnqN
pBCXKhM8vQdwllWcEFIqFuOPACj7uRIaCP23bbYRAu/MdLV3OWTbwUiWek/Mgbxe1a/ViIZcmNz2
nP/6o5JZ+rXA20xZCsS01rMptR+7CfRFsNgLWCgjWjD3Yaqtqg7CAN3JKAXjP+eR6ld6+Z8KT2bg
t6Qb5jk2DblFYQFfMsM1B1Us3lojiYr0wJ2cA48OfggzMQzuxUg1HJjFVqXblUBw32znafsTjJAZ
LT8/ynASURNB6NkbPPCwplidm/3laAisjfDthnjV/Lh8YaN03pXvNQii9Hx25eZ+ajuilDUnZcaY
TWhrDTe8HHhpPHyr3Bg7uwAwaMd0Wmb2Nyvyps9R7OEO1jMzePyDelACfQM6s43w4iJ/oPj2WBh/
OUljP0s5yx14MYt89pEiBqUMOLdN5hD+taa8jbcf4pKn/YZjstXZ93662Nzrn//fMZgk2U+W2FVZ
GIKmAZ6ZSE0VbgM/FGfjx+h8kPFzwc8HphCjJzpoqL9jfnBUQmxHHUYyZ34ROcbPwvGJuGLyaa4h
iWUAYPkbucRJPKPUzMe96/Z2thGqYmKtAKfcFHhpg5DevHKSk3sCO9ugn6lBR2Viw+uaj85DQOv8
VSMyREKpD8KVagZzafvZoO1hljxmwxY2MLg+5Dv7rguOesfBb/mGtYxt8dx2WwPKOnk6xr63qrBd
sYItgLM0mM7BVjE2lXaeEx7Cg1HfMdmJ1hWZoxCCGohdJ+HkBBn8d4oPLmGEL3YE3UsOjh7VSayT
YSw7BF1nTe1BIb2e/8LKPmwv5DxOhZDRda85EckfWHbTqqmK339kZpJlqoQ7el6I9sOxvt7C8Rc1
Nv2Gb4vAl42ShPAmWGNXIuBf+jrhpmjoiGzeiBYI1oJXlJR33XjW5q4Yv0wPZ3si1U5zaZrZjfOU
lofS6Hlb1SLIMqKgd+2Q8kRV8MMNVxgXGdZhsc356kQK+xy/7NbmKyAX71iZAxHy72AUSH5yYqJ3
igP0x7pT5VrrQEC6rdeWFM8WSPd2S2qGhGMH0f3JcPsy49sWT0Br3y9k2NE9/F4s8Wn6jQ9V+bfU
37vhKbuweOXqRWWcC5g0k7C93+TX35VGBWlHgzr9JEIwbFiO33aPtsFIemIsWPb2WdI4yaeAdjRH
wKgSNsEnwX3nkUVbRgQB4xCGfrOLlNXc2/SeDD/BrL+jlgOhRaHS08YJnRzdqP4XAeWr3ZOykh/c
pWfpUDdoRfucjlsGn05ifIFZpFK8XV8TiLCzAk5CJqgo0u0XioK5CEH46JT9gVwh/PJXUcyCkj4a
dkoT9pjwtG5c4Vp6HNeLhQ0wTLg78V7NWLyWKWiDv1VpUiHVk4KSBF7rTgviPgdNekaFrAs2+ljt
x0zVS07NLPBa/knJOaCG4a2h1znT2OqG/tBcNLoxbhxFpMgkGPzH5k0Q5wvd5oJgFUhtFT2ADF6V
noVseyKInnyUrzZ16u3ziIyhL3ryKel8M7y+iMgm7ETcI5tCDTW423r+JCGza33zUEbf4hE07SLc
NNLsSSWXejjv1i+2tzcTAL3RhovHTxSKdUNFH+hC+qYKy8K4LTsYMtnGymjFwVrRxu3mIJgiJCbG
3KaxdmKJ09QJE4pDEkbKxdo0eeviGr3ddydZOy6ehvRZEsTl+o4Pn2oe5emMJ7MK+s8BqVeRoXY+
/JLFFag9LMr68T+7hE6RwMbNYzPWOHNk9VEgMhcHIMdVRPJPin7UTZXpsZ2Ew149YBpD6o3o+D8S
aQwDJvahXVKBFO8WdgIjBRXlaeGaIur0Vq0my4rC7IQi+AS9iR+1cgHfAaq6bTZm/WdNOuGS3dwv
7aMyqIxW0EZ9XXKwhQapX+NF73dIFSZ2xbsefWwPD/87Ip1zvbjYCfGJUQa9R20Az0YYlL8RPs9V
hg80O9TA045dFN2w1G/jwieAeqBSqT8l6HjOirViiueiKAuGa77ige9pOmHJ+UCgWAvA0hy22e1+
dchRBYtzYN7hKvJN6hEan+DNwhMUgRSC50PiRKOrJUN539Zb7EDVfVh5grlDsD+EWavWQ0IG0Syj
zEz3syW5IWIT4x/wnJl3xt3vVkHZlEFvMgGRg6KDMUgkddlEgOgcNb4tRmXnxDN6XRBVX334+ugz
MtMtFcHCd6OV5yLxwszawX+eGsz7sHliTLlTNGGs6tHwsIM9yQiqDUuwEwGAupyhZwnUKCT7bXe+
eKFSXf1sWHjfx4bl1rEdUS+GQh7U/QgGjUlDm/SrJAEkQBDSYmswuCaRW0nEJJkHd+LCnEJOnBCU
eM1wYSKLdSJY12EZBP9iKC27tLlsPsl9J7ih3uyvbrF2Tu1oaVnpYwSPDxcP1eCH7si5bsRJnJY1
E3HAtMxWllzVkIheRdWatQQmXYk4YS2wFjL1zWZR1JdG9QHB0Hm1mgBM2GVRqM+eaGzug539Sg0L
ZqSGLec5Mw3aLv31HYuHMJJdiX6jPeWLocFJqu+J72TbiMLzDUYfMlqnsa0pgdmS0Smnmz2N9IQn
QmSfz/8YzBkrT6rNdKXNlbRFJx39zUs4jQ4YChyjrzART7Q3QwOVYvMjBxgeEb0PezHRzPD8BnWG
CJ7HTDG+/aBSVT4hgn+n21bOUnwgMisk/FshhIrqCCOHhBZrqnVZ5l/ApF1oFYfXfwStWTCDHk0m
lA+Pg3o4zx1QFnt3CJvqYpW+QFTaLc8nT7uTEEGM0z7oPcLXjB389SGqyyL1ESZVlLt2A1y1CNEJ
drm0frS6lR0D7masUT6bzDwAbLnGF6MsJvMDJayzInVDLnPgs1varcgcWi2v4yEMPNP7JrqyEWow
KWSaS5NAY8fE1BvSFrOUQKjzNqleGj/ssDzcq6efSGQ7/oe0jkq2Bh6ACYiPxOvAun8gzkjhyA7n
Onx6dDiEUhmdNmyoJKUUQ8xLzgaidSM7Mnvd4yoinGYC32EpTKwMYGhpFWJUt3jz7zJE57B2OeXg
vZNiaN0KMGVQIXRG81RB0DOkbmLnHjSi84VvMkF6OM2E1AbrPH23DIvpjyneEhSAMAslwLdrBJ3q
0uFDhWwsUwflmpY6htlQK/7R3LPwKOqRCucxLbA/eUjoUwFolzohOkwm11K7D0WmhbchV9dm0BPF
jzVYWmq/Y71GNRWXWuf1y81lUVBs4Y+nKDeyuG51Tkt/Vhvh04K3G4V3KIrH9JM+i3FPWgEV74a7
kpM6aReabejfN+u45gpPb6w3xfI1sYJjPcW0NBCzNkyn2kXvjlQnv+uH/KTi2ZHe+Z+v1qYhhCy3
9Fyj8q2XEUu5idoiQYQQyaU6sCMZG2KYvKuDShmySuV9kd1O4qv32VvxLe0tQVoDIha0miGkFXnb
qwOwNCHlgOhqNNchLVP1W6MHPYOUOEZ3toA06we1LBPwt9Wg3K6sQUl2RdUUEwjGQWNCT1hLP35Q
5AsSUSQXPRs8rmFtnuVm1sE8zYEOJwp3uzxgONra6sZxyOW73GZ0EHf/nMNghkyq8I+G44MAO08v
y+fIlL4iqNMJXtJr7iHeNqc8KADL7Cf45GEAUEu6fBVw4ZbIAQmEfg78Ifpn4ywLmmxs6qNep3vS
SmcGB6PaVzo7qf7EFr8hLX6sYoviSRaQz6QXa1+EAZyyZBkKRLoZ9J/E35AAgvIk1ycMI7pnv6gb
+guZQ2OIRR+K81pcQ2CDILwmBjWXqXFADb/IVjHOjHJUqM/7hC//T0BntRBmabf13ciqhP9t0dPJ
xTHX9sspxqmP1n6SJYe+5eq3ikwtqEmuZYqXWLd5xgNkDgSxv7my6Z655iB5svJ/mPglYHWE9Ui1
xqIVdVKccEa1wHs9iUaOkxPo2aO4Sbuj08A24RtM7XqChQ4r4Zir4d49wH84RsHZ3hMiFcCUZJsf
zzLxnaS6teYTVa1E06izYfRWdWVFtNbQ2QbC9imWdGmArLoDxLLDgSuGeEgLUfLefsqxUUpTC2iq
J0Ay6kCNV1Wd0vmtN3ZZ4wfVQUxZqGaBRETX/fzput7jPK2QP3XzrTR3ifz43H1/ojQa5QbxTACw
8gpDAWUzZyvshEyUXweaWqtzpqEabov37bPgzUx441Odnwcz+1RP1ARqaU1nEW0edH0LIA1SvtDt
+1ewbgavV11jPbH8uimIlWgpSJwWlcp+hkdhR5SwUdrqJGZ99wPBVyen98JMZdnafAN0PVJSG16B
LLVgKDOSAQoy91RUy/RA7HIrVQfOLCKy3JfLRc6TDCcw9wa+Z9gikduEMdOr+Sy2B45OAehkf9LR
Ej/oJMg/ekCyyOoxSqGRJKY7SEYHTmTKo05RyEYTBdI6RYywMjGP6Smyoga+2TBT8mEPkWoZhj/F
eEgz4mtFFVFViU7ju0rhTQeQ8icGI6RNKUKN0ndr042A0FbBV6koKw8KOhNrPuaO480CaphAy1LA
2eqCYfKpfjEAk9tGcxOCpi5gBLyN6onf1z1KaEby/0VR4Ynu34eiEaFGt/5S96HTEzSHsDEuPrDj
ttg09zfx7/uQm71gnh2FU/oTvGGIjFITjzG6gyUVKq/PAVAamyGcWl26R7EQ2e9rTU9NKrR3ljqL
vIOqBMKaQLLj1M1nL4JS1IGI/kZLyTxReQ2OgyTOcQleAZLWGKi6T5mb/P4/nHBsGOFKQFAIFyoZ
gau+ddzwZDgoCIQ7ViAyjh/s9F+o4jJhBuh60s8RrFgzzdMV0mp7paABo7tKJK/dexfqSLWpzQa4
/1SINYI+jP+Z7lzyRgAwJj5Gy0Dvpbe0QvXZr2jQfZmog4jHznjpg+vees+Yqs8CEohFVquHAEyu
hwOpSabGgcGxHF20mVs/JLf6R3AhHG3ooq9ZPjVeLY2R6oIdDexaccPdgaqrgMUsPbruPptWJ63E
2EjFin62iiZV/LCQ7D9tIH1IIeVFZ/REq/h7cucNFPYNIWqEzIArsusCwOGG9jUMCZ7wtDqlX7dv
W4Rzq2hnpBkPx2F0eINkdzHCRwMBI2piVZgyxxYcvRKnziob/k5YFFR/1ffcT17wAoCipEZ8Z+tw
72Dsc1nAbyPw46HhCTVOJB1T/K5jgWkUB5YT2rD74eliKBAL8QkcLG9XtQ8bVKOy5xLE32VT3FcH
2NOjG2CNOB6vqMOO5MeHwpQ+AnCejNvZCXZMxm/ppaN2CSleEZmR3hpybrPMSxRrr/De6u1I73m7
0Zx2kmI9GfBcElW31gMBSAQv1nWIGmiXgcn1fOZ+uF2CftN4D3SWSSvw3ZdLqF1yCyjvackU3Ux3
JaGx8ol+bSo6p8RLj2qBi4DjCC5b3iOyw2sDrIeeKsK1c8Gh+N6G0irXOOkBEAOnr1G1HaWmlVov
P6IiEVUbzuKLpUQHgMZkQx1l2aO4rALsocJFYNXvjWV+ec5pl10Tf3pZoiau+zzPGwOZgP8yTRAl
FdtD6OPPpjfmWEQKvdjB/1IKvLShuPT/X6oPUoqGHJS4+5Gc8ZejHAErQ6Hwf00I5ah81J07fKNO
GOab/07a9mEbFLVr4uDqffnoUI2rrAvK27ifo06woOHVRNl/Ro3dgekfyzFL0qZ3CRSk1sC/OOk4
ndMpnqy8MZ28CeTKNxQA+WHzs95p2rwOfQlcj3Hw4+/PTG2j5cVd2PexGkR9XvG/lGEDNAi30T1R
H4P7WKCjTNnv7txC/+9SMgnqT3p78cceNZrnHxHNdxRThBas6LE7fYScjyY9f6rcR4s69aHqmuzQ
QNNs02mjYhikZvegzhcSSo4K1WlF6pR/2NCcnKjz/1JUsWrGtkc0gdyK/aCgLBmaVD32EF15Womq
SiExRrR/0tjlbnp9vuLx96fWZBdQfUs3LeoIN52tKsFZtskgQ+d/qcB+xS1RgIkW3AFzfdQiSYvX
rnfBMY5ngtCMyvlAbGwd8WXjece8VUKMPx2zRY6vqwA1X704d53qYNZ6S2ZXO9DlIBRDbPyRS091
H0N+zekbqRn0ebmdhGGBAS9IPaqcKKoxu/fQDvT9j3tP7K1XJ9hlritRfnprmg+RDk4PkYDKAgs0
/mPnLjtlbJv2PVfcDPwDLsJt5Dx0793MaX2SLqko+Q1pqJTZ/Xyb/+EnoNV+bYpOWzEFYAMvVWtY
cWP2BFFXoA1sY3CpqpSPPqu9nQDxr+W2Hx2jUk3y9Q3ZeDBdyfT1x3kI+B9qnzmLusprYbq29zTj
CgcC8sgpEKYWzLVy3UHjJFJLqUSUbaA7+wzRvtyUDAy2aikEDIWDJ2ysZOHkbyd5eyp0mzqWlE25
FYUSfqyl7liFNTL1nNQc5li1kmX+mG1YtNCtXF73c+usYsuJTMSAnzNxp1T7FOr/DxNCNyW5uVGa
41+UZszjKI6KdV8nNvtNNdUG6R15Iu1Ovu8AwECsoogpXXpZ/OX8ngQ6LJtiDpAmylH78BBxz/o1
5264W/TuAKdvGPZkRyOvB9+RsIGcyK936clscRYVDjNlPhx2+iue0g7JA9xapu5t2mdjuOG6Oz8+
pRlRIefyqI+eebY/Z71R66KENsGy662nZVEPA2Q0eP0ZiJc4hhOi0mgyRXFRJHCwV6eU+Az8uh4m
qf7HteJlNDAYhAHSBRVI5REu5IC/m9Zl63HVFVgw4cqHtJqLW4mpenWHQJWGbUUW/JrMgMDu/yb6
jUsTTkuHirjaIqZnVWiTrPfWmiVsXKhmsvwFjq5wEY3Hj4LPDeJYyNtyCGogwLxt43CmvYSA6Za0
dtHPldpPG8DVYYw6DcgSBCTP/iwYhniAqY+iCHseO2C/em6cCYL/swJV1cjcRB1wNYYxZ5f07SuH
GE8x2CGbD11B5SpF8i8E6HyB3Qh7ILkbmVBqG6KGngnCeilRQTJQT+NMD53lMqZgcUAAjhBBIogj
Y/YNIbHRTwAURQOL36jvDPnVS+Ybi7Z+o6FypypVnDHzAU5W6jZ+pBzTOCZgAhyY9cJNBwLvb2pY
S3PP57p00D0Gx6D/kMj2AVqBlxYpRLSuAHjXQIqsGRU0YiciMAEA5jNZAJ7vQ0V4iCcD1syPxz6g
wdkxTokx3ZIdJpeMKQMrZm5FrNAAJT8j2HzLs/nhEy7uUst82FXapKNOdA6byOFHT4JylfuTjqyk
6357uQCW7oO3ic6J+wtKAlr8a7QRzDAUti9B8FT5sd8dI1qqjScjiP4+2k2j6AmStQqHcxVy0NDq
7UdNUGeK943Y1daHDk4fe8XE+u5nd6zb0ZqRozGt4O/Jj0ydcIk9Ex8bQib9+qYqt5EEIYyJen69
l3G8G4YrjTCGF/un3God0SP2rmhy7kvwfrJfmCoAN3xi+5Dky2IVxnETKm5GzAu9IE9gs9/y0czb
dPxhgNWeKvnCLytQO7lttVwEyll5X5c/TEKz+sRvuWsduY5A1qImmQ83uGpR4QCTBhyVnlCAg5h7
jum7jog5D+xu5JjCbqKdd4PgZDuoPnRSBrF5o+WkW2c+8fTO/h3cdwlGZzFtZqwkM+EFuse4klBH
MTYj6svoJfqHTGSx9/fPo0dR+RHzjwXnZntnOIzRAlYKuHjOyOghJWfdqzDBU3Ayh1JsvgfujKNx
PCUlst+JZjOqqzHswhn0DRqa1/o0ljax/K93qaw8Gee5yhO0lcfBRZfMBQcsqccgfFE8kwGDEnXW
vrv9ODW05jlrjVJjnUkGQsSQYPW/yxJ+Pt6wh0+2sIxc9pkdS3TYMgNAfxGRc2/v1czgn1PYcTKA
GO/eWb8uR9YL7yn7T/LBcI0IPKG2L0sciBd6HvYdT3vvW/aSwFJpHYfya7J7f8tCAnujuQ0zC6uy
lYtRNrjle5NUMxhTuOzmTNWjIrXUq9EPVpwiKn9K8nxYEMjVTsYdyQjvj9FkRkmuvgqzTjQDPPoC
y3/29jVymLzfjbBQLdtPeadx1ub4KNaELUV8aYNAy3LOyGsHgCSf0+4+cNHMPQElM+CAi0ciapmG
EpXYnhIhB1bN+WGDbOnf7Hu/gGMJ5N9/BLJB7tDhpjoeLfMoeZijW9NebneVLRxjml9q3IfUzEQc
6r3apuylxlbH7U1KpwhpmJkNCsYGdgz2O2InkrQQ2ZOHDly1KcDNbbgU/gkZnD+t3EmtrG50s5q4
XPIe4wOTE8vhd8xy5JT/8KEFIsATLP94p2mS1I+xb1q4jmQOluRMxdxwrv/hwch4Jk51WWstbmTj
xmw3umrRcS4Rukx84OB2ywWcRBIj6EIK/QvDBQnFXbIAKXRnOzdr35LSfEvreK+peR0u9APqpIJX
hj5/9Gg+VmcfVOTWqlP3CHKY5KuVEVurunXQhbiAHRdPa2caA9OHBqvFnfkSLlnyW4rVv7v+JFny
sT+YPnlMHzfWwmQV5TJnKpEmoGsesAHZjenUl3f0DyQFcY3CS/TjsnJnYmsneUTDd5B/mafmQ6yV
rclruhFzL0IZvMLfQkhmhxPRGaTXF3i2V134NgA2Jvcah3CIKg00BeNJyfwIFA3CsgITBcsIcFv5
VbFXH/+Gb/9LX5sUL4c1v/sHB92D3FUbp4aky6QyNbb+PRETw1ZceS0LdKdt8YFBdA68yem5Uvh/
CUtlX63UYF+Xnn1iBXMmTYx8EqzIGqb6agfpBnUhY8GH4Gq39gYffXURINMpZFt0UMhQ1VEILP10
0sQUAbPTmgWRGeAVyFsR2cn2bzza6o3PPCvfro7N775wca5LAiumRLezN4QXqyjTDmOpncOTT0/4
nh+YJRdqcWxr8E6LFWuHasAJuBRCtcr6wBRk0k/WTwKgFe4e9GH13f2kyM5b7iRD1eMhAanGfogB
P4VlYH6ATSDWvgQG5TQqvBa448ybbRvmbFc89EVaP8UmUcUq4yvMmHWxT5N03bFdEZU+c7ylASnH
ldd/aBPBIqEW4BxIJ6o0+bkuc1c9i4ySyxDHnps26hQ4Om1VNZeWZdXbg+s5qJ32HHGGAKpZ/A4f
0eVhShSYWPqoeuIcEtKrgKVdUDP+5zjIa7L3M1KKmoDVN26aBQJkqY+EA+nnUi6aqZYPkxEQj22m
L3KosGQGJaU/ILSk0dHgaggK6ys0+8TIprlugkFLS3sL8y8Ptqq40Uhn3/tH758nQml62FGUSBzp
plcoRIRQjWHNfjRiMKb0kvuC9z2yHZI0XwM6IDMIjezJE7b6oyR3fiA0SCgr7+jl3KTq6SDwRtA6
hyBxFwwrDLRwU7Tvw1ncgEdAgk+7ApRkCOTk9Ce1Pdx/dy/A+I6WbXeYx8I2HNL2VbmW59LDREwc
0Shp6kOgQFkyjExiX7Z09C7Rgm5wmyEDD+54KIRvfcFDeJrhQkTxb61iSZxTjcRBZS7aso45MC9X
Vjrm2YYKkWGfLXEhQrD954wBX7D4ZYB31N8Pu5QVyELIFjzA3VnJO6w/TV/8b1L/5sds3MC7aq6z
zr+javDL9uJpkwB75jBh5rfgz+5LqU7Mwh25H256Gd8ggVQD31SRYUM79StgzkJtbQ7b5UT4FKgr
/j4QNFE/0Wxc5NOs5cL0SDv0kemH90hwmYX4Mj8Ln6jQoJbo8ftF6PsdzB8ymkPvnH0LZnvnPoek
UGeNDVr1G6+Mp+ZXnyJuIZQVQkUmZO+HTw3zy77WzoSDQkFmziIkfImlDEwwP1XUA9PUwEqbyxfC
hVJsfAmxqULZEprL/F8eDqX1Caf/7zfJXYatSW+CGnug/ferJptD1BPl/Sd1mLj2XifuZVYO/Ial
Sba+qlLtVllm8czI5axhh6ldGPm0FTweAFwexT+slxQgCKVfuQg4n1wq42h3Je37G2BOaacOFlv7
TrTNQWnZA4enORJ84zzJvs648ysdjN8N9Qte/SanzGzb4czNo2TztMnoT1Fyv4+1wDhWQsA32mcf
2Pzlls+scPNttoNLu5pywThFvtV7znkciEb1MCQna6TEFm9QpxzzlzDXKbAMNwcpndfzhsoh/KmK
kToehLtRFA9SOOThyqbwjimks7WCowBqlXFHmm8H1rzDGlYiVwmCgJzrfrGc+psSTzoYk2tufdIM
PsuW7KKpAI1NMd6mecGT/nquEFWVsikYvzu/eG3LiGRnxuflclo9tFDUDw6sCOgSJHmAUCsrKwZ7
5afAWJpbxTLKJWdSPB6OlUdeazWGx2lVFUCx4Ffo1yA4Z8TEUz0IbaYsaXQjnDE6x7WeoTomZFrN
JnEyTPrDHzelaMhmckx8m5YYRZGZE8j4hWK4JAaVV83EZWz6Bt3M/uTUck+vQQkfHRCdXNNLxA6x
HYGuYxqKO95jirZj0JSVEzCmY60wWintxhLqnIyVBNbbKWLb9B8NeJuf6wpRggklMXH2xmWyvA==
`protect end_protected
