-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
YGUaNMcqjHTm2QDEimtuVnYRETSC8oPMvj8Lrpc2tVNA8NAEfn/PbDKkqSFamwFY
n3H7lpQMGXz+8m/qtMBicVcOclGP2+YRZA6njEk9674v7LUPy1GBzfT0aDDpHr/G
RYUocjUa696Zfssvp/kVJrznnmdtcukXI5U/dNn5Xhk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13635)

`protect DATA_BLOCK
r54AOv4eOKedyP8SvfGqORNPuSr476pZkUJdKqBEy5kGPtOqhr0PxlM26IAM3Ej5
MDSUd4T++oQUjNMwfAvJ1+hN3o9dVXZ7onsyhS/WMu2IRHVXQmj74plnHh/dsIX9
BrwHhRGhQYJyBzIHoMVtU9zRAGz/e9Q1HXvMQotsY4wfCNv/75d+9qtKlk+95zGU
Y1KRQZXEKbaC+6AY+R5VgXkUqGabFCYIOM/wdNv8u5PksqMWmAVGArLiplRQNrtt
SpPyvFB6nuiV62OLGl41UCwsYPam0m432tN7ANYYJfyEDj9k4qxQpJu6Ax9tTNRk
s0Rzl99QFfKrF8DXf4ELfgDhARMbaBDgC2o3Lhe0nEYF5cvmd/JOcOcWKJx1rAtt
IsGDuMJGR1kbrFpL+xDbdRu/x1Txjf5jrvuKahnc5v+eIQpn8SHw5wTAB9mRUW/o
4azYKybzzlV/gOX3VjabC0z2R6qynQHHcYEzk0pcHKSB5pErlz6EDNyelillI/Zw
GQXuChCxZPOGE1+X339CZmf8BTFO1lpUXrTNvcj+Ki3eCXM+2c9JQVPM9JT2rjlr
/JkcMJ56zFQpW6UV+dyTmPxaFqehFH9UiDO5MkDnS9xcct0bpb1MYcZ+8pdxjNNH
HtI+qGOlJO/sEC7eZWfDXgoSlKf7U7+x6UVtqbGk50M35P4oVXOHLXAOvMzOWDob
j1cZa8XytpGq6nPyMMLSVjeMSSBXGjXJnXB+5oWNg5Rcqv+PFYaPtXSGJbvQyk91
oaNZV3veU7l/vd6zspFFadV8t1yK+nKXf9BaLcW4uQMljEUoOrhG73Uifxi9FTPS
RjlBG2dPjiX7PSOoUheFdLqX/+5fPqe2tgY8pMd3yZFUfKZEWy5iq4FBJJ8cPzYo
WkQRx2TVEto7oj+SEVUp2scNTZrJEHVPF2PFBmDGWDFpUL7LAsPwSjO4rbuIQeka
Tp0yZZh69+wIhEktWQ7lb+AtB364MxRuWxfgwKy0OZA/oBRCwNW3hTd76xappRM7
vLbXq4Ok94hNTyVyCZf6Ox1nD9IPZdum+ydUQJ4Du4UazAcUbwbTitixajxkANjD
tGIWiEqCTo6+UDyGb4NqaquT8IEwPJgJLOwwS6YSbi7zTqKlqZHfnv0+COxBt+/H
uN/lM4IAaf/4JJEVkUTAa0N/R7EYJ33aZuSALQozsi/GQGLSGmPAwpE6CjxXP8So
qUNIIbiVeyGGOGKJl9amYepasGFGOoYeNFuE6FsJD44nV11fbOEFlS0Sw8fAKLOc
0r5xvX9d0bC247caKOplzTEm1dvfCdcN1WXknw+puUyhb+FWOFxNUy+7T87F0Lms
GSnth5XBB7vwLKtvn8YbKelaAIPorFsKWOp6p4ldeHonGt7q4kRaHpx8JYxt0OWK
3GWxGodyiZBjZrvtX35dOtSwsUjGywDjFMKVlDmbLvZgo8PZWH7Sr4wXuuFRo4af
WrDjDiD3sVItXryAFXwUQcPcuNQdh+cTKQMuXDt+j/802XJ2bVrpPPXxwx9WU2eE
wx8cWkCHMrTe4/xqHwybWqSi9WvknAG2xNhTyLOiT5UUAX/Uooer4jZef0kpSrDY
aCPGcIH8lUe5SSRlCRGxYL42IztVvnML8Tu3Dtp2qRHh+tYawRxAjpoFIZBhKhNk
o5hV5XMNeiMzfDjPHHZpJmelK4RSbXyf4id7dYIoM9hzXYE7QuXAPWhELRTR6bNE
0OctBIwdTSp1xyP+lkcGcjKEOFM0lOrxgBliKIBhGx1WYAKzwNtIfSKSeCiMjKBW
WH/01lQAm20wdl/ws8Z2oa2W1xpH9K7WG4Gh4kgyTaA+2L1yBqhplabvXWGWtiQP
cPfx2cwNZxA1y+WSSpvSG8DceJKNXkpqAt6lrH+g9FhhXvlLpMcNJ3925PXUR3+w
79818KVURzrengsJrr+Z7k+OfP+zLWa2xmP49X7vuxSjhk80fBZ1JDD0qVOyQkrG
fQU/y/SrnLyrWHX5hghNHQ0wZAFBY58l2QSYY9EJVKZ4ZmSG325FraQK8TM64C1N
sZnj9yVI9yT6WY+tNMaC8PGPWrem0c/LOpQz3NGh8pL563mqhX4p1m//k66fqXv9
Qhdk7KoNJsTn9fzCN5CP7OxylJccGPo95KD0WwuGO1cdb6PZrkV2aD/4AyC98fSh
FkUaB8U2v9SvykispYafEGAb+XXsE7ja3xS6OQkefk/YG1GwGdipG6Ta0FcPNnb/
qvFhACY7lgeazG7awhcpXoZPL66DqqkH//Bg3bufwc+nKOgrQNODnmAauCMFzfzn
ASQMxzdEdWaR1eIyqbfQXjMBm03nCjSrQbgDYnC+8uWdgu+4cas4tBktUrer1C2i
1tD1204+DiyaS1LJJJa4lM7nfUUS+VKseCRK0NRNm4f/hK+U/2cd9YlLoo5qXB+t
K6slXUrkrXrTV1FXGNy6cGO+QmzAqeTrpgOy9zH0ref81wiXFTERXrbbJGvh6ZqT
TTtMqXLS0EPtmCQTTaudEmiMCiun8a66Ztg+A88msvG7iO0ab5T4WVEK9RSKIvr3
ioNfRaH5P3Cd1OtrkyeTnvUUCwXq8EMjd/Rq23fsoeOV0PtxkQkuSQjeIKLImCZ9
A7PjDHJUrCwGAJh0Dc//5FUpAS93n9lPXyYI3DVPWPoItu8V7iozvV+lTSp1+aWg
6UX/SuwFzvWm5cdWWcPvOB8grV8oGME9F+VT0N0AnIXHvRUCuicrsjv7LmMKMXak
85lCMOQcQ7Bu7s8SRRg4E7kBMpu8rGalcJUdDX+T3MTyF3XlyAijeoEWD++WsGrW
khb4lgZ2aqFUecgQU9BSuHolhyMn9LuDZNwXbgCGFAVFYTdYHYrUHlsrpLY5+Z/h
AYYYEW1E9bhGb/7iXtz/igU09vVzCs3TjYbq33ZJ1t2IPZba7RN+cmFXKlcOHdL9
WvSYSy5AKtDmysp6B1o0rUqf1gRjwOaWlyfrqWRLXcV2nRjn2mjF0ys+fWjidcvc
J89CTZ7dOfZJ6kjTQIModabCU6J02I/Cca9gIN6Fd4JLbxPCZSt15W6LLRHgLwoC
3zgdmq+pEv4TuqwsQiyszLbJfCHg/C5GhzX0eqbNxl7Bbe0JKjmuq5IZtQEaeFSJ
TbdOJ6dO0cdc7oD36hnkxmJ4BjZfZZ3TaMMkFLhs01a/cp1BeRcfSwAjQQ/VYbzF
YYzGgP3+sbD5J1w1wPf0ku71hQXwlVu6XPg4+zixFdPAjZihaB3FPbvGn+447Qbi
dvzLhNvK9JpDviWx3iJjLgWx8FtDbLQGh8h12fd6LsibzjrxHyWgMh7+hP6ZAozU
7wUgjeMAZs4cBUm1ZpP0rFntAfVoM8AQL+DEUKu1NtCttTs7SEslvGO6QDqBf9zD
R8YXXo6rcjohMOdUvVoLiFAvANySuCoBYrSPmiJryGw/xMWUGr10/d/i9RamnXh7
uLjYugLWyalYHNiaw2H1C/Wf/RPam0QqxrXayNlOI4HxurajmV1fv3VQJGAQeSfs
oe0b4kCovB9YmCJiCLpyBBBRYAujX2bknOmK2PcjNLxDil6f+/K8ysnZCPiYx0/3
hEvXI/EchZHUONGSI5mtXUOWC1fZG1xEVBM8jxyGiJgfB0S4W7huYQwUdC7EZbM9
Fx8XLo1dC6KuNxyid5dSBIeFW4IRC/GFH6/yVSTRd5D8AatoesEdn13fTwQh+5+N
giR29qyqni8VsNK5M1yNEqdlVhA8miAjd1CN/9Pj8BzWus08Z2ixGaA3gk4u2r96
ywS/5N7RqovgXMYqMBsSUUu52HzWLCNMw6W7Wpx1TdigdZt8qPrf58XZFELORVr0
8iCpmx/RPD/+BddcSnW9stGO+1fkcKP2VMktOA3mf5nAtn7iF9j2FycvVu6Mluev
Z2cxwdXuGSHPRAk7ryAjGMaHPeBSMMHmr0Pa7DfACtBuQR4vBS7VhG8WIdXZKQCx
2cX7LqPNX8xcpcujbEMhhS1M8nnfBjOXg2APYD9cOu1p1QnpcNx0K8h4XS/8neOc
slhnt8EeeLt43XmFB9/XlhXuetwSNr69k7soMMSEeluo7sos+nQQc/Y+e9UUDO6z
tcHK7ozlsC3uKnFZ0YNCLyiEA9vL6EJYkw/6AGB3e0+DAHZ9tWG3/1GS1ezNitix
5Py1lsmDvwkDUIKzshL8x47OZY9N3hTLq3CKwI4f5boV+BjioAkGtxtFTxLyq7d/
ubRs93wSNHVk001ght0pBMtOfFQ7r7jqAZQshEbAMqsZ00pBY8F3+GXj05vYitCj
hgaDDd7pn/HqeENUEcj0wZQ9v6UhqX6lBxnHRobnjT/gWOZBDsy/TxPRTXK15w3z
fR9tHgIHz9vY0uqxOEcbZOT/2TQa5ajJbW3woA3afgtlLeLAyzZdvvjnBpQayES0
P3uvwe31rIyb0pwrYzxvtksbshzhLbNCBx5ZCKwtm6CBISE4vae9sqwoqFor9g1r
XkCPaX9beXF5Vdxn7m44fGgYosOcCrBbw8CpKiBouDaQ0VqaX9m9ptgUrNCOKWB3
p80XWqFbLzkiE9rskZtunZPlUrSpznpuaspiEMflN85mkHVDE+q3SV6euKM3ipx3
ciHZQpl9wKZeIqvWslBk8gc7YufmJu5jPyTSNRYLUHddEZjeQwFsu0bdrwZoNqM3
SiQPE5v/1lX+tlfl0M62660OnqiwJFg2p8BM9ZC4EoFDebJyFOo5SjVSCpb3wIL+
V1js4wHc+BK5XJlsm076Nbep89wIRoDUXjng5kpfS9s1OkettzOgsYftix1hDBAB
dleCqISRRkRYqJsgSb6UwlEMYB1uRDwRIjo5AARZ5afjsPvUUQvuW/WXQ8jKcMig
VjCenqkODCiaRExcT54ftMPxNCsqABPcmQzCjcnG2PJTER5fz/0hxOuO2hZobyqO
2mZa2CF4PzsWFdC1yL1JcvrMfALHXDD1PtQzRP9TjMbRG8t0u/aLooJjOrG2pk0Y
p7VE7OAqexrKKZ/l9L5NaZ2bAxYNnuK9HVGfHzMEFukhpsXhaQNl5DcAirMFYELp
T706zO58J6JjXGFX6ZjQdRBjioxZ2FWHRSdy5DUcA+e7oLyEB9nM/y5RUT9L8pFO
6GNRgWbSbfuzzkxW37KuYNxiGKWy2kfFp7HN+A1p/lX63HoCYVBA80z5n0WAyGN/
TETiSUHCUXi256GvEu3OinYWh3ZZ4wJoePqAvmP3VPdrl4RQuwo/2vNHeliKVXin
6o1p9hQLbQg9UTnFnE2ixKFr5ILR4rTgSt7/zSnjMZjY9YyH1j9pZn7xW0SgnaGH
CN2KjPzR3ug5+zKZKd1/NFJ+ECLMX0OhmZ2/EhScMlCKcjZp2FVrASb5G5V3ErVD
09JbG4UB6JydEX/GuNRWwlASYWs4oTXgALZOnOrQCQUVTHCRXQfIK0lWEsq58uhd
hSxcaM3bQhnpGRXDh648/1jGyNE9nL/wWs0cn+j/WQHYeu72xhvGX4I26HeBj5iT
LajtbwVhR1jW21DFQELXdvhzp5/leKunDaAoFPvHF/4U3qV5yOIFaUxSNNkR72tp
7TGJPJ0WW3LQWiJt6MEETQFIdCOKTIa5PrN3Wvs4Aecqm49Q17BoLZjxHeL9uPql
PsMSq5C4xVT02U0rQ+l+AEHpULFFNTluZR276PHA60jeIXJl6g5ynwzj13DJ1kJl
WDltSyYo/iwGMQaQpAl1OAS39tdBU/eXEoq7icRUZfYk75OKXdDFxZ3G+g1IcHvm
YWrahrCr4x8rcOKn9QHhE/d9vGSQPBiQx1zrGmOXtp2R3cWtALqtOLDHLz5Q1Ze4
+W0zAXt8Sb3VRIvrpHCtoE2LuZd07Xlue24m47MS5Wyp9j9uBxD7jRO4mHsEC+6C
j9EwbaRJmsxfHjJz3JQMAJoMBtNpIL1q7zkJuSQAQw4m4HmG55kqFa/MfLp+tXs7
720vi7Pr1SBIHY16SPZHeEaWoMq8+xJI0Yowwj+xzSRTSKxCXNDPgldBDtGUi/cH
pntCQPyNhsdH066bohsMbNTTOjIK5sK9oD1FgXUkpRNvBQmLxCD0ldOpD+BKz/Pu
8tGuXAvql+IwmECRHB2tofJB8DE6hSPmGdJGVo8Ge6iTS72+EqVwq7L1SK1AfwmG
KoddA3OTW0WiFezmEim9ElHpu4fLjcQFHvvoRtjMzxwo1nHYElnMln5DsmITn3Sk
Z+sy6IbUq0vCFZLjjcpqP25vh9+vwArDHL0uZr5DdvmneUPBYrdKbE6tU+cirWJY
wxxqoaggYvABOrvXcYq5KvyXEL8WzTCXYDQ5cwhQZ03R6yiQrc44pOoM88HlXmP2
3zmIdsN2yRUz9NR9yaPXvpIcFryW+n0GUeLc4rar/888sH1GhrSW7FmVpgRWwWmt
5y4Tb0RoBRgA81gO3EkLUwvaUUVtzBbAKfaxcx8ePr+aRERPz3NZRNBT4mcabTpn
jFU+ezJiduQGJLlQqxE6Z10207ga3LOg62gS7y02bUFAHalSjwv3i8oUnTq0MmYb
kG7RDLVRsjQCI/tNKZGVOW9tPyxlfs3TX82j6ZAsCh4FNjCpKRgUUD8q/Du2g0Zp
r/nB9vM1O5pcBs50owUKRtztEA4W4AUhmCpYCUDwCOhyH2B9EYGp8BRxz0MW9KS4
uat3UHFs9XXamS02OcT4nQmnOwwa6FYOW54xGuHMG3eUPs0qKuO9jP07loQWes/C
paFUBDGo7lldnPD4GP+wmq7Btwl6bDo0+Ipo5bqcVOUqAHnalS/iYVT+BAunlVnu
z2+KeUo4R6wIUWdDJWHDqywH8ea2lE3Yr+rQPwyOMiZLuLu5rgPIvasH9FdXNqT9
J5aVO+rHWRscf859ZvkNb00AGGyyj6Acgb+3AcFVeywt83XbZsM4x9Nh06t1mpyy
NYY/0uew4Y/Tp1KrhIlfgi3WLxyzke8ugQpM9I0VkHoq+C771eR/1TBUoixpoOYr
GmUwBTqz3VzTAZ6zpVtl3i8wMNNwPfKETqShkbjJuW3qkPWTVGdJftMdxE1jJNpm
IgGMdGjPx7fb8nFgynij2UfOPbX+DUIJNcTiB3MUXaFeElhCarmQcIuTIP+3Z5l3
/8IET5+ajKqQwyhgAWSD4YsqdeYSyXjzOjDavGYRYRlqDlhnmV8SXMLRIDD920oU
97uNoUCkR+5c+7zAS2yv2h862lNYvAZlGE+uZJenr16VzmA4L99NoveV8WMSVnO2
WH3Ry7a+vhLaCZ+RlrOWcRypZ+utRc+Wy8zfe97dKFMZ3WmtKCpMvMsV+ckG6Bg5
1XlPTy9UV/8YMkY1dj/PUM0bX/s0H2DbP3EDo2qIZ1dIRyursFnajHP9Ng3cp6by
XJZsYOIfZaVzYNJueYovI/ZZ4Lj+HA5AlGt9hUVdehU1yxzLSnfLssXzxvjldE8j
I5qcB4iCUb1CbhiD5rTEmjB1ZRImIADuntqZtpMj8u7C50NI2SXX7JMsyK19Lm5L
fOpKXAWpCvDmWrtd8PZE+c0+wU3yNo5Vl7zAc/EKecSqRmSeOw6XlqGG4U4MMHae
mX4yqgEjSea3jaBZoI0Ly1pa/k6huJPmHQNjBDGh01T1KadiZERKw+K1mM+T7Fn0
wbJRG2xTZvP0ofG31B8KrAxec//scOlB5VCcugK0C7yg8OHZjH5J4YLor/hixGwq
gbAXUJNOth7ZvV1MuP34Jw3QdxHeBr+N8V1fPTX/14HP1/5dxbOq3dlsEkaUdlUJ
MNwA/l+SPRIZEiEGqG7tcw11xgyvopoCJaiR9rE338U87nSwZRWVpgfUWoBXs81e
+BRp6qXdbqAnX4Q7JFxu6xSH3pXZkFKqdPLS1VlnDn0RKZUeloGUUZvGKxUxe7kd
9KloWMZnw8xUrxdlx/SPE0N5SvBJ3auxVYeSk42n1mE6IhX/yYrDZIJ9gP+eERQG
ESDsEHGd1yIg4DjLvrQpAeNxEAGh5cSt7tqWIwEjy+KSqHGDtgYehZxiM/Mlc35t
hNvGwG3reH8PYt3pLc0uoUN+QPZ3dmPL+wpSEiDBbZorL8XcN+//UPcOqjxnKN+q
fTNkhOrEcwBTvF0C3TBaCXhyktcL8RVZfWEItTSsKe+SFh/xe7FxkutCxmJO/4AP
gEbJ6WinjyMdePtiO8zZrO7SkYr/hlU3bRECTRJPyPPC5BrkVG3RwQfzedcIoyCs
iBwBmuEMVhVpPFfF6LtAihXLwS0pxRGnvu91tlvIzv2egqMSPDCqFOcKsIeXDC+t
AIsIEvi1eHwiPN02JbY3N4T+r3WSD5UvX+pELeqoDcMLtaDrl5zDeVV6pfWQQj9v
WeJaHZypjNq4VUll0iMHZCB6ATlgTevK9jIbmBOoOiYQSDynEpC7ZEVQ1TJMSsKm
fu+Z91nu2e70cVV+fAljbTId8XjNj5AXK8dbzPo2BjGjVcneGyZS2iHjj8SQwpI2
Njn9jKUEceTQImVXUXyQrDE7PkfOSfzGZ139HIuXVpKvG5JjJVY0NAIyNMhkCvOu
/cHYqaUIsK24xmLd1AdrBsoqngv1UxC4Uyu979Z49FKxXdEuQ7uAkifo2o+It0v0
RO8UTMEbcsEWkc3D842I9pH10HkTKxKJDJbb0W7+IlT7/K5ZfsS7YAkHxJbQtACG
0BYX1L6KWChIIM7EndTrVTdTyeYc7DhWaORcDoTekzFpMNbplpltsocjI7Qz7mLQ
Xmzs53WpqhSSfTIHpCAnlx0LZ1x9dRk9Hk2Ypjv0I4tEkIFQwbeTpb21qTbIxBs1
padZxGym0EaW2mbodo6n+WeQE6FQuiPtE71gzUb35/5gw23yyde1KqsCsEudwOE3
ZdBIeRB+lY4l3/OBuUES0PwKM4EuASq1kYewvLIKQDSCQwVxU99Y3zfl+hKOe1ai
tc9d5hm0X36SFAgF3S2FbUjz1h+qLa6gy0cIGd8Ztg+M2HdDNNK5UEpD9hRDAH4M
Fx+/zvJ4dkrOBAloIOkmZu61y4YJ7OzsWLyD/vbgra+BoTETIB9gYZf/vhwWSgAD
+WkZUxSZA6HH9scP6e2KcxkHyMmhAQnlMzm+K3t4UKBBpCeCqkLli4opNyZQYXXq
uck39K4GkeopxFRZbktwhABhiwtcrsMbsSY58WDp2TJzr/c9MCHczpdPvq24s8ZX
x2J/+noF2ut50wJB+PWTsSF0hMw1szMs+9x0sy36XxW7yTvPsZ888MkrT8w4CLYV
mViepCLa4UYhiWU2fVUUzrqCocPT2iMFatfxGbVsyx4z0P75FMGs/YpAY1v7G6BG
v5T8PzkmSgvQVOYBSLbQLGq001af73e7kHEBfDr/2tI/QxYC5ib7YlPTztmh1sb4
kVIJaurDEpOhDuhNU9vX6aea+KXV/+1p8ycZ5N3+GPJOJO0LE0dBAO5CjpK1lSM0
2DrfNbMTVAHbEzSm5c30HhLidjr7baOZlpIIaWj0LcnN9cp0/SFCUFtXBguzYO3A
PdWZTqo7BKVicqfwN22ldmqdLdgD73T+uixSCdOjVxb7mRnncmcVd1v1929leMiL
aHRh/dBcNSY2mvchbRMWiNLxXgzFRiqHLmcQ30/g7wy0ybFgzF4UgXlViUUCKY98
3ZyeedjDHLLG1iEYSzlysSPD9+SsV+FluWkqeihzHW4CHiUgkjsOGgzcAmvYZCkh
qjuA0cvwSoilYeA2krKUigvvRQVNInedFfPcB7FBTeBJ1pbHGRxPMOJRRQQlVeCh
E8fZPimdJZSAHjiDkkmOYju18/0KavddQQMSBkBzDCNyzE2bajz3c5KYMDdUE6gL
zxikzF0hrAQRddr2GMdI6EX5mZk3+bxQT68AuThvcv3DrSLJFyt34gCniFiWS5xy
w/m4TQTSKj79byEriPg9dXKxNwJhZhFQoQFqhISzt01EFAaCaGhb829qJ3xRv1Bj
eGWevwgb8tBZpDTC/AoSAYHDGvQ88vXyGMSyzawpeXX7ZqEXY2FNastXyoDF3FDV
Zc1VPS6Clo0YxAJyPLnn27q0WZecHKz2sAkPHNZocom6ty9rMWhm7gW1VG2tXhit
Ulk+wlsT8QJFWSclDs81f+eCk7CYz291xHNhY44LQRnNjbahz8rctc9gXRbXnulb
imsDBV1Gv29NmQJmle9vxcNQswwug8zgILAzOfDaajqqZVDHdX+SdJrKrXgpKDWn
daGFAeZeu78IFfXgInPc85yC+oy7pi06xl/hVtM9K5eWwxmIeCpWoKustck2LwYQ
pF1yl9WjDoGQta+3Qd+Fye+wCHgFEUfoi98MHyaWxinMwOVTQ+Kh1+HYhFhWeBN2
TZk2r/jKcO5yN8dbx6QEiYeA8Bvc7+LN5TrLRmhM0Jrg6fNmoXp0YtlxF+Vt0fXq
Bas/QI2EXF8iHX8GoTxNBIr4AYEbEIw7RxHyUEQEVKhFUeQUoL48W0wfQQdC3OlU
fQgULIIcy9xpkQbSemY9n7pzI2s409Mkyxh5VrcMYM2xKY/Ku1ua+ipL0onR+bDP
w6dF7hE+MKj2V1k90kjDg1bMA6yiMeXGgg7YIA3T7F39BwC+d5sYsuD2ICthfT/S
CIc7ilBM4iY8Q0pZOyPKibBXOVwPbjo6oKuJwqcQU1/4HS+hkC9qwzAZ/6G5+kSa
9nGuWywfRvYtYkV1YXu91Q4WyvS4NmoPHsOhWPEBeiD6eA9dtv0MRzQUouvlr7kW
gB89DAu+yShiu6wp21YjYizTWt0LKBRZqcF+OySqzP9jvoO4irXq+AG1fGhskrXR
5+O9gJcIa4WUTu2OWLEDjqA3k0imqpld8zl+oq7o264mOmtZLaXyFqNGY6hYNCTp
7tbItViaOht61SQiK73uTxmTvbr7FlAIgVFKXffZhUz9HO7M0uY6lvn4N6d3fbLG
TYOsKJsVJEEbDleJxX/3cOLMwE5/8w3o2X0L8+QmouvrcsLxCO+nVzzxdSsCkjso
iWJQcWqTEJ4TcueHLRUJJHSptW3nAKtwQ0PIL6x01lNiHI5dWMdHcomo7CGpxf+F
mOrYl9lxRRwna7B06ytKd+rH81pMs50cv/Zyb7aN0LGLX8MngvncbpPo4UhVCLDZ
MMEDgSDNSgd/vFi/zInb8piQUOX3mFisoodFh+oFSA0uIU0GM0T5FWpzBYmP4le7
/pnfdAWSshHCVj59EIofarr7htFdWBT8kSwCZoz+0azN2bG+luyWDx2vrwk89PKT
JfmMXI5sIQNMLdGsX7TPDTbaFB7NKLvWzUS39lgexqphD/rZWq4im9iMlKV4WC4a
c/3V+D/Qjtq0sc1NImG8DCw1tZwD1+gRQJaWY95WFtT0hUIswdaDTWZjrpT7L697
ypJxdzW4dZC7SyZl9Xsv2oGBW/e9OThtxRJ7NG4+PF3x90P7RFQwxYbO0JsdhTd4
tlc9E7DYDK7K7IoELabeuwXNBgJO5OlBOedcfW1HsU+rnHvgZmngvWtVuX6kKOlc
RHMULJgWaNNF7wfLmpvLIJDUa+oO4B+u7quagGjmSRDjiRpqcWZ/820up0RYhLmV
K7ogWe3aX0EanxCESe/kBpOAWN0bvJG6k0XopyhP7TGnEt84dYXdmaPNsKWJU8GO
Bxl9ca21RbLVBbEFcl95t0XKKOlsmbUihGdPmA1tfxEWwPYQhD2R0RY54w1C0KyI
SqoCRlw9QyDaNtXmmbzZhsggpe+7AGIeeTJFRHTpPg3eXilznFLpRvkNL07xDrVG
KbwIyRSDIqwoofrQDzI8p5yj9M/YkIS6GRZ6xjS+wHVRErBoaH0rI19DF63nicJl
G+2HhQloC5EzxEA41rZPHvhD4U78gm9aX7fqHxAXzvnZEVtps5l9EHnMPiipInzn
a5/o0UHf1iDE8g40QMKaaSVuTWc8MIGEpR6Br47h5q0GJMaAT3/KQ9QzT3EQwry+
crmX2eVfxVZ69x5mOu1UNLbXffH/ymSd/Ul7ARO78m3xh8LNzAJXV4ooVizfRff9
yvXc51Vb2szzs9ljSJyibTwpYjpQxrcAMKIrv5eog4aMEJhPpceBr1VEYqBSgW6l
hAnCxIFWwiac24UWzcihcR3XUtr03O+bluzJAa0LG+mkJQIeKdzijhfLcWFdqY2F
7piQzoVl0gFPLx+ByKSHHE8fd2Vwey+rUevys/8gxtSF2YFmsQavZO7ILggFFgp0
rWwwuMJK2e96LLGAlKPl5L9ptacgHYUzcDV4rc6QTjZd1X6lZ0fb8cYO7cHrXs2V
tHkluZ5TNieRD3B1gBA7fFxGs9x1bd/zjoKihpoX9GPWL5erEOmtTHBYWT+wUEUw
u1JvYqNFIUOq0FIQw7tPJg1Fis2+aRIiXcV1ppDxyF304old8aJJMrvRXcm6Zh5o
HkhEQES+1xBOOSkCNH6WUUECwLaAvH32R4xzfMoy3xU+JBC3iv1NM6bzgXJ1pC4j
ODGVWnJZjRbhHK5KgyaGlv0NjLMNrFfmdGVLGoexI5h3k+17yiFn2cdwctc7tMmV
Bnnc2xjRbFDrq9CVHY6D/1B1PGu8VJ0XVglCroIzks2QzOT2SCZQsobMrnEOA/eH
v9i6w2wi33fihB6i+lyGq2WHVZ6nq5RGzfXcbxhggOcjgEvwcG0wHA1IMPtKAAet
HbfwUuot92Bui1kbRSiTiVOGcG3113bju0XrwP5oKWiH3E+E1V8Ebk2FkWLDHpI8
+H1PZIH+RFm0U700AGUXUuRBQ3iyu/YdZJzqrsaxx+7DJm+0jNV7MG1+lxsJil27
GA8czKYCSj+7e+wovXCxCqgXFTOTyxx3XpS57mKB476VPa+GT+86Xhs6c4p94kI6
jOWiysQTjSzJ+FU9BQeyanSCVYA++p0Eu6txxlXNJflGXuo+hc+S+ptrgPpRnqT5
qULCMQeE6yfzBljiN1af58sWkkWyls3mzk8cXhvWxzIQYcmLKKt+DivPYBvf8FGH
M3NxoGq4CQ9hwYCCqGpbHrniX2ZLfUw5RoxyinBf2c6x/INZKuQw1wl1FIrnRGki
7G/yk3aTLcKesnl2Sqh9kNiP2eCBU25ifUz+KypjXy7ik87ZTwgpt1WzxUIJ8Uge
T9bkAhfuq+VaODRUzwxaX9e/42QC4dCXpMfAXnV8y0HsGlY1wcf3jXxNSlby2osX
/DrI7+x1mgHtZViWM+RUiM9vNuH/AQITyfV29qxcqHjRRlbS7DF7qwJ5oK2+9aiP
bkSaik2eS3Rx7BfFF/VXqZw33JOgDzda+unbFMH+3XNJgGTPfKAIjDvR6ZZmR89K
4kj/TP3a6c0tZhXH+2q7cS516G5evzUYvh5shLo+r3yQV7SEb6N2KaYaYcm9P55m
QxNFoejmF0w7pLOp5V7aqi2q3aigOzjBXZS5yFskVXH/31vSV7yL64NBmqbAV3w4
HfShkKhnluCSI1Jqw/dq0UZ8idSMcpg6c931FbhoN+6aRh9TMxroMeee365rAEsc
HnLkztIRQXuzZlnmY6VoWQcrbSn4HKVs0qq+8AOv2UMvZLLgPFhtA1SkBOSVz5nv
SeismT95boSr9c71AwO3pzLfC3dlcNdZE4/FXcy6SAwZiP/kRG97IZkIQiSJgvth
3q5nyuVzwuYqMfOJNo+Pmg5WgC2WiM0bRCF+9uPHWOW5ShFnlCN8T9AhTx2HJ194
FX0n7c8byOWsfLQdxrp6v/DMmi5C828SUvuQ94IQVGeWysLhN4z167CayLyJJ7k/
mIBhJYeXZT/2TP3DcDP9w6lddnI2RbWEpM4l+UlYg/yCEREIpTc2PCR4T2LSeVJW
D8ijlarIA3cM8Mu53fSkkGCYzh8rx1fk3Dl3cDrnS6ZEeHfaPaFC8cFto9pLVtCB
k1Vnt5crPh6xIINrFn3kuF1t9SBQNrmy1hEmJYpPQayIFMtUZ9QpCMSv+hU9Xy91
4rIq7DWk869fzaj8O2NjpXpuVc4nYJbLIFrhLhUZFNVkV8JF7dZNTTnYRxS5N4mr
nTfhq6x8sbKIlqNPlubUuXBlB4+fEuWx9PWPdtxnxWi5olyYJ0kb9H0LXoJAEoUX
5jKJfmwzfBHlDR+Cl1CNbMkMIIYyExgVyv4RRYKkbmaUxXklyE/GktvWz45iozSw
zAP2kTA7hOoUt4dv2wLnPhvmFw3InnmoaWOL7AD2aL7PjLjwkJfQlTQorNKjKaKd
uVFFQFCb8pW5gP0PGAr9E5SP9OrvMX/2+09SejmxjzMYJ46b29mwkqYB5z47pa6N
bo9LYTi8p2mMPjsERMfDf8PCaaXin43eDbWfzGvGzxiX3b9pORdPJrXw2LzD82AX
w2f7YaPCLSv60od0o4nJeyqJDTxzLnmQBjULjjYKlQCyMaSnGSEPCsjtS1uKuTSU
hSHvqc60hpqk4qwJLQcag3Ty/pOzNSae9y0ZM6AliC09WUfY6ds69XVCKYryr6Eu
umeb0+5H0ZBN6KvO55a1fHJrqfuwCxwfwt5hHMWYDk47YEU+4ONO/bZUNLguvHEU
pDcmffWI0sU59h+pSLprJVVpdZDnfab8eCu4weT/tWZcmUG3IUwBcqT6vRfeh+uh
HvqPSEk+Dk+61IGjZNBiwmXUaBqzAJsuuG7pS0B146FSafi1pbNFC+AUKrPKsN3D
KQYIqY1apAL6zi2uyfdkHrkJGyFIVsZD9qa78q3ZQA4k0eqBnSwgVIBiq03V9ZdE
7A+Po+8nao15AHn5/Mr/BLndhLQjlKH+ScT5UwNKaYAzx1w442AWY6xro5DgXFyN
VSrKsi8DWRDUkASklegXrX2C9tGHkrFhQNWmk0w1ViZgF3z1ZVCGhu3+j793loW6
/uJqf0u5kd7epn6dIh/vJamh+s3wEj0DfRaglYORK5yDq16+XWKzqwlYtI2TIcGY
una4z+HJqsGqZhvr4wCCVZ26CHr1SjPanbfmw0Q7Suut1DrBBc1m98BRRfmM9/3I
unn30CC+b0ZWMYVBavbp9esTmLbvsER4wrJBAZE+w8YGrHE0YiBTCPzB7hnL6XSd
YM8k6luZE5oZiYUAb5da5adANVvaS4Znxvgcent2DpykM4/SyU+BsDlsjpAe30iT
JupgWKyqmEzvXLh4Wbu5Nbcm6aWo1iheH4zL0fJuH3CP666UlgxBZ+pz1usQdatx
BTVQnw1NSu5XX/TScDjIfbFli/zMPiq5SmOBBMNxku6mvUgXf+pnZPOADQCnKXk3
yVGjMGnn5PTIu6NuUHGdjqzU+ZRoM3ab3qQlwOlGwxRRFR3Qm3Sc6BVcin+D3lGh
X/n4GUwmaPvNs56/ZwBr5g5FBpoAMvl9IDDzcSzdTqN7sYQDjZev96uG7u0zG2kQ
22rrKMlqX9agsK97BxHmHDp9CFTqiKn8EX06EETiaZOA1yjXCjHzqq6GgqrUmuHl
CFKMF7A41MAuqXbSnh77w2bQpnl8dTs8nrpKJqwsWoh9I2sATcLwOvGCoQ9jKr4c
j7U88iIZ40E3K2tsYjr/4fQMsVVJP5I8aljemwoDqTzX9PEesuZS6xOzQoeZfRbR
nw79ctdbfKBLfQZAqqSsfw2niRJOQFdEVos1WRe0Dq0s/KC0h+/3rVORk3k2Dx3x
Tiaib+RhpN4QuUS9iNn0nBZ1jBoEJK1M3NAVQm/zQpqYsH5qBo4dPfvvtCnnXZYv
adBEBp/EKWMr1zJI2Y9EZvrtNyK26qqdRnzbDitlcAG2ZKLgcTjmURQm0XHFYv5w
BW3bJvKqKzlzcyirtgwj0LvVamzQDF6jtqfcmHFlriphXa7VaBZy279kzSiYPTjR
lwYp1GdCSspcd+v/iZ/Dpolj1SPgN/6vZGFHOlneEQ3O79MXDuGY9B/cbfK4lqTE
95KpNM/x+FTvhh4vcPcdVlucc6xbDF7CMSyn20j/lHO+2sG7WRHdH0C9EsOZnFNe
foAKWinTmEYUz2B79Q89V/E+yRTpklR3LArV532pYRJf8GzXSKVv6KO8rFqZMCYL
1/MgTGH+lYxvSURN0RChjKFLaUhpwG6L4usgLFDDjAoM7QajxBmov37vo5PpA85x
HxAvgQsSHfvBmTFV7DUY1rA3BhmnZhCfOuFmbSg7YjyUHvf+Rz9rpz5ZncV4Ix8B
SMuFri/AhukTmZEm/73ma59YUHmeUFclB4oeDoYF0S8M25Avnet4EnGWUvg0hUjN
uMtItubtu4vSjzG3Od2H2RT0Cuz8e67nmD1vyobwqOsSXKiH9BW+Nl2N+ANCLaAE
Bs/ErC6tyz2C/F+M0quiM2YD7Z23sLcGOme7RS9/CGWIHT0TDZWE7AclLKWm/ujI
jd4hvmVuP+KrzlbujskQskixMIYZOhTsiaJaKBS+HP6ztpHbr14mWJjgfxeKP1fT
WZd5gMCNlgNbmUna25knMfaHB+U6DCPAkhTXwUh1qjHImRQm7E3ZFsoirsMgK+FP
JMDT89AvjEz3uA1p1d+VvZHp71M+wieHw+2tA0jykuB1k4ulh4BEMxM5svTNEaUi
O11hgqdRobKe/oYUcYPCszMhhgorxODJkXRpfoxXkfL0SEiCdmA2pXbtkJl/BQeJ
OeOZcADJjv8UIutVKlA8qirLKKa8NS+PQnyi4MgCfqxQ676/vEG1beWLnusY9Xpn
hEsNVjBaW7Hyp/6Lr+lBUbdfh5u0lsVUYZlxMDcDpFLoL7ZI0yoqV9fX2TZlx5CE
3SKleSiH6RQ2Q93dyzeX71BbzOWlToBxDOon263HXUmIEqc86wUOzmm9e9xNeB/P
zvgc6W8l++fvDHsrCns2+I1XJKMgnJ1dRAf5TtdKbutg8TVtiQs2g+f7SbwxklO7
FToDigOWGsKMmE1beHekn1UGhwyi2KOVkY8XHrumNCSxqejEnGXWxfuRyoxXiTzG
tiWARPg844RzLFQ7Iyk5T+hIRSpBZUPMCLlpMccNbTvYlf+SeUeavnXHW2QeU8mL
iqIpHfya9W6QA8PayNigcySBjXThx5vcfBg7P/e3Yp8iScfyXbXj5O6hxwg1S/a5
WsCVP0fmuiLqdC7ToSc3tJbwy8NF/r9+Am0UXduTPOmI4riaH6qN1ulkgHtNmIwc
TKZ1GaQjvqoPTpwhCFCTE/qtCH1tKcG0CuW6/20o6hCED/0fuO/9ssfL3IG8fiW+
CQR6pke/bUQcqex99X8T5tEKHMmO5BQX1TEqCZlCGBBUUrCfyzwgxnjoZXGUkEkt
VEzpuVlMh2X1HHMDZjHYg+WSgYvwiPf8Ew9Vv2WZF0s5htC6HfW81VLwRyz7vwN6
7JHoD0mKc82zJiaqy5BfZD6gP5vwSLh56G8F2omOihDlc2HUMNVVI8IGxrAcaxvl
IcK6hjUwDw+nfC9RAFVhOtHE6lczOTqXHtMl8lEHo8eOet+Z+2jleIe+AsWoc4Qr
lYoAnVg535z9cTTIPsrprT7C12AEhbB2JIhtEknICnUoOu6N2J6t3R/l3YQS6eb7
lR81jQkItzAcTAcqq5zENUr2aZybh0ZJvin1nNCh7dA7Z5SlEvRUUej56PZOJT3F
tM3rKdqiJbhTTJz1YildEmFuBvH2Vo5/Ob7jK28ASpBp8zitbvYRPD66SrORE9F7
4BO1zA4Vopg8R3EtDdfFzPtSZ0dwlxGTIu1eqKNEaejGt5u8RGqDMN2o5JNPTn9r
1ZhYhyzMiqfonkFhg/KWXsswW4Cu6DV6OhEjgEJE79m1TM7+CZgipufsrrX96IS8
3MonvvMvjDhF/xVXDl1140V9khMpusf8/iL5FKJWqgXlHvAqekqEK1iKoCCzz3cT
2xS24tmihBsAKPdBU6yAD99au+LNC9Ve4FGIZgR0XPMsFk8ubeFSHjxpiKzdKh9k
bCm9ILqNjQEAIy8iXNHkD4PqSpq0CKkqSeVK1aYg1tZE1Ivnhp8pTGDsZNVchCaQ
6BMcsBf8swVPjIndUxEdsoLV499MhtrP4s89IXJ/p61xNC3Bjom4DXEF3lXuihq1
kGbhO+1TKy9WBBxP4AfYhnQ6NZsHswEXmBSVqq2uloi+r9LrzlKB7YYinFLm5Ms8
tVDblml3WL4f1D78+wvD9t+wz5wdi5M/iZtSi9tjF4JzHXLy7lAvhKIgYcenu9OH
Imtp6f0Awbd69jOEKwgSPYqhP93ixpiXT1K9V9ZSvuusaz5C43qmA+mOss+vhfiM
+wfN8U3kLmFHjDVXkMcZvDhLIz20DjgHwXTCmiWDKTrGsLjRs1MSXPBLDEk50M0f
2PwP2szdt+5kTWGMJjt1+yFxrsCK0J2tdhuGwcbeuXg=
`protect END_PROTECTED