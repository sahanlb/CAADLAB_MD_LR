-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
YAkhbRM0eJrhHkwhgbxDJ0HGimoUut0QskQ+wuuHjO2GLwmNE5LGDyuQZm7wS5EP
SRc6XKzAgnAOfEIwhztaSfmYeWoh0OGnji6e/xFD5beB/0zYEW3/08eRavmnDfAq
I4BFpukn+Z1qk/rpiSAO3pnjuA9LUevi0kJZTQrJ94o=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5472)
`protect data_block
UTBiBsxwTr5xqBvTqMwm3SJffohNYBvz2Ygr7+2lPK82V8meX8r3e3fCKtBd71Ng
8zDuWdxmYFfS2nfwo07XzjU/UoTXWEMC8QVNGykgVXdWQ+ETslObxtOE0fQsBGGz
MQ0JSVk8w5oOrNmNj3HAONQQ+wF7e1eTsLs73n9t/1e1T8wgkd7TGYreh5+wg4/1
pFDk88kwOTCJQQD0epII9vlU9kItmFLEo7mqQ2qsBW+B8HKwNNZKZD3YJBetniCO
gDMr0BBgzutfy5/qKoJJdLJivaAtaHowWTugMhE0dkHSsrt/+mj31g3nSSJqET/T
Mvdx8tWBN/2pHmgWlkEhAAgW9XUjzrSey8oG5hdYgnmtb4DTGEUTRC0mtyy2Dpit
OfarpmXRwx3tJvbu9y+fjnb147BuIikrjY0F35kYmchMc/56f56R/u3AK/IRNH2B
HKycUK6hspGhBJYeBH2CRr0w3NdZMQ//vXUwIWfAObi834tPcf8nfEZcwXnDxCeo
e/enNSuHJPs5vKB/6Z3nh7oWpdi9Hu213phpZqsapMLTEVhgNXB6yMBAjAm1lL7n
NjuMhwckFa5FxA21NwhbGXyXoYyND7re3K5HiZ4fflLTV5kHh41oJM8YOkzRNN3C
DVUdUV5r86YO1hh1u51j3DryllGLsezQvApDCFQuof98TP2f11AKIZxLrvl4NCiE
cQQqoAC4gHoK3dZX8jV0tXNO3C/o4v+LZGSXHjWFy17Zjzy+TXuZsQJzrZliDIux
Rc4y3DhgYhHH5s1mX+1gBdhnFG54AOF1txvAySVIQ7+Qr39hPv1e5z3Wj9hyRN6V
7mHqSBZbrEN6KtpYibc6VJT8ih4jl7L9n7PHDgoo5UTraQQO1f+RWL14SL36cVMh
06ITHu4j8l0bzWGkRtO3HF0qSJbMRAcY7LyQprhP8yZr0xwOOsYq4FuFO0SiwH88
CbBjBMPh+KI92c+arBdh9qlNiyKtpJKcqUrsX4QnYp0i4yoPdmZ1FrpigXYeXd2Y
fUbvuFvx1EsjCwUGE3GtF7dNRgkvqv2UPsf/bAlb+QKIFnuL9vPqrc8lsb5gSlf+
miFJt388ykUjtA/2EwVOJlpKFpffgSaonKC/ukv/Vf12psrFpAslT0Yv4pudzJOj
FKobCf8aPeO7ZiGsL2CLZBHgMqfSqpgI+3c9dqObaqNkT/8PYGmns8HJrupe4SkM
eSbBRRxCR+4tCW8BqBPjWIseh+rrKyH89ayhpD0kTNEqFtahFu3B7/so8/sAFqsG
eHm5v0TwfUdrrefFZWN8nacRJ+w81Amrjx8lSQfGRfLLvh5mBqElZFOmOWq49blt
OcqiNT3K58c35cJygTFqidNKTioZvJN1cQJlKZC0B4UPxNymAgflr1bB/mPIzwDG
UWIhhH+tVjabQUYPBO3l5y00fRCQWCBvCAcKXCtgCB6dtHl/Gr2DO+P+bhphpLni
2kIyBD5oMdn9t2zdBm2SG2ErFYLJndihWmfKdnXZ64xoTs1iPJXjyxajmzYX6oaY
/gkC7RGH9eabAgad+ME0baoSpgsej7grXttKYUxaqmDzlHjJRHMQjqOow6cvH457
QXJKJxLfS4HBGvjs1J+VvXL1NlZPZSiLEqJPvFiQu+DcIeg0heiXMK3y/fClnEos
cnvesM5p1ivev/jUiE4WcJzdT9+tFk18L6tMbkYN6bMFj27vHCOQ8SNYwt0PxwMK
bd/0RdrivGE6j+rHK/wSduZ3FCaXemBA8/wHZx3QMXX78G0BiNwb/faX/RT7LVpM
Q5cRQo3pP6ZIaa/tHgpIGwynZm/L/oPmFUkqLhy/7Ka7Vtb0KYf729GdJV5tQmft
k0vhrj9IvqDc4/xL+dFAtZV8gbx2aTagR3hZQfq7V5wDpfqnQ7Q2pJKa5jAhK7ar
OJHK85/EFgvTkF9P8RFvgsjPhxwDiGRYga2mAs3TKRnRg31To9uQrzpYy9z4im/i
hCACVuVZFomZd98Jra0/7QSZqY86S67AOqA6/d56bJcg5zXX8rzZnGf1v7qAGUe7
DfQMtvRbDmLGw7L9+0aRRa2ij07RUVtUurHLtIYYQSxrzsJrTpW70zSSNtdGUO0Z
RAEcb/NvP3poDYnpF0yYQ+KO/KWUxz0xqldD1nx7m2o9g+K55TIBxW+W+Oc8lWHR
LJkTA928S93fhW0SDXp0jNzGNa8m57bPqki7h0EvdZUAYEkHfeJXVcyYPqdNxdr0
F8nT/gaF9K7ltAw+FK0gjrzCOcnetuOmnZmGp0bvi9xRdPSmWn6Kstf6wfi2HJ/K
iWlIk7uaFr+Q0IKgJK4LEPAb1VuH4J6rgU8acXiU8WiEprsSq4nhsjEPXljc8VHA
URVQBSvdnLEFrjbLTO0CwVCb+/zE+0WVR2pv+LDE4uSRCAELjvm2nCSqF+jsV+MV
7A37ertWCbODNLv9l1H98nhstPKSzvsWF71eaJZbIw4yJpqvYzX8OoeUXUga2BsS
317bYgNp9jpcUwaOB3InhfmgFPUFMzgg8HVj6N6hUEWRJkfMgRr9NEjT18thi9Lw
7Tbtr2M2Lu/41kce/XxURpUVzInjpcuw7OZu8bXdcIRNXqQFSVAaGMHv9x/SLol7
vrJ3J3qRph1YgfwmjBHKlzezKhHWwy76Ly6Wu02QEnCU9Eg9nEUFJaYFnbV/jd1Y
63NcJywwvN9VC36cyGcq8OWFNGEkL/YAwpV+Ob1VtbWFtS3B3HI3ooE/ITaAZcXl
abCcakglBzs7CyBkmKAtnV9PXOJl+p97bcpN1INyHrJO11258cppOw7hUDZ8V3W8
XN7ZaEMjgqJ1uv0bTse95D51UasuxVhTWzc6mbmF9NyuRJWm/dF3bFavhJ9AdGa5
Kk47G7k6UhEQzNa69DjLGIAc5Bf93lUxOkEerV3vzHSUz5iuqY0xHcMIQmyuwZ/U
3Ab3K0lqGxCNuBN2EWVFnwpKDSHVdUMLkvUK/MHYQEpzu6MQqLl2Qt59l9zQwPat
KGulV2pDM0KRwgaIdnWg3zT0U62PWas+pDXXsc51EHJ6mW4TPzV0GMrLYm2Cz77b
GeLKu1rWCaDufN7T44XznY0Ho9/EdJI5rExDI+TWyjI2WFO5yryiljugUcwlqIL7
8JCpCHrf/MfHioPCTwHJD4/WWPpdm03jGfeLbeo8Ni6lXB8s8HqeEyn3Lz2bSClA
tk+sUbpO7C1Jjy68Dzmk9qD1aDPu6Rh3xwIc35xhtmmDFjuAEVUTeXQKmQdL7+M5
Us04A2ed5SzRWFAUwxfuFrVFdSKHOPIZaiQQF2U6bmQKztwfq/ado3q2yNfrso3y
TfF8JF4qOVN8ikxKnA6ghTDVuW6HXjOyEt9kNElIQfg9fiOsnSkwpAZmfUfGAy72
5/mSE6ivQBUPSx0NRGFDLaXky8piEQuiSs5kC2g4RFlcu2WT3x7aroLAv408oGhp
v48yC2JqGhnjAsV34EdUvJlGtt7X0fn7XU4yhW2NIhEPfTRLdfqFHbTsJCPiJ5F7
rWxqTIwdrqBBHmZTPR8lHFINTuLoquDjs8OSZ9Z9ds+LUvw4zIEoYlg3Qn5k0MuD
yEPv2807qWIcSgXvg6WRVRiYdlH9DpM/dpunyj7RSbZNwa5ht0Ke/nDOcNEcRBiS
0iJFEX82IV2onYQQtB2d0TnFm7ar/R+EkU0iN/Fvy9EaXDKZ8GSf1qVaZmubAv9S
f2R6APj3fSdzz7k4wgXCJuBsltrVTLQHcGXNp7Vd15TAC862jhATxa9/Hm+VM/yU
VEm1wYbedZcuQ21BQQePrGAqBbxnV+ThS1nmeZbrHupRIvkMTObTnePCf5pk5XNN
wSD1nYAwE2kBqQjSwALnStJ5Rtja2wvvOBIK5X18hkD7NIgzVmVALes3VikDXh3H
I7sb8mloV5cbVzcX/SSRJac8KXgw2ql2+y9tINovfQ08sQ7u1EScICel6Ucg4z2O
g6SFTsg1FRgL8VG4OKdgDo/NuSXqkwGqCLUfW0TWYnCoF9eX+EaPeSlpWJNF4FIS
QphmwLY6OB4+6pCkN1w3xFhuBIU1V1caZ7zho+9oixqsGbEj7bMfoGuqFS0tODjq
JIrJ9fc/ApMDLOKhpCDDGnmX+K8RXnB7NV/pGkOZlR2663qw2vT91HYiwDc7PPEo
5RzFcrtBtV4LnOKJAmBcZZCHya6j1X5wstPPQQIgfLBIyyAr5SLJiAA3EXycE3uZ
ORvtBBQ4BLEn2Jmw/RCGqAOw/KcDeJbJwxBK/Dxn5Z6VnVQ1o6ednrAMVt/yZaGL
a0xwL+No8akXjHNZ/meQzLj4ntbcUeGiVz1fEo39083YErbfS/643wfbxLC6+eOc
lwOS4ayZSGWXWQhzFqDje4U5eT+Pdb37ByAnkqvkv2z87JE8cW5xcvLCGSjTYaY4
6nIgyRov3yHTltQ0lJ8A9C5qO/j2xu04OfxjZcVW20wpCG/XgTj5g1T88VQ+cHpb
85UiVlwzBOEORFNijL303QGnMtDjEDjkhQUgS3QWvOozIYE3m/VKaGSokDUAbC5v
Z/+IWbIC2pGL5nzubDQVD6KiCmJjr7gNA1sS3rZc+6x61EQ1W+Zf8eRMUIEQ2a6+
h/LF0p84pfTf6qc+fUfR27W+OV7gLsleizr6cuuTahcYSi2gz/xI6ofiyr8wUoYS
wz7f4/oRin0JPK+hvR7OsAZcHNEKQKtMkyC+iFkxlUZjOoiv9I8Ux030c8b+FBUY
JZMW9fw4k1kbj5a8yQKzAMmg4/ZkDW0lEsbFGZYIwv1HP0MiyMaykxgDx7csLj9g
iP1v2EnJDKRNu+5wLA1Urcp7T+MqHETnRDXFRLATHIYTzVw7xCXBne6gT1TZB0Ke
IySQfc+OkAHx1oi5/KHgSacFzZiVwIkkXP6aURqpa6N0W+MJHzkPrKpjVMZGI7qo
OFfI4lUHRZQN48+Rb7qP1TGsr04rnWxRKsSs//iG3EUnd5WCgxIdQsuY6Oiz9nUx
W5c2c8Nwm/DfDrXwIq37yvaej2nc3SWq9yrE7ob+n+EmYhI2RJ/P9HTIRs95ZHrz
d3Y0YwqahRLRUsyB0UJKRtgNymtql9N4RRQc9NhtsSWT3bHdhpGDouQ6wjZgCC2+
3BKSN8NVQck3uxOuAqsHp0N9ukQX3hgbqJI+65nGsyIZTUhkZ+TA9JipzER7U7Yy
/uElbRcCBNrrl0UlQ4LGtR2Tf5mW7s12nrb58FBEYDt3v4+bUygsOv/O7dH97eDo
Q7tA9+qcNSnMFkGc/qjx4zSKf7QCRiJGI5LWZ+ibbe6bnlgUaDpizbNXz2TJ9wyi
F2HuqNAYCN9eK94jOqfynJlQnTtM1kbW1Cunc6Xvm8HXg5hYX1lpfC0Ja/JmYx0J
JR4PVT5qF/acNOe01sAaeDebtYCWyOCF47XWkYCpSEsp/sRFaZn9YWxg1Kq6JsPL
Qp6B8a1Le/LpdMIGk+KGT2tEgEoNJ01Oi8OPaZu31CCmT5Hai/FfF6/56HDF8wLZ
9yyMgNCQW/WU7VGuyC2bCCTZ0TUAEk8A0W/FS/OJxHj4i+PbjgdGpPqj/DshVOn7
uO01/lIKlBmSCwszTEmi57tNpEVnLq4XFO574BoSYKPoaaUIHKLHdLalXyRnE3hG
VeM+NdLLInPWn3vsKpvTxzGg9VLU8HAu2JWt2ohw77+BjvNHRe51UVrU7MryhCyl
eISngboBBbiCiXc5t7QWaEcUDRpR2aHzi8z19piw14Y0NwuwOaVxaUPqadMYJ5DV
o7zWIQSwV+2FsG5iaL5o3EeCeLl8UTBu39QmUbHApghhKIJmzfnUyUmz15eEUDoP
hSSMJK0LSZV+S6FZHPnpqKw5uTMl07xsoSkgqtCFy+OgOKhWPjjgp7tIOZjXl2x7
lQ8l2G0Funkx0s1TvhHIrf6uAaNBeTNgiCWjxEH2JpT81VIyuMIYAummse3wiqPr
u53ezYvsWcXMVq8mQla4Hps9Obo/YBXCzmc2NcyUaaFM8MqloJ5LrGQi7Y/jXVys
PiPwrNZh4XtYcl2rxbNRapa394SDshANSFtsOrqTFu+UKtZNa/37uzSdD8sXBhE1
GRfPD7+MP6/PI2k2BmAJ38P+3lT5MdGAD5CxuKYBBMj/xUkSXNLuI+mF3cBXTuWR
buNMO2SgCMRZ9mA0417WuioK+jMIIrUphHt3IekrnqS0HR58n/uuK9WZHIqSE/Lu
ESUkWp/qiw5hRqRMn8ACY7xB1XBQlDtPhkhErUIeqWjYMZBqfzWCTW1+F6C/jZQb
LIXfYva6r80mdiYl7c675K/huBff7ENhbGILGPYwj09KGYQIyaxsVC/j0iyI/tTy
oEKag0kr3dzh66spinZ3YKhB7gMTXSadvNk+pocCDoPplvJU1fdneCpjq99GrFw6
7TW0Ey9TKg1+5bMlNPlzRN+HnY4TayUkgeqKcYKMPjqH7YOaWOeGR+eDnwMrZlKW
s2/0tN2d0xy2SiMSTmTOmCyv/yCJW+Nqjpc5JkaTHeklh5d/FrokwFLWqw1VYNP8
NUDpBlIKyxgwKxJ2QOteKPFt4ydgd6GtOR9T9164vuBCc7RKOkMJiSWq3xFPpJJs
YrdAYAcalsTeifKraa8W+7i9NZMKQKU/LcrkpZ/PzabEuCxQQcIUkEjVuPfoN5Ks
0VdR5pPy19kq8bRY/Sc/yKy6F3VvdsymCIOWlRZar8AXJrDk6VqLOTNZjatpttcU
82utmYxvYP1A4dB0olRPpc3sggSfU4YZlqL/y6dkWWSLuLiJadHgwRv0QP7iMTdG
FkcAecvxKF5ictQ1yi7sThsh96iLWRwQRNPQlb48CLUI+9sE6TVmtV9/9q8xYAc4
1VT9Ub7LLfxWBhSi3zMKmi84opY2vuxVnl3ubbTwrsYYqlp4c4nJz6VbpBwUVvo/
z/4Z9/viNHQetwtGhARlDZR95QlQcbn3O55PyZ7U4XDwvVUVq6edUXNj59MVOeGe
qgLAZXhbssXUd1CE0D8QkXqKZwPnC9vGAkv5LK6BU4TF/taTjbC+i4+/E1sohIIC
ZZHPP2YXk55n74DB1J3mFgcpkJ2a90HTHyyV6QpXpg92ZuxdsQERD9zykao/zI0e
zr+GIznTJ5+G3EdajtG2qMDH/V0YIwdeBtCLxgQVGGGBls/MPgzC4U9gc1NWVgX6
Tc2Er5clG3y4Gq2eXDJsxkND5htJv4YB4rOB+6g0QdAJhGDz1X6eWUmCMQMyp6Tw
iNOJ+h6VwV0rLvuwuyA73A1Tz5s1zKOIazGNrQDAvpHXMcuXrl2BOSR1FSTiVMYm
`protect end_protected
