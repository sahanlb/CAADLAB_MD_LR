-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ruPNY0B3hXdH24rcT/fmBuT+6sYYuSYB0Gb9y7YTYyufRFZvR6q12uZmpJHXbQkWzoNrRXez4SeM
KmldD86VsgPDwlBpq0qUzPD6Yc/nFcT8VJFQuc+KEGbmWfON5cxP5CZpXXuvEcshMOYh8lOek1ko
jtatLsYGI/akgk5rGujhuNej9Fp0NOEjDArDuDfWUtzhx81HOlojGeUPW+d1es7tbep0FftyjhnT
nddfyrCt2/aP4qQPMwbXX2jE0TnJ/LjAVY1H5WbYrgZ62ykDQ9D/7SebCqd89nwV+mruMMk1Pfjm
sOnPssmx48EZjXAZWf547UNqYFpYJGhdDE6mVQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1680)
`protect data_block
BTPyMvIYUUoaiiR8Q/rSpL+kdrcUXUl6jqJA/m4MaVaL54ZYDp6nmPG9IgK7+uTXPEGCQQ47sUn8
AwCDpvzx5rfBHWjrOHsVOiOCji/Nl3t+UVcUDDUBxV74FzNj9unCO7X1t/zRc/VEU1Ewxf5jC8EB
3P/GDj0C0bP89dyim1w9cfYhUWg4McPr67axQF7dTRiMFcdbqVx59yWLJplRzWpGK5AjkPikfrJN
y/T+q2ji5i+Uc0ewdMSQG/ikE7kIi/4P+K77GMYO34ErnUqB8lf1s26a/5tye7pmbkPe4i1gAH7W
2kbJb/MBM9PAV1gStsgJNQ5Ms4XR2MLzGIlNZbBuotk/jHOTCcHTivKR1OU3q1Pp6UVRaAKGD5tV
Y+2e5sRgsk/z9xgo/lWR/l2TZgu8PszvDmoYqksYmB2tYS/raiM5WW847lVEk2q1W8x9ZhKXxIN2
XTYaJWSYb4HrFJXvNSVvalNboL+Lg7oVw0ChUTq9RGqt6JYBYOxddeYhwcNAwEIz6gZs2m1qO534
4uSbO1m7rAqpT8wTsdPcRNm1l7rJlr1VQ2hk0GG0jUPZ2S8lzwE7wJEin2QjcGwlv+1VAiUb42gW
p3qr7/YmUf0rFWN7oL3abz+OarWfshlFCS3Ok0iZGZ7VSNpvXxFLybZxiI3EgJpvbKgoLP0ovyBH
qkl/Bz7yGCHwjMvhnIBd35xPoReL/cBZ04qP5ftsXC1c0O8EHGBkZccJ+h7K8Ah2LFuzRWPVHxu9
5OwVdfRaNIJqlRgJcL2VDLdwBETDv/zbeilZdDklPPcFdgxDaM7Ccw3jjrn+CMitce1+CejzWGN1
y0WESDaNr1hrQ1cwZYclJMUuXrTSQdOIhAjSrh4lgH8oncEl0jCcNmhxStjdnyyOKmMlHZT0wflI
AOTgIaRdex+YHwZwzOqFkKxeTbCriiHdh9daW55zkJJ8T4g6+aajGtB7RieDz38IC3XraGW02JzT
Kx+CKfjbzQqKqG091mXRAq7Ix16ImuOIlAOUzL4+q6crDlxP4EsjUOK9BZwOA/peBYLVhIuf1v6r
udffVkNzcUehhExbkGZhkTB7hypCG5IMZeaDq3iXpqmC5hyx8sBxTyvNVqbUpf8tDkesAhXoJyom
H4Bwp41dc01UExL/qBcNVqIRe1TuL9zU9k0Xm3ty8fz7byaqSE3iVUaIYrgyBM85tEbOq5JDhJfj
d+yCtRfu8kn7tAEht3ti4RagxSNPTht9IIQ9lHzNCPoGkJ/gsBb8PG+6ApjUQsT57b9RTq5i6Fg6
/7WonAxvocYJabynAcEe3OWgmmmQ5iWx2c3968w4Cjz2XBDXw1YBmVAtJZo1YjYylkX9Qo61vpu+
eLEurNDMkAxte9lciEyuoRtPReb7qqIkEKa3VIYgnfP+kn+N6shPYFQaHiafFA3Bkb7S44fXUuVE
td9IuKzvkx0ox2ijob+axxYDwBbWxNEomH0thlbiU9X0kiv4+TDuoHRFv3UT94iOz9ABQdDHZgI8
4JSx4av2UrzrcorPbcUnaMmGMNz/rjLCf5bawTgJY8w9HN1pH/HaD6HWgCGc7AdtjVhMEjQe6YIc
DDJZg1c4pA5FJ7H+R0bMpVz8jZVWDmC1QAosUF+i0019GSEhnHAkBzcZL1QuMXCNXji66tq+H7jU
1+Tmt8sHP2GCHvLQJndI2wo8UJanOr/QpXzTdlv6sP8WohD125P/kp42c31caPKvTSsHKXYMidgr
DEfSFdRi0bIx8kJn9Uuk8v88dc9sYtZSFO0vdWuQovLkADNy3lC/XjOBRPA81Nu25WHkcgmsVS4f
SUILLebl1o7AyDyd2thBPeXaTfYo95//lpPgb0c+Vm2hpYRuKxsHbAawYCHYVH+aYQHOmffWQfts
dzwTVZxDDMKdSEhU56X0tIW3E8D+qV6vF7UzErM5+MpkBrP3Gl60JnqQt55s/2ESsxsJmYLSiTuf
zQiHSIk6+VBLPhbFx+QOM5X/Iv6QY3ZsNFuvm9kWQVE8p8ZrqmAHFDlBh0FCif9Cq7s/UYSk94Q+
sPvTmm0YTZ1KOmlPLk9rzRxgFTi2QWdSfuiFo0r7rtny8tUqbi5VsdtlA2Vj3Vmzqtv/7NKTsrgb
8qZvurUlGtg2eNTGxMo/wp3LE57331PsBQ8xYEMKa3DCMvZaIb8zh/kSqWC/mtbjqfox4Yxv4oiN
IIUuuh2t+e5jgIFZlHK78IjQ+XXTMzmvXtY3
`protect end_protected
