-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LrlKV4LR36zEjmDO+O7UJ4mUoD6mViSybFJUmHOy55Wa7Mguu5gR1iiSaoHzwVudi8nPes2t9duX
yuZtRyAXpkc4mcg/+LLQ9ZMxkvucfEFT+YcDp1a42HFNHeL3EtsCCM6ybba9nkFV+UIgGsMcV6yB
fqJle3px6ygTDVnLPlq+xLkCijmtRzF+ohO3q3jBb9Fh0B00u3byW6Uut32Up1kOQD4bKv/PWZgX
Nt0Mng9lzbW/zunwcbCjxkKzLxLqnlT0EysNPvF2U5gqlRe4JTS49Kg9RqFYkfGV6VAWVxAbKB/B
KTdC5z1x0kt//BlBZyWghJzPhHDzHChixLQvtA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9488)
`protect data_block
lFjpYVOaWWBFHvcYxYh7tRIWFK4SVd4e5Oh4BOjJPXMgiGsooFxkfLuGm8IVXZNn9wnUsCZmy2v/
WFZ/h3ja5tyW7VXnnkCx7rqlaJtWiGvbe9NGdaPGmPtBNYtz1YPfbV4s+xt7AkiFuxN9l3NYMlCt
Vf19+28ODYtGQXty0tOX1s/bo30gx6QhQMQwbbU1ocWRaQziIfhnqlXrp8adjv5uR7nQLK9a0fqt
B+BWc9y57Ig1WE9BHGvZjXNC/hmY+KOiS9NkPeh1jcO5qdMEz29cVHSjrkUjdQFuqzm9SLJIfLdk
9wYV0/IvXJWotMCHzvcmeNy0Hr/VpvGmAdHKVxO5MZDcCOBmQSm3sbC7Q+46CIetOBL60e7hMA2g
2SkyobF8LLr1mDgvZSmcztYyfFFEo0m8pu6Dm5jngbqDj9Cy0r7DDCRHBstdEBRmWG5GT4dDu0Yv
rffnH3er2Dm06uaXsqjFY4AdyW5QcjkoapHzMfcS+dIJhBdKOL3UxIZn8rtZwxuKxWDcR8JGhgH0
9sOXBVsSqSFURH/w+0hw4HJk+AW36NI5fotqDsnNHnrJbW4MXz237w5iZIpPj+QddOpzKip5sGTN
jBfpEvIJ4kzVWOHYR2y+bJjEovj8DuRb0WHOX5sBsvX/m1r32QXrqIr/cbGjCIcMM8xvl21sLThX
6Fm/nMwAD8EN4eOtWZpUi7ad/L4xyE5wS+SB/dg5ieenp0AXPu95rk1Y4clgFVvbj4Ng6hJodeeg
gMZzIfDWiZQEqLjgMOyBFiO1OFK8MXjOWOXa4gYssqhzv9Kz+ZK7Noas/WdhL30zEMrDjgxiDl48
epL5iOYO9Mzt0NFCiGwSWMcm3SOsl24txUJnI9xFe3HVfX2nDhdm3tUlVG7zI+lhkKmulJut6aFu
mrtt2/XCZL8M95Sd+FOPjG2+l5+3SuzMXKRvneS0aEci6Np/CjpQVnEImKzgIQb964DuWlV0Ru5p
0ntuwejTGp3zFYEOibNzP7RPzZMv6Qx0ZDIFz/o8Sd6nc9XckHuA4UnNk/l5vJojucKdK9HqZvRa
ugIjbUOtJc58KjCD0ssm6kWzVx8ejtPm3QG+3+MEGbVwtKJe1cojtMz8eLr9gFUE54/lklOg+ydO
Z2KSsUbKms4BxXMfizq+IC9chVcE6uk2Q4vzg3XoUMNZWLjdGAL6cUc+B/tbJcxohKl3r0vqtP9P
tYR0rnpdPgtfXtSO72m+oZnX0snt9KPTSFFhSZ3JBtoae8H9yhwvev3Ussxlk/JHGdCGxUhy6JAN
qHUaPmdVPwtRjqP85jTXXPA4Kg0mJVAW/WBrdho3dH5oXh7l4mgCjjdSFXf+TOQlEuZncXNCjFjo
2RjXRIT7nnjgoSkx3/QfaSUUYIoVLUxBhujiGCJJu8IChpcl+c41yc9cUyqLzL6eedMnuBG3zLfl
FvLG7SOtfVsOYQzMovFSmeQz2KC6NKv0FP5KVBF3NVegKRew2FLImOdQyvkOjvk0Aqa+xCO0uPC0
Iu9R1DK7dd89SqtCvO7wbB7V+iWlEcUPSWHvCsiYi+iLGWiwrfynLn20bRGCVpx85fMkkAVRFp9/
6d1kMQ1Uo6NToL4D2lSyUs1MbTVjyTJ+EAHu5arHStC9cE16OlRUqvBF6NEB/LULg7MAivG5bYce
2qVUYPsIrcdEtN8D5weWmhgmzpa/35kfvX9Swx0y3OcVDCtXYNAWcXoQljd2mVNHdGvPJPWkRDCw
yw6He89j+D1qbASl02st+9OOilVas5sEJ12PiYopp16AaDngCBbZk3cRrZFBy9b3FESfErWuR/7Z
aVM7K2p5l0/GdrEE6HPmc1pFMHCfuS1T+plXSosEnJdHCToTcka3lCtzSbaWH6mgVKGaY2tEdK2t
bbTE+UIq9srgvlB5Do5PKfUt6pb3Xt1qrJbsDmcOMLsvO+JPjje4C1RHenmNbpAipuSGleGbCRzI
luOz0vPm2DZFbf3HRRALrhdyDf9mz6JkCSWam4pI6H5rRRq6O8SlfvULOL1fKuPNiXpOsJceIOg3
eOr2SZEC7pb6mbkF/RmolwbKmBtR+OZWPnEqsA97x3fKe0B0FsUGBzcq5+79ipVaiLZyVJYAX4Yu
ujbhbU3b4hswG6qXs1RwevBYBE4D1+CTeD/PlRUBWI9hRz+WNgTXHWCaWsRBV8NkAl9UqZ+teGON
nAFsCuxsIG/oIOzttj6fyJm5eNvsRn19BtXM6YlQC272g0n+CqqYnkHDMN09M83kE4wr8IzEYikz
WcsICYcinsS6j2qFyEJ77fRGU+gK0Rf8zAFqg31HgsjmB17jNcZzXcrhJmntmsCKuYulaebpII9R
lXdK3+rzATqToAFBzZkxW6qMiprN+dSJg/XS8Ed3mcvOHSfW9lD3ICXQRqwDCJEvX3hKAsVUpKzP
vOk+2xElZE7OdLkTQFKa4cXuYfXiObYfainGnvQ96JbEyMlk91m8yxfA3WDKt/BeGbX5HPxw/kaN
cmMQK3fDPhKJC7QSk6hr5gvHrrXsbxMJ9uJZJlRaUnsaGqJ2nh4k+I0EXOMZe1WKNgTwnjTisegF
qJvrsE3q8VBN/euuI2g242TYLKYfquRz7iZER8kgGwO00uO+olItYmv3w1OC2xMKj/CjCTgCdlbq
e5owET0vc9bqhlzwenhrQ3uf1Fd8Vw9UWZQ6DkyipSgc3N2ZKAyjXKcl5zAaCpppZ2p3GxD0TFg8
nSh3y0KR+LecHZ4pMIGyGGTU2Vp0QrNaJ7Ka9/1lurY5O/64wjn0b7oVMFp8xEsWB9FmJEPb8/YZ
+E1k8EcqM/BnHeZA3jhqbzIVnaRPOi4u+fYioNZCaFyzYsOBTmMg9KIfNMnj+9/PSAzUDcMe8uqf
ubF0dhUov7qjysD90zYstBgIqZOjUXyvVJ2aMvsKboM1FIP8Em+vYTdFxqut9wdL+EykO1AqiTgK
3zPb2IXfSkr8Fdwt3mMLiCf0OQGxpqFf+vJ1DP7hAl7TkBXUHtqmRqMtpsLx0k//Idf14gucLc53
TXNSpYEOcwQcmcWNF9YZDQU51WWbNxZBM6c8L1NdhKxGoa8lAA6DyGJ5bSyXlirOC4IQbDXSk8lu
X2VoK/ZFoiKYRb0O8m74I21gdOCBfDU2MXj49zw8bPeLtGZ/M/bE5k54JQ31M6c3otrVxjv221Jj
6umc3kq+99itWyXazA3wuAgpbYc/NWT/4OK3pJxM/bXqERSBHFyj82BIzO1AIx8824ue0w/0xvhQ
WqdMileEUeR2EYgwEBGdUD8RHwH/duPtJxOSVtS/nMhSg/MImVUzaFl4U3RdpLeBsm7Pzg2DviGq
U+C4Lk1EUaJflZpx6edkffjfe4d2/qrrEyuwfl6xaAtXPHv1yZE54DAnkGKH/xSTEMkqFgzVEHtL
mwEug/CIxKz9Tqi+8MO85n8n9cMW1Tpi7ZtysIrbb4unWjfvL3DhwSFEu2ScJpwAobSPc21qJpGv
O0+NoMXp8cpjHvosR0qFQzQ8NdcMEXEvyfON0tOmlYpS6/6oh6BSId9NwCXaQu5ULm80chvQ2Pym
q6JAnfoFHCejqzZ5Ls8uVOqZqdNTPk4NZhILVFDTZ5bUp8P/JN68Zx2eUAMANqs6Cn0wR1PAprKM
vm4Zz78AEFkTbah8kdD1gv3scEoM1nm46NFg/hnIDbemeOg0ercpPwNmLvjvU9kfOg6Wp+pRC8zw
mRq8Q51ATuo5aymAGHdwMHiHA6n54JeVvNMRBnG0Rmg8cnrI0fBLZWlb9Bs/UcXWAV9ln44NRRIx
TCKeSCNh5SGaEu1CJeZe7pKCc9wsIj+mSvZex5eS7037Fb/zTsV03qSb2n1siMx7Bl9xUSOt14GX
F6XKCmSq8cJnRozKVwLdhE+5BcgcBUMi50/gR51bqHkM7sg+dJXGvc4iMeOwQFkSaxq1TzdCedYR
lExetN1f+ZZeYqHrLaT9CEP2tJ43Lryr1HLNmu3olQWVEErikvr6R9tGRYmyRBiwXQ8L+nCh+db0
bwwpqRRdUQbTofV330IriZNmlEUXLEQu1zYkpWVqcI088YkaHJ2E5oF4Q5dm8rhVzmnIUMeux0BJ
HWSVAexRLHFz4jLKWGDx3ID6uwBCJ4/WVXxCFZ/pBN3FdwvjXeegmzDyJU+HeAd5MyDEIZbJoMdJ
AH8Vm3JAiXKocMpsKtq2yY840B2i3oEVQFjOq3Jc7Ca1yc5aAMXLJQ82QAJQA1wojfikGGESa9Du
ZtSASoCQyVpvsKzja+8vkJjyJruIsydWRzLkl9cdHC2HcU4QUgi6yrSqODF30ucjG+vfKe0y6l3x
Wkhs5WZm5o96cOUqHVRYS8G0kElszXzzMv2q4eLuf2+LHr7iTchoUz4HC3xvvFzHd/z3U4fMr/BK
d5GUfuBY/Kc+ZI4pIubweY9xJhccPyunR8rbMRWoOJ80/lyDXZ/ePe+Dvv518RWpjzepSKF/KG4s
1MV0On8Ia6QlM+o/TlnPi7Cwx0LreF7MlF582Pxu04YYEsGpZO2Kc3QddDS1xBzlc+igMCAS8pNx
io1lmchzXwHxpdG5lgqXaEBB62jyIUGj+3XoXhgOHr0qXheJzP1XzWayvPD6lqp9t5hxn7bzeSof
vtjKL/sBbzAgqa1Qu8oRsu9WHPBpQ6QRdKkAZ7yaNvfO5yri3wXUCd9d5Tn6tmyp25aGx8Wrk5BI
4kzmMoW1CcD27Dqak4nS9CFJ5kXKDIML6J2+HMfYGynKV2xD9zgr3Cea85vtzjEyPw2uqc2Nw0aU
IhHL46moiDMizIS3+waW3L4uRrZIMZTRGy22m9ewHCAa7epjqNlDfDO4Bjz5Kqs+FX+tpaoUfdaa
iHcFKdDhRFyzAMk6KmtSA4rcv6YoIcHyk5D6zyDKuyNt8/oXXboZgLOVu16AV8T9uxCP+dSG0qPk
vEkES+JQC4vweT9hMLPN3ZHjpEciMPo+n6jF1Wt1KDJCr0yFobaFKXCa4wO7DR7zmTxFhq4kSHDy
nh0MhaO5a7lHAH1dTLw1ZEev4gjjxvAP9tv3FwWmNUVF2JEn++tHTp5B+BMm9ZF2Y9BQZDz4g5ye
WlyUKa8iVguBQPDt0ZN95mRmLqwzvpXtw0g142PnkeW/knXjm4Avi/kCkP5FnacWe7DclkB+3O4n
1mnxFjgrqjH7zZIrcwbKTRaRUawq9K8jBMZRYgAd7ZnZRPBO9CnXn7eBt31E4C8I+ErQuQghW9U7
PbD61zbYjCCgOUQkOzeEIAHuHcYSehdj7JfqV9h+Kcna0XERKTgq/Uu4Na+A+v9gxdDpS8vZCcn1
NmX6ZeL8udm6lQNrqEvbXeE3lUkbYRezkPo/sLCGmA+hySKJVhW1F9KdPUUp6flcT38+U7IU88a5
hOkekfy6jpamgo6oPqnnsJMp2ypXgtVPa0MwFhV8IDV2x0IoMpQ5DVaOdMGdMI0NoHWf4cvdnYMe
KsZN2xae9eS/QvaERDuKKq/q3y3nK6WItHu24tFPJ8jkbvZ7DFfpOWbyM94DN40GU9UunlcGBeAl
yEbMgAP0inqC5mWxb6XFDvYFBAXQ6O19Th9Q5RJX2apY+xCgm4INeG9tD+gi98CDZjg8YESU+o9G
Nt7ZDG5U+dq0lEcF8wKjMq7FGpKNi1MP1MS/mqyKwqmxf1hSNkB2N8TgggtR5PQy/d4GxdIo30tU
QGFifsqz7gYkD5r8og9kNU90+IFhAmtXzP+J31lvhZGRFrpNYhM6ALfux/O5o5gj1bMSp3K4ugo2
PIrV4PwtpUANf9INiW+Pba1qvyrGvMkEbw3Y21IqtjwW2rhig0gJQy90ISkblRSMNd0HJpkQmC0N
5jm5aHFhIIC3Mkyo45JKV2WSBl9+wTJ9bJXXIrJYQnJMd/4bDTTa+6s7e262YTw5BBS8NCkYJORQ
5r+DYAGwBxj/76zKcKtIM+HvcxEQGEmxWd1+RKU4gTgajw8QOKdZWIfjMC1XLQQAbVD5RQuTwVK0
xisYM1JYMUC4luvAc3QegUItHPkaEMLU2nB0arY1D5ROYotQi1mve6eJg6dlcjkS7egTDYG35RsX
VgFbQjcpCHgfMVU07PYs1mqXgsU9SG9gRZS0gA+JcoG8WUZhQTVutarmzG1f4nz5pnKw5z7pCBv2
ggJ/qbqK74NEo9JKPK0apI5wfJ1ns2MNg6Mzrd6rZ8U/warUM7SCCuAC/jTVMsj8WaPbUs62lI+h
Q/dcTNFj1S/XOrmEOMhfVrbKbkXa4LB6lR5EYPU2a+If/ovhy3PTQ2Xc9gBeq4TXQdIC/MDw+ztG
mLSlZEQlpmMv01prT7SA5VMxIbp23WgyQv1Yk1j5oGKQJ4cye4Wk2aZyi2nhK/wQhcMJLWACKFqt
S7EEXbu2r9LB6SQLbSfd5oSwJichBBoE5ndh5MriRQ08grAL51JG/9/llXg431gB68h6gIHAbxP5
xRO9h7HGfc5cppcJCsAc3kgpnKINU7KwJRZwv1QNaLRbFdI5PxniKHA+0u3jt0YTx0anzSF6MhyG
Fw+MpSz57hk8UY073kkJT5uzz/0nRjXMqLZNxv60Y7kLvjwp4LaFQUuiMvekZgJ01fZCEEt37RJb
SXL3x2zGw3CjbiFqEeiLickCtZGvQ11CxAnwrs/CXqI8qNNfwqgoJ6k6olUWNVdPc37lKVmcde/2
2aNct46uLSTKwaVW1zZVqzVwxXCqrVux1InRsdGMz/4uXtG3BawWbB51JBnsOGbBH/1+yBe70RLJ
hv6+DGpCStuLEpICYEagAX8B+HRjMPEAzNNjvzDKjK0cVhPgpVWAqEqq8MFi1pRN6YuQSe7Yx7G+
+SEasZDl5ooKqcNNZfHymWtr2aouqnwb4uOFyhCEzA59GyfvaF75WMtd/Hh/MXSgcss8bU9KrcOV
cmExNCvswxvhqXIUANsRH0gdJuxW4xEsvGGzq+800TAAlsrZocp0IE2zZ5Z9LGKwKyZRxLkfux7m
yAqO5D/9lfvHu+PaPLpl4oQq/MKtqhNE/yKO103s4r1MIfUUQOCLEeKMvRbxel0xmnOZTgtwd9su
C0Z4cs5iS5ocg4M/BtLxZfgIdqRblcplvK5LuLZxKuHBgw7ektCdEgcBkn5ykYfZu9t+6UcCFvPT
180SzzKfSKEWVaS2eYYl7BtT8gdM8fgLgtnM8aMY8NiqScjMeIKOi3pLocAI8G5N27qWjEekbYC1
YNc6XuElFSYCEUNBxtoxO0qf2mgPCQbRBkUTv2fzDZMIlixp8kjr/kNOKPZfr+08lsYViwC3UDXL
1V3xq9Vx6XS5tgp3/o5NFAB5q348EFnVIutILeaJy3oA9oQ7WdlsIc461t9ax11OJJgGj+71lFFT
gv1/Q0KpAGNze3NY8xTZvWWPzClc7p6OAlLpI5koz3AQM6yHc1R6t/vnRK6/CYAy+j5xesYUdgzd
fujnbQv5Wr0B56b6j5y+Vmd/0rlmTU385+hUcom93D2qT8x1v8rGV1GcS2E3U6ORgDqCTRCzOGab
2rSULgKCDio9fAUANKza1G9QhZc6kAtNr8KupTdskOgdwId/Tm0LzquN1Oqqar1xidbzq3huwhoH
k/CI8AMH73bUaCTlXy9OO7vcsi50a/2c4GC7SNMEvu7wN0PqgWm8SC03JqdkaJRBVg4YN/KbfBDN
yX8duI/52QfSR/pybUq+8r3YcdkyqvkxOkDNpyOoXxcMxNHpP4Ny3x2VBc9kqqSeYPOKr0rYSgEO
EFyS5DieQKlhbeG44ZCIbwWDPOrpUkvvbpgc8tX0luOOV0nOSbZwd4HPqWU2BSxN4DaCcngRZ2mc
gfR33Z0yU3YKsWrXLM7YHg2HAnOrUX/VY8LwdrKPk/1l2nurtuHT3e/hyQrgJzrzDkkCbdn1FnV9
iWpQSbskqaaYbrANfRSTOCAnR1wiZ4yAHo7DGtuX6nEE7CcxOCUcWG/GdjfibADvmbNem2l7RPas
dUrz2Iw5n5mxKxx9730xMMHFz+Q1mp0waP48yo91LguO61NgSXdYDszVT5KgeWqfapjVHw4ZAn36
2e48qDFHo5LSakRzC6YkKqBVepjppb88bhSDMtjZLWcu5dSzW0NWq/8+cRleigXgU1KmACfbYcNr
4tPnpXI8AyXgwxyc5nbH2345Oe0CSL5SDzLO/wv4mQ6jECp+Voz7R49TNqbXOGkBIC45zXXYZfUK
DglTU91wmc7TcTVQ3sfT3fuYdqE6f4t3lCXoLujGW1NkreWTvnvGUHFnx7dhHR4maMguKv9DPFI2
ejjdjjLwPT41JjHSWYesl/3kk830msvP43kt5MxZqCq0gjsdjQYkENFj3EbBvG7rjDtYUyubjYuq
zNIYDARBePxRcWmQwAZKO8f/uRdWb6lyv/JzJ24sKWvqwPv+wlt3m05JGG0DLmmVvn/XIEWNt/xl
lVL7T4niPSa0nJlZOqwgQ2jXqcZGzpxwX9F5b0BrLLiW/Zs46qIm+QsWqPCFH/9zPjIh6aPCnl6k
scaqNhd74fStaNyXdtbGGJs4ogUxon6PJif3M6rPPFio2J8moatA80ip6v55sE6iKBVLdfm/s/Ay
pH3SDMjU9UD5boWWekDHznrYaMIakDnTwHBu9XP4PA9PuaReBofSrPbS0+MOfkFGDvxVt9q/woRL
fhQx8nAbza4YVqb1VZGv1kCXMBij6LGODhjlN2MWs98hZAS14v5vJoq1lLJF7Oic6fXTnCkBfQyo
/Ppb+3CF1ZghibfM5ViucdC0lEWdi01WM7yt3Wkqd+ErtYFMt09wvr178TO9gIWAQFaqKCGosUwD
DWGekzN8HRvp/BX9n5SXhI6r4D3zQsgpJ/LgaUhZx2hSPu5AK9f4BNZsXhPoVO66E7u0PwYWuU8K
r0ocdy2r0TJnaPdA4GB6FKa1ctp+Er4WeD12VRV17VaGUW1NOxbzrURlqR0+Z7BGzqKDdSYci9uv
jMrE0wEdu02xBdic06NoKgIKhaiWDctubMRIS9+EI3AaI5dKlkKyDWPpd0vVfI8bOkZnobpADGtt
f0btFIRR2y1BEdijcEX0vYHnLUI3UlIZcqODCskIzkl5leO5ufdZgVkYYigDmXB60RcMFq528vgr
1wE3bFOGjwU5L7ptWgjoNmK0/AGpPw/wv6Vrz+ONknPVkOJKl6qevoYjsZFSh+tRDllQ/e80xsyX
+jTq9DwhYqitYhjGbz+5EdAZ1TukpenJ3VQkUaeS6i2OTTVwpEGWXRYotU960fvvepcJfE8Q02bB
TOr+568u5BQfX76+6bApsEElfteFxuPBRBUsF7l0CUf6Z5Y2ik3i5kezjMspRR5Q7NfLtYu4LDA6
oTD+nNwpIZhm2rA+lB6r7DuD+ZH9molHPbBZeKIQUOqG/iIL6NxVrFuBujarimKqgjybe2bsjp+O
qY4fE6A+NkX6La/3vlz6w/gnmwTLXdDEhGD4Jc3/PHyr84UyNbtPuWIQJVUGo7z8Zs9+HmErS6Ko
3yhOo9AmrN6sR0DaImbNWaMYemb0Hy7lk/Bpkcsi0ALVyNYSbT052nsLVQ1kugX6Y2MIgpYsOV5V
NRaRDfYqfJRD1Q4kxNFN06xed3r//rNY43fdkppMK1foyblDb3AJrRnVEOIEQBlPTJ8jCSsTh2LK
ah04GsPGQ/YMnfDZ+QRlmVjH18u4mqBXFhZ/vnvs2CP2VtPmvOZFzgHzCHjgCfsE1a6y+X906jnq
r7jh3GmkPKawOQLeY7ICp5ttpoTy70TIAwfidvSzK5/G8BoYYdnUeUtTsSyrfxVYgZOkEjlkQvjv
ngm4oLmjvDrh7g/4+kXFyElMyZNhmairnniJCyzWwIncL4XaXcvgmY/r8tzQQP/o+UYgu/r7rxHO
ZesMcaH2lAMDV4C+WAMX1dFCGqcEo8ODalVDN4942un6DVl9gpPnEThLdIZVxiwFYo4YsSQlc0js
5eUX15cPsbtX5nF5Ou+PNmDpH5W+yMde1HTHt11mt7EcLXv0iu27I+PE7cAC8PIMjYwOfTcy0Qun
8790t/P3q2+6GIlDVUUSaocKFzOivWYmNRY0DiFWC7Oj8zqQd+F5cXr09BUTA7AAw2zlBK+Dzlyx
mUBC9q2DpDz01eZKFiUyDnciWO535e3+cby+uB4fu6m3I+iZiIh3B9EMDv7zXTYs/J+ATlg75a8d
GL3fQWZn1xG9dq8S3H/kYOuf10mcYNUefdiKA4HxrZ4domZOHTGo9Rr92KJf3244+YO8W4vjGK9G
6ERaSvXwDW0+Do9i57Wpfw/w1Yk/4jprv8SFjYXSTdbPVR7mFhlGCh7LlEmZBU6gdQv9bRNzjYoX
B0KBgyaoQgBbWS20VfSpgkYgmyHhDhLZVDYgl/eXWJ9BblOrpfuvjx5X4UuLxEc/suVV1QlLClK7
Vi3c3rjyIdKaMZyLbj19sG3z2oLPd/gYtbmePB+kn7rLOaAmS0Zx4QdWIPXeDlWwnjVeYYs/mY8h
PVynetWdiXxQ6VTgY9K9mrjL5+VHuc/4u4szXPMwjZiUki0eIHt/OANSieJFqyvARh6cL5mfdujN
Zvb29+bLRUTxNQDs9DngSExhTexWUlEGrUJvRfrcWx+4f3RQzXS1RUO+oUF//HNX6p2ffo/ZXCvO
H5uIXnz8nArCIPAy1wTzhGzNFSba+eJGMEfv/RCb0VDqbL7YZba3MVxOUCSQp+IOIXolFvxF1pO3
RxLqdMdej0YQsi8DQtutgTqGvW87WGccW9RkJQGVz5Nx59tLeQARorTRUnrK5VxXCiKOE2DK6hxP
Y/umRUvMyKyG1otialeVvsh1/GywRhAilF+5rgzExeVY2mH6MHygut5R4pK32fVaQhPzNGO2iMIg
X/DdhcgaYz+SB5iCJ+2UxQdm1ar5Aioelg7xNITxhNlCpV3hbu4eLrduCMQOn8KUDS4HrdaZmF6p
ltz1L0//EK7Um1nx07p36lcdsgs9A8rV9/hAmrToL2ucps4yKbz9wzdf/Zo4sly2axNP0rZC9CJU
241sw8D6PoUXTE2DMMqgm8GYNPe0tIJ1PkxoMwBwxgGrHuiz1GibKEq/Q7xbdJ5hAY5SV+H0PDIF
iNZEEGUy2k0lJOnTeQTIB7O2BCPcKB29+hMxaSqOBe+nfyB14+OXwMMMPuKGnMpRDDNLWImCCOZJ
xPR5FB01VF2uKfBiMLFk48JBznotf+qw62sd759tbIbH60AiE/C8LUn1IFNFezVFp48ywHrgBXc0
ehbphsuwMnqfjarlpuLTpVmQUNIukkABB7WKzgoPZHZtDj0SPy+Pt/w55RCVvG3Kw/rPNrKFxseQ
eD+bMGQb4T/4TaiQZFUNosMNixK6AddIrpAJJBjT/Gt2gt+KiqX1Sr3/DVkeCS8Flb+w58lgYdhk
wDe57azfE9yPWXephM8XMqTUhkX9qFnJQkK3e+InBAGUT5oOQvYo4rO5Gd86HJrrX6x3ze/mKMys
AFiZ+HkUC28uQuT14xm1PGNq4REjgLeW3B6MaOXHhJC4sUxDOOjBBh59bgTTpX9Ezy6346L2MDIa
oFEnUUlw0lKrj1ZFwgJI/pY+pNtugwO4h0vqnPY5TT4Vl9+so/HatcM35dUcdMN7T5ultzgj5UDb
2CQS+LMQcZDgHHAymMXfc4DuPowZXDqYZnR6ZRluhkeFGWRu8qrQUwsgcpoFtZJdbOsbO32ebfip
Bo6cVqM5Ga95kWFudx05wqq6kicw7hdtA0UqMhpstZhG3r2KO9oaAohReo8t6VbT8+QJqH9chJ7l
hDF7RY2WeZgWufq41Jx2QYQKQK/ZxcuyI2Wr6QP84jS1PBBGof7xDe1RtrKxIuuTn82mRBFnzMcQ
6dbTLkC9+q0FXUZKy/7SyyEDISNI+0ELNwT2O0Kolk8vYd+LVnH3QyPItv8vrcFQvau+WuhODNHO
ABQ2jT/5Kp6i5cNRjosmk3OUl+5/PmrookXmoEy2peAjVJEaKGeTCTWkE9H11twA4h9ODMIHOoJg
VQxrbYlTwSKHaNpLsnaraeTn0jomxuElpnigb7Dyiu/qeSBv/OWa/LxQrG0DDq67MJZlEHKKzGrc
asUGPgK97r2HghcDeuMJvv9dym6b0WhftxizfsHpWL/b8v7REihx6nikk+mvw1LSnpfl/K6XxO89
1+OJtGmZf2kY4Hx7AKwpNNtOW3TTLU2O1LSLMfINjW0FXnQ6uydWMJjDgc5l28VTLBdt1dEoyjOT
pPtebbt0c4XBpM57YNRyL4mHe+NzZaoRbM3vjjQsl4f/5GUGGQgJC4qjPqVT7gr71P6ZyA3tvtka
YyPsS5L//ThDvv0kciMxkHqj+pMpWbH7Boc0vk/TmsN3MV7urbsQoS5UWrAMdv2EWak6xARqFSUv
1VU5sR0Kpsv+sxjHL+HdD6YpNK6a3DBDYBfVx0+Da4097bPCGvmL1r60K63jm5IjyLorRDLLjjFn
eJBv96LCpgaQbeylnNXEoGi46EbG/8bauy4t2QE30QValNF8n9Hu32lOvPhMVZB/wnLXfAI/5Uwm
SWAFI0rnLifFq1jh8As04pojUQii3a78TFc4XnpkXUcPCgVo9fVXVmtbiUe5Em/cgrwvOai7Ie/s
GLeDWcsJjSF6gj5+HPxtot8BhqohvYVutjs=
`protect end_protected
