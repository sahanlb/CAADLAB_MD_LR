-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vaZ/hArZGX0RtQ37Lm03Wx3HAR0QNJL6NqACHVZmfYjAK6m+yH4krhsKs1+QGE0i
5s1WsQq7geLjRdVkGsjMGhbyA4SRU4Ls3S594IuZwcl0XExPgOU20GH2Oa6LyNX7
gYUZ6Wq8zyFdpP8Th1dpdOM6i/VL5gcQueFTj2h8bHQXCTAg0sne0g==
--pragma protect end_key_block
--pragma protect digest_block
SUQtIAVJHC9uxHgPKRlbWW9QXZw=
--pragma protect end_digest_block
--pragma protect data_block
mtAl5gLGjVA4t91wJyY/Md7ll082IN066xf9PudKL/9ySPZ6HlIFMEqyCkdWu94Q
hvLG/vuUv4YdaDui9ndq1Lb2Aja7wJiQpDv6F+o0sWVPEVFbHyizdTpTVGA0vt0y
l6sxnTdNAyIaHHpKJhVroZruVi2SEinNDX2lXxFVVhZk9rQMPZQbRGXkACiysHEA
Elme9S91FcfL5C/Qh6ggl02cOOsYO7J2+6g57r9KayY6aWtdIbsgQQapJwl1fv//
uPiIkB7wfZyj9SSMhYHO4m4TzO5cfoYrafOi9kmdTJtMJrW68y5eLXqvSWRR9505
5pK2dQZPWcm+6jcEFRMGz9XPTbNJ0N/jPnnkvzoHEWDZHTPgCvPUglcusuLGNDdn
hGdVbIChpnQJy5MtpM2JkopCSsp6bX/WGEdRIDv6qWxDz/j3KkTTugUjolTNK1rV
eExksF3PwLJAM1YwAfmK6j8NwMeHImMKT7br+Q9OSMY3atn0dMa2bR+KG6L2bSaL
bgQo6htxgptRL7+/fjWfzXnY2RSWAIt9pp5sxvcDKcXpraDZKs6Lmg/yTd2b+E3n
+onOk4ueNkcEpde1rurku1Cv6AAk5+9i5GVP4qEbLTO6oHXQSoNueviYBKBYlgLA
Y/vACztLoBT9GOBjI4q5Rz1e1nINbdVevOVAUJNFMTYRKD90x4gZgpM4SkldDBoI
sjLna1My9+qRLDCFIxBuqgEJP4J7Ox992ebOgfoIfkAjA6mG+86KnmeQUPRTgUVb
EMVXT6+JDKfGkyKKkev8ES5KIOi+pQCzQSkVPYWzB9Pv4x6epMUQcarxgsBv9toS
fPmEbmRE/W6apdG4S6QVpHni39DbOU1Fnj17z5cC0UCflujFZRbHIWAsnW1mVxpl
z3uCFKY7YOpT6p7F4T9350OL3FOzstMNII7VSqbCyj49//IPJdCZoHDaosf8BpG6
1+1Hq7Ya8br/J0v7RF/6O6c4iEf1liAnvtb9o4EGNgHSCvNqe5NNkvmlyQc81RLL
WINhbyDPexieZyhduLGvlu3yBBQOVfm9VIFArgCsCXci7ycmVssprO/4wTD1GZSn
e+EToRJYELzZwZmc+VAuLmqVJyuiwcTztvhTvdNKfR4X2+RZEw7rm1ezU4K8ysY3
LQD+AdUfQIXec414X1ip8xenSXPjHxnZZJ43ndneWYlcoK0kWfD8cTi6Vp6cvtn3
eI1ufSlaY1xrxzcSTEX9w9jYS97LnhOBLYtw+2T/QZsYjOItOd57vb0+UPeU0fAG
JxP4IKrC3MJQAGd/6216ariPKplkThvUrdEJZzcVo/Agia0Y+OMrpclaYwXPjELn
Zs9RchrD8BqOhjqWJcFJMXsEvMCS3WEnDE+YMK5Z+jgh+Kl8F+WluyMOaeHdMYLW
7yf0z/INIVIX091Jlvi9PBprC8gnbQ+KbTfvR2k344TaVxI7N205w/HQGYyX2RKq
NVtSRR2Bxrg8hckSoWsMZGuUHYIy4owAHJxRm2DpU4QVxnznzvdCkrRygkDuEpoK
u0L53Jux4Cc4hHk4y3ke7uz8g2Qh3OnRTzgVf1BMDSSuEQ3i+f/smF16QzzHFbk6
tKYJmCXFQ+bnktA8LPK52U4KD95U3CUyagoRufI6LfRYWDiP3dyW4V55q548X6n0
KtlJjCqEXC1+LSrZP4sfF9kQ2+CA4ooRCJ7PR3L2tTTmsz6RoMmeMBoWinVAng6r
t+H4atCv69RByCstYLVPQuI8dCt3OYoyrJI1ferwXzIoJbhb8sPDM8gVBE2iwrco
jAlp1/jfJ+E/+SpCzlAFzJ7hpj0afaoXjrCy/cCddkYvHOLWa0n1NiMDW1N9yI3o
uR38jZUkD5kvQtqJ4Wp0vuhiZ4hA4wKeMCOH+uceashpM6pz0shO0Pp2UscLnsK/
vkx9Qcy401IgVOKtBkl6jcyoR/fGj0eIWdUJnwlMr2NpqUdVE9fMDSKpQXlGhFgC
MRLXVtEix2HYHaLWHwmKkmPWDLqF6mkmTgDjo1JFo56bhVY1NIWTUZqkmMSeg4XP
2RBvHQH+V4CfhTJCDAZRs8J015m84nHWqbljUHmlX2Bpr0en5+BSaA6uq3eJi5xl
44tSMBLiQPI4kEHIa6gpmdkTxE3e4wZrHO29+QdPOwLtlH60+L5Rjy7ojGfato6Y
Jlxw1d/OzBss7oRq0PkUqPRuI4nCmSvNkox4ov1hFRMSF+4hl4fAne60R4gcqUJe
kIDYDeEXqiNW+JidIEamN6+0tXU9bczUOt3Atjff8WrIVMN7o6wFrMIdUCslJp/e
nr94lxJ03V5mXbMYjjD79GvhCJtNswXLCwsbG3iAT04+T4+G5GqM5xVpZu/epspA
xWYSwyLavOcXpLGKEWKH7oPTyy8rCePGcZLDIp7na+3LRMXQNp+iFQQyYKv2U0LF
H5rdNzbGnsnyW2tx5SH5CgswELbLZOPCGZCsQZG444QbtIWGTzs8TYReQBLIJMEH
gjSzwiINxCDDFTQ1kVZi8BDMDvh6i2arvhKf83F0lhGchzVMdjscpNFiniv8uyRu
Sd2faxUSyJkMJrMReG3fUMNZxHEMzbspPWEFBRsyp2WNZVXO8ISZohZ+H3rto8f0
/jIhAGMBC4K8bSKiwNbEOti+Xy22EVxhe2FE7Pxmm4e8GUwZGZRiZ4Dj7voMRvE5
2mbdqHjUaA/N6SCsCnm5NceMpKZYfOI/Lo4CaymWUH1SYbQUhrFA1S0oPCL55GK/
JaxBSspnMq1+VdOAm/VSV+/zwT9dhWLvZKzdDSYiBuniQ6CguYSKk4eim5vAwCdY
TSpTQyA4cOwJvdcbhK8j5mojGyUt7EA0Wu+VlPtAxJZ2YlYMhqiBRfMvQbVlFPHa
oxFzcRG/5i+9z3IkG20pQLgDKTKaJH5HC5e85TkI4kxRAgho8Y2HPgDzhMyF1l7I
T18mNwiRXM3gg0MqnNzoSGLAMfMKPjUm8c8/+2AkOA+K/SKimoM1o/pS89UL1O+l
Xui2zlrWiWYaK0rhZ4vnoYbTB96tzVHSazI0jOsRkdQs6wBnyVJQidSbQM63SP1B
fDRkwPPp5wi2cpIu8yZojml/3YEgaCevlXp0plpFjGt2NOKDn6Z6t8qD4B4sg7h5
5H8FrPpkjAilurKEBxkP0Z1joT5Goh+wz5VhyKyK5EFWHtJIH9KOEXJTUN3ubT28
DP36M6xlIMAWBG8xobVzvFgfaCbWsLMGSIAc+tRotIGYgE/nEXygKnGU+vb1uqyy
oPd43G3U08SwMUHnQamcZuMifGwWj+nIlbdR63i4u/JBgM30xPLMOZi+NgGjnGJc
qGPWPsL5z8m/p55oRRUks+tPoZTyOqK20jipTa6vZEjj1JDI8CWw50dHY0796qVv
eU8rUhsVBuOmCf96ZtBywFx2KS3auP1Hivz/pbPfcsLuVnNC5gIoTqDNjD2V+sOT
AVEnA9Gc7WlapKr3NjpY6RbL0aQh9d8LmpOGP5q5vyTGZaM2rPk62jvQmh7HAOAF
j02QbtchO6uJFIzRrvFLwqV6X7+bIgCwwe4DTN5BQY2Owt7jtFpiWI4ZE2/dhIg9
9YT/8ExEr0y0gvqc7sgZ4Cccd72jz277SoICiLQ7s/4AM5pqayhj118c5Kbip/50
BVHWaEXv/3HR7pvP6dYbiI/7KEWTOBc2q7Csh3tMC9HgV+b55KuyuyhBPwEQTN76
slCQV0DtV2ftE37jMJS/WS4tMmXx3NJs66q92xDCZvL4SQRTcpsV1H0z0tZL+/nc
nyE4ePaE0XEDTrVWiBxVmeqfkwnOXTImXxztVz+HrNpH/QQ3DB3Eh0mevPEH7ulB
nntjglefy+ZYnW8038ghLdzkGIDcOTmqbroYHwlJnP0dqxrhUXPeRn64VrlWItTV
18OOwfBBERj9oDMy3f0l3dwjzgS3DnWllpNLBANflG/rHQdGCgnL/wsdywdrc/jL
MbAxdPWjINvYkKC6KWY9Wligmlc4GvZbpX5bdHrVDGIWly4yHAqP8vMEN95QGqRu
wVYeEumIcI4brjP2or/QbBV63KeGYSKIr/HIVSas+UOQ90/x8kuI9sbYhnc55+lS
g1CgpI9zwCH/a3ELznqme7LGDVav4M/UhDClnw/We72+tQLkIwTSEEGLs9+vXfxN
NDfGohg9vTynD1lmt+7HcFKf16SNzGPT806Sknlgk3UTW0QW8WgXiuMdGaWLNQ5B
JHgJZ83IYEbof/XoHBbUKdUSF1BgBE3wMjKYC/GU1bqkO+baZhxxlVolONjthoqG
p5ECsrb22f+9LyeHcONsr/G/xGYxuc87F/CRwIxsmNmBij78rnQ1O6R1b/1GhD5s
6ZgaYkseEv/nhtDAsiNIKrjggHsnbeADAJjKIXli2wu+4AL8YJcraFdiCKqGybJG
56rkKUS59e5SxxUYpXPRTHDu21ESv7kodVmpHufEvPE4WTDrZ5LdtGlAsisdwBEu
WN2eeAkXqr4NTRcWHpQwim131g8LiGIQQO9wwZnciP9MFv3v+AKf4nJ/xkVr3Bt7
aHSZR16Ny2uqE2j5G9/T9MuyzDGKM3DfYjV/V449DNI6aZ4T64kFl73edOKMzDAY
X5HaTcA726E26pYT/PisbpkxCvK2UWcQkUtV/o0wDKNogH52wgxCC7zwXjgHiPUp
gFBT3VbX23MwZJ0iPzGTfaay5pcSS2Sn40CDS/fPRetmnpObFtwXCWPN8uCBdSnw
3yMXruvIzaZ4+PeO4+hUE6pqTh8W0zg0Oifb8xj0bfYBvlQPPxWp+gPuXShnGJMk
No0ApHWtKAOzlzhTOGDcLw8yjI86Z/JphqUZZOiefgowh2wKQ95e6I3Vk5c//KKf
VAZIkUPyV0qU+obKwlg3Td6+8FsIalbf0ypLyjYKSeNFBlwcKD6qtmm57cMfII7T
H85v9ssCBpHJJpWV8U41HVw32XGUmnB155R4QuAO/0pR9OoKVpPa3LpwlXlaRREN
l2cOSURnySYh0q17Qn8A+iIEfu0XKJdUtTN22SD0e/+n+oeiZdSz5N7sY+uifces
6gpZ4HtizVyribjXflMjxW0sUhNP+G6Aq9Y7SiWWnxOWU/35SWzx5GxgZ7I8JdN+
6DQS7uWPWSYApz2P4YjuuClrpqMDjEWQs9g6smO2OFDobqRofzApWy0hE5KK2hqP
rG6zh78pY/LBNX9eiFvHpT3KROPkV+Lvv0nntdw8iKDv9CfWFJbIgEZLbvOZMCdq
DDVk2dZX3Wzr50pVePyai6bOZWAPCP5G4qCrdTJzXdxjUF0N2lz5hCiDps68uOa1
N16bM11a7j+EFSWO32ardQ0SpFtNuC9+fKU/L5ei9mjJvQUCDPVAfFTPTV29YXk+
NUXUbI3rluJ9Qj5OUVwSqw07usnQXwXnnZbrIFO2rwrMaDs7GYIA/7gt4md4wpY9
CAxG9GpmyjZwIH/qQwBXxftqvV8xvkx6zuMsr7yjxJ6CCAHyQPRq+zf77l8gHRqu
MVoqB8ox+90fJivLHEqGe1sSFbp1PmsYf/KXrrIRsImSpKP8AutNE7ejk7B3TEOd
HbWDvnjBDU0n2KZqm2Tf97YATqIWyjwWdwDHQjYS1PWxG+dBp/qigM5N/DUas7Hm
z/wYZ8lKO8KhXL3WTn5H7Y/Ggu5VMdmPHHYnjSdr12XYVLw1d2YnTYzjM+XW8P2O
kqs/lyJJ4d1b+V7+qFP4N2tcRO50718qNVpzh9cY5A1ndK9mmKvll/5IY/HUEoA2
bqqtlPkiER9hkbI3Ir2GRME4BYNTg3RQMo4o3M5kz2NjHOAQ2+4LRD8//Rjsp+sp
hFZucF+UEheLYEkwPdTOsS17xxmO7EUOtI/SmEsogPZ4vF59u6Y+siVcI6+zKimV
AxOBEhHpemuhu7T3wlHXGeRBRXtjkJM96ENFrxHzs8WN16mM8nwr0EdjqIQGYiM6
7PZJjVT944qOXisnadkF7jBluyvNtFQ60J5p/IIlaFWi3ZVlZ7c/IQCO8n+bi1Bu
ZxAX1SPrTGN58eZS7hvqP+ZMhcdfLKZqE3VgMTMTbQ1xU7rc7X6Z74I7pPS9k3dY
e82VRFCX3truLFcJBjhakeMduQXLEcvkkG4Moid9ogCnJxE6PG/bc6mRx8qS90e0
UFGHMp37wyqbo5byVmtzZt6Plfeqx6v3alm+K9WMEoNzrIO6ElxBlUO2zFwkOVA+
4XYacX+TnMg4IwqZbqlWJGVmqZIxPfwutZlv8DtNUBD5BM7txoNV4T7kqxa+lQHz
koKkA+ms9GtWJnMdi9lXgip7w59d6iWwLDdAHsvKSfqNgFDiuffaOShXSGg9dv8j
XZCShj7VgcinwW/WFDeRqmwW4Y8xfS+TjMuQW4U/QnO+HSF9WDnlX3fvT1TBbqmv
EFzrl22js3Rkt1XWJ7ysgPnZdXK9kJqIJfx5YH7Pz78eMtOb3mmGID0eQ+T833AS
xJdFdOSYXwj6dRbfwAas7SWUgURAtTOvbtZzmGnRYhSrqffrel3NFVNLU3hHX6zQ
jF8UJFaz3tOUJ0x5hWtHoljP+Pbr+zN54ghBdKEdH1ZO6smI+sxAaOY3P/8cAdMF
u6A2k7kPmhLfgql6a+IuOUbSUhLmA+uT3Yu9T1rBUh9zxuDKlV+KJL3zegRWMvNq
ivPU7Ws8NNenhD6njoxJnSxEqK24izVYVC8zCG8IKQV31jQP746uyOXsIx3E0EkK
XFMPWFIeeBI/VC8u+oHi54/wRRI2Osa0ifU3kZnUd6AiTo12pTGyjbOxse7w7qVX
vQLxH/74HcG4FKIO/s4A/OYiDwH1ynsjUSph6BPqC3Lp7MhgvYk4uIUOy5K0GYB2
SSKf2IOIv83B/8c3hQXX9v6YkRMARuInrt2CuZDeXc0uvdbQEn/hzxf5yvgaW+Dt
8lu0NdDVQDpmq0YwnlnnT7graPwhAApqyshJx++w+WulDfO3zXkEOow9u68ThSIc
njbPbvZYdXR10segEAX0qQ6sibS4Zwh2vaP/xcwn8uS6qhP/z4Fek2gQpqtx3CJ3
HuR2sTpQ40vz0En/ZqT0ArtO7w5PVD27CCjLmAB2mg+r/pZrOY3PsbZMfdasEqmO
wm6IfBwHCkutPmCb0o6n6J3pcG02tjMgyzUarjWM4vJiEwN/pJY5r5VHvH6XaftE
ENsNJ+Bb3glaFDOF6ib1EOjdDfVcDVeIwMzqe61UjviJzo5pOTrSCOscNv5yOUzB

--pragma protect end_data_block
--pragma protect digest_block
wJ/+0CwKM8gHXXM5LTbD/ogN6Vs=
--pragma protect end_digest_block
--pragma protect end_protected
