-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WzUD8vDRo94YqdCe/tVzS/cSVQppAU5mLx6NhNdOU8ywQ/VN/Gp14NqUWowQjqGglOMwfhWWoRCP
PrDcMDaWYLFpzkStiUs8bagb5VQ6OG8BwjE4Lc3fzqPCNGtHy0rmFHzgsuaIB392It7NTPx0zRwx
iCzztJgF/PG2qvgXt74cewywhqCwcvk8s3TrgpT7cNXFQNaAw6rjS05UX9s8ZTqLR5DSyhoz6ck8
NOgvXH9oX/hPWin0eSXGJzExnzvmiFW4BHK+eeAda9Tnx4Gi5IXsBqSoVucvp+LCs07cJPTTQQBv
5XFWW8Mavp4+pkFyiVpWz/px9l/MTmHltvtufA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6832)
`protect data_block
OHdTchCsmnli33SzkdE10JLal0DwBAh1GJIW1AYnuA27FZitdy5xhhv/XFqTCqtHm+Bu9374v//U
BypPT+gV8bvtD88yb67MXB6mimGcE3FnugiD0Qjdtr/bjnt7u0K2z3ga63HIZOI53Lpx1Zx7PFMZ
P8dAMfG/ACkGM8Uatzi2HyLwet4UdMO8GbFYXOMVqkJ8udWw/uaMn8Sc0ktWPTR3x/r4MqJNrIw3
y2Me4hCl93TmUG+1YTNvxfnbQU/UTUh9m/m+RYvDMi4FGyhl0L0Afxp0ZYGnz47I4suq1LEXkFAy
HPuoPl8C9+NgKk9Lx2EXqhMF2Y+9xEHZIVkIjalBIfBv2m7L9Sy6bFnePyW8LVJ7Sc9VHmuKCza5
xua31pI9C3pxqgvP2uwSIQ7Yc2x7MJIPFW3cqtQTwXV6ACADx81FpXT3Wroig/1NDdWSPs5EsBLX
yU9/jbsv8aX84MEOMSBpznqLqqiLiLqfgFHU2lgkB7B60ahqOtIvYhXUHHEL+KhMataCtTpgTCkJ
i8W2uqM57bfHCrLpA866TMoZO40w3+ql6DCQUe1WXt00tx3qTX18ZjMHdFAmnhPwFuPHxZ/rn7C2
kUjqecaCUB4BGPtP31qTue+KdpMbA+4GMxV8K/rlzhnS240+lNhjb8bYUWTxgALEQxlBL75jKztj
w1lQxxp1FaRoz1SMZGFfT8OB/cnsl7iz+P42KDJKvT7fNHPRJ0VUuowRu73Rad2Cw2omo8+C98fw
f4dKSL/1+cQ8ONOO9VSgPbMU6bzjTMp18zN/PKANpMKsKVZy957/9WD1tZprWZSOucHn1+suZgxH
95Y3Veh1E03PkG534aq9w+RyBqlUKfUC6onKHx1pJ9Xr2gskC+aS4agdgv5oJzSgfOgTZ2d7o6as
Qpa28j2olwcsT2YBodkvYIQw9t0rJ32+EXUVZrrBERsOrLp0Ng3p3PFJ7+IpmzqLnT2jOnlcCpCL
nvb1kPneHfK/XcaUTPNvgFm7c/v8hlX8Mm8fXvsERVLZHwbS8EEDeJbzPHIANUT4dRi9/4hX1kIj
uTf1j3CWA2tPKFXLEISzeGPZZGdshuZ6cNAPKrn19HOhUOp30mALz20NKz9E+u3fnDPDPE7pje/d
i7TUgGwgUOW0SupojxyKZ7QNeo9+shZsBipj4WekMvz/PJ3BubzGdK0WEKGlQbcG6XXi5Nn2oMRv
y5avSZnwnobuiaWrrE4WYDAGvu5CYgj6eOnqWFkGCywAN5UdIiuviMwjA32odhXqY62KhAijoagr
yQ6lRd6itW/j7l0GDy6Uv7L89Xr9On3+PaSFFXjCNGiBzO29FEOpsnH/DzMqdAhdMlA3/rTM6RLM
5sgvKnCDiNYqdHlIoPAP3d3xaBq60yuT2uifWJYm+Cs3ji4A+xw4W2K9U+nHXFG6I8S1gl1+3upy
zQcGgZrKCE/d0kX/Hks3jhbAre0T5ybtYAl96mM9AO6G03ZKRyOb8jgcTBl4QPJC4XEWF1+Es9Z9
gVTj2VpXp5ZuhIA676cX9M5PwkSzXfrsQJi3O5DKJBXjEO8Uho3lZDqzas4+myFA+/46tTSKdsCL
EWFYI+tzeMMWpaI80Vxb2/EvUcxskppuIAmo+sn4rTZA1sxbdGJsm/UqDY0O3ciMLSFtWTJ+rDJs
l0hRSEButQG0bjlgHINsbR9UE7EZsdkPbzAB+ThCYeDeVTTy/dJjjFgK2mvJtJlcWH9U/ZXGHHQV
jn8mL9Q8yC5ODdd/mvuzTIr2/NG4zC76Xr+GtJJg8zVznjZfXDOuAcK4npK5P2b90T/1oPcLOsDI
VYml1mRBij2BkF+o7lAFsvw3G5g/EbNJyZy7kjcs/g2WWQ2+P83jRTQiAdCjw59a558LEqISRCCw
OhBf0Mqyx9YA9r3oAqdU5JAvDOZJ8HSG1RUA0R7wPBdSugKqrr6B5eTkC9ShdCyvN3RUZV+KfVPV
uSMeUFMGQmTFgRboesb0CqD4clpu4DrP1flMuH6C1y+3Da0LqYXfx9+Ue2+avkGTmBALR/yxITkt
jFIJQkbZytHsse9W9lgggjukzLGun8GbN5AHugFCtph9ilPgr8SS1CAlvwtB9DOLd0MQB4Xbgbsd
yk6hEc1J9et3E0mC0hW79/xb2EqgbV+6Piof3WCx7Y9B/pE65KDunmZKzcL39gy3eUPcdtkCzIUk
pSW/5p23n6x7S9/kBwNdHCeWdDqyVV+5gzDyejLMHc60Ap2u/UWgQ8rdJBCshVX3Y89YrQqcYODu
draNG5wCki++bNPy2lcwNy5hUTKBia2FE9Ij/0BLXtiC87/xyGgYR1GghggE7wUGN+wPHSVg/D8t
0OvcUCTzcFWd1RArZKuwPjtUF5asoov5xBXW+iPl4PtdoPcP10kBYzgancMr4PQo6eqD/JKbf1+X
wWsQJ9PQ/B43F6hpB+39A/QAl6WPyc6VZztSWLItlj6+CaKpzUrrMelr1XZLa9neq1ItHKOtV2yN
LiBMH/2OR2SKUNiUP4uVgUgUzyar0w2gFYQ+8oXHfFSaB0uDvi3qhA6VmbraHZwisPdet2XBsWFu
1OstAPQCDfip+OwF8heMQMAQyKy77gDbnnmr+Juk4PLeZyp5LRGNeYWXvZIYqVPLF961z0I2E3qM
v6DDG9J/jSuUPpWdzgACjRRcshIQv4qzkmzWdvG2PxOJCiv+m3ZeT++x/6E9Nd9LoAUwSu5F5SkX
LhuSfCUY+IlbeGpSd34BWyrp8UCH/e4lhSafRxY3b0CgSUBA7guB3ZAgINB7oWrRqIeayI2BN7H1
4jETdja1Gi05peTiZ0n3MAgdLlOxuEF/iih5W8M3+Cw6b6+DNEVGSJn0ZQWcftb3XytM6pe2Ch0V
/U4ktYoL9d3qHoCTvsv1czMSYIbHEVvfZkU2dTxlWqz9c6DA778mtKN1WIPBZUxgK47dKfQ7Urkq
RP5iq80h1x/3pHMk71Sd/80TcDrWZ1PF1I1DggJdqQjyaTDhyR3wIyDrDmTTOD5PWj4xLQRuFFSm
3h3nD5wpMqG8E74gFey1mcnr+z217S7wW7kXsj4cuklAFKD6L65PtJIYiv5TLyz9E/uV8xs9y10Y
B1i/Huf4Nd7j9zW3H+ui7UX3PqcIO9+MA+ghZp7twUsmTsEcoBX9aOTjKKobQaImBaVd9CIDpr5P
xyBMJf0kU1xaj/4VDxMshSQk7eCBJNwv3vIYbAYC4Srci1kD/w1BZLdt0x0IUwT9xzIDXssmO/RV
xemdYurUcPPugR+Ll+7UVSqd5ZE8cKkP1lMvBcOKaHkkdbwYw+Hf9CQ6snbSLUN/APvQK64CqCbw
PcFCAlkgungRK3gV0D42m5XajIx4KA8HxZ04hr4XflQdat7QzJu8AExjXUG4AybkP74BY7MFNSks
SPkuo6Ok+DRe4OcIfYOi1OTxMdLW2zNosu0EWXp98X58dKUJU0/rg4ItWVzKVzhfqNcgOk++jsQR
0eZyxd+fLK9is6OFs+PYc6xezOP9WKzRL+tRHYGHkYDsFPW4l7uK65KBCxxrHytboPos1e+e4RQa
y8yhQRRPTX/9aCqg8he89kjZBxlYUYNH/kDa0BedmnfKBxOrZs927k/oC+e30knh4A3mNt6R58iz
+iEOJiaB99CBPHtiYOo6kSpk642OzwBYPBNwcR2tt8CC6b/sXCEbd8hrYZNN1JIDOsjOQoHtbh0q
AP/OzLuPvPeZ2L6kq9j0TfuYW3pCrULLkwVNzbfIRrVdM2vLvK/LGRIuSqA6lPYZ5H0IyTZYj6dW
bQw0TyZqXsNI+bV76QqEjzZxpj8fYhobozQbqIMhAKPTtKLsTUf/O++aPpTXSsfKe1jaUTkwz2cu
Xl01zJAEzMQHapibocJviHtDVnyA+jGw4798AYFvjpfND0EXdK+r3wO7qkEUVtNuYcATp9cRItx7
hRvpaJrYISczcMzat2ZGuAFAElofIK/9M+XTHRToZZOsYe5sRn7F7AW0G8Fh1efDTnwL2QszZCC6
/rx3cTHQgkHUy42tjKvqk0zM/yjLE5IEDpsSz4xaS2BoIz7fTYyKIl+RkPBnyFi410pZ9AcItOSm
eP7mbLIYqUvNbso7LmGwG525sd3zaOgtlaf02gnxogdip76aEHhR3WnZH4r/lD3qeVK06Xa+XDpL
IJzwKxwujw0IkPPfvmNsXbI0bG0zghxpRme/TGRC9qFoIZ+2obKzToHjeXik3FM3zJvNiI0tyavo
aFDzz92YdRWen614EFwKauHaOp97BNNLnai506IpJ0E1oa7hpp3kEU7gNz0LrTTm5tZun7i/uTlA
+l+bPEAI7GX3/MVmi1Df9ihll3ZasfLXCcInfUKeWkiAggk0fMF8VbeJVgLqzP3TPnDs2yPV+DXp
9OnOKs+GNNKcnBUTDulbAuuNxjIRKsonK1YKhhRu26ccqDwM71xJEyaLfJfFoNRucCnwTMfLgT1B
altrBdn910VxpgJ7xyEm2Wi/cjBKFQtA+dW2Hk2MRRLL9pbn4vhB2FrrZ6MOYfOato8kCyDBlU9Y
S8hLmszwvP4BxEEdqWwG/4xwZE6hhjSFRYWoLFHW/UvNDx5C6P552WWGMBdpPiYU1pzBzTqlaseu
gEWO68S36w2axl+9nlm9cxB1QFqtDVCl4cycQy0HfgcHHku7XRRniVrnIHxtzsSjKRhEAKIlNMDS
HOwXXbzZ2sSQaFTkcTIi2bW3fVqWhzx23rZ8H/lOzUI38JHQjEeaEnkbvFDe/4lEyY2Ut2bOifuP
fQY01WeF8mFxnPHeaMDwJfejxAkLoPwFdJ9zod8+NRcY+AumWxm6kW0NYtFlABdHtjbtu4hdGvYj
CWHRQUXcYJQGit9NlFuyJG094e1H5t3tZPyxkjyuUZ0Tgp+h1kKc322L4x4hL4foksna84GbA3cZ
ecporyZzwpFlWW7DH9lJgKBc+jfIhfmP1Q0/w2M9ATO+JW45sB+PaAVFE5UxHPRYJRBoRt+HYreg
i1r/nxxerjcqOS2ptq1y6Tq+Qe64DKQJ5dKYN7Cg1x9CY3aVOO3kvILYfDOozWNJKXdq976g5Ajy
S2uhoDJQWFrCFMURGWnPQVe9/AqBi9z929C8vuZlZidsEYcwTdeIJss3f9GDa8zgBZELaN8kmgPt
5HMwvv+/WsyQjqZT0G6khMOUNx+oLD/hILVtnyO3KKXGThfIwILHt/nAoSVuXUwY5UnE2/UrUWwy
1nDXoW1E3FZIILEy9LumcW342sid3shiXe2BCiaZCdoK5KtpvwuBVyHEl3k5YsdAhpuGiAvd/zKx
9yWqT51xU/yMJPWDRSFsF+V2j39rW8nj93B0SkBoPl6OJNPi1LO/1+hVWRJJ7xhQjQZ+UOa2Id8A
08anh4S6tKF4Krw506U20hMx7L6Cohp/vlRqRhe0N+L+lP1BmF6jEikrPU3prXhFZVs/HlAA3Vnd
fujkuzTldbNQWMTP19zqGAh9Nz/XG7902aMQvn5OiAhG3Ixg4zAxThefJQxdZoIDguB9fJYaVMMj
y/6cs0FyC40TDsznO96TYxEfI4i+oT5E8gQp+BzPEz+KP3AQdwcNhKEsmrfSapR4dw4MjZ+4ivWv
QhBBIJEUZ7QXwnOc4yZCBYxux2rNbqyu/uPFRsP4LBe+ekVi8s1V2dLczL50e69oBIGefNrRPBI9
2Pb9bQ1kGzTiKzdtx3X4ejGrt6uF5GLYziHT08gyqxrLX1cvVBtEsOVp6FEs0VZwQUR+mtoEwSAR
ig+iwIfzGZZ0jtxYOqY3rZfU5AFs1hmz7TUu1YZCIdBrhcfa0KziYYbaRK1GGlNzSq9IMQrQIduk
hlqlkcKhegpbBvE6zHUYxXsRP7+5Bm1ltRpV2fR5KO5agUjyVhkPhi5W647cexV7hJXbGd/KTxoZ
8PO78I/U4ZL17qWqb/S54NQc36QT9gy9vN1Lkd0t3oz69YvX34c9L2m79T1CRnFn9JdQ8CNvL5kt
OamoP25kU/yfgl1I9P6Kf2CU0yxsfONy8GWaru80q1TroTa3Ey1dRzDvtzYTnPPA5N2vvApdFlO1
kA1nA/LZKQVad0nW5pH2HqetPHqFe9ub5Udl9PTMtei5UKat4Y4/4xGNlQ71AVx11BXhtJlOaJq9
vH31raKNpJVAkmBHAONBh5w7IcgIytolkxmd8FVtYndti7Yf+ez+1GWjGAdE/G26885DLGwuMQUB
ZSXOdtvli2tlz3X93dLQyIgogujILrbTrp6Q2+7YsSZvOxbItyuz9mBTnJT3otOClCH5B4HqzRRm
EC9oinr8EzuiuxffddrPeYLaYb1h8Jd6Hvt32Lf11duu3ksrAjpgYZTU7kuEv9MHwpnS2Ix08sLr
xqS4cPpLWHk61Pt3QddBZewAkdEPSUrmPW6DRIcx918jJSZvpcadAiiKO4uyUPxbFjHr9Ozt8DR/
1Ago3cuP2pacm+WjzdEP7AIVKzsK1RKzm76wig+UClIfEfGOJwecFM5nnxOQFdVFq+SOBOXzH2Vp
oea5DYNxIAbnO0ocUcUm8NP1dTG6Ase7iK7xZfB1eIVE1mI8wtlTPEAV+fDSeLBROFPiJr1eqJ2a
hSUy5a3CuhD2t0ooMxJpb/6Ux5M1oNImnWBaE1gw/LexwkziTnVI26LWprhYcmuuOZ/2OQ2HVSgi
lQyW/kS+2naT1p+gFmUszks0QrwyM7OFH0IxW3THGmAHiB/obN9s92mwEbsn1B1n2vCKeevlvROs
WfVl8ZCeosVh0aZiX6fs+yjIVVRsNV4HlYkxbk/WAOtwr/s18Ju1WQrY2sA+upFByWts5Ms0sfXj
AyhCon6Mxpa/aDLCkuQE4F7KKKNrXfUXhBIiA+0WOl44Z03wXvziJhD5NXimQTPCSGdCVNyZ+GVk
TvxgP75PpdiElk1b3EJMaNPBMP2xZ+aBWPkUdLSxDvNCmHa9JOsl2Rp4CWJcjy6T18J7Y5KLXW2X
2p2dg4EjrCFcQ3h6H5L693nNZZz+O5btoW4U76YtyLVGOTU/b6Mwdt0oNwoZwb0ZqjiJXjKn+Zir
IXwYXkoyG1bE9HqbdzE9vMbCALdtik6EsetLbQG1K1TPcZg1agdz2fFF6+AQqWV0y7AH+l8+ua58
OkbGkhRNhdrZk6ak9IjpiChPB0YM+v5M4JTojt9BDgro9VJprXkK1RtDvKi5jvUgiktRmHZsRCxy
P0FDkVQr/zy0VjMIIMp9EHST3S7dZ3E/GoFnotWwUHuL1le5c34OfDaqNuXHxFrofIbO423xACec
s8bxXD/VGPc5mLCSNTB9quIbqDaFvDCkuZXfcOGJxblJYW0HlN9MAjk9WzPZ5IsbdeoMeyrmxIH8
DAflL1Kj5coBuFXLw2PVRbQXNpms0Tv18oy1epA0Cz5NJDNmNOlucLQTq3tf/HmT9b1LdO+ezKxG
RxwfUVMmdTuVAXS5XQlBL9QV+YSRQTwqOX+rKNzMoyaixSY1GbPcDl6MlPl0zKxsOoXXIWW9i9mY
nZfqg1X6qQ4+6JcQLJhDBFQ6pnqGA7Vv14sxXyyWhGxgz9BmbJC+FBZFc8pCO8yyPl98gh6bQS8t
JD13RIuzk/1033JTJzOZq9/9ks0QMR8iH32nkc+8nUC1dVjl76eIBCf8kBMgRS0/SreckJIablPG
0nel9Jlqn8d0ckA/t9d1esdilXdMmeqPxsQ4G0gXkGtZA5BovtvBRdSvifkPllhwll+sIzljN6I+
qFtmO3anorrvKOgQgD887M0zuDffmdelnySL6vAykODWywJCw1z1bXc1jBgYfnUYj9XE7TURNHlT
wRgrEQ26PzUezt5btyx5rBleLQU5VdGEgRsq7BRqGz+5+UX86T7ELAqXbeJvbbc9IPKJTsJahxMx
y0lBva+kmkawcwg/LWn0GGpddSwazGNjmAnzNAY7KO5I+kHjSXVxxqrt9aLpLeAnM4510Tvq6gIR
tb3g+aKxsD+JH5mDZBD8LgbUUwtaXSzWm6JHyYN4Vp50V0TAgc11hEZxxZcEQrj78uKzo2TY13D9
jR9VV1Y631Ttw4W/oANM3GTeN/w3QYwELK1FeowWQ4PrbPa9oTOV1lIQZorDm/R5RHbRLeAOm77L
MnVOWf35sg5BzRLZLNWyi/m5hLnSq8mDzmtRt1vClEVM0of7M2Nh0Xzrz3bgFavc6lzZy7molsbl
ZYpJ8k7K0r02Akis6ECepD8Bj/DzBTXANsT/tDijGiWjQLBYt8V95vpXDv7YPkCTEUhvIQ1FYPBx
/40Zh3+I4S67uPysYFx2tVVMwAJd6sGm0axtcJt74I3vI+ws2g+WGpZBmIfaR3mzamxm4G8S5yDe
vvM6o7BpNMpzLO+7NHAl/woz0XdcGJhWI2WYRuC2IFbHct98IRiWFHmpp/he6SDQrOWkZZlhKa6H
S+lywQ8DeO3fUcLTQ/DuGCzIGmHTrHCgnHJaHfF3UdZEfWasRX/en2U6qs4jNCUrQ4y5HLuXbxT5
GD9QW/TcUhUyYBnII8sFeGm5fH92rUh1Ta7NeHYlL0oFJ5sQfs98OEj3d9bdNbXwXueukjPK1qqT
Lakpg0w5SjAhVXZLm0a5hhu5DvGq0na8lF8CnL6NuW6JicS8UYRZlrY6AVKHkm9qmtBw1DOW8vUu
G07GWv21n5Omh4gnXTKelcYc4yViXMJkE/kgOX3weM0uRxWORipMqbfr7grz8dya30ceqJ6aoMPX
o9p5aEFbLXUiL4UDSwjIi6bujjDtD5kXKzB4ap1rBLV+0IcQyUiCiWa0wC4RFfdHPFFaV/3TPqOG
NxeEjL8YBAByVAA84azb7CgkdGReTpp5K1kPriPGaNgr+4GW+pqf3OX+gzWZJPAxiK2AWWj/LxNr
RhnxLYYMafiT5T5jUZHMjdWIzIy1rkOU5XCFj+iVvvU5XxgfFUHzhF00Sb6EBJxfTLjNuyE2jxe9
Fn12Qq3LMBbOJHMfdst/RjHoDgivplBnf3GY9hgF5f/khDqaIAx+Mfp/jr66YSyN2kOIbMZcibKr
rp3fCkkBBgWi6HCl9Wr002kkMY2J/kZ05u6rRNz0kk0ItQMTh7A61nVWE+nlK6U3Ug==
`protect end_protected
