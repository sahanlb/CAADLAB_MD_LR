-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
yfR/w0+nTWXfDwevDTWpqo2idiM6C7UxNFXc7C1+yZcgr43J6QQtSLmYBkgS9c+e
96qUjNiZCqAyqb586ezHdPk1nAC16dj7+C8YS28sz+oQanuiexSjLF4d4kLznDF+
hNyPgnJDypyfD2gf3bfbwisbC4T46gOsO3UjUf+E2EleSTluRHTI/A==
--pragma protect end_key_block
--pragma protect digest_block
6p9EnHns8P7mcqFM399+e89L+eY=
--pragma protect end_digest_block
--pragma protect data_block
fQCyoSp7RxEE5rBL4+zNkFfKgmJTZe79Omsc1hU/RKUlwEoEnxfPQagmF25EN5j/
TO29g6PuQ+wkvtiqU6NHN7WJ/bi4LLPl5/XPgFil1kBj2b+FPleBoK4YOTfnp/da
tTYtKJ4MkYSEMWkopq6GDoERNXOqaZCDpPx+TsCbfQtQDyiHOzYlBPcJxl9ZaohN
eGYDrWmtn5pFDqO7jwrkQaAWgMyRCdQH7ietr6P/g3zURiUQL2CgoykPbePem3SS
6YtYKChP7+GX0Pm3X1EY2rbYPWofhpGjiVkz2PqVt3e0+tK9V09+74nn70pbOoyi
hErD62cdYW3FfgmSzoz6FmZMFdqXp19E+/mU5pLvb2auPxJDjf9GEVDIxHNfjG8w
XILRfn1CB8usY/IzXU1C3GiBLPkmmc6/9ppDSPaQxpZMjHiG1wYhP8QAiNTghGOb
sEXJoXDP4KKTuQ4rpqIDMU0ALnvMuBv8Jx/eWk7mkk49fS64eFGRl+BlqTCwuXuX
SUu2XCoUk+vr4myPfTnwYwRN12x3I7HWkgArnEFC3av713D9Xiu39wakgJ9Xaybv
7B+rJzWe099MULZ9iMFvIKZtE5N0GhIXzHIny/ZwPDIjEPt1aPJrIXcZd+mrBJdg
Li6wTkFLtAZarsGZBW0uqlzAt0qpLhhnfz577gV4GsLHc+RUYeAl0/t2NIIqH8pQ
8uKgFpChdJYfK4KvVS06I0iR1mSLyNQZhCBmDwWUuXpqcpoRILMHL2DukLD1Kr8B
WaR+xB6mfNT723PTD0K94tTtctfnwJIdAQaMTOZFh5Wk9XhXfhq0v4oECzXdB44Q
qLzbK9ROey/VC0V3vurcR4BEqFxh+GNpk0q1IdgAqC0Jo2VGguosh+ioMmAYsTko
VBB/3cNRsEpbt5d7DeyWeOg0ysl/Bs/Ly3L8CVrf5VwC9y7/BCSRarf9Wo5RKelZ
iqRELCzvgwpiKzM7T6n4Odk/4k5euVejcjYJyInWL88mJ6IHRukBt3iDtJsZFZKX
w1CrRyZ+PBjtWfPxU7TJ5R3BMKNTlhn9PI8zm8pnXbKAHH+pWKqAiwJmE2LzWQkv
a62FfUkj+jGQKBMxJTZh7X0BC1f8p3r7xup2W2bw1BCPMSuVn552jtQ3A0ejopqD
woJ8VymtLADo8RSvy/Eu6qcZSqzfA3g/JvjzeltddC6PmErfV/lk8f1FJeb6rbjB
iRglHEOPU3GpIY0RlaZObnJxIjEBXoGp9rmQcAPuvgYfzGQRrquusTuRoFd0mqRu
Rw6TxBzQm03IIJDmmCx5COAi3oxn/lf2FkKvYxEXwrFCkkzs1kTp6E/2XXoSB7dV
veink9Wc51ZVzUZlPDXAbfSZRRVWLLjM1Xbzd9XzZFBI/X7xN5uvy2JP3/j2LEGC
S6+nY1gCrqaAgl8szbNfcpiDTDg9D5/fEwo1gDXOEdQrc3WZogf46v21XTzisoVK
JPucTnLqJTGqsEb0/TgQqaDWhEoLumZVfzqT9XI/FY6BvNO8YlPtybpxd3hDkhh+
7mJKVV6S/zqAnrcWGE3QV9Qtx/msWmgpsCMgxANde4P7zMRNnn33CTDNdMyLfHOF
TbcPFc2QyR6KU5eFKzPmyQ0tix8Kd7EJxLtX8R42J4X/cc+uv3toCU3NoWIm/MX1
7nr9XehaFWTZYEcZ2vs3BMkuJ9f0RqV42hSyiHB2Y/YnU+d3+MIY0DrtpoMRr0Ro
i8GqpZu6FJoP+D8cM18/iJYyf36bmych9lh4hQ3dM3kPMAZs6dQjFV30OyLPMzRF
Ksq3jtXK4/aQzWNsJXwQsy1bu8vGUxejVKR8VhFBD8VunKBuhkqv/TTDD5vY/11D
0vUPnh1K+Em9qJcPK21lXH66IMhX6GtlZ8EUz16RTEhJpS8EWYIAZ70EBrgaFipM
uMXaRXfxhS+E2jcFKCK5CXJYwe8IEi+R/GOv14P2Rt+2lDBUmWw7HmlVkXlO2JnP
8Hz2UaAHcE2+IpJlXLuN+q7NYrwo/XqRT0wPPT0hIj+RSHbgBB8oO9LYNYQySPmX
LICZ7CvDqTh7Fa0bB2VrRdZmM6PjL1piYhd7Gn83q7ERwJKqnwNrBrb8R2ASaYrj
SXjP0gqQUPuMAg1C4JaQ1bF5Glju31Hcx/8qXvUPP6MRF+KdadEuTxFJzUX8Te9p
BCJSOwCjGupvuH0sicavcpMkK6GpKZfKetoVQoHuN2/CwNvDC5paLP5ejpZ43c6o
N/5FlKwQepANImIpY6xOawZ7Ab7R7DZCiiy6O8HgjT2xNeNANU2kl3qdTmxhZ4r3
B3hzfnURgpI9xJKF/OcH3ZYD6hbhQsQYIVpI2vw2K1EXEjDK0jqjtwHVPe+519Rz
SUOqEbgpDCrDg68vE74gQeRlkERx6TjZlL56b6+geQkTjZOBqFYMoqKgs/MFWrUq
1joCfI6r6RRY7POXLxf42LOiHxBxx69Q+0Gw5QNipPkzkd78pkJ19e5xMqbG1Mz6
4W9ct30XmXpYmcJJL1q1mK62d/cenQ4M1S2nvZawzsEjCMNjmj4v1Ihhkc9eRKBc
V8lpOsNpmHVzjTk4E6cu9vxcFXakZt8Dkn58TS/RBY0CubMVP8hyTGMo/BI+kdNe
i+zNoCdhODfeINhAkXdTPDgk68twtbOfzNYD2Cp5ejP49mCF/XT4gzFwwQAzrUfv
O65urb+DWS299GYSdbvL4jrc2x0O4C57GPzZqY88i9Dt+YUhnr7yORe4T3a8gr3B
JfYsd57spHbPD8keJpnNKK8RnsWErzx61roZ+EJcGb7cEZ4smLfYKsjHVnbefASS
Q8mZRQzZPk2MmQWDPgsqrfaV9bA5M7JxYx6AkXAr/Bp/bZDSCgRlI+H7158reEHi
RoPqi/cuwUneF/E/1dQB5MzZMcMvZnf9IsS7r8Gr90ELYXXuUq5uHmB9atYV0fst
0sPOmixow8M4aIgqlxzdhVqVeR1W3GLqUDVwgXiqeAlJyZi88djuCo4wNBoCUKuY
bhsC69aRrcavFXqsDBksO67GN3w7Smd2QLMRa8cdIrFsUWtLjO1ib+I/ZLuJCAjP
AZAjRYFjcXdvV2FbxW7L2bRGu8pEjsUyh6dgC3aDnhiNachidY96iHAaD6PV9E0p
hd6yW58TTwxBVQMzqd/+vMbt+b1nuZQEEUbduoMB10kuGzCu/s8SQ3Pamleqdw2O
ItnXthOcyOE4EOtInD4I1jyzVa84iWTS7N0cM5PzLZ1TnLXmXOMxtT2NDuJdvoBk
njNh1umCTcpdSVGgVAmjY6DXp06L9dJkNNR0kRNVXRCUV/8bUoi+0PJLpNLpyvkc
oY/BNf8uP43UB1m4srvo31D7BBmb7PqtoF5Ru0uQ3EBTpPVAaOmSKUMzSpbpCaOw
g5P93xWKr8Ue2h+8UNkf4u9BatJoSQBzpEGBz+pGDmmwClxsbnJpfywFM3Hf5sJA
maj6NAFzf2hJDsrHQeAX1wYDeVP0x6sK94vDxXbsS7lxmdgjC+Hya9mn2n7o6yI+
u24YvyevQg9tI5Xe0Ae+RWaFQtFEB1usRtGJqYnW/sWlRX5vLOQip8ks58sS+ssp
WKUh/6r5dsmW+qIAKweL563jLiCm3OFPsWsk0/BXjS7zYsS7imXerTwDkI6rrJ5s
zwSyYdxpeMsmyNUlDrGzKS5FGgzO2CF294yRyFrPLr5lMxyfcJnP4DJ/pEaYMm81
aD8nSWrp2kbJsOLlXR+mNjJ/iaUBSLIlxAAYfETaYQN+UnsNaNRgPBf5x0ZBimDJ
J6uAE+5T3dZUXaCXU3UE+xpGaXLeWfPqSdeAWtkjPAYlGXiA4lZbZ+2mmD39yO/f
VQ0t4bjev53HKgo/j7DKKv1Kqap2seoNfEF0619So+3bsCoAA4fU/8Szkcypv8nt
jjE3IzTkalyDtBjCoVzdxmrwp//PDNrMKSQrKGdqJHjkePioVX2MMexUbv2kcgqK
ASg0IPQurWbjlvkRTLhMKyRTs5yS3c6LKM6RmPqjlIEXOlmiNq/US3ekXHewL8O/
Zi05adgAXglPDvxRc3Uttd6Aowapw9anQxcRzWnATw7ERtB2xjJuZPym1JiUptXp
aLyDvjzx2EI0sf93e33XZ2Z5lu5eYNPFec98gKP4H90P7JLcTuWLx+PTVsU2FgNk
zqP0ULErSNSbm+h3kqOnZjs3ogjSqBHIJ68e0CZTquUEgfJrcLMJQ39x6aRjIXu4
75ZYuEhB/y4Y6SbW2bSKkLecO4idDFqNNq8oihmw+WvTEj+x1mgJ2msc3RQb2+ib
U5sCWjbo+H1T9RKCTZw4PUe2FFOoxAac9IRJCOMhKIIB0IPlk1sZwlbe9R3XtrTa
9JSfslPwrmNXyY/qtp2owzjtydZNP0aYnXmbG42aAulABiZrqpYG4DqyaBiuc3V2
LUkPnhix0cVk5OoCb7zJjaIsY68rGfk0DgcMRqMf1lb1DOcTK0yCN8ZHxr3WmwUe
cSH8UTtBeCzh2LDGZkoEFte1tzbgWIia+QvXQUgPrKJs7eQNRxhWt+tUNj4+i9ET
1vstWN0wEJM/dfLMzthBXsubeidvZPDoH1jmyEtBc3uT0mDYVS+AydBJLbD9lAUc
+SOKmC9Qu7/gzvkkJ6+RbgyKj3GWmsTkO2Q9+l7UOJkFVTBOZa5uOtdSGDqiePJT
P5QMCePdScuIGSzWokIbmcX6tBPVJ8MRfqdZem1ACC/dy4FKpTSDOus2rbdSBNAM
thxGHKqGkJWM95+UZSJIbg==
--pragma protect end_data_block
--pragma protect digest_block
achpRy782i3oBOEHyA8f9TMejt0=
--pragma protect end_digest_block
--pragma protect end_protected
