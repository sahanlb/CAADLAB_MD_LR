-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
nxoQcQvwLvoFIwWXT6fKOhwesmoTfNTKK8SRlhRaQTrkHAPnF6GO8WGrzOw07oDQ
MvCbF0EtlmU0iO4HUkGiMua1aSYwVo21UokGbYLAueea8tU+uCFiFa7v1iCu4Sip
a9nuwent6aAW6qKeCvhyL4457ZdTGogj9TdpRJL3uSw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9856)
`protect data_block
ys7kXy2e0RtwFC5G4V0ovjXWl9MT9x3QGytXFeIYN4wDEADTeMeRHPio91KXuvFC
AIllZuv1RmVxTbA8xZPKHZE9eTolLtFsfReZ3yMOobhy6GIbaZmxAUylVQOjf0aS
6XlgPLWjwCweoVJGZGP6mwxRgyUYblu7tscNSXh5K5sDjjrWIUbgiF7Th4f0Z/Ln
W1PuMrtqy5JgEhiMhQDQdG8BmuoF10i9I7MiRJuPCFDLuzQ8zhHz3YxK5/ML0DNy
VDc8g6QlL6CL6EtIk5l0UMsjI971TtmwhU9x3LjeOsqEZWpMY0tH5qSu6zrMVRpe
4wPODIS85Hjy3snaramhsvU7sV8yz1otDOP73aox91buB6HF1sghWhCZKtAJwej/
01EonuVfdSRyM/D0342n38elxz04KWTaIVBVUsD1xJlk6simB00UzD8QZoqN+vFR
01UymmAdg3yn7Ekmxwvjp5klYPrfR2jttvQjpIKoj5Hjv+f5znSNraZVhgmUTFPq
/z4tO1HdsB4xGwi5ljkFiL4PfyjwFiXxWjsGiDSP3Dlw4SgSmkUjSc0/jyyw4aYV
YtCEpCoeCf1f2+ImIWCJ8Q5BXMJCU+D3M03j15/OMCE8w6yg47v0+shVCVAqkDnA
LJkLyxqKBJDo+duyEREY65RGlqM44FtrnW/RjsgFV1U7Rftcxj135d90S7a2U6nM
mBmZb94P4sRnrIEltoa3Scw7iVnfYIDtAo0DMRa3MELKK71nxSjzqAkL/emGmwV7
Tdbx61ik1fSXujd6PqC2n/stkZl74o6YsPk10bAQUHxLWbkwOTxyBuUzVKeiDj4W
V46ulwlfUEpSEmEaZvCv9tPonRvJt+VOizknH9J3wCGPia9KaYI5YM6BpAf5H9s0
GzrG24keAdiey0UHDGTd3CqzyPT9s7y3IQYmomNl9nFjd6dJzHt9pIxT5q6xr20Q
++VgOwgktHqTqZ7lViKda+BwdJhq3xBlyCgYJ4xhdrlxDopz1O1WdBf12dr2Zph2
ZZK3za/4uMJNs2qZW4OVxnbBNjbedeoiONUbl25kbMyoP2x/slhtYzGIPJ0u3wgI
UFshGyBGk5/Cgkw1AI2/gcrnnZbbjaia6bz9mLnvvELzhKsgbN5PuNIECL0QcJ+s
6hYLuaBeHnk0gWkoIrke0ucLIisE70/UNoLtgGD7IDkLri+DAhnOMRMw+WgbSuZ8
7/2AMnU9HzX5QR+fm4m2QujPIWfwuyeKxAF/ceHIeA50vEZ3EDOSfyI8k0VZrLYz
ClePAZrrNyxuMdx1J8DJre7B8eHg/u45Tz82HcRIPBE2w1C/Wk0IOZSxBSf6jEDF
EVlJGGo3c7kvt+Uoskk+RT8Wo8X48pSGXDD1E5wryoPnob8itGOLKO1pk7W4QTcB
67SUz2XkpQ1xTUchY10Zn+s0ZH7/04x6po8NT2A5hxbtocpV/yiGA172nggwl+A6
ci2J5oa8jLuQOb0rnbtZ754ZLpd3hWTxCHbrK8sY73lsSSxr+cfmHjM4h42aJnbn
Wxm2nWOjMoSKV+rdwoI3NuMCR2SvEXtcaTa5lYa8ULN5WgmT1/bGPZ/vLydTXNKz
leNuS0kjFOpaCHCLZgJUIkuSTaPCh7a9hHO7fOVIMmbpe+0VmRJ1dfTUxJ2u5JG+
6IBq7w5Q+QHVUzezbIsLjSKTmMPBRTOBH1+HBjRwPeftPdIKWp2lLn+kNTMJfHe1
7FL65RIetbBhsiDAkAwje4xHVrSVIi9JKc7DGyIcFiJZWA2su+m0sYnTZSNBaxWD
fa5zQThjF0OkBsQtgNWebh4n/pm+kzLKnvqbPv0qYfp3H8jJxJwtJx0TsroqvfVW
9Ro/IfL7felooi0RFI5GEXoNop0/ktfrdjUGD04w+EXxlg2HBAcCoi7NFW30YbP5
csa164Eh7a5/A3vX+L94FRJq4fdw52ay2f+KfmqqWpGqOGse9rc4uO5Uanc8OsHp
FOjMOrTx0g1UPmcn+fSWmAPJ3qDzQmm2WVffKFHjQIAPK2Fo/nd6/VrXxdplLfyM
Gj9MQbCF2wqGjzycjlRGj60LkCTOJeVi3/yWT7ukYKRMcTGBXvnZ0NOwgYiGkdEj
d0bJGhlprraGsdc1looV/ptwrf3QRkI/c7tfOgd5s86LFFOWWMYRLrIgAFJ/Dwjw
TVCL60kCzXuzHsJ2KvuqSUgQ8eRVGyDA/BX7pVNl3b91/rRRhehDd94hB0o6svZl
aamibKIJe6SdKpmbaTZpPXLLy3ywa9H+Jdf9vCrPiGB0/rObHycqaxW+h9dVtiWZ
0ZawAb93pzdhzLI0NJHvD4yBJ6VfA39IQ6hIRRPqAiD8s0F0HSGseOcbQDtckq3t
GZz83hUFxPj8yFavbRPsdc3eHFFSEv7l8O6qdIDUArUKiJt8NdVLv4zEeLGUUfIJ
X4C5YlJDVvXRZA9dShYDqURT/LI8wfzqH2s0cO2OgWPYlud8W+QQeJEoegXsrCGl
W0vuYWFdIi1+MBt1djjdUoAOKLdMeEWzWq++KzKHMx1zJ3lSCGhhV2CmUh9BflIi
Z8H952J2jL6w6Q34nXALH2QhyX4j9XZbRg/PIalIhqYfjljtUhw3pyzPm5JFZv51
j5LFwMiljrD3hsBYkP6EUOjhZMUVRhqwHbL9tyg528JTmpjxhJDx93NaDe8lVig2
UQakC8ayGD88FH5MhHMVnF7HFV7rJbBoowrzCBGXJaPK8g2Q+ZMkV2CuvOQUzXVJ
1L5yRctR5pX1Hf1boy7qaU44FwBFEFDwv67PMQSMyr+rH9UYz8pD5/U7vJo4ao87
P7e3SGrtInS9PQQ4RgFf4d9Nij/GaWtl8qIgXDw79JwWpsQv21KHIe0VavDFLa+K
1S4oULql3Vu2jNoAv5CFcvqjRsZLCaWGRKKMKriTW+aCHsL8JrB6d+7Knpb1+BKK
rzG4BSSz7VLYnyMpFGfLeHTXqoN1DnVTco22LOIzle1hQ0OBzO6sCqSp65awqGU4
R/BlHJ/zLoVbfb5VI9xe6Oxi4sblec8Qu1uRjFzmr2eZWLWFOvZuVg5AuqVtodIQ
yYKFadm+gZg99s2JQGlvwV7cGWfrGGkdE6q6MozUI6CVA+IIqmkcS1MjiH4hkynN
UvSJnBIKGIO3StgzNc7iDeBA5nIdYml2U9SYSKAj6fzXF7mF6/jCS/sX4O7vQFE4
DIKSwUedWYUu+TFTcjzmtGrDx/LedyG1PRgFwLqLJqHIcVvj7IfkFuXgO8/bvrpC
sCN9o9nCE9ClZF1rEQFmlEsUYbBOi4duAo7ItOTrLzN74RP77szyVm1AxxnyhWsf
9EiXp+LC/DV/xre+I/XzpuQXfUXrfSjIbf8tU29CTnu34Uyl/s7lCFkyX57MFLzb
dq8udzMmjiunOesB+FPboo+k/ILladCUNnbMUSiQDVM9Q6kScd1s5vUlHMq/2/Iy
Gg8hvY3rcHAyXsPBpeKjJmCzkSvEmNht54cyKgdvqNLfryx8cZ4QtwMqhpUeHA6G
EzKj6/Mil7MbFLQuwCpKqH2GFRokrd6xxt0klviwmsL3SmsUUGCtQ8CKrzAhxlag
ZZfbI1FOTfu4rS+9MPAIeeWeAev/I2bIioDzsBsWyQlC2dKQg/cbuHE9eOdvW3e/
D+Itl1lddCmU2a2YOJ0qIeCL+6diGWWDQd/vNA6VEStgah75gHPYSWG0X2UOqn95
WdKrWnWEJacTjAbKNHR7FoOfYhs4YIyWeWc5Po2H6sSmOfIv2/oHCBnlHiMO9D7q
OgaKz432Glq55rDFaBKY6gI+HbDQSHJYY0V8q3IxijxpUSCw4KHYm3izsTGS08Lp
Qogu57fWb92El7FH6prDfKPpwzj7FBq9yorzCeB1IxNpRC0Ttga1l3gmhUNMNGkd
fwvGIAkwH8noRQQHOz5JmcruFAeQL0Wzf38R4Gvjh8dz4sm6IAsZ/NxC2DU5smBx
NvTZVOISIElLBnkY3YIypXnVaPYCDfSRD7JYuiHkxaCCPKyXuoxwboE22WPLJ0z9
l1Azmb5ts1irmN7So+4J2l+nCZ5E8LVXWbqPJs1hlw1+wEn0HjOlcM4wsO5dYjWO
WFaSHDQKbEz1JCU5mLKxopE6d1WmshOfKRXoGH6hEmGqFQ6+aAVxfvdQR4KkQ83S
XkYm60gFzMpQyF1NmPXd+EBTQ2KH7uFzlN2ijhtCViVeYsTeFI8QJ59Tqq49GxDp
A77CRpgD5qmuU1zBng9mUMrds9a4+y+rrFCzB/mPlxFe6guOEPy/90CINCc9WNu0
AZggEDnH/zd2ALjRAu2Rz7NEdXXVS6yLZrF4KjWZfPT9qaVDhp8PPk9e0wX+gquw
9xO/zzDiE86/vs2SjRZROoxB1zureWAMf/q3fIBT3ovGG53AduVBBTsAPWFXjnIL
jG41R7/JivQV8sdZzzCKxFxh8fJUHAyGyjVWYJCPDALAIQQSiZ0ngo7KE06GUy8G
UMYI/rGCta0dlkBkT3h0xlU2JMyW2paC2jOlPagfx8+9/AI9g+hdij3mI0Y7Qafv
yEkeV2aOH33DRjNRRgTz6L9yL2Md5mt0oP33EZKx5mHyEi3dvOuieyaeFBu61Zxt
fTrrfwV+QjF2RkmzqhmIs5+tQeYr9dMqFlkXZW8/WlDS09A2znK2LNjfIV3zgZj/
ljiRZqptn7sEBM5WMBWratoppYRX8LH2GaWpPp3E86vCxxXawPjU50P+8Lw8CBP/
GQ3hBwl5RKTbyQWCPkATx24nP+lT1Mi8qaoDb1qrvwAEYz9SHDWKjTQSSFxGB2uK
6hJZN7SBdtSVrp00xNcUp15ZeNDRzYlxGmufHaXMeCT4W4r1ewDMFRuCeYThGoCX
m22LbJd8YuXoPdfv+PegO4vQZxrjTRwK7Mh/yeF8pdTNkcWe6xWWTDLQpIjNNkvI
90yAgp7HgehKXVM++FWruQD784lb5BbVEu8m5eu97MmTyPGo9Q5SpJd79eTgfu0D
ZDsN+N91w8ZEddSTXHeec2YH1UJhM7SeV9DenPGG2D7td1bAqGxSN5gWgR3OD2ds
DKZg9/BKUafl9gBOgOTvCi1XGkkGeIqqGJG3cEK4J9JJ1k3xy1pLDltJ92cBoNpf
BzcwWE6Y/H/K3PcnOIiMrUrAjdo9z7g3XvS3LovEn6EWaKPhtiTrQ6WK3G+3HDeA
9EQzJ+lTTEZk4fuBxl3zBmKuAqJw8b1yA5oDvezeoC3SQBrx1rY2Sa1mfkFF1N7a
/g6PvxOjHv+YjlZ6Zd2+0u08p1j5eADqiDK+luYTCSwLg9J3LmrbOc6v7PMXG9rs
lJWiH38Dr0PeG4/WKlejwOx/fjx12q6nZFTlvsOp1qkdZBJXjvyFqw8Uh2U3X7AS
WsdzIWuIzCNnsJG/V+ASG/eBE9qoJUu7Hnh8O9/x0H7aJP44v+G/3KlysGn1RT28
AigGwebImzd8XshRBE1seiOusTulj7hFVxNcpGwFvcJq7xTz1PoiI3Kp6hHNNnEf
wCaofPuA8/c7wwIsznmL8/e6VVlmUCnbMducCOgK7cRPbUtstvoofQISSr13dCnv
9qB1sfqCqd/9FGj/4nrI0UHXYyll4OhOaT6ZzKalgwor+q5bbN3FRRykJtYhocj4
E63wAnkbO11hf4IkG99PzveD9zNMrEEZN5V6XU6ffCN8eQsxqR482sdk08dCsO4l
rfhcg6Dk5KaO3lskCCNALtmzQwWJyMlzvCQYJhp6lQfEW+eZzm0q/XDG3wqD0Jmy
bpZJ3r21qgK6NbLwWbXKCRKfbwbyTSxpx1XHzsCM4R/3gXt2jS16bBx/pTzfcz62
holQjp09GdaPGeG9pLHRCnOmof2dj+IXV1jH1MJbXS2gbc0amgI6WpWaagpzWBFz
UzvLPCl3IrZ9SRL6FclGulppp7En0+bhw6w3QrKzmn0CqiZ1DiQOTvqYOoge66PI
a/Ydnue8QtPbPC9Fbh5ZOWttHnmuhsZ4UEaduxVVWhJHKNw3ZgfZRPwBGyyXSjui
R+WHlWqpYS6NG1agioboictSJgeeMyzWN7UM5D2kqRp0Ed5gWd/0TVHUs2WzjUUt
MEwLSA5Xj+0jganSeanEL9XgNkgv9AMU3hpi1GKx2voA4gNuScOZNwBCND6ylHjF
Z+uT3xR/DVKJDy3clqW2NbxqcUkINwSkpQkGNaNArj/oyc6vORzLHxeTKPt3pVh+
McHusAEvoMSDnkbVGb+ofUMwRd59fNrrl7AK5LWjsAspt/bvkQVsa3/fYablndJZ
LveEmcMtK1zU+uGqncWB6h9KiOiOKzDFkgylVbqcFpw5dvMgQ2cIqNsvfMmymCos
53lurCixzp7xwFgUYnQZDI1j/CvBoRK3VKK9NtymMeYHGQBk76Ky/ae0yDeI1jEk
Y3pWa4NxWwGuztSTTcHpTj/r78zAb7mDFBtK3JxzqTTKk53aF9o4c+AWD8srcwjz
5aUGAKVNk7MVvNi1y15hmCDkSogpLERoxiP6F2d46S+H15l8QmZsstfbW+VREMgD
EXxoEE1LQF8++soiACCE/f0qKQVwO+QsBgvQUo3PQy9BW1bG9rVc3guy/sSdm45z
LTP9V5j0uZYE01KQA09KwvP3Y3Rje5WiyJ9INglzoBez27ZBn6cSLw4B1ACJChP6
yyij5XNeItUt+5u85iS1pZw62WUJItPr5ZUJKxQBjdqY8UrGFfPkAaNZtTlUPxGd
KDwfxE5r8hsey+EgVhF6SpRsCGgudeSXG2AGOtLW2pGAIIJcWyC6QIvIxVJG2Qhk
HDxoDkrHxhketrL/cu60RlQrAZTiD3Sw+G6p/KvY04fsFdqxCYOUMR7okdG4iDDM
ZfWg9JWkwsXAW/5sDr120Lu5LnqdGVHEnbzwKZ3w7iMwFwSnVic9a6efGopR9a/t
Fn1yWeSQsWpbV6m3PXBGjKOl1HsGzpf0xl86z8QL5OPnw2fZjGFwgmxuVsVgx3cl
STmbYcJjksyGNiIIkRCTMKbU89SvKfqkpeNjLXjboRqw2LuLxT54ToRB13EHc536
qZQjnR/cUqtOK2HP1oVXkKVknbvFxUTLiC5/Et+9k58e3OxmrsAfsNCPcFFkR3IX
6xEUz39QdpnIYPwrzCU06ggcjura7PJtMjzfwXaAzRqY9hX4AproyMVZbzvLQP2F
is8JL/x7KFJnDxLceCcqS85V3FO9CPFKR+Gff+/w3D+vk81xpHcx3lATN5FZrpGJ
HQ1D1u3MtybgpeniiUOZOd699Tfkyd5M9WpixQNQWLwKcqA0efV8Yc6+jBb1OY/j
5zw+0hzFqWBz1DK9aliguB9t/1VizM79R+b6ihFcOlOs09CTUiEtR1t9D6ihYuFI
oYOZjVN9qdDbQdaVedLh6N8fSuttKp9jkqiQp8QqFOTl4UEGGO25178DhpvUcFw1
096Qld5FenN9NDIZ441t0ldqXOgpXLq7/+DkanNWo5Px2odKrzjAogGHignQS/IY
NbO2COhA0VS9xHtzYKZm2agC//da4CAmvRmJjSsxYMkAHGXp388mbtVChXkYA2zp
fIXMBFpfQLNPJaWPc4Csz2xxAUCXHKPaBOOyDGY0D1WNSu1pYoHfyG3yItiWXZvc
oHd9b1tfKaPDzisf8Yib7AEBbfUeXrNl29yA/E9TuJtONe1KGFrh8mHjqIWsJNhw
rF7roKmEx5mte90jkAcLM83TjGHm5krkgcvvv1FJ9RwTXqxHgowDIFsvPFVQ6fqK
Mvz5vY67Vu5ZbWZ9E1/dASw9qVDwYy+n9ZgDfQRz0MV2DpYwVTeJdgBLuey4O2i/
X2QYJCyQJd7jsVBFk19GHImdsUPo7w3n/iuDNDAwwzUVF9fszBorUgb2zoXJ2TNW
HegNdSlEivKq2n5IZUdMdxPdpel4wazgrDT+r89u1d22vXyvsu123lNzsY417cEg
gkp1lN9RTT2f4FI70MuE4dSoC7XWxf/Z0lkXLRzywsAaSlTBU3MnmgXqDqqksQ/b
35GdGNAsNCEFk/t0IzTZZLJtWTJMH55umGYFTm0ctHhm+sm20nYxn/Qb1fjTYcTP
7hMd3erECwCBDlCjdaAZRYZ+AJt8l3/+U7QsYn6erhWD1KC2xZU04XCknTQba3JH
Sj+sM1pAxMeYqA1pFpKs77S67SWfH733fQQpOEOFO/D6teTJdtVZ0F2hcyIKI3o7
Jw4xHls0r+mlEwcZOZ8okoTINO7J0Dh67iGN+68L8jDQSjR2388e8q7I8OW7/l1B
UTJ4N4KKuwchm2Uhm19xZ33Zmd70r9KRGhLKdUrwAC6wU4iiGof74GUhQEl9fQiq
E1UDYQ+osqus7Zw8FiOuT/c3Js8Cvgr2FCd6N9iC3VbH2sy+OMU8x9MoTk8hUEyp
WP/PHcXJB2z0IGQrXajuLUlooKDl+zPGoEP6OywNIenf4Ed40WLgmvMIpej2O1CD
BG2M56s3QBKtvb42g2S9JTaqUAnZwm8/7lDHeRgArQjiF19IVIe7pK3NavCMywjF
nxcXpQ9YGWs9tqoe6k72OvQ/FqzfjPYXhV8JcObjcAdIQ4RgCaXunvH6eVOVHrKR
BiOJhdF1BwHeS3AHuwAFrh4eDOkto/qGu1U4qVd+28Vf5lYQNPww4vyBevl785PP
oyUPDsrAJpHZcS+XJbRcIW+AZh8ETQ8NXr5hSBOJjMT+WgXWuYaUoBQo+gmgbf1l
gr4v/KB6XhzhE2p5XSOSp+7g+KqMNBfXuVUGhMsVjiHVRMX/aIV7qlEgJaDhLQ1x
zaLb2RdOPL6CtROtG27Jjy/8+Q1jGHtWC5/8UVpYFn0ocYKm66kkt101rsPTNh7h
HzEDpHUinYE/d/PdIc/cVa5CfeoDtogkUGOSZUvPnGU4WkbXzREOmy9mOqMaHy0B
cPLUNO3wheRKWwyoimcd5OWRZeCfxp1EOheIE7HNSP7ThIPpCw/hyduXQU42Bwgt
yky/f9/Vase+gxzXu+UbHG0Uhrj+7GzdLh0lz4BrTR97CYVHWHSATWgtp+2EeRrD
wIKl4Y1zIKuretgCaJVICFM0kdgfWKn9VkfBHWEBKxIlTkCwFlSfJnskWFNGtKUY
XKvzZidoC6RvKvaMmndktSimiVefHk4GjuW/++rnpEZs/CIgN+zfVfv06IsETgF5
IKFYYzjU26YMekAHa+BHpgqBO4yD/OIt/sY5X2zKOYqLuj/L28oNCBAUT+p0ZRVj
2lC4oma+qH3q62PC3qHeq/ivGv/AZPlovEeE/nRP2vHLph4MvcqdlfbVcwxg0a/e
0cTwITBDrj/CHvAPu2YhJbIbnydAjy0XVXmkDZ849yXRWnn5c97Yd1K+P18CKrP2
YItA+PW/P71guu7RUbh66juWpOi4WU3SNNVDLFOHKhRhqUkDb8Orok0UX09/GPiY
F1UDLh2/upMb9hEF1kb/ABckpcX0Ja1JRRY8MxmeEN5XxZWX1ilg/W49A+HM4UXm
+8mgQPpw2+DMZpOqc7oWUkmB5hOloIAtXYvao1+LiobdFQ1EAbV1Yn97Id2+b7u/
gkCItueUG/BiXjT80yKY0g2KMsxP7Ac/VzvIHEy7hffv3j00GjzMUAcPudHDBfaH
bBjq4unxl5gmT4tXU3yz7R5Vm3e9Bq0jD2daJDklusTNijzgX4b+Nv5YyhzZsuht
an2VkCe9IWqnl6WQOvXbqm1VDU+yCtIGeioIV1OFQq0wFEn8CEOsPV5i3hBwSa4V
Ob8mzmqrR9LGD4GSAAkyG9QU+yLcku1jDj94BeD7O7tOiI8ltOgaYFSRG1FN8CIN
eHoTBAWKQ9bZP5bRCyU/OKIPC4rIogE0ocD+PoOx7F7oCoxl2TzwVcTlmZfAH6N4
NNA7Cp8p9uyCg6p0rblPHRPJxbbimNfvNYeuMVqYSUc20I0/cQelaEpSrl1dCvK6
1vLlF6ugHCskVM/7aTHcuSi5O0sfBVae3ttNkl/JGnS8oWInKOQGv18hhgzMWrEM
sarb8EVayvsr5WWZyc6nwnufqFnL6TcdzkDlLXNuAyVfWa1cmcNGZiV7jM3y4ZhE
RILP8wqPR5wBAiu4v4JVfxNKriGTRj7Gsmzho0jbIUKQOvyv13mui77lN/RwE7Ht
TidCqUaZqdQoT9CBzQY+Vk04ZPu9s6xLBxj/lBt0DsDGTKSL0rhU/BBN8SWJS520
DrjSLyviiM/QahEVqrbl4e5GkUXWxTR2FaviKgbo8XHWXNaVxulzEqmIhlSV4l6X
tccVxnGY17DIYijQZl02tX9bBJEA+cay4RYiFvf5jBUisQeiVkf9r1pY/v9A56pW
uTrTb4vnKKBgDHkx9JlMcJUqRQs7cWcYpEuzl02ASHTCAkGpzfn675EgFuy4X5mM
MRqpMU1aXgxVjcXTAGTeliWPmgv8SG3gnAb9kgH0803/ZnPVOMokqAedSX+XsP2k
49bds8XnnEvTaV81fzp3fom+dIrd4JIHEbl5T+C99oTJIrlvCi8QuMJ0/xT7AHqh
o/4vT7CERVzhD3LGXI1gYLnWsZAB5FXcQB5ydnFIinNLP9dcK3WDGDx+O7JZPQE/
xUQXme7OSficHiyB+mcCff7pGWuLwVIrg2pBSHHoP2UJ0vhMmQIZYBgphywaAMAk
SB4rDVM2Fp5R5OBPgKeiXorF7vYbvLZroRU8Rj5CYd5103bcTh0Ey2c0h0DpN4tB
wNfp44IkbS5seivhJVvGqK/T9pYE9aOsAaobXBZJrsX+t8204gqqJ9QSwYTARVqK
JoZQzlZAjNtXjWrVRrJWYhgf6VFyjs8Gif4YGVV6Ep5JtKgPHm3U4DR02sLQSoGt
K+E98PNqOMzetDKNhprEPsO1+QIjJo1pyiKZlQG0w6CJl9PKFHDTJ8I4blwzGOc4
4/Hkye+VDcyUVKUu4ZJ0DnedxmGKQN0BnwjzokT4wjmrxy+1tlNw0yuKqYdyxxcu
B9yGCvy0VV071Ue4erCpeHgW4Cb/SqpwvfDXouDDHqSUB7tGedKK4uU1BZE5G8rO
oVuAMUBPG2oo8sZaLsvi+zIf+VHscslVY+gkXBvecRy8E8dx6DcaXFLJKsTcm9KC
VaZ0W9MsT3JrHWtXY2VD53+tCLlKTbhTFaiIo7PikNuHUVON564MuW4RveIjWKU3
IBe49vUwjh04HMr1BjNs97p8xU3hmcXD4GlKXVFzSzLJRmNWk9htmywxwAss/oCm
VpwS9kcC9SnU6RF+Ab3jttCk5HHCQXn2tXkIAYaPwzgg3Z9pZDfwdubvnn8PL4Rb
rfmXwKPzV/fKa9oMTa0PvoqU8VbfcCWRL4HzIktnukrMPqCcsUYQN91yXSGnMyl1
UhnxjUvMdZYMVh/8aJWBWL/Xeqcgl3peFuSd0Ban1whZXwuURy9GIpqbtiJ4AZ0I
BD6PrWQf8KpgDztiuVJFzlBdsCJ++n9x9qdud4nldGt0Rdsn2YfEAlLg08pwm3uP
OGnjWpxB/KHlKERofiS0tCADE8GDLUY+byNCBFzIDGGAlnJvh3gKOupdOZbvNPqM
zxbZeWJybg75UiZy+spIXQC+BSgrk4OR3pSN+Cwdpw+Sowo6/LvoaDwIwgTekv5X
a7uM0u6JTpEZ3NZCS2/RY5nyzAyL0QDSzSG2PIF1O89ue716fSZJAgKwMVkonR9H
7xNeyFOXP6puhIH6311P20GIMeCjuKFyQOQvJqu/JSd7JhzhnknuQ2QkrtllnPSK
m9wFIpru78CITs3I0d6ndA3m7cIZlneIcVlrUjfVftQT2VQXUxSsv7vkB4zox8aI
NGkxht9YP2Pe13+2REIdCpcJZbinbSehoDHlLk56d9Ncg90ExU62WHOguFrvhx3p
EhLVGfE/ML2dWdj/DESvFP4D9rlK+/tnb8H/JWkSqalQEGv2bBPnGAnyo8E0f4uG
4BzXA/I3GfYgVY66TMFtih1LsfwWKe6QZMh3Vrptprk/IknW6QZlwvg42PmX92m5
0I6DpLReVwO8IjMtjMvJmXDFov07Azd3hl6Vt0JAmDp7c+/KzgvfzXF4I94MUH4n
/qFztwyNQBYdhydnrlfKGUE1mmZTyfx+svTkHfcPzQHjIRXn4lxtDUsITXIuxkia
J8FWQb39voDR4HIpZ9ss+LCllVa2NAYb3Px5/IKLXmI3Um4LDIBRCqRcIvFE0ysA
NXfzu3kxtyal250k8Dj0d6vM8EHZ/MQ+tVIY+hgX9E6wYze0w4c6RcA6TxNG4wJ7
MWSs3qDDsMsN9vidUSHQuZL79Az1+4JXsqSBparrLm2G52X9veqB6zDT+XRMbhz6
OtHiUsLr7kNiGXpQ7LzyBSLvOyyE9dezLOpKS1W6zGV4XffbBt2HBa5+kKcOJmkf
2vXhK5tIdgXXDbD3yK7YCpPVXVOmQtmQgrj7AmMl0gYjIKVn47OI+6EDeLgVi73W
ZkrlKO4bhVLT3kGfsSPLN+aAXCGeyrpQteVb4HU9cyrzDyx/wI+DJV0S6sigZCu+
BGqasuystFkHAgzrMTvz8HG0ea58CWwVg3iLIqCMU098aIQPMXEfBLYRExFQAjLe
UNYyXYWnN81MSMQ7BC69k378MF4nh9Aqj7kikfWpvim54tdcfY1/I0lh0kwI0rTU
Wd7ym3bO0YO2I2tBT0v7V6aOgJN8OzDN9KPPRtMLfXTrLZgWcdkTtDZrUG0zAxDW
4AY5OWvMCtHhkBshEZXkLij3ySdELTTM1U09eIUBLwmCWVJGdsBYY+6yhaOLs0zH
DRM5Nf9+1TKr1YxSJS0SBq6CbRYCI/6IfItIrU8cEMxo2Q23FVOjKJ+k66bNi2or
J3M2Rh0rlSMIs9WCNswClGJJz36ACGH59r6Z19LgpwxtLMcx/+dsyYb1SCzmPMCk
C2JEOaDe4LisFbd5F4Xdy71Jwb9yGY9lAjvJUumu4eLuC+A5ViGt5u45uOMERrcb
0s9K7qT6h04Dbm/JNajmiTubfuU+VErZsxcnatyebeRRvxSbcRus92YA8ibwadSy
8IzwWTaRtzs7nJzfVy8J0Fq0eYykmc5AyRYur9S0bZstd12IcywACiDuwjMWFQMp
JX2PrEytqwA1qpv1okEGCf3DaNJs/4skqn79BeasPWQC1nhsRmkcmCDDA0HAM55Y
nrZI++gI6AWQNbN7GpjxEw==
`protect end_protected
