-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ZiajMxy5IUowZPXNNofkY6OcCyKj9Jd5Bmrs3f2EMYfrDo32LUSgYiyAuUMPfyq6
8KnLFvFzp+wsHCY+GUc6uk6twmYAJCrGE9LqPccpuRLwDWs5qhyFM1qHIyDsBhVm
ENSWCZRiwkHqh+JFDXQbcBigmaxbjyIieXFXxZsuMp0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13549)

`protect DATA_BLOCK
Ok3ehXriVtpQJimWfPFAA3zu/vKBsvhxncdGSUXkn0MOn/o4BYxrRd2iQ5iITjLs
05FF0rYPDKoKrJ/oo23TR/iX3J72HPMMAafqIErcpCRi2/7yQKerV7Cf2JM80F2G
r38GbibNPeLTcvu7m2AiwKjzoWjumfXPdyh08+tfuCn1G7NRRnifC+p1wprWjldU
3iA8Dc9x/liiogfxnYc+bhXro5evjetBpF2MdQSRSr5X6D80ZikAI5RgHj9XD0jZ
8Yemgr0cYtMJyjkb2H1CbhMQhHjI9QFvyYKmUIULlUO4dwwHeFKEzJfs5/qbQmfN
2lyAtqqOQtC+op4LvBRFx7OicIRDS5LLTEHgKvtSaNAK6MGDWbmOYfNdf8lMAunl
YxX4FNUcSHkFgfufznVp4ByAVJXsRUEmH8qDyYrgLN/OLsV1//aQyeW4Cp9oBIxZ
pXUIIJ/UXUCU4Xk3XG8Yj3SEdUCdYw5PO1l9fHBzThGtN4Se1ckGbcN08ideW2eu
7FMTbA1K0UIx58E8RyWKgscOXMpptsHaW5WjlcR7vZx8hfG/e96YI+L4/v+Effs0
+/2AM4HRFlwvRWFmD96jq3nOWARM/fwb4+sekVeqkeCrKMXCLqsEeJwSnXhZtnnI
dkUWwJT36AWcP8tEaNdbKHJq933vGdPiXeLw8ZG1aGg3L7veGGakWvHYQtr0gBoT
qnBpnfv+kgVBG8tRZgZ9tnxfvE2cGGjM1pFSuSJZW7yES5gH4/vuwvnu+9IaDpQO
aV/m3uBHAVEg3fqsrAmtXYpvnhEvjfRL274To8p9XdBbCMbKcd4xaxpONJIUrMDi
UIijMeeZR0V7Fe2xsDkAwZfUu7RqIlMOwuFL9+gopDpb7UNXMFCFLL9wBNk8w/HN
bTs3n9otJQ1Oev0eNrpS31WJ4OU9w8e82tmD6mkA92HSOozodHOvYRiUqfJvIhaS
SKSw45sXDLwAUI18dd4Yak/22r8HPSNf15WDMJyycCdBzLGUgvhPr/mjrcrrncOP
ElL21DAluG2YiTTvS48jpvnANGmXsTYW1x240IkEN3pYxhJOQg46Bhy3+TAjynKx
0qxEBqRQ2y0i3V6Pra8x9qfcvRZz2VgTgYoccnip08XhADo+GNjCK6tNqrYnN11U
0IEIh41jIhtY0j7Sb7YKaAginWFw6j7bOz7yowB2Ip3J0TOVLgrAG9ew8BQG7GNQ
CfLiC9o7XIeffbI/h9yBF0M0mQjLsfv7Jd5pW8Udo3P+eGt21y3mBsi29Qxr9Cp6
nUxDGYok/qrA6vEpKXUvL9yf/1kRUqB7MvdkNQ4tV1EvyMoP7eAFH9oDqeKw/KAN
QRr+mTR+Q/z9njKvGyl/2doFaHZD2HNiWeQ6sRAGzqJqWYX6B94fjw6lalq2hGtX
64GBDZHAQuDyqIUABwYOQF/iaq9SK+axwypd+WJaf4Q5mg/MerlOXCK2R9UkhuSR
iE6yqjbpAS9c0Vb8M2+zNuzP/jSaLkvZIMaevJqlOsYQMQ3HfYQOYl3b6ggeIn+o
IgpD1aW9yhVHgH0Id0dyBF6k4CKgZBwMKIvBq6MrLQEzVtIChfubMdTy1BD9NQUn
NvXln58uVGT8Wm7+aBs8vii5Lck/iE/ZtnwlC2Nn7UVgo0rWH6nkuLiavNQJohDn
J1w7gACNBuxWOiCDTGYd2Oxvdv05L6c+7P1IaP1jMyxqSCxCOM5uDoE66SRjtL+t
yzhC3RDV5l4rpcAVXtJP0XegL8l9awq+Wpm8vmjtCLI+0oIk5o3Y70CIGs7j0mtv
DwpuspYFLRLibiXrT+0vDGESFIYBIGj2UiN595QbwhuWc86yhVQfoFtS1QkJwojL
N/jEkSSSwzWaRoOFNvZo74THoMggVDpPP7wCGckyKIQOTgSVjiYOtGPt8FT9S38J
T4TRlcs/c+efZPKpUlJHu0+XxX5BR7KZYZIg1vw1B/Yx2uGBqTKUG9b0WLcGs+Xu
oyMcC7ZOIzDpgERrIUxUZLGdCLqRrYgaUzJsuBicof87oNDs4+/vJyNCIGsDYLZh
QtjyQ+WZx5Di5l+wEz5EA/VGdmryR5aBEnfDI9LCtGSfWg4zQ16+sGax840EzQzD
WWyQ8TC4Z//vgGSGDAS+OZINtPRedwljw4aIMZrWkM5Gcuys7iqLDqoNxY1d6iVt
OFG8qI5Ri6XacR7aisw19MvQIQAXKYHdg+6FwNEerxUcr4MkhK5MGkwlJa66F+cP
8IVmA3mN8MTMW2vEU+swlDoXgMzuRRDmBaRoP8pAoY5EpHazCMPPfzbGMBiAZuO3
xxYvSrVL/Cu0wvmQzEzwkiaNiMfsfxLZCDANMK8+Infr8UYx5GQsBDNXMvQQ8/JS
Oo/DWKx4YBtC2Q8fHPcZq9giY/RohkWz2A5cN91U3k6Pymtds9MTnV5DLu5J0aHl
lcHlVmHaosO2KgOUVSrDDu+SGFeiUArAKSSz4679lSNSdnoQ0LK+gZ2IginejO4q
oRuJj88zMrvC8tBlWlSLUuIhxzBE1M/DSFgfQmliGPXx5dPanfIGIpb9Z349hVoA
zCit7/UDlL/ZixEGNQqiPyuXqgAcuWdOaKR816izRIkFqRVAU9B8C1/a+aKkDOD8
9i6UQEjMwjGo4gvj+AEKa9UQ9WNjwD+usGYjRN6r+kRlAbMhHFemwZJitpQDtWYY
fqLIeK/M3cMOEWiF9clFSRt+oJhB0Rm385EEPk4VFNhh8xuhibZBUfQ25/yQwVdj
hWrA+VLJ7PQ+QbRKxVVMcAWEKM9temxkBmZrzS3osb3NeARtENRP4FuFIpMi8i2f
szV+evf6bUbrJzvbYuZLuhb8t6dCxqg+Yq676bci5Jl//wNUzhgvHtyOFMN5D0AB
0picJclQ7iFti1LGsvIe+vOStD2mX/DQWB23Bhg96M+xfKFYz8ULpnqnPhfQQD05
Z6rdjFcpX5fQDZcM/S0CrPevY/uCe7wUqT4YAO50W+3ntgBVRGRJjOSn5xoy6Fuq
Ua3zo2QQXwpI7/nGVxvI3eGwCM3+5UzaVXehrBA/k5fgDTjoYKYV4v4cDVPivWh3
Km2AidKcaYsM8jZQB8CZw6y/NqkVBwyiIL3GZCUD+3CSuW0YcNWeOj+90bKPltf2
TVqI6/IbKVAlIfrE2ZcbS5/fxUW8I5FgFDDAVXuQVKMPaXMDlB1HYQLfV+xu45IJ
s1Sg/aPwT4TVhYYxTSbVl3azJJ1osqQexvhW6nUgNFMgm11vB5pbc4eb4bhEYahf
DdHf7PT8J2XspGCttrUo8ROaOPnQidZEgxZZEBeX4IVFWWIVUphjAqCVOdAZ6q6i
EVwFOCXYLcZ8R2se1iMRALDnHkYmLPee9hZuJAVY398GOCeatwNtfQsdqsfXxA/T
XShxUslhG4WQBI1OWMrjSgnUBWuZc642qznqh+AT9mZNay6uDp5VED7iKKvNExAg
H3WHUFkWIivbTH4FutufAaiY8WjyON+flfMBpspTIXLBfcrhI5McCCtOK9pZXpq5
MaP1xjxIzPemACTYEg1XH3jyvlRk2/coqQDyIQ8dpmOFFpOlRVFRCAVXdCugv8p0
Wk4Vx8v95agAbDbfuhizL5VHAiV0ajkwqBtzsxwLf/URoALJ1FPjMIdUfI9w9CjA
6VUEUU9CjvAbROsRuKjSut7svJbsu705Vi9qJRWRtsCn2O/okTvbYntsBoaG23Ba
cWkmcR+M2InbYDTiS0C+Vs2+UDpIuJAbff/MKfTwuQ66bIYDlRNmraDwUjuqAF3W
Vpwp8iAb8Y1c8vXFBPNwrTq5fJS4ToF2PD/RG3B9bT9muDa1/Cd9xiAJHo0ENVp7
QF6F1wWcsKCeUrXNuckLnLcAsX7nhh0JSO1RqGDvArhgXIRG2d+Z9IJQRxy7g//5
qKYNWeyX6c8lxJrk0vtlz29EbQSIziamBS6Eu35vwhXQa1dkAXlp2MEqSqTmWwIh
jvq+Qh3eZZUAjEaG1GoxrZvH3fS/iO3Tz4lWczqz0ajFbi1gHNcMwIyyhCEyDFqJ
mClsWei3nLp4dNaxRfBtKNPgeqBUkQinSEV57AOA6bsTftr+6a/j5twjhix4uNAV
MOt0ghfuvuDtXew8IUebk2oZmzKEBh95gIvw/VKg7nruhowmRlm80mvkm9wIePI3
oll1hTbQ6eQS+AdFLu9YdHIua8d6Zzi79fNVuwzdffOUCBMJ/jWbYNQkk8ZBm7ee
WGSmlfW20lNN+Mu7kIAjArFiYgAPgFuNV0e7flnbJmSlN0BMD1JYsDxhxizIDNzF
bFM0ULDuEmJRK1ki/U6Ou2qUBuxAomBxeBxpoIQed9L4TiEM/1ARn+hepvHsB93T
8h8TkHZU/avCWm/9Xi1LFswdVErBnuscqxMeVh0z73V2dgFSAdPPEWufc6gQUdXd
+5Y2nd3NXa0JrcvObHpLoJUfPfMj48ozPsbYeWoXnGO7zAiRN1uWYOHlEjDSeJBg
yN2LvVq7SLO00a69k25m7dP6sWZ1vZKabWZ7jXYq9m2XDBI0QHUPuHAfi8CAN9Ln
AcE8ysriH8fDNor+9Im/Fc3MjmmD6Bnv81LWGE50hObq7h5mb6PR4E7oJOmTLVPw
T0s46yncyQktuDIygND2/M2tEm61OR0VUIYIu8PT14WEXxNd73AwxUeyRPVGTCnH
kD4Dht3Kpd6sPWa2GpcfHzQM1MVeoCxu7WCe6+stUYzC7k6sbyHmBbM7XFQUemXD
P3yodLztTPyqpQwKBt9/Z25We2K4XpisiNJWNttW+RZwbkhEcky/FoJNFovgz0Ie
fIf31dgnznU7oOIdY0sXT6DgVzccJcHqBxbjMNCmiBQtVBd4fRZW4w1Ichz05NL3
cvPmAmaAU/rJrMDPN+x/x7T7FvHNcxsS5NgnRQbVsUAC9fdgmz1TgvYago5rOOkq
OGWxK9vPbwM6oJauUwJVWqOh4ajo8bPNxKsD3bN6AyD6evi8rvs17NMewhS0mbL8
5dNhFGgDojP8r7URpXG5Ngxv74OqhpR/OOW48jkav/JxwyVKLoc4cZIjXUF/h9a9
JzLuATJWRhfnnrnC5vYSoibCSw+kYNfkOZi8WH3gIeiP3aWZ1z36903js5wTlZAV
EWZ4aCq3X5JdSqH8UnHmR1FVpnEMXryu7WbcZsDYxJt048YEylx0Eg0AaRIUaJIB
a6RwDwVBOV7Yq0ONZoVrNaGkZWOrO2i8q7E+cJsV/vChkxKeKyfyuTOOxenLqHN9
cdByr54hur72Q7NPH82FGC4w5w+4sExGOsOgB6/3ir/xgLaEBysz8RUt5+zE3Kzl
Y/aD4iHzPcNqYyujC9bMLEgjibhP+enc7CkDOC2Pt9m2ySluy/g1JmkL95ChBgwE
H842zlY99iA1krgNFmuCD2V1A9Jmiyy17/sBne9AowpZWEl0yLSWAF1rsLDmgTRK
VnUEVinWZevIaNMOlYWAzp+EjXaDqg8x4QLHqMgCc3/oRVOc4HR27+XYiFSYbOtI
tOuLZ/UhuVoT1pd109/9l35t9VF+bVzeJh6Tjgp4KdKA11/tu28GPfhaOEATJ0uO
6KbFR5JmO4H6DKEhKsLxgAZx89SSbFmo+4rDmVkavvEKOXUctjgnOtNvf3Ty5Blx
4E35NxnIT274EBocbWzvj7hnJVELu/nB6Ip7iIpndLCYAZ2glFjmaWV1Jy96NQdS
YmA/O0ifXIZvlMiEzjr/q0PCRBWH63zdaflmTGCOAW1zoNtx0LY0q7cv/h6zUKoF
TWNdnSsxNkgpjoDzrKr1ohApyPJfXs1wkIWUGVIgs76RVP5S0H7gtUbrk8nsROzk
rIm/t/F6sSLGcuI3uxaKBrYlGgYCs/YPU8fXzKE9ZsoNePOzrJPyBgP7BfypfYxD
dlNEQRFTJW/8uA5e+X4dXDopQnjacKBb+031gg88EuXOc7wXt1ZrOiRqMaafxFMi
riKxAzORYyyJti7aS5NrtsTSfkc1CghLmkNF7TvEHV1KSh1//PgBKAOuyF3S4++C
iZt4VHWepkFkz5Pje9dUJQ5zgmYmA+tpZf79OQurXF4NQQstqxOb49pBmkFSktZG
tpE56oxYIfgbiBsp8PkQU7IBvF5xZcSIddUllyupOoC+3TKzqgugPAfIf0piB/BC
bXw1LtH5b5FVI633LaYxx44uqq3oZiXVS/aA1RYQKAU9R9nDl+/b+edWEaFjLp7B
ie3Z+gwTZILM4umtyPqd7XBq1xv23DPrSAWxF9GacfB0i8M48PtmMcXLKJLN5ZT+
CyAHlIaFjLd6GsYEb22XiFoXzXX8TOUrUqkedlpkgIzoLRoKMEgyJJyIl/8ITqx0
I+NRf8lOqifX3meQv7W7D+NbwDPI99tYOMNi+yJo+viYc2M/6uBdL2PEosO2arxc
/bI64ItIs/6Yj8BP8vFY+AcVkpJJZDiii/wvY17G9Yh5Z4Tc7Rj5LPPEE45sg2e0
QU6emCud3V9QiLIuvdGLiFEsCl4frbkPzoAbZ2CCuNeTbFAzoUKvEv2R24Zk7QP6
CfLeUQACsaPP+exbChM8FEf9yxHdUjaYhNRc6uhQeaz300gaYdJtykLaVm6cZOSd
zQp+nP5GBR08HYVWVFGJlXIcHwh4Fe5YsTU4X/VUexCCJ6xZj3xPy5XVpjxppbvh
rGZTEXKW/0sHGN+AlaoJJZ7D3+l32Bf5BEzhgaTtXJta3lOefNxHbdpf5f4q/YJP
zQJWNS3rpYfTPPCm5lndTdnNdCEt2ib1OPIO34lug1GL2b7JcHQWfttrGVw0dTK5
b8UGhaZeq4/Hz13n2h4y5elskSl5Pyl7Y1YPneRhPikfAW4r4F9Tes1z8jkgPrOE
axyeiBnYTn6vqpvdPruIDQ4nFNXMfFyZTAWeyt2pFwUYEfbvxll+iBOf+flZGuCi
kmnA6JZ5gFhFvv1QG4pIJN9rwzYR+cte4HRfYGgBx9Kl2Mj9BPQCSl3J4asmdcMo
rV4iBokQB11nxCZ16qxiQDy+dsDKo0ek/5N3z1GJbL6KitbO+fOrpfWUGKrVN8Qj
LuIIvGPH926Ho2vnKKUWFgXvSbepSZpAxPyQoACKOE3pNa62BkUVPjltkWzK0RBq
bpEzcqsPeXg7Q5B9rjrQxA+454BBZ4C5Zd3ibewGe2vXIQOfzu6/dWm5JaD2oJuk
kVko4WcM/YSab1intoYq+S3ZDkoH/DL7lZKfe75BOZLbWrFfH7U7RNnPWw9LmQAl
0VbzYgD8cYjEFo6v95NSr3yzfUeLjnGzvNXWkbmlfYuKxY5iMKSzy+D+8QkcfF60
98ZasVzk87NyEV61WxXzLrkRG6bkOiYzfFFf9Tfpmv/lZU2z5WIqjXvSu7+D1ZXP
UDHCFfqSQ2NcfqvyNWGikl5mXLn7+/PT/WSmc5bp5ocIUfaGDXwNjavEuP3brx4W
DX3fc1x4gt1S9nrb6OpfywRrOPMhxDGhg+Ro1YsW08+U6E2BqJb8C4WwW8XN5AgB
HSAh1jsQeik5eudD74pIUACN2v4cIMb82Htx7KFHf5lyZATfcvnidSV/fs3b9cLt
5DYQQ/q1MLnj4TRWKnnkqI3GTRV8Q4X3sHxorSyT9eGByt0W+rgkiPZ5BVudHDE5
rPpkwDA6txysKznuF/XUpld+q6/JIIgTVylthSc+k4eH7fngvt3k0YtO+gWhJOT2
AaifzYdPw/dBHTYwJ1Id2mSMlReKaZ4/F0F2/twg4jV0PkudyYY8rua28uRBzs3x
jciEIouD3MJ+JzUCyLZJo6iFeWiFADIJI+A1myw9Jmle18NLWOKR7B7fRRAGJ480
Dxsr+ozz539UCgCBqU6VyvnmR1Jm9C54i38HJuOZcc5H/GvhYCsRpAw7P866agi/
LHqL6Dt7zalfmUpl2705Fs/nkGBXYB0SYoSxR5yZMf6UdCL0kW9CcfOoZZAzq3OM
i+/AQoIjjKQ5JgrAlXsbR4oBTIs6oXCn5JfRSlmw9JwcruKAqhMhqEVhE0GC5t1o
EworHstjmmk7/lKx1WIApV/JLXByoserUIUWkvK3peBbQif1osca5E7xj7nxQHIY
t7XDfn1uftoco3mDnXRXqeTHvABagxNh6eJRoSxTLlBh9Qt3EwLVtqOdA3JPwl82
l+tBU5hbgqB+ltsRQCIN9/UhoRWH7em8T/O1Vj3U3oa0Iei89LQVuOxwTbpXBbJr
Q5RbO6qtetWeSakY8VFtXmKFXtkoe6WZoHUDkx77c3OZFe797phXeTvcr7/HWzmc
hn4SdjEUEhY1RbhskG08lzEab1F5Bfq+GJcRAbDe4E5vRIZKKIWFOWf4+R/hbQkz
nJYxHyiLqgoo9x1V7ZsEXwazgsoic9OV5mYYPraCm7RsvVJ8A2PE1ViFzrB1f6hN
8AZD5xmwz6sKdn5Q2E8nqiICzlL1j/LcnU+RIQqJtlmsMHzRDvh6FoZ32Ws2mPco
8fvun6pRMnLFJo+DXidN9z1m7WrVY41TMyhFWTzgqK0iImHgNSbFAkmEC4KMlmCi
F8TWmhdpMKWIOR4Pzm8DTw9+YtJmK0gF4vxMPy3DTs5ouFCHIbym+hLodPA1AaAh
eR5Rk6t7NpURR0SRaFo8SxlSsZxWgLrr2A8hT65tYt4zaZErJyoo4wBQ9PD6GJRD
cQsE4wIgHyjpZN/TG0aBJ+GeysidXsGoEtkdCeipNObUNXYq77ak7FxjInQ3pKDe
521ZF2DYcClz/rGsb3tz+beDUHs/KgQbqxx6m/Lrh+Eq2sJgTHsAfSqCTWUMPbSP
Zhrl0hieab36PlBz97iHePr9ZIfPzINd92plF8Zk2nnbs/878+0tHGBSFAeUZoCt
MSw+FSHAZzoP10wtOxKJJqZjM5GyE9Hv4ee93KN3F8AQxTFca3ZX3y/kRfvrguDu
9Jcc8mzKWGtpc2UNdvYDR6N6UnCiytqbKHAECqQUsBew6fFJi/ZA2BPy05BwdqoJ
cxtkznWfsbZY/Y4zkxDOZvZ105zhLbwQenLsVeo82N5fi0hwypT9953vSifX2TtJ
M0VXOm/963I8sCr2JGXa81QZEDaJJDr5Od97HevuHvgSFDVww+1WGxIuuFbZsh92
jW0BC1uMr66DG4HcT08c0YzsTIyKMt3v/2XoDxPhD0ji49ZLJ8DN5Db6axkP83tY
hPGboolEdA3m2Uwrtkcgf9v1ThzhAX/GJEnIInI/F/juxie/ZJ/KqrKPCb98CwpX
IQApa0hbkwqXbTC4C85RJiTXbMjdtSeYbaY6FKhJeAQS8Vn3ZOh32C5NObKkK3Qp
3Cl4xo6fzYA+bqo7+jkZt9RNxr5iKbQgUZbYuVycslNZNy2vL9SYycYs3jzxAYxA
F2tVE+ozmzgbY+P4ZqIxzoU55pNTv7f+Lu5xqxNF8VoVfDLOCddsh0N16N5rQjJ8
/VgnK9GTzCtJWB5g9oKGEZxCxq8LpjI2OpO3aIXLW0Se4GPdZyrIieoETDO5/F8J
48ZF2pcqwFJTtqB7I5BW4rz6+qMuVq1nkJjgIANX2/41rXxYa75eBZcSlshd6ZLU
SsdceGyCsIeEQX6QEW3wUSgmFd9+is+gX/PMZC+XSj+67gtZpdHghIdYjQvo5diu
e4ws/GQ8ikIX5rQbQdSJxwwfLxmqjsu9Ye1agXoEBbo5KAfct2DmX7Oly8XF7Twf
FhBkf7Sm80Tuh44yM83VsVN6I5buFpsYIhaz7pioepsXqmXq+X9hSKBkFHjwfYG+
bLE69dSwxoC0lvqfjdEii6rW8+MKKIp8wjgGlKFCCNZFEhB4D90NvwmQWoiRfJKw
KTyalW/2wdPmXIsrEOdGG4YY2ZAtDsPxCxfCwrAVNRzk82vtKiKYM33up5+1wNMH
vG1FE3X8C5g9vhiIkfyHQyXjl87WobyG2etYclERKg3IjBRyeVceP0rgV99wfC40
zRg61A2uSRcygkXyeVNRNIjvoz3Mvy5xjuNjNu36gMP2oGqy1NaIJUxsqZtJj4Q8
S0qQJIjMxUdsqeKEbLWpwyYXrBbBf0aTuUaL1LD3/5I9vp3yys0Gt/GiizeJn6u0
dVJfXEXc/SAZK03DjbgNIHH7G9cTuFZHCg683nIWZkWMs1/drbLtfZtoz+1LD1P0
pwv/Dcn7UbbDzVqtEi9V/0QhKGveLUD2PDqvZgmklwdJ6LaBuk4icPa6/B5Byf+9
tJbnNJxi32RQ6FHu6WXFoz99K/eXkeBaEonrz22X/YkuzvZR7/fSaXIaE36kemHk
RrWNvVnO/jKMlw9Lit0/NNSQb8ZB8oJCUSqKys0Epydimp0Pt1JYjobOlthVNaZI
sqFNyvSNPWQni0AcNmzM0G+gqTs2zZmJPB1HvPotCkf7mG7PvJpYiEQck5envbOI
YkW+I39LepwQsclFRtdnUmAz6eoU8P63TNVX4eTaE0u2ANGoJNk1F00Obzdcxch6
7f+f2mfqfXXXvpmo8RnODvKpTW6S8jo6ZyTC2c0zvF9LS/8aIyvVCDV0nft9ag97
BBYtmjMJHuBDaU8Dk7KEKeawkwYYW+53ycqzHO7lCfmldZ7lbSc4mz76GHr+QrYc
Z0CPK2//OBXB62iLM7Ncc9juR3KXiv0ytM6etG1a5to51Y5zv1C+zL0pQYTUrNi8
/srmFkf20FRea3HNr761YS157S9wV5uusPXV7FEPIQIw0tUvduTPYvPUMt0pSRJ5
R6JDNtvcMLre0TYzVGxvySfXy1aTrGVJckBLyX/2Ecz+Op/j+aqB6mlPtR/PhUuT
LBCRI+tUKkk1wiDIp8oBNeCNL9sSgNtgNcxpJQikT+GAMc27S8XQouqpA2t6UoNH
zcgG7KUa5mfQvBgmoNNnHKHWuXxk/0XqmsNhHgnHlAp47H4F0DKnTzrnoheMa4O9
9KDxhPqUi02Axym8XooFGwlXW4me4WOUA1MGvcTsPJW9CQMmAndei5xxhaFG0sgN
oT6NpZqoEXrryJm1MlClnzoMZ/+e3FffFQpz2e8OpZGnicaS9mf+9DXXO5tekg01
gxs2MG6FlBG07LRGSSqeKpAUeAmOX6PZAtyt5sfFXBXyItEga18Azh6FdRjfOtoG
s8oIsB1ZETX/o3obrgA9CvyJpFVKSq1HvBJSndOpGukZHvJIKIbNnHRghqIznDsV
aa0gZZ/85Us+6IujL8+N3wULdD49ZKNBWu761dULVzS6mVaOcqC2E8JteFMteNj7
RnmLb/hpb9ZhV6MNgC7qwFTg+h4wlYune8EKszFe5WuBY3TtXiFbQjtLYk2VyKR7
YB0BzdciHaqCtUcwgSiBUBMJ9TVHFXklr9HpHaalod8q1SSAqPh5VLTXKRVCqghb
A4/Fsvz1LEUSZDTslbaNoqlgLAkY+cacdWtvcY74mXicW9gh45J7DopETGOs/lbJ
VCVLqMVWnr2fmTKFSstQDB8UrMsD3b4IunBD37cKbhFuex6NrpDy3gbm5Gdo5hTn
xPVX6ElkBcllF4gamQqDpYTncobssr/LCbmxYuUpXPWyhF+X8EVorvLeecDWbXb2
isoyr1NZB+18a2BKwfPQo3NA5KJGkK7azZnsHYfX59ASsJ2CQ4lVTj9W1E+MQV/X
SiBA0CFlQhBvhFluG8i3a8gsdoLD2rKgUqUnIZxRfPATF8taG7mx1W1aWzYcwkMo
bS98Sp4BLCwDhJESKlOfgZYqRYkql5G0fWyBdGTx0ysB+RR76Di1v5/9YwELl/2n
nNou0JmXgJQZflc42lbVt/e+K31n95ej5ulCC/GJHxUKf1gRc6q6tzuVueebM6Ab
AE+8ER7EFfhWDscyJU2cAuKasmkHm3rwqU5HGLHYOCwB9nStAl3BWQxICR6RtnMZ
oMCGfFmjz3B9gOQef2UMxRhX66sQNPECJFl74kNc/S+jiWUQ5T1FzE9PvyG98yXt
CoTBLoqh/fBw1cl7mOH6VMdF4cVFE+18tuQpxNfeD7WBFE+t0NDJYkSwYM4v+Jt6
TvIOWLOhnOjv4JK9brBpmoUY1sXVnl/IgfRVWDYi9c7PoNWkz0V+fbnprIHZwjTB
TY/gX0DcfnB78QyC7h1Iw9KZ29cPTNczfr9+HS8kfy/fDatZtqDA1H7aIhfmE3Wv
08yBluF8sJmati0qMkCflZsEssiOH+imay8yHlaEMsE5zNrA7Bo8Yo0AldIwSh5F
Yf1ki3ZWbwsq7ziLsISUdjs/3WXuu4rT7+fYkXDkMGDhVYRI2mxW6NF6Vp5yeDTH
mja7ZrgRL2jt8rCGoajMsFnzpFeb7h4imSuMqDrRBV2UTa6G0QzEbBFvBrTIz32T
Y7cxu7x1oYvI2z/SIuUacSwtP+F3lAwFuJSBzPzlpIfWIV5Nvx7DqWMcNXoZb6K9
4+3pOwzOSqrOnjiztOGPfeLLTnuSqhhpgkoxvM5z0SXSjJDVEbsr798R0CLdCYz+
PLJ19tqGxPYJQwfg+80DhVTu2/IC/D28DipYkRd5ObckXhWP+p2IyX8O1YFZKfmx
GwcFqdBnI1UwFrV01DPdn8iKq1G5zjNAGH87HOKIJWfNTDC8dcDgk9U7Ohajpk5p
nuiXG63cHPZ7HAleb80Yc+whmrkib9vHh1QoyRWi7s9ZRxM0XwYrzSNirNaJpax/
ZMVui4eYy/PhvT8RHOsU2Nv5U0bhRlg1m3YXrLQ8OVyj9z8J8tNAGFVO0kAu75fc
KgBPxBk+2Q8Dtlzvu2WTEQadhBaEsfTJeGq0FoD1fW0vaymadFoGxgrA0NEbZdJ0
VtqoARV6rhZZHOGgpWdrWxoKsCyBJv+w8a63bXyvAw6diEJcGRf0hbbLmBF6qCyJ
vk19efUti+Vv7TX05BxrSOUxHQAlFn0IvZZbnoY6yIHlv2LF8rvNYkcRLUHj70Mc
MZ+P6tXlSr4g4voTd3z5oduR2awsV8XFBhEe5zjkohxBZD1/gYnQS/1j+pwlcPFI
ZKn8Zj7ZIDyHcvGpigjvFD9yyRQFZuZCB4lzRs8y+0pRrHPEUHj05CQrBvoCPCIZ
WEJz7Ev521u201LZoiA9lWVVUijBNC0rZGYTK3v7c6FIf89YPjAaBaivShHUF5NG
Zmcesi6evVzXpigEP9duptgKd2MI8dSX8MMzpqAxzF/jOQ63hWzRy3gkWqFtWwxN
tMGl8SF8xVsbwFPYibaOKRh1TiOnnJD15b++6ximoyi84uThYR1pAhX9usBFMfjf
PEcZGwHfdKtXQtnfw5Zi/R9kcdZtWuJanWGkIg/BqPhI09y/kHrXYxz2w3Okf+4a
Ml0aGot6wCsZ7hxjHk0Meygt+Z/fFct1oGOdpCLvJtNqZOSLtrF85wENOjOmb9q6
HLsqFdOvcUeClhhf713xch+GuGZOL4xDAdzOKA4YOp1DAeTCq/ufhwZq1V4Z5pbG
F376K4Gk3/9TxSBS9P53QujGXO5I351/NwrYjAt4A5//6+YnRjLOy6ZLwKWHfVWz
ui1ZFEh53XhTrM0zFvy0MLV731ciBm6kobBgUy91T1vLddJ4IiM8yAlBg+V5+LMp
ZO0/ToH4BzypEMGxEtSV8q2MKONDhZb0RgxVxrtbgYeHV/CrL5IsOizhMOFHNiXS
Nyjq0GhCGzrHQBcEryghdGWPxUzNZ93SdgSP8ZfMKdeRL/j3A4einnUKvNntv/Gz
VbSn1SOI/l23sGfyfEqGU3ZJci/zG0Uhbt10wYntQhFhK484MXruZdhhSTfLYnIi
KAw0wjUXMWmkbEr5mjGdxGc9HxQqBEtwv5njszP6baBfZmzmBVEp0DvJU9NaMuPw
BkTBEb9iwIJIT668mXSeyv/7KbOrFZThMci5+dwOZymqd8Vh/TEfZTgi/jzg1rM6
5FNGN9WGs9mrOOtsgEfwggQt8G3k4ILRbqdohuuiplF4c4qtCvc02o44HeWsJMHx
pAp+A4EUbF4pzQWTMld+cpD1KrNuuHQYEb5BIx+a3iX2hlCWdyfM01pXVspfkfSi
+U63VbrSBHLLaVxZ9Mqk1gyu0nsEVEpF8odeqgkBAjZkcKFS8PnSysueON12KOO5
VKe2YmfGN5X3ftQJMpiZbt597UOj66JklBMDbn3+wo9/faV0kcWENawJ9I1w50rF
x691A63UDS4v6q8JDl3XySB01P/nDeoiWjRRA/IjxIBv7uSSUsmJokLsqgp1GFbJ
LF2hb01zkw7peE5mHxOopV0AxZEzAvdMFwcOADXphWvGkY/9tRH8ERC1VYoVKMbD
MiY+C3WEspcTa2a4wsBd2ccSWEhCPxMVDQQ0Wlq75yVWbc8asmMhkMla0qgwosnd
duCEIBDsed7oCBhXd7pJNBB8nD7G9au7g4EKKEv5Gm8ntsp072frApvDCKhscpVT
4jTfc1qM0JB6wpgVbCSFnRSSRzQ9tARqan0mLlAUntw/6ZXEPlh7joM49Sm67MH7
OWmp4cJrTV86eBpusDddaN5xrhfPV/K7+iNCjIQfryq2UTuq5nUr328a9rIMTHdz
K7Llb4Bc+uX7UCV8nRChMLP2ryKgALcaL0sJMWmwJXFYm+tTJymT7C3g1VzdnhDJ
hh0KDLC6mMkuaMtNaB3U4ipSMk9Y2BZO7myPBBYs18IwMnfoy8wNWzSXz4UUU5Dy
bUDFbf+Lb5AjB9KYlUs2telYv+Qpvab1G58pcEO8+DWNeqgM286UFw7Kf6EUakqt
D4zD87FfMkOmSAf2fAMbWOnErjbev1VILxWYZyflaPDhaaDiaas8/oVSoMFHWibC
Ge4WyfTY2Zf5oTbBJ990YOyWvgQJPAXf0M7HYtgWxb0tNh4q8JMKZBCL1u1JsSON
wICHCXDsyixx9y/40uZ2OUwHp5s/0xAXBLf5VQNSofoc7ysrIF3y43iSwfaZvKfj
Ovk1//reshLLPKVR3znVQdbuaevLX6ODlecdLQ24KtrXz6uSwapbF0YEXnNhsPrO
UHl0PdYTN3z7GkuYL+QJQijJgx620eOeYX/Qaje2eTmAcE7SYyQvvUCY7i0AFzcw
YKrSJfyMfju0usmmrv5E3NXhDmijIGFCeAv4flritbWe23vCmN4YEf0YfJoy0LEE
JEYUlKdlSuoy9BrcXMdUtFveUDA0F1EvAZCDxe7+uHQp1PZDzpB76WUPN0rQPVGb
ChDvELsKVgd4aSm90DgyYygQuFQGC35cGNhfXp3ajGw/2f4z9ML/xongWj9lJnZA
RHcAYZhYo8BeXHSZgccNatz+rPFFq6WvqEqr+9XekL5vsVqQBmIo9mz9xRjjjRBW
W1AUnyHWQQYiWlhxHBlqFpUXEikxmLf5GcM+KYin5cya1R3tIZXb7J1Ll6zLMUyo
f8eWoPKqnpaMKwS5GjrBdPAdBp9/CgyBsJoZSib+vg14T9g0g001OrIGKnlERCx7
eirRIsnfLWlXP4y5HH8iHkJb9QB2gxP/d7/XrqwqJIn/paxkKECuTfwefGVk/Mzn
w0AQr+iupsmOiXvvHUPRD7NRudJt54IqiJ+MuHvgRmluMli/rTLYXlJoGVNxVlTc
uueWZHx+Z9OwvH4W7Lcco2suf7N59R7g5vLXzJ6JIFo90i0GHkms5+5fSGPzAtJC
sJBQyLCZdFDYvXvNMm+GyR4tFiMd2HaQG0vO+2UV+g/Ltey3Q8JGcIXtYbHoP2Rp
5YJMEx848SxCbslIEB0FM9eO8KONls9a2rl5yZIMwQmEJe+kazf5cRa9zNhN3bIO
fpddWBGbXfqx656tTu7O1q0YG5xJeJPpqFTqcaFbK1W7AGcyGvwtibUaIztDXDp5
MEX6fHxM4xRjm3AAONsW+kerkghyIdvvx7sHcASDecXcgCjLk6Br7Vl4jZsCMAoL
AZGnli8gGDPEwVt+9cO+Gt05lf0imXQs9SOatzTy+NLxL3XVU4uz2zkmrSzEDN+S
Zr4hMC3rh/cKE352yzI0dcQuRZZbJMQ5Q+skK2qfUNEFwuoJAxgMTBJqKzPbhB7M
k21JmsqfM9EGiwyKwLZQZpoQWyF5fWkoYR+bOy8J5fFsRVUfRdNCuQpwEuFnmKlI
qvBn/X764fD0b+shjfJx/eGF/5Gqp5+HPLF/xqwzuen6hTMyFs+ZK1SwxCWt/cfP
7EMCUspE8BCc4knczdQqCOoKul6La8u6qKXruoq66IP3vP3xywfXPJ+uz3062NHU
TlpNGc1xO/lQC4GAQ0/EWVD446fGXRTYROYSfA5HhPwCK3UuySYTpWTJliRK/864
Acm+k2rRywYcusUzbKIBUpYfKpU7Tc8SZGgPQP7UnLcrigfEeGdadPDdUQeE/3OY
biYSsqQAfrYP/J/4uPDCp7Z+6M9y8P6WP6ppRSLu0lN+2VBEYOB4ZA1vY6yWu2lF
oICn8m86Gb5hw7lzxUp111Bt7AjQ26FEZPCf8YxgPDas4njJG8pHcl0AotgLOKve
EVXRpUS64gEeos4qJj326K7gkhwHaux8BuivD5dFyfKD78nOfXnKKuodY2Y0v5pv
r61TegGnGQ+EjpqdxDv5a6kQ/PT8tVKyMGEISTqanjPBITLo7l/eWwvsh04OLFtf
557ecYTOK5C+UMRvimV0HwUD9FxFCiLQ/eOd8hCbwuZS0rlzQp5uY7Rq3a6SugzG
C9e3A9V5As/gFRGXBbPHmxIg7yDE2lg4dr7hYK1zwNekZ7c8HqzwD00DsTakhETt
XqdRI3NFZBF5s3cyzZ4apDmXCMzeIuf/62rzFuF95M2FDghsa7Fp9hikibPtp2CD
rK/2FCP19QiOobEydnM3HCNNv/LDLMS4qRBKzM+N0t4RK7S8Tspj5jsF3hce2gTp
vXjtwM+oDM6gtz2CgxMBARsYVoYCBgkwfL+72LGQi05ztsxdChLRXZim7Kss5Ml+
OPQNNCS+VBmvoLyHcRJ83wNWtn4viqoOCjH+A75qAp1/EXHquQ1Nc0jauN3zoiUz
DPdYkfpYcN9hvgHZhf9LEkHHsvxL2GlaWbDUYVoJ9kevwHI0wXJgA3FFaEkKEU4X
u5uM6NT5YuAJWWuWevZ57l44GkD7wl0xXw0AANf9CnacLjhsk7B+QI5v87nhS+k3
U894bAZjD9qIBGgz1JjuSwMTvnHSEvQITcchq+lB+IhGt+D8igOesSZCvLMEfcDB
7hpyWDomSsM2fElzMCIYk+CR3vPyEWI0hs4+8eOI9Ub2W8V+jQc+AmRGiEmpdUEb
CzGh2c5JU1as558+d6nmwXydpMoe1iEVbe/GUHkzvo4WcHldNapNF/Llhdl4ZJWG
ZwwEncurxWH44QaBy4+wnWilQkqWPyOkc+dIf4JsVBFJXxgemp1/VSnbJUXDHXhW
7KUybRIcrcBfB6tPdDHYkh8TWVwodBOeI9pKlIHzNzbgp6ng3V51dhZUqt/UvHFQ
J4d0Gg3ozIKa93CmwddnuKe+Ol3C0mV5HCmZ3/ScMJxOxdjsC0Fj9mcPXnvuCAgs
7xGHSWeOuhYXaNf0wPp+MyNWBqh8oc68s4XyIOd+t9CHbYELUqEVIxT9gHtTZd4L
YNdSz+4GuTVj/VJrL6Q+l3TeN6FktQsYfVXtdHcuY6zO2FSimyFGwA7GmDfyeGNu
s1RJhYX6TvWyowWfC0hbu2f3sryygAKK1TwotJ0bgFg4+h/XxlDVaNHwZfOKp25b
B29Mkw5TOb7hOG/JrpdiV9B2bJ6ZTPK53DU+lf9VRFbO8483AcJvJhdtrPNBZ3nq
Arvj4H6ip3XZeJLx1zEuIbkThKbTq4HG+6N5uWYhE57gixP13RUvWCwx1/Bjcay4
fW+TjrIdZJKDH4RAdNSUZ0V62SsqJEpsdiPBjfP2cKP1eWZOl8ZGbJjQqxw8SSPy
WpnOyZlc1mJWRb8mCbL7NSFc5G/bPXFB9emDNMuETQSCjaVyUKweJjUtW5ZgD3g0
DTAap9ftMtx9JtU/wGAUuBXmYwfnYQcVxR93grViGsyZ3KGXxNUMn7BCin1lCZWD
gET+RlGrLvSD3qUO2dmCBNVqjNYfiA7GLCkFSp14tcZGLQt1/ONj2RtbD1bD12IB
pOzKfC6HppyI3DScXNPA4jYLyar42fRJ9Xal4UXda39PDnKrJvNqjk0SWk/DS1YH
lc+2n8ZLUbuslfoNIwBU/FaJx0c4/EygZ8Z/GIrfI7Y=
`protect END_PROTECTED