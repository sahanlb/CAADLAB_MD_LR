-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
AiAUdO6w6BiDOjLTH223OBNQWUjeqin+XG2i+k+YuUVFbcne3JQlI2m/VcpNHN6g
3um2YKegddi4d4IYcUxXkG4ta95HWVtFNUTx3gHvm9eWVMaS4MSIzxkHnU+rmC7t
ifYNeFgfUN0xnjwxZXaj4JJjr76mV51eigvqqp0SQDU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5447)

`protect DATA_BLOCK
C4u8qxjRZ6RWOZ26oq19KIn2vfnvm1uQNKchrIjMA9euU4a+iEHHyhRGiEzcP8AW
DzGh5y9G+aq5WAF/Oha37xUOLjL+0IPWORQVEeKO/5WWqC7eRjsVKaip3JLcAVnQ
lixN1U2rBqM5io/PX0g5NslpN7YwRSbbhrFANi8Kxz/+GT7X6HE9vjxrL5sbXsi1
Lpi8bTH2/hopiFMX697h2en5hbcWf7dz+sTU0xxq3eHwt5Le/noA/Ox4DgdeXAls
yG4ESqJeJvKf8+oGEJXW9DimbFBiQjl/PqgiLfMEWBnoGz9mPVf6LxcdclImsLaW
DUzo+9MIuZsDHc6gOECykgGIOU5ZJfagGeAU/FzkVDpU/BBfhkGAVE/w9g/6jhLk
DFsPt7EYW88vzg3mCwVS0nNSTUvcdLJPjg9T6HInOP3H/TPPPHwylFEcZ4eNpbyd
3fuWKJ/Npgvn1x+YfZ1sncJ1kV2SKQlMBDTuLAy8IYlnIg018Ynm11Zbikta8h5s
ar3tExb7QL67WPSDBHelQquBlKDnSmEa/ydskSwn1YfOZAx2XyZZzp8whv/DeNeY
PeQDXiAN3SNiGrvKbvjNyUvS5DEFiQ3DdpfpLYkfn1eXAuNnpCHRy9XN+rtl2ciJ
73iu8S2gxLzBy4+lj/zO/K6o7/RydCjFAuly+QjPYGcdN7nYaupR3Nf4LRF1jNeJ
Kgyjo9NlIy8xRETaDK9f83wQHzO+JZDob3aloUHqBbrdgVNsDzDUSc4OJ4TgWfC7
AEEctAFksbPr/aji+BjYJcqgdRyflQ618woFdxmUyX0+/EnyS9Q7wq3D2zsuKbzp
8lVVXQq1cLmGF0IJvs1nq3dSUyfQr3FWs5ipw3Huj/nnJjMLFx+WEtHnnIhMaKzc
N4KltLsvO1ubNZRw1HkcDhBAOX2iwowtDa8I2+Q0s0nRChZ+idAsmvb97ZBsbmuM
JUrzIrPhx7V63HPqzg5ZpclNu9qubHCNQVxs0Iqx4IkL0WtPJ3O+6DSlhaL3a7ke
6jHL+cBjfCnLE+1Uw0QechMOomGXvAQpgb1wgM9h8PnvT5oGFc42nZabS5xWVZh7
z61WB4LQ9AthC7vMcCdYhbrBYvY9+WmlHyOToGxCzt2gGQegHsnYKb/ev1/n3UNp
s6y5K6O6Lqa1BWPOapDJUnTymDRaomXeIDgMZHp88jMX417H/z56MQZqE+F3Mvew
MpsfiFvhakjkC8okFipW50JQ8ZOL+7Syth06nEkiTmflPNmV7VxZ0PvjxCi2aU74
JSvK2szfZSRoSC9wm/1zQlJ3t4ViDHmKawb7/imv8UlsJqiS2G0JnQ5yXLVn4Rjy
piDNRvgiEq4/WfuW1mfCY3lIrMQed/rnACrgJtqFscu9Z5AK35nGcboutdqB+jqF
ckjsSHSGI5cSgRTVPcRTlCgWfFrkQE4G/SO0+ncnnNP7oyJ4OVa2UPWPqXDKPgJp
mNAPib/UHOFqp5SXTT5w0ug34B3eCfLncLvxS79gsnY4rLdwkG/LZL9RK0bavzii
JhyCZG3i8W5J5iFZWiFUQIrny4hrMeyvOEfOiERBFDybYYC7gPNe6CoMpdY53RYN
/dluuAFxSHrUux+ow7IinrbeR7owAfEtFTdGLmj/MgaF2zAIHesbzl8h4JPHlEtx
ZOMcCr+sFRCIyjMdSHgq1tjUkIR79nDsuGSZ1Er5JyzBRVrWcdSkYSYJ3eSIEbqw
TaUTSf5rB6KEBSkKHmnMOaUesoaPI3WznPsgog+Q9tzTutIO9o5VeHxHJjz8uefi
HBnqtlqQPqeofY7GvPzaZ/xWClcj+f3TIgYLuBFMP4e4gFPL2tWRAE8cB8vcpVkn
+kzlclkbW56gtLRqlHvv6EuF8Zs1wXqZ2Ceo8rXPM0zkA011g/Ji0z9lrNnMjW5J
ynvobki48pnpau+OU1ymsfWRuIWYOwqIbk/PeQrjJGagWUTDyYeGQr0ZFiC5EPqQ
avIkgEOyaLJqbYFquRGuwZvYHH+rjKeG/koTtyJdGYjxCOwMxWe9rGVTknSDtgaX
a1Hys5du/ataDw20Pv+rz5FPR9yG0NJ5YF5mmV2QZ+R/+H3ANiS3atBz6QCKioZS
FDmeYsyI9vdPL5+kEfk3u9XWaCWlYfiJfS7ezrPX2vwte6FoY7W+KNKC+O4WCeR4
QBZptXbRCmFVYnGuYzpMer6lymC5NyPn1cFfDW/ZAR0pyewCUC2h7/EnLYuOcWsQ
uhXn4ObejofpY4eRnu0M1IeDRRbnd4PEbmdCJjqp1Nq3dqzUJbdPy+NkMAD8bYdq
PdBqH5m2wxxZcLYj5SO4Yh9OWz0CjGo1XKgYVCHZ8ryNPXDp6j/mASl8VkfAiChg
AUCDW/iIgIS5AMMQ51dOH+Mc62n9nYY+bH1G10UJHxb1BY0f2rjKDCHhUT1AJ43f
rFbDxBsX47gH3NXUN5ihpm+Zv6WQhMh1PTPHFFw0GhA3wxSKupM8Hm4CYUrov6UL
8il67ItaV0KL/X67eoceVzmeMEIQTTMxTvLaSOcErJRmQ2EpRc4ukPjdnMjWFlar
p5XSS3cICkXDKIhhGFzCAE/JVVwgO9tJkpCEEh9ZFFYwIAohyQd7RhlqAq7wsgu4
/GgnwfUvxz2njPcPyaBkgZkLlOpPKkICaIfZ47sYZ0LQqQSjmrAyDu9Pi6N5AgJd
TYCTi0/UcaBFngNq16V441A7wYo8pIAA1ivRz/TMmJsn5cS+wnliN7cXorLKUY/T
L00RwRuIvxTRaV9uJEyjvP7u/0Zs6qpvkeRIUudnJK/oGas7+CbM+EsQD2qn62yi
s28oL046MoSimK3BxFAFX3lCt8wTmwGhiUOue7UQmqIDaEr/cWZFom/puR/xbZsl
ZUFj+IydxvOdaa+eNKP86oAIJabDfkLP1FBZcU+xBxiaEhnZ5F9ONnOmIqJSB1M5
6Zebbo5pDpLvZzoehim+4Fhk+RRqUqJkdRiOq3P06Du6hiRJnwc6SHlB5REByJF/
uPNA/NxJAksRxLAzySyUjC8YwAEd3DL7uAttGNfCs2GSVcrqVk9FbZpVg0Yb6cCt
jnskKZnV3v0u3LuyH9RnYIqsFYHwkj0Fbmq9sj9pqEXNtMJSIR5CrKw4fWelKV6G
nPfryrAy4xJW1THRyyPz+28iZfbcoNUiF647TKcT4iAh1BdeQi2F/1gzpHFrPNld
mKqugRAZIt0wpQR7D7JHPa2lG2kZyWUyhLtrgDOWTlX3GRLa044SKU9QH12C8y0w
UvqCnpbaqVYoiNXHKU4Fw7/EWzWueWQ622Gu4rJrHdGXMbwtdKTcVXt4YxVgunh4
+7/Z1np/3/2a6cKZc4xBkvCT6nUpcf8R2N0HdugPD+H0DlzqzuVy/Ywj7jR34FUs
ca6e4PjieEO45MRwZXp0zaRhCou3ES0vJMyeMiSry6qgLq6bDHBUP2j8VppPuqoP
3o3oHSj9Q1DOE4xJ6L2lki+ab2gufdVNqLzq89A2aTj+/woIP8AvkY6ud13ZwfWu
EOUovl60rDARdUoK4+/stSb58zMJ/ZPQ0byrlpbN3BO7H6oskr9QIsNlLMG2KKnO
f1weKMwWC2kF5DODw663LgGZjT3QLjDVT6VDf6jMC0LXuNOf/BV4atlK2yj76BnU
0btqTQiQvskKG1eePJoesCRMRH2JVZhHdNBaVk+iYPC/wX+BBbFiAwbkEi37Z+mu
zZ9MW64hDn6E4jsOS1TKWdC/oG/T7vWObUQ5wh90XDsijAuazH+nmAoV4w0s4tNo
J3FI6qnmHX0GbDwEePr+kolVhE0d/TDG3bG4T7QgKnZSH5uy4QEUfzDPQ/YRhdV0
Ach92MiVXPxucU9PqD2egKrfj5mJ3W9wV6XyHKMfUjwmxkVCTQdVhpDCoI6OE2Qe
ln9Xs5A2RzFMEHB7RtIO9GHLeaZGr4Iiva+Vwh+O0abx5uVRCU2Tps3d08iRvqrO
FJAzzFKJqUw1vEKCqYZx44fh0FhhRDhiUUE2ZHL5Kr2KzRFaDxvGsrXYqJYfYXla
5K9jkdyujIADcV/yOd9NTpi4LS0ejs4mAJqqXRmZqgFFY7qw6oYq37g+7C32c/V/
Tcm7FQ0y+K1IvyaFKlihI1sAa+uzryIi23VF6R1MgTFSid4+Y/77dYCaNniyZSKc
4LZaeX6YMvNHvEm2FSdqEHdIjf8cB5CFLA6A7cjF6CtBdRfF8MMHxnD6u8JHctJz
vaSMXb3nvJB+SuyDKqB3Au+dQOt9p9SJvotV3RRwgbyruf3iWLge1rLdRTJMKOiW
93TKleqbZ0XQtEbe24uPg4E5u+wkuEQrtOV9VijGWrBWqg1p9jRlMizM0uY+qlht
8BSK2TMhzb84m43Cew6JsWaHPjwux2t6q7XilODGisegi0itWillP//BLAAmR98A
NOzshAodIjdvPTguz4HTzFq/uYMpYyvxIfSve1COoz81v3bCJGgtjVi7NooPy8s5
ynyQ0inG34Q+1+dSE7zYpULoinKOvOoxQnPEVaELUIDG73/e/M4kBrLaxvZqLr7N
UJwy0GLgkeruVEX62tITjcS4Jux1Uxv3+BSpPyt5LAP1NUsECsVhHMk1zdMTxHnE
hf/zB/UjuEFKPqMZJXpDK/dAzjLfAVmYT9TOzZsX02KJlrPZdxT2GPzM449xmB1u
I3MFrf2slGKOq5SdFWV3QKbGHF1UzQchrafTOBq0IBj5eyuyu/q6W3TWFaAasRvu
2qE4I5d1a0nSe6ZwgdQQ4Bbe1qLhpB/AqudgU7R1VpbmL86xSW3eG74+EuH0zayI
Aq88ylUi1nTXtSUVnTIVCnAW4EcFsJ9RX/pm8SFeWShaW6GGw+n6/PHFHsL7k/Td
iM1++hV8OGGrZEAIexnLmQz4Q5mUo/v7T4wfTgXtz4hYMvD+aXsXXaHj3jAt/p/6
dwFMTndhByMttRZt7AbeLGysEuxvKasscFmPepYw7dnT8d73R7trEts3/UPiNTqQ
Q5cYs4I2T4DGKLIyYIfuz9e67TlgGAf3mXH+iVtqlfdpXPnQvv5HUGOu+wQCsqrW
KaIEBs9Y3ik71Yuu6d9e2Ht7fH3LGeEoj520LxzD4+P2f40CjIT7Lk/X7fZk2zmO
5o6wR3uOgOiNdW/HsfLdwbQ+U5q6LSfKdwHFxYOuYv7tA12cvcY4NBxHMyX5g+po
q1XIdsPjDYgeH+UyGtZ80bnRa0sJr46kUleUTNUrGdv3T8nWZLHJu5aIEthOzfA6
XcyfQFDg/3lE5yt/n8UjsYb/7ON+LgmjmRwBTHmb7WSyyFNhC2tgBZd00agp4ioz
36W+K8vWpdP3lAsyNirvloTIcGiEvZKoIC5QDheaQdwvXXX0/f9rFm18BPd9ZMfE
VyxMcl2XgKMHCvHfAHLtLdWU8tZ0q1JscofEvGJEiAnKG4SAB/qphawOGxYb0SqF
VGtN82jHbeHVuIjw8Sra3BKXZtkxGxrsspnMGGG8OzC7KQ3hrEF8KSqtf39vjgTU
5BJRUNmnbww6CDOzhaO7THF0xyplGJtr+RmBonMF0116LoWC2ktdmqrgdKQIw301
a93CIVNxrM+cxRg8XMXg3mdGiphZhl3bnpe0Z8aBEZuyQqOQ1HIpIrk9MhbypqMB
DBL1STRJR3rDtDRHt74NGmP29ZKfVdNDQ1buqzTliuo54glHkIj1juVuU60HA+GC
ZK+nud3yatqAnfQBotG17OuKQHECsvBmFPX6Cb6avwnQ1r9+q3payb2SbxPqjszz
IehEjElIqex/ap+/JKK1WQI3f8rOQTEeUbfTNp4JEaEQoITxwxT+fMbW4bTBwjtS
ut1xHSDXVKI8QKi3xUdqq/VVD0qnmbAc167M95LkCJCEziyek8er01zClYVTwoT4
PdPEjHaNZ4u3/p3wIR3JvcKY48r7eD+P7KbDYhqzm7eatqoqoK6Xv3+C6Wf3gqbI
6r1ku+D6+V21R5eI2o+V+l1qT/QfH82bY8JJzzGPtyGOXkyHG6V4VgKUc8bRzUUn
QUr/ZAeTUhhzrSmSu707ksXmL8W1WZyRWWmdjNwBrURKtC6KxI4BBcI8RNkdvMcZ
5X372v9lexFNfoB+WZCwaC40KP3xBpUS4OQq6t3jls0+m4l4jV5dwttEPzt9mhoU
Wmu+nMP+YGiRAf+a5NRoAP2YKrt7uaDfy6vQn68mHpZtbkFzgG0iY+he+TlHVfvp
UgpMqPpdBafDZ0SrZw50ZAawqFLz+qG+7JGfBIYoznEJ/OxvRujKFOhqToiu4czs
wpVwrvkEtig8vR99DoCmoWNCx0w2pd0/SGsSs4gfndLkmoe6uWxA/RadW7R1pMsJ
nu9M0kXni36v7MexJuFr85u91LAywzTPWP7iNnjuxMkiujdCu1ViDZquGHabEyKK
8a+z1MXkdRfTkdN6fU9vio8aSooh/pl+fy2xpXWLWEsjxztPg8+sKYQ5++wyZYxc
LsZ/fUxo1yblPX1BxcFDWeSGxlC8qdOTO4Ai8bz4gMnp0TdtNMTcTCk3ShAdrivq
ISuL4sI8rsCg/vQ/+Xj9Z4QVHnO9JqYujQwIDNRUacPO/ybQ2depdfrOvk86zv1G
PbktlSajIBJlOIkE6oSmLuhSr8YD05Mr4oDUPSaVmn4s7mt9Oa6HOu9WF8c8ydAM
enAHXra9cXkcFZqov0ACSbdkOgHph+fny8n+uvrlZdNmN0yT1waSUH77imawPdlP
ySz+9QupAbVgmtmsb0mmsUQp+6ql0O9R6NqbwEzTo15f/H9VS04zQc+Xq2mDGqxK
ozgHlD5J9C8IxC92mOBVdR5g3+TGHmU3KHQMFeN1opqZFkb1vnErI6iq3MSsEDij
RhqCfsskaXP5mxofwvjOxX24TiGTtGp11hyBSoR3qOwxQ8YQxB9V/9b9niIGwawV
SEDmJM32ml+jptgWKgASmCw4/VVvpfukSdNujlmEiS3ZMMDydu4koOq7iLT3NMqv
6PIAqzV4NxXyvIO3ypUN8FGZZZJzZLa7U9wBN6box2V9ejdtjekQXZe49zjjyHF1
iPIVDlEivedM60EJpFDBvyJD0cuSDmyzaHhgpLwdn/ffiinEWcthSUWyhJ5tMStz
9SnAe8/nKJM+IBjRAZBfDlNgKIdOMgLGu1G/PhZ7Y4Xd1WoiO65affKYCe3jCBrq
1AAYLslclvbZY9h9lOCOx8qDeoSe2qPZA7IbklBDHreaScnoeX2td2x3vZKrmqOo
QB9e3JBcZiIGikVY440p5HCcsrqG7lAMTYXmcLzyrJh/z+SxDQE9nL+uUC1e6J0U
`protect END_PROTECTED