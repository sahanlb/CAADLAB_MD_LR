-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
0vJSKQD1dFHW3A3+UD9YnaKA5wDhGOZwgdhUkHHE8Daofh2ga5ggVzQy+Zmb5zl3
Evt3HgTbeQ4DvTcff+AJW3e54KNUXr8eMqRaF4guB9LnBtAuXNurI8B3JZhNg6Xm
kMHuDa+D07Uc8fKdWemymA2XgXrvz98qPtJO+KCHRcI/Xf2N2oij+w==
--pragma protect end_key_block
--pragma protect digest_block
Q0vyHbXvKBSWywyT5Es846TJgBs=
--pragma protect end_digest_block
--pragma protect data_block
buk2Ssx0fV94Mpl+EfpTr8JC87HanWOB6BrYaDpRi8k3iOPWswyWImLGne+EgAG1
NLjDL5KBv/T5wiIA+qTrww7xMs8Alf2mRN5Zft1zbabz0lBpN9mYnU/7lLQ1nkZ7
NezVMxw2CxSGrRbBZJI4JXNH+xWJBqjORcsR0Jmp2nusahX0sA8zwcV0imzbHniX
Z/mDFM5dMPXUGnrDlamvS4unQPHuqG5tPWsXyefozV1RAfJUmLxVG2gD2+9p1OWc
N5IJxtH6SDlAsyjuHbnRvvP+VQuiQgsQ/vFBbyliTmrA2MDe4nCnZ2f3zxkJ2EzT
r6+PKRiSjSHN9DRRZcx9Bg5m4/J4gfiy8CQjJrXoMlpObWcZerXabYrELyRcoYZP
Bx3r58ynsUr9dpKgRMYc0BiuXIjki7iuTon8IkJNIBuovbzUs7ySCuUE3IsXTSFi
OI5LOjthLLyRK8Xabc/cDrHEzBwQQtKSaCHca0KvirHESj2dvjdqeR2164ZEs6XQ
NVaJyIAgB3hIQKYFBS7Y9irySFSSqMvWybXTNLEJq0LnxSO/eVGl9ualsAunipEU
Y7DAICoImfFVhsXmdIdGuuaHYp5oYK8bzyMOQry6yKcYyh4Uj4nmqvfCEkgB849C
xze7hv67HFKqFwikT+enl7iy57IVODZB5KfYulg5glIb3J0yXw0wmdqrRvoywG5O
K+4Z8NHsmUVAFTHBfYnHpOJr4b2WzrN+tv1brHQJ/Bc541gh53X0mJr1NdgPjj02
b2LbvbFJM61d0ka3QfK7NfcpvFHy5XsdMMcKnKDtBZg987fTFN8pjJJu43JZcd7e
OOxht7h+RGc/Ydpb2ijyibDncZQIcdrwV0t3OY2bveFFjWugs03cHfZWlckupwtz
pj09n3Q94aUM0te8ID9+JDB+JTMKLXCi06Oze6xJVPmPOf5cI3x0Zgki/WD4IY5i
YCW/Bx9Os9UpNfdifmU0ltJd/t1G1jZlyPL+HcNb5vHreR/hXax5tCScJV57ax38
yvOrs/0K9GwXicoImxEodD/RL2iNWo842z1mAbaauaYi3TPOW9Rj898fqxAVDTO6
UOl3aWkXXyWfGHs1P6C3sl28NnwaLO8DZ4KzKuOzZoPoeKY9zGo8/gu0kieALkeu
5CXRnQ7//Z8v5Zm79MNR1QDSDpbjP7R4a/p2LHMN39ProhQN/0GArah9mI0Hi8m/
feD7vZ/9/UKOieLeMmMyUhOutYUyTK1hM0gybOAnG7w0p9AHbkrsqOe4FOrX6Y+q
graW9Qtj/wPDZKyFAmw4CGSIUJk15RTZ0zT0yJg0xEYkm0uwiuW3bi/kcSsomCoS
2NG700gNtVGIVbSIsuKwtwZ49kXOewGVTQKbuJGqCS7ZpQfplvpWuIv8X7CAFgYE
TYcxlE0mFcUyWyLz0VnGWrVqoHDChTMWnD33Cfk5f+OxBecpD1XZ2sn4+Xexupnl
YCDIaFZpLT77FwxAIhxaoEN/l+MxVt7IZ7+uYZuvaqDn/hHL0YSf2ywteVhr7bQh
13rK1moNsh5UBp6STghizXkydiHHQlyxk9zUF8AaFXMFiCXT72IGUUi97rnVoxRw
fuqOhelN8z3m88gpISdEHYnnhVFFHukjF6I8PT6ZuSnpWi28VQio1zWItStw+B7v
L1FP7a1Ie3bqA7boOITzbmmXPeVlRAmtA8J3ARH9Z0iJSYVMGKOZDbZSvryumzxs
Kzp+5jm4N2auqWa7TZ0hCXsC7GUYHe14OEpL+9Fk5UGLkfd4TwoHMzNgm1UATrH+
6VBzAFyxBvLVNe/2tPVb1IbhlcslmZcnjFDHc3552yKpsNOtWrSSEaY5Ms6UkOeO
uNgnRyoa7YZZYOLbjGQ+gcj35Zubfqeo6Siwsfa6Vh6a8c6XhaK7e1Po3tFy5BcG
AhHd0urT68QT7PD7RE5JQlSHXVrANlnxXvrV42fRkXvHGbGNH7B+0hXGQTCelUXn
c2TVmzhrNYP+YPpH7mOnnSpeC/zWHYQpVJphzTGyPyFamSR37Ni/ZsqIW2FppIml
dCSzuS1uiLRmgza1blJnNRZaFgD4uHl99wGTl4ek38frBEpdLb9J+tdPHBcl+HcQ
wOKthOc8mQzrlNLWB7GRnEMPYX4PWSd3IykRDXWIMD0Ko0lKhSYUgjHQOT5Gl3Cw
Zd7QeEa3CuBfwSpjDUSbphcx/7GDipr5kig6q9QxnnjZkaI8Vktut3qDyIn2MsLK
ey3CvBzhjeTjQYjvGqL8euKfmeAQURSQUnkmPVm0mC3qeetsyOv9FwWS8XJfTH1r
rP851R8jicP+iO1Jx7Mst99vnbsTVjruzFC2W56hKTfYcqclKMTLXKqifolZubxb
oiDbAz6LyyRUqE6lcxrDP+scQGAfdDbyLixLUZ1id0R/af88sHw0ZvERFlUunj3u
/qzscwERWfeBw73/C+AVqtfsroY2oLZYxSZynx2oz5/+uZDyCLDyuXjK9Vy1s31b
v6yS0zMVuIxluR+dqHQb6SY6LlGkMqCTJMJQR3Hk4BJWSVGo9/TegTwYn/av1gGS
DCDtuoF8lL+8DacVKiapF4wgE0CYmTsJKLDRp8IxGN8NAdGnGnH3i93DW7bfQrwA
lQJQu3OAQvwRHZVlS32KrrDocXVbPv/fmZW1eTo/0PMOtfDRmrgqdwzanJmMvbE/
wC5jPyGMuBt1uplcfy3mTaFZrYmX4kG2TLjYDIfWdckV17V9Uhkxd280rzqMLhpG
pVMNS0D9bBlbAf97CS5qopwJpIgYwMjcivf2nGOsuzoAaThYXISa5t3vt2ti2lPB
blLA9GiWi9dRA+NOI+/0xsJoRnGFrNZMMdIHThTZxXfpHELkyiSz0gIbrS4DkaaB
Io8oS/zbHJKQ5g9n7F8Qg50HshxF//6i1gI3q/s3wDW6V2q1Fvqi33Pf1RicxtTe
c3D+NmY+2ICQ5Nxcnzr2SxDOEqxC6ALNcAD8gBLB4yoyMLYyxZEOuY3A3VwEd83r
10YMmgwkRPYRcsu3+awV6nljFDBYopiZasmakdDjs8hesWKvgBlqfTk8MpmGITiN
j2HolOOLDMzlTCPXuHjDvKv6nndFzAgC5H9tDJSpMJw2YMJSGHl2wDYtqcij1OnH
Gyweu6Ww9ATmfxzr5wGkUY55AATaVdXkTm0GMe6j34TGPYsk/E3ki2Z0nj5fkmbx
QLQBNo4b9i1akm9V4C3XrGJEbejvZhVEo93+3Iiu90HcIKmSGpEv7k5KzcB5ssvX
V44ia4iMJ4UngTyeClpAke5cKTeQDDju9xDgnQaujXW2VMBiCX64r6toFglZQh5+
26IWmWBpnOBmGt1mVDUBKryIMjVZatLfhAYHCmUTmUMZRmoHqI2lh4kGZEGLYTtl
gRh20YqCvl4z5xknPUZ/oH4i/5kAlslo+4dzFntb4Z53q1Pk/3ijwaJzb8TgxImh
Upd9L654R02Ur4OjF0rPjM171+JmCkpLw4D5euRgpyoTEBd0AhSYgRcklsEiNnxR
K0xhYVM7HIW90HY239AxEhmM7Vrlz2NB9NwvfaKO+CjJywTr6SGA5p6H5wWloGNR
E9lgEheshASPF9BdG4oS1TfpYLYA6+fP8RX6emFdKL5CG3cOnfzy3pM+AIShNesj
IfX9vN3dalpuxMLOCY4hsBZNxxuZjwKojH503HHZwCKwt4svqWviMIN2RbIQe9s3
6JOHX114SWF1O1U+OPTFJJLCXMX9MPYswDsXX8iCscVtbRZlTL9GdaGQSoVYs4cg
JC6R83LNY3vbSLvcMRK5iVwvHfefyOeqJ3Otewz/P4YRBgGXQJAj1pPmJo+lEiIw
sHHwq70kuCB/BEsLjQr5Yl5fzWownaJnzCZLQqUPozzjYvq04w7q71g0aYfhxiw0
sEGq671S7WsuaWBJIxSEV9Xs8d+q/0C1ZicJ6JYOxfQ9pzRX2yFVEcC7OsuR9tMk
cn8i2Z66rn68ANeYravQiJQcl4EKrUaG1FXy6Nf/n/J7z0noF9oBKgDskcHp85/O
u9AyfKERIIn7HD0L4mdsgV1gSxnQjwjbNhoTjZ3gPbRLmxUUTXD6c8WUSx/GfTes
eQwKLkT8NNpj7raiMPr9l/7YtPWv2r8Kl/b4t0ZRpFDuxwLWTfWYrXAz1hDVyHkR
RSpV+Kz2ylld5JlEyg+smTbeCA2+Rlh8sc8r7PORqpTJKB2Sg7HhzfppuhEjOhr3
LGqPCJgQRcfjEd424y5ax1x1wq3ll7mGGnwvzLymu6cGZhuQJ0amS8Ngzneghtt2
GekvNewTwrqRo7a676YYXEK3Co/DEqUbA46uUucaHyzOC1HyfEUsfzjUF8TywGdc
vUXyKUzq+CBaTGLyVrLYsURrh258xSteW8UfDLVs7BDkdH+vM4ArgBXd/32JRofn
kWnaJS5F2E+cREYmbniEhl2z0AsUHhYFSXKSalGoj63PeKdU9S6mRi124mw+IORP
1KLYH3d6r+tO7vwRV7z5M/8UUeVRkzV+iekp/g3P/EhJR7lfZ09BDBGYAg4pTCwB
71rftqEjj2GWJvg+z/aSp5ErC+OXkbACGQs/S8P8PftKWgVulS27ountDizZxeuv
lMwVpa0WxJSvQejS+NpJlEoAmEkbY/DHbjbKYGekxlaxEy9tjr9JDBEaQ5vORyr6
09Bmj6LWIzRd8o15G6Owj5tde2Prdh5BDzHxPonisXXGDvFkgoFecD4WBppPFkS5
s4J1xUcWhDPGZAG3RsdhZa52FW8ifPRuwilp16YrqMNQQRngS0vJux+AjINJLcCD
7l3g3DHJMYk96Drn6gOudftfYNnojxvL01EmZ2/RtsjdkKJAWcxS4WnOpsCZfyLH
dOCZPsolC1SXio+Qq9Js/cwWTXE+6P2/8o8i6rPl644fnTsagAr9emFtZqHfm5Kw
yRaXR6pVnvTwVgPkMluvKWDaUY758Am53IDNDoIoDUStILfqhcipcF0Gnd0S7xDo
BQrZ/qwZEa7w++QRabp4OfjoLmoseH2D/TI4i8LixWJdXvo/l59ZytAhn3p70YAQ
E7CHPXLDuFd3FUVwo+ETLXhCJv9l719JEg+wLRRroEhLhJmja6vM1UtdWC00MCBk
xtd4KeYz+bWj0B8WBUzuurIofN+a5AgOZfs+JYnO+iFBYSCPc0BgfV3XNVUNdShF
n0jHFNT6sUzOBE0vtx91g6EQEdyDnBEjfg3YB2pRYSJsU3VYHkhZHRk1NxKsdsmZ
jwtCt3KNi7Fy7WXgSfcc4yFDYbTLKzDBt50I4ApZ2NXXPNz5OqWow/cStDjDMkSA
40TI4oniguwsNuvcKivkXOQk/FvoaaypG20f6i2YibJHEbeqbHf5FEXRpRx/dsWL
vJWYvS7XzNWrcgjMK5zeOaLRr6hR+L5nUiu9kCwAtHopcFcNVeDBtRDDH3YiIBcj
ZdSACgY/K7SaoyB++FM/vBcKC1Cmp1bEYOX/TqZnHyPha/EiYzMVNBtiXqDBInVI
4YiBhsdPHoCNqBVNJSHiY+b4WcOYk52ar2oISy/qYVjPpc/xlXuCXFVQHmy4qyB0
ja8loxQjp3ialm8zwFkSvH3IBBVro2wJNHELLpPwIPkvON0fGG8/cNUvi5XGmcMW
XZ2nT4fFtmMqcGaL4pXteXcSTCx8A/F3F8/JkbaUk2y+tQzkRmvuzs6sup+81EXg
LUezQUAC0MOlkn0bVNX+uHpu96wNWPg2cE7KthD+TccbpM1+gxZiUGPeoyVXlxN0
07ybRd5AAwAaLQdPzutZ8TaMY4ru/iBFpRTKF6x8o8+q6fzM/ZyBDy987977AXWR
sirQLwGJD46rHp4xpD6b4wPFH4KuS9ceBbmZQpyfPNS/If4nW1IghoGEGbKPYFHp
kkpdo3V2B7lPgzVtaRAS4e1rTMHxq04G6n0FtIHqQ0dW3D5WhnUOBUZRU48gF1q3
3GLU4Bem2X4iB3edmodIPx3E7odRTWZVJcdPIzCVDcn0aHJrjbTE/Hxm26h1HKYN
7PfWhwRvrI2xR0ag/2888PhP7ISC2vw2hB3O/oCdwJywds+SmXQROw/ITRASrrXh
OpqOljSjiYes5p8FlfgrbxzSNfqszUA/thBXKFdBwvnovEjK+FMdCF5oVXkdIbJZ
3HqAl6EzWzL8qFMCR2TWIwrszz7V4DJnJAJ7JWq2KpEN+osJh4kcg+TDTlpLUCxu
4iGe/l1buBqRldiDQrGqVewjmU3hQJ+gyxavofjWfJ35knE6lt6hn4IamqEs2lYj
uuFARyyBqFgONp9NuYJgAQtPXgpSPBTnviSo1Sf/xYYZT2J000SFzmV3+fYP4YAw
nS+YFBbgh+pBFwgGcaq+iffv7vn1ZlzZDekMQQ+U6vi9bA9E2pM3aYTNHHacfY8Z
XeSBf0ZqnNT1mj8Gr841wuOezgId1NMBqrxhfLxzyZi3BRC54jmNVd/CI0J6zPx3
4pgzAw6hScOvkqnqrBNMDvgJXfYYvrBYJbarVyK3ZsmB2tdXOAyk08OA8ZrfekE8
2SxvnAVpSkEtH8t3/IVYes7MTwyZZ1XfRUh5n5YUJ9xjyQPL5OQN5+nGDyewNH1p
bO4N28vwhlL+F4G2I4IpxA4XOCP1GBfktVQuQMlZMuf11r4wV9yIhPNksFLAOUUt
+sSBDcvsY2LGvYdolo7jfwVKuc0tv34c++jf4UnPzg6nig10LZLGOkZNgCEwCagu
Qsi5gmvQA+dTNYVQ/z9vAlJK1jJivvr9bu2Q90HbbBOGDBZ3AAuoHPvosCD/VyBr
eXdt17Yl1HyozAwId8SnNxgSlFh3700Nf99uME7k5PsoXK5CcO+6Dvl9x6cJIdyu
lEz6xnJTTgh/mQzUxOp/nZmdZM1GVayR0e60WDHvCzfz1VqNI6/x2iFG2o3aD1h6
pe1iPCvPSxO2ctJzmjVy9VceB/BPN2nh/S1VXc6FhFpJSglHOBr28xkUEjlUCbgZ
aNxUynRObXTXh0zV3XFJqT05t11gen1wV0sOVjvAeMMsJvq1JLaLBRhHMIV7KbFx
Yc5V+36v25FQrP6BpL7J2os+KbS4dVk0Lu+v6NvOZe4XojN+M4+4JHhIWn0BAcO5
1cYQA4E4AIk/nIAcrcSnv1FwSLirZIOJqjSjzH1LwUcKfGn5xMuH9LGFMdNVeC5m
bEcbc2PA0RlxcF+VvsdWaTrTWZCnY4nEupMLZNc/mqN3MP9wZcbVKCjyK7KC27dH
iNFfvmky2hp3hMg8G1N4PSsfBhuxdxwFWo+6jUTMi1kJEt+wgfI+a95yX45J5Lg+
pxqFxHEusmzfhWSi+PEqNAaWt0HHTYFyVB3gRqCrSyoebkcBAwkF7BsT21V7coqn
aMasAoscw/W/uLqoW7l88+Am8qDwNtnL751lJt9oFadVPGdJ6XVkd8OJcUIouANC
TBVRFW8BKQW3i/Ri5vzFCZ6cgdFPj7dl7i444JoJ7IHRAQ+33VnRNaUTnAGOQmUN
kxgRy2vIZHCTyIDu1cGfKy0X+bzMLtH2BAmOSfkp2YKzE1gOhbEGdphUXDCXcSXy
UIZ1Ae/M7Ozr3mMO1/2Vm1xtyADDHWQHM84rvJq4FV7nZDAJk2+MEnnvjHVkyqwT
hEyWzN6cee8snsOVglmACfSU5CE9aZK2cqDwAZgk4oS2ai1RBHdqfcsivdzrri3v
ocAYXkmWc5EhOU+brT/pMRonVxXxjf8p3DdXesCdRGZ5rKzT8CJvrQCw5JblsQRP
4+WJm7z6vcDqRR9l4GZWSyeUgFNhNV5Rmx41wt0dNkZkIg8Ql09uMSgEOvT0ftTi
PlSwGsmPbn44HobAq2ZUYqCeDbiA0Ki3kUxQkmCobAkgMJYybWIxl3KQBNLt/A9H
fyL48PaBOn8g7/4vxP8Jreu11bIuJNcZz2cJo7fjws7iigSvcBv9oKptzzBHrtUo
osH1PMQ9wGt22q5HVzmByDzB1SI4SUAlIO9jZHSNa/kutZlBsrAZmNJ3pQutuche
cGPaHUkfgcG4/Nc+0Xzp8D2OUyczzwn+HN+iA6WdavlAoJuicgkWNdwryYcjHPlk
BQ+AJiA22b77ptmz9vJSptMn8Yu8qEQHGM7RR6aFfAqkd/uRbmG3mHlAKAmNN/WR
S47aILCSjMiSeqfQmLrCcdbwV1I7NGYJPULGjihkT8FKxNd0kv/wvq2q794ain4B
ardmyUW2nuptxJzSeYzO6zvuvyw3G15j/gC/9b0+wd+OydPpdYvItFmVVwgSt8PN
f19h6CMSRDYdRn0sGA9kNZgJnXWL0AQZSbcgF8V3gsh6040fAYiq7HVyohLZG+P5
R1zZxVRvwkpkF2DsIB++074NV/USAyYf3MPAPahA8t6eZn+GoCWaJzrWb9q3Aqu9
1dxLofrmTu32rYThFxuUIU5TEm/d3+ZCpa79NdHWYK8dHGbjz3XLbKouGvfnFkiK
/PeObp1AAOUoo8UIC1XApvUw1y1Jkak5BIG4E0Ebed+wWH6MxXxB7G4tSsXyvLsH
Lkan5VUzArPfum9iHzluSFu4lrXpbBZ4zLp30rDmzu3zSrUFJO1lpRSO+5fDK1bf
vTN2shlYDlWbiP+ElcFqM5FGm/9bIzeu2mN8B1uQbrmx6CfLeFcmhrFErgp1FpnI
2kqKWwiH4ihr0pBRxo7PhCcrbvIcv1GAG+v7c85eSPcAll11jhod8gzIRCFd9Lic
a/xAi9+WMfZfpka6N/smS3cAl5FaGnn2tSMAWy3zbsTQU0RunAa63hW4xubVwDfF
pnj6S/aMiIBQQk8cO2EO8QNLsnvWzzkBAqHFAmTjtksodeagTvhDCduEc9z2W3IH
5sE+6WdhqOxjBZC35dBWFzaBFxVY4QNw6C9eEcCXWyn6CJNdImggJw47CoJYZQlJ
FgXya5XR+egNwZkhL3SMoJKCtmJ0ygIJpQgmAl3GFNnXYGhA6wsWvFtqhPSTZaVI
z2DDkxvMFsT6RWXhFTH0DY9h8KlRLUgI6GeMXHVl2/w8bTerd1uaIPU0A4qnUd+q
/2aVElW+U9e2oiJTPIsiQNIlswpKLyEmKJuJ2MDqqbhUFT+nM1ZI1NDdFfPINcW0
rQMsFMYuoFuEcXtLCMQpAVVeTPGFMfVkI9ARQp86cIkrq8TLdbwssWVW9itxmA6E
0br1DonB6IQiG71cV8L4BECEbVoa+Vx4mFtcrkW0Za6QyQ5OQqNh0CVgj/F8kjmD
l0oAUzWTegwtbG7+Utm94WZY2q6ult4X4xIHZGhuXUYePpnKeAXzdHr7Wviq2Uda
mnz3wBgrW9CZp6QqaRzjYINsuFh3GNEcJdEJIlwh3pwxYOiVYvfhG7E47SCUmDLh
JGsMWYcoGugMMaql575jMiR6aEZscwMntjnS+zmtx3PmX1faUufyf12JBQMq5G62
S3DFJSYkd16Itc15x3UO3Jof98RL/PgdAiWd7z/2aVERJCyxERt7y1AKGUPB0yGY
gEmJYfrOuMo9CRA0TIhOGWJYIwM8eKuAxDyarQRqYdrhTWURpUeQsijOj8KZ8SYL
X2IvQvrKvxdPvPu/VCqhEfrB4HAh9XraOdXBu9p6fOuIVnzsIwB3eJUYAFWdeHcb
tTDfuo24/cTtS4CRQAKHs56vORvuSDiBUL3wcFVpQwR4w19MqVEb7Evq6+EMbeyA
IvUbfFOFwibkLRiR/iP3mO+bP1hwuXyHXx4bkMNRNT24+SV9ambZCKu2A9nAtopq
r7/SzfcKrtnGMRVtydnLlb/MNFKlkEdJWni5VWzPWTEA2Sq1l+vmL2ILx/8rW2AE
SVsGMjy7XmOLuBdcS9heIyZNyLXlF/FCIoIFYVWZ3SVvfba0A3AXKPXmvUouEYT8
gO8Om3mTB5YqoKz0aGA5BRoCwZEaEtMwaxl0SpVB5mA+dgXlacd8TXP4CIsFI/tT
NmQaY42rIEVzAXqaCp5G5/ya5pIP31Odp4BzGq/FH1xVJcgh+V0G6HOhfsuOv3F5
82PT9l+gxe8+J5p/EG/BzNHEZVULEpPolIVwX5NLsgmOTFqKQyOcYHLM1sRpjHu/
jVbdz0rqCxTFY/BTKQV5prUgmC1m5RcaeMSxTOVWx6RMEeONUSJh4g/uVsrAF3BA
cyBQJ6dBMAdLDblYOtO21tMG1QVBHcLv/wFMKDZWZezYA8f+o7L/0o4CWSC3n+HS
MildZmVR6AH7rCGk2d/zC22VzDxGazQB2QQXpQueZVQbhEVqkN9xuwUQU1kljlX+
pxhV3+8ltAlY6p8K8ylNmvy6IlMe9WWZrgLfzgz1X/+vkFRrWzmpP6RdosxgPRLS
A6gV5CZ0mdHtfPypJIo/nw4r1vetMs8x1O2rMEo2xqs05Z7Oax3aNnkNb02/S6IE
ucs0on/IzVBosHbJB7zZXbn99eSPa4+2qOOYevHCEdIVA9wVleDaFg6u3Nk98tIx
JQMyFeqjzlFePzlHYhi9zs4Fic3i+dVo8Ns6AHyXX6uyVQPtUc7WPyOGz6aiN+Xq
UILKOqHJnq+uOMmVJcT4rehxeLOpvDRmVX//AFWI19jmQJSjoJ9ehjaGgtVvTIcO
4dzX2sJJAdc6Asxo4FQO6CUd3VNB2rNqoYcxsYFKe5r3Oml0/9ShXqWaJ0YgYU+r
BdNVexhUkouPN3k1CUBeaJ10xOH6GKMLkAJg/J/xV79N8rdlfXxUXdLv/gImFxEN
u+31xINhIeGdkrx8bI4UxQw234poV92OpyJo5XY/Jp3IpGwATJVyFcSPWnJqySFF
VaM4Nqs8LFP4CMiAUHWjrtPGnsU9eLJTNQ1qs6qUZND3OOda2ZznG5eIUqpqthsG
a0FLXuKSpxyt+c1rrRyXvNGS175VKcbjosKBcYQzjggLHEiYf8eHmK+pT2bmP/G8
2pwMdUjO0n1ZvSQZo2puHLeNf0jr9Xh4bSRglFxJ+hVOTXkqXuJ60zBtDe3oQvCy
ZqioEQAnSdrnmBbt4wwa3s2VQrxA1tsNJxu+FyKbcK2K7uBtB5GGVD5Pova7JaYi
1AYnNfaifnNksQ7+jr8la6u84TBwyZUQMVs9Dfb34N2VfZc4pVYKHwUevqoUAXip
VUepQqHsr3uQGOYc1CHUdXhxUyqG3T4EVFKUBlbWoAF9WhV8oz7OPy/hs/q2HFB8
q1F/7YrigTz4M8Vjb8h71eGXb9xEHGMuMGAYZEJJrdeKZe04tMOFF9QdcY92zQau
alYkEWm2iOQLp1wa8cPJ0UlXXpLtkKDqTAKQFKPhRxEgteO4gfaKbXl50j2fwB82
F+mKOS3E6B5Mw+9DZonRbNflW1Ja0XsIFfu+9rsfTZ5eGfFq9/+FXFrm91Lpafjo
75HCyzJT0QkVujx0cOXVkm/ir30p39kP7sZnKjUm0hRQSTw2tEed3N/cY9hK7sXL
xWVo5rKJ2JT6vFd+YiNxWIeocLREL+LFTdRmkq/qauVREkQai8X+30zuDOoP6Rqi
MW5zLdqtPYnaJS5nv24c9MNUUUewW36nFN0hzVu5aJEiDi8BQynWqGXvLmQMrpt+
E9UrXhy1pCTjoEnyx2k0cN+fZ3gE3nBKQuNvJt+mgQHLXuuyCsu0bNp4Tqq9Sh64
icHh8XKiehePHAGM2IGKEF2W+ZgDVGaMPain3XoEmR5Cu0HypKezwPwuSxXDT9+W
SXMlFkfNR/YYh6mQA+MG+czAHSPBgPIKfHgAd8pRwdtQjstVV3ub3HBLlqtfJZ6b
eSUbCMOaANPvLxNMJWGLqxnOeEhsfZ46PHHmzy7xUpK58FZ1RPJ/jzELCQypGuKM
aNSgrzyrXz86NCRG57Vie22ZBw4gheTyP1i0i9A3mMPOO3WYslEUIAz0ZjHgXf6r
eG9K6fjtDBidH97NfzCuZZ/PjJq+eLnc+RFBs/5Ixt4+/hu9Kia0/RYP8pQ9I95L
XC8kP6/6pnjxwWkXGKOGdI9m2ZSwKZNP/1Ol2GVNv5UwW2gawlGOwq4u9Rz4JesY
GO9U08PaeaXc9UktviTNWnXTlGqzCYZS/P49cAGF9X0XOND0GbpO/jHeq5pb5+SW
e8TTZuzcMEaAY1bqzErFxaTjywuxdi6u9agRmpjJ+sV7hdmPWAMlX8RM0J180NXX
JDlqL6oZ4sR5CSrZHd0bIVAvW3xsmojaZq+CNYQpPE8PavK5Gdsai0i02FQYycdb
rsfJ0d4Wm7qYrcmJVwygwQPhWhK+4TXopc5dFABcYmj5Ll3AZ5n0LYFWd3TvVYUk
vAyfLiBvePkOUjaCdJHeqYUtfOYtvRe4HcwkCJDdhCKNN7tOVCXUs22aMWCY4azt
Aah99PHMWU6I97J11H+dkQj/FOPHepgQcEsW/vTxKou9DCUeN+7vcxm/IPulpjcf
j5movNXSJAqz6NWWZx9b4Edn/cyogeGlAi+6DDJ0JDqoaclZrO1iCPu+DtxdwUhK
QgBIXLp1A1KRPyp4HANVHaT9rDdrH7a+1LnJo646VW+HRfTqMqA2Npwg4K1TN1NF
Waz3DGDLbCzyy0bWeZ40I7l1nYJhKn3rJ66Libvv4ETntaV6xGOyFFf7oGjn7ioh
4cCI1c7zOhDoIyco/6cRV/Vl+/ATWGE7dz20NnIrnw2oJn/kymXLTROWoVY8Clgo
rF3dvZaoEpVFQ4x7ddmOgSRU1Ckqf6FdyT/C8UQhkVZ4KHJws0pYFLr0u83FzcCI
9OaThSLV2r742Y7jciM+Te746E/u8UcmxQ6bYhNyXEGr/1O4DRHa2OfRzS6EoyWA
9/HbYYUWEw/FwGHXB64urkA6YfCaAb96AxjINCqu621MXWq6NFcvEFCX4o4Jol/h
IQaWHpBfX0IddUz8anCUAhZVED2pG0cjpgrflE0Wy3ytCYavr68IUf8Vo9cFmEsh
oVOsB3JQIpEz0uuVo2B0t6bu4H3gQnAsLZsCUKqH1eaq2BkawbOakmYp2kl198E+
YrXq1f9ey30bVnB8FxFJbgaJQgX8v/jmpYFhNu/sy5KGlE4sGXwrSGobJnB5Y+jU
n6Mgpfx++RFbqJWNjuNzylGg1unM3vpP1WBkUbLSp4naoayx5x17JvRJnkFVoezc
LSNfa8dA3EGp7nE14WKQMidAs719fv7dvvLkAv9CEDFU3LYNcheOg7c5BjimaBH0
1zLl6baqamhgWTY5ZVIRIZyVKj+tbB94VhWOXdBlo+wGy7v0omP1KXHSXLe1KlNV
7DOOVuZhLxu+UgOMO2DtsvpNgjZlHL2Bp8rBAxKRXeLbqX6iKkdbw3W8QMZDus9Y
qoOtk9q8xP6g3Ztv1nlVNVjdHHj34Gbf6acnQDGz2GJXdqlc8NOJWgO7nURoVSET
Bt2C5pHwnWRt1lobspNsncZnKg3IwFaN2sMMkR5d8S3jfDZNR38EnaZHedJmzviZ
osrKw57Ka9WQZuiO7j6plCHSjVFLwelxj8FEj5pevMtN4LDU4e726h7vWFMtKu37
9iQMs7u00brxAC2ds0LtT3IZBatZqJ2YoDP6RBLfD1x2oNPKgo3UmMhGrOE6gijA
6HftSAIfWE+tbPPgBxaTLjejyerf8pjO35WAHbe3Fqd0U/2HySWJTuGf4owg1K0j
oYyQQv/20FkzaUA6hxl5JHKnDH1VVvWzm3GpdnOrQ00l3Ore6TYvM1okTXaAnc51
M8AHG55let04b8uBmUTNRSiu5YtmjopFxysTS+jRnDGMPGNuu3bK+PEPwV0icVS8
uQyf6C46Rn2lYxsVv39Mee6cZGrMdWEb8PUtysBvPkz2bsBostAf+nOiii/eXfNM
SOtODUZcDgF84RxMq1ISajzlAzJTzbU3wtZkDVqZw6UOzH5yclx/9kaZ2WU7wDiA
5SYrhOHox6ElR1M8rsi1pQi8guXcEQJ6WQKUi0gRTMiPXdXN6B5+7J4UoiIM5C/C
KAG+AEQv6lEhbw0BYy+lAu40r9X7qUq4eOIrs9CBxpMtjAzZPr0R0I9DSJI0nSDi
I0FQEGXB0J9zQOxNajq+1vpIdYr7AzhzsPGb9ICWj7/xDiyAOTlxOTBPU27x1OYN
Tl0noaYhI8ncqIQwgsJHlQr0xfKlTP0Kl3y09DF/nGTiODv3inS6D035+qF/iPfL
yE6DMtND40fWc2JnSKBFjvy1P+k7fx9Xx0YmjhFUXIDCcK1lrWG+cDXdgy5CCI8g
ztFmSY4+7VeI+EHsIJTo6A4kfK8hgSm56Y4J3sxFzILSgrHWX0zonLn3EVVddgKX
MwA7SHiEx7QzsbXJ8IKRberGn1uJEeYsrE6cny7KhD6S59adWbODq/H9ECLNvCMH
WymprMPRG9jfA5lNapztSWqo9qQUP3oIGQ4aIH+CjQ3Gz978vt6JFcd2QG4bZVS6
7CUDUk7eVfnLyhQDOkiWLV0xOETau3AlP38ftQFZYoeCSGMLZi5zJhqfh2cPk1+o
z+Qyn+Cyq7dnPZq+UGDrp9HL1g6LKnBoBudEo8DKYjeo6gSabqalE9qzjPAbPtXi
gyquNW+28G3P9S6ZhaAV7eg6qMACsFOC5N+efVIB13ModCWz7uHGmKZcXA6NZySl
6DN/ntvPIfFnOw48IEwLanuaVPqKSGVQ4wEwG07wtEdda8XwQyPaWmV8WsrbJxQh
uvom4QjQWEgK7k/tnjiHcgx85Un5uid7Q8CMY6IV2sJex+rHyVjHZub+XPDeT69k
Kw5/kTCNC7Bsy2i/vBylDqpRbdNyusyBkXNaztme/2NKLnD1xgj2lYEdZvrZzzxG
QY72Qgyq3R15Q5UVXdDDOVNZVdOD+adnbFKtjGhm89e154497IVomM9UXlmbwPyO
oapOCNgEgM99dSW/avqNM/PqXZlzgUrGPl4VWn3pHqG0hKIfuOnWs/USnhUOAHtf
Os+qdWdTceGPYlg4PurwvAATTSBtozIwlpMiTfhy843RDI/RTSwbOX6oC6MYG5eO
TgocwcP9UYjVTNq7vXPhjad9Yaj9hIAYDtiy6Y1J2PjDzxetcyOk+PXbZD+Ez12X
pVzm4KCFWVo7LNXyf3vKL8Cv9K4odrhonBczuGPw3yNCaHVvnRDveIDmcnSjAqhF
1jSLeVXFsI/QoKh5cXdVJ23+ZJ4ilNE8C5A9cDzZ/NX2gV0GUxC7L9uce9BFCISD
bOrdyxsVfepETqAhcqTmqOph8qZRTfQKutU8Xs7wbMt+UGSoDBU0lddROitiaQBb
XBQrUgFoyOcH+VgGoUmzbFjUIGouKBZ01NqldHnFlSQvpWIvDy24f8plnsMPQEew
Dl5OWjlil3eQmRJjfephCBRdA/7jLCd0fuOeVi/OPB9SQuZTnBzgWo1lTnBTLpsE
MTyaxFdf8TIsiKJDJWVvG92dcPqRy0EhUVrn7t749yQzzqo88tMMj64bFNpmzNxo
TO3BpE5EoxeLuzfdXHbtUdC1cSEmfkgbYFH05ZnW1+emLCtMnIpC3YhT6t8AHMcf
gp7gsErSvujsnUPrIJjpmUJ1eo0uVlf/bxMU7BZMhHPs3YYdrjoPi+bQvkewNU3c
sem1oWeOyA0vYyB+iDHDt9e694wmSAdhRAJ15alc3pha4N0c46NA8oq1VdTDS6cA
ilMWiNMPtYaFBr9upEMcUyLEaEMpTmoogS4kdtB1GcBaEZHj+ER0LbkLfdRrDZQ7
dCJSYR+zEuePxIPIkb5DX/hbDVjoyJnSgTI1JIjw8b7+JYsHw3oDEBOTa1VfJa+p
swU4iciKBmUVH6sRIVRsgtMttKSPiUPFvg9QM5tuhL/P8wJAK5HN3sMaoghy0YVD
DYEa0WyU7ngY2bp9uPDVrG0zKmqkXmNgGg/LN5Q6/V9my22vkuKPc7hdN649p22R
RtPOtDLaJz+x0gTpmVnstrtTGIjs2YqmytDaYb3y4DPjLwz6ygTtNh6VHsCfii5s
yRZoPBCnapVg1Op15NAK9s1sci/kaqBIN0Sr9j2Z8a+3+iLuLEPU4rCPraXWgxYd
Q6Hi2FjtPe+rzZLSwPelMwIrNINBx3nMuKCIYo55AGzCSOjMZu/cZEXLpj6FRhXs
pmHH3R44Cd2EFjyBG0G7Kv6uJE4B67Enmdj4U2KH0Mp/qb/HHJ406oDDr2LbvlBI
6VpQZceIwUHU7YREntNGbG+JJMpDVk2QZxCQgUnOxfyRta/kH7tt1DUMyod6MIBR
Dj0AEYY64ScZ3AWvgejb0ie+jDJEjLPv6SmyMAORzxQD3l/8LLuoWCBwot+4G8H2
v/1dmlpDgVZ4dPmoxucr92ailF2qRBC21QVhei2jF6nOxh/57InvlQMq3cl1R8iw
XoL5PrlmN8ZvXQa0+kvfWRwbxbvgjXkQRj0LWdYfM/LF1Q5iTl7lK2b0clOLaWTX
DFWOKgiG5RhczfaI0qaeqokz5DUrcLDSyAO5ZWPsiTo52k5BQcKpE5EKA5iKP3Y6
de3Y6zPR7lHccBYt601yF+9YNHvbTvZuYZq9vyuVYsZLOLg8C2H6FOAEfgEcZtqu
RMRNGbjLswM8gNm9HOxC2lyHjhjyNymMRJYS04g9zMrCGQSFW0Pu2uavDXQ9Bt67
CA1COXK56RAFRb60J9uhGvYWKGJxCb1U9svkTPSb7/HZfvG/0XkV9TBblcFb1959
p8e9U5LeXLNEkLZF2+krZUdi1YscDUOlTsKYdzhOT1/3+wzTV26aoQ7YXeKzWXIg
AcwZ990wFz0fnI+xQQnkaK7ZQWxNw3eduNDuh6nYvUaixwim5AUaJvFjEotO2Y0Q
Ccmx5FYvm3xs5TYg5cIdsXKw51WxDrjehhe4o2LWxKgWH++LXz+BOdJwSh3Q9BTV
oUF3xMcHeiV9T9tJo5dVJcmK3r4D+z1i7cNr/1bXyXEDQVY68A0vjFIgL7uoSPUF
yrd7r3MkXNHcrgKeZBm/qDAUKnJMmzPZgrrTMIAFdaFW9y1xeXzn/k7HZxcQa4fU
wgkLnaQLqMSZKLkpJRaajD4RwE6vBkcnaQRJptfXZfmeDd87vezueCtPJrYMYSDY
AWv0Aq7DMjnhf4XE/zyIaOVNAoBxFwUXT9HIk6zQnCECwboC6qxy+4PnCD8iafwi
txHtrscDI/DEulUzgNZy8FheagVN1d6p0RUCA3OFBeFayst+h7dYH8XoXRO/iB1b
fZUhJ8AnEXo03nUBEaBvxdi/137lsfNNp0pOiRYXRUpnK+Ryvzd/zKhiBCMuLdew
lX5fPNs4wH+reRUYsIeQtHCbNHZMXo+qO5r+nPH7iQ1DQ+Jn1sqwH8Bn36Sf2F/3
WeNPE6aOd22FGoklrtvcMNEA3nW4V1WOjXtiYyDbKgPbfs8EYjiho6T4O4W1wXbJ
y00Hw9i0mFeL8DJM3HEBdS5nfq0HHMxwaPwS7vlBaYwTPa75lR0VbewnEQ2g6DdF
L1ncnkZavdaNiAIJomAWOS+QLX7QooCLulogSJAXiWKwhEWimxMPsJEGu0yTSlJ0
6ImPl/wNoNSzsSa49maqgAYrkZHtXvjtfdwVwsIBb//Tg/8sOXxPyxIPCuQcNtWl
Y31pofx+xX5+4rYcvBJumjQpLTlZV/DoOs//NOBDcIoE5URRYZxBZoY3pFegBgZ0
rEx268i9KGnhxpkcfkSgnRG6NeI8l+kxtWDnVHVsPh83Q0tLjelIdBM9tLGfqE+8
EDRZ7lu0DDZVx5sYVFIld4cpk/CHE3Rh7LUBRfmOwrCOEbhT1nZZEVvQ8NzLWMNj
DT0xCEIAvDKNX2guoCUVx55mW2bl3qD7TFme0UxZNjNuvr/zWS/t6GZEH9i/CMmx
ZP9ZnH4qjQtVLBhndAwoYH6tKAPq/qQwqjSSmZUBpk9wVyYVGgelqZIXqyIiuQX5
1uJwJXb8KRm4xUJghOGGgM06njFgidNeSvlgkYPG76ftgr1hI5Y8gcDQiMnc5Dqm
T4nBkRH4yagVRkpxSJP5UewiTwGQZiX/s16GRMmocbaRQ+g7TnaaM+g2kDY0m5SN
z3ZCz5/i7AMRJRfJfL/Eo2QABQAqs9lkM3KkUVhNsj8M0/DOV97ipFaQjvA3bbt2
Trz5vnp/RqL5ky7GSAZW+DeszVYsPbqat8DPotGKVWYVA1x8H5dR8eek0qeqW7cb
20I/cH7j/6o333zUkdT8EA9JTZRAcWPU2Ous5d5RXygiEWV8QjJOo+1R2iwxR46B
vK7awl1sghZFfo3bliFsH6tSNQ24csgJ7aDr7m4eqCkAczJZRGnnO9tPMnJskn9w
IcTUkKBEGr1aaR3DcERm6YNkNnB7hsgq8y3Z25cMt4Zg8Y1fxSrQWLFu/qWqItKU
Q+hQludq8Zg3brQGbIGElQiZz1isOELkFXpOeKjW0Ppb6Yo+GYskLIhDleT56ibw
0p4BpZOxHlH9Socleifi+8WG9/Putk1VGHkJpe3PZa4+0O4MPxxW8RxZUfwpgqiY
/bgDA2pHT45KK+zYod7TxtZdJV/TfQrd11dVWFTltt4Og08zqG4puY6GxCyUWOBG
URbsMZE7k+ShtebHQTeotSnVWasjHDNl1/PRlLOqJqsC/4oRDO1abbok/rTPuFt5
k/vVwadnVacLknAUFImLFYHg7zDSaRro5T7ZD+xrQoPvTtc8WU60otqpGicllKAb
fe8UHP6qABvYDnODO5SxE7JqGusJyhPm+1vOaOCJPmKpZbPwb9fUofsz4ib0FKTG
LNvzYKIc4PCL7h9Q7pH4dlhZgDLsCt+UTpnySwN0uMgxmvQ/eCKS714kRb3dwwVB
uXPhB9uYv67/kUBHbHrGric50DWFTdNgNkyI1A9Ldxqp9NvSLaYM5mPlbOXWSRlP
3RQjogLIc8Z+D/FO+JF0Z7RYag85YmAHY36B960RVFzqirH+FYZcpyyd5rPxEoKQ
swi0ODl98PkFrmsSo0bZjUUkfrZwYM0xwoF5t9kI4SJPpxQnF8VC+GIv/NyPLMrB
RSiC7+5x6n8m5hCEiy08AhgGH6Dooz2a9isTA1+vytwgKI0ASjHX2iNjOSSbix8X
nt5POI40aLynhTZxUD3ZbhUusssaPQXjoTlxP1jaBdgUxgH5KgTcWxM2FNApnA8L
DSged6KApebeI/OCgQTExReQy1bQFZpLvqoqMoxSpOqLqXpPcAEcEaNTci8sYEM7
3zbPePrLel6t/YFFzTXwmMFXbJAkYX8+bYgn0CikTRGvRfTNzkH1oofwX0OpU1lh
dkfmI1mTIRl0xQobwS6ZQC3UBT2cu3TjONhTtvDK7sDsWFSfEyPWjpjqJ23S+nj6
dCJo/HJUYFgb3uMmetXVS4HAG0IF7MlDZJGF1pAnCsgtmlzSz4AJ2Q7Cm1+DQrca
ME99Wdmr7mrI0HOJgODeSgj/LiXlopvfq1aVCUuNZQN1CZtxBt8am/Km5kfgQq96
F0uwbItBGcXSii3FNz14UQjxVFT2Ms4wdrTridrhCEDLScNG3FBUglK2ww8Ixym5
3oveR5wdRlbB+39KReLftNW4aB9VA9LLUFL6Koj0mMrzTdmi7hjaBtws0L+KYOws
i8Ko8i5CXtIofPnUgkX9N5sLYhEfJxJKeW8h53HYbHLCZmpt3/xJwK/WGSudeEaE
v5fJgRzE273Mlb/dEU5dDxMtGmpQ9Er3Cfw/zt39K2LyiDXQUPsjI2QXW3c9ENYr
0ZMfS7vUbfLczxskkTpbq8squM4940jOFnUTtKflDF+JjW9M+H9ASAySXAJ5asG8
oEWL/g9nPiSnNXIURcCBz1wrZdigZrMIvFjo3/DYzNILl6/U8gzAdhtPxZjhXLrR
pNf8V5mG9bTLYFg9YpeT/aD0lvCdSHJmRn0zvEhKtj7MgL9y5tOXmfwrhcJH2v+R
ST3XMDA/PKDgzRF2OIU/5JAPYQQjecS2krJuNAjeeuTJkzM3pa/FmGFh3OXvf+2d
A0ATK3eprS5uL79OwD24wHnlFmYxM4c8xUmR+nfCCWz8OTrW2kEGAsnAQY5DvDHW
gnksx49xtXrYp6NcOpdYNKQ1GT0wbL9AAFw+BAIpbiOOT/fwXYM/sQ12Ee45FyuC
uuj27JFR08nkQ5UFr7X3yyF6fL2U4xkBXvkzgXHVsR2OHsn66e0sFKogr3veWm2k
3GxQty8guJySk2Uqu+6AunchuieWbFy1ylbMaK6AsmJ7+9fpxmd2sfOFYzhKDQl4
3VjKZgd5yfbFaHgPnDTkRSjE2DR1F9mCz8xTtCxl17kpxYU76ipqV3f3Nh/eJjrQ
fG/Yo+QoLn4O9iGziK9AB0gj/TRJQ6QEsNu1LZFVWiY7ZW8OGjCjppIaytXmqSFz
OOx7OxGxlUB5H9LesAODMWYGg/NCL18pjeZRv5hnxpvZhSo+BzUGokqUNL4I8Ewb
okW/2YXSIec9EK9lS7VDAo6Rx0MGuFswWLN1pSwM2QlssebGijpojaWy3r8Yc90V
+EMNbAZAXbDl3DvZi56gEVgaioOdxAXsPH26lzZpJwHHmT76rIMfariruGPeFf9q
jEtvRJ4my4gf0Z/4WLINoPHWMEWfHFTSeiXeE6WO4qQf8mrfEbb2MwBW52mzSdMu
BvWBtmpR3wYUP/6hzuJLiSoDxNe6YDrhDpjQB0uRedKd6Hcxd2mKp0j1+fepAo03
pkIaqwaMxIWbcUyCwjfDrd/nqXV7lt7CaHba/577Rte0EyE/lNQ6L+L3iF6eEkMW
ljH6G+d+bojmhtqr2LBFbsfTdW5tiZ1aEum+jwj/jYxx0TFXYc7TLbGI2hdjr0lq
U6gCFadqd6eLcgQrIlvCb7QjAFprGVvx88O3aBqHXYxAvboyCFD8EP2ZkG+CG3r6
EJ+en8U1Qk0rOkUKKh0VaIgj7z28QdRCgXrjN1fW90BrG3vlBBryLxJ+vWm9KfFj
1pN1+quq5i0ASUvzq2FDTeILl22nEl9fO6aYoXQAciu3TnqeK4E91jh14Xed8HJg
cj5DBtqFqom2xUKNVkTdhdV7vxnfDW/x7NkxRhvIsv/CH8rvqTKaiGsUuvMubOfi
Phk1J6T5NQUDF5e7nuWfnXqtLNqkn7o66PjBE00drrTIXhtROoUbKmHsrjVwuP0f
LfyiFt7jCGQW8i48EB+u/cdAl+Frtt+6dr4UqyLQn0SbnBSNmLuBbljFgaOB+/Zl
x/hsHKLEdLvdRHdkh7qe5+JufmXxkojVvL7Xr6quyCNadzIgWb4Qa5GCFv0Afbuo
VDfvQsjfboGGcykfC5NsEtdAL2r8rhmn8KMk6qzmh1EvAd2V/T3R8B7KoSKTBXLP
Csc60fE0Bd2l5Yly8FEe4QwD5ZyVwy7Z3fHKs0bGcuprDsi3UpzmdaEhGAJOcHxy
5NEl/z/m8R6StDscPTdsVp9jD3ldzHBaqXhvn4ZUN8xidKhVPCAgcj0Gc+FYWSHX
dBI7Qkwcz0Oxe1/U1VerlKvoW0lD3g3hiZ2UkU20/uXS5GH9XQOGjaM4qK1xEjd2
9rad2G+AnxQwVEwIseiyHipKksdKKlWkX/vmj3ecVI8YqLddD8G+NfTYpGnJZOmQ
gyyQVCT8MDVD9dO9SkNn3lOlUkMOKkgoOc8tZqRxv1WMttGhcibJoyobMsoLV3s7
bRqQPzQx1RwSFDHW+B2V3M/bapvV44YRjpGwVXmhscKxwIw38UdVGn8T240XXvBa
qGd8IS7THbdkTOzZzH4oK70HbR/1+vWCBTACTdcwRcl9qdkdShipQ5aDzb2LJz03
kQ0+Km/HltgDk+N2d/W1uFlBiVFvzPfXu4kEAEB+IlGTM3bNC6osl/TemyeOjowC
4JNMVUNrT/RKu8hNAztX0lqXT1LNS8nbTe4r0A/kGVLlY4o+OeQEWDZvzoK7O4YH
UpxniGkySza2VBvjlUAecpPR5jt54OU8W8ACir31XlTE3WFurKmNg/lZE4x0DjWt
8BQPNbh6IVBUSpCWMwPmYnwcXo9jSnO7PH4m47kGuS3IIl8N18mcbUFN3BA3num/
snIj/BYP+dIsK5O7E7boWvxBCEzvVdQdIfoAaJ7Xx1Qebsdddh8wYVtnT2i6gNAs
dUMv3JjkGWivk7muStjR5mpnnBzPM9QoPJBM9POGbV/uBET0iARXN4uNCdNnEwpW
cTIbeQ5fX6NJU8SlN3Z5gywGjkfIqk88cP+sPGnRGbzNu/H8TKMSAiQO5ZJ5419m
oR3oTySJvR0pP5Ewq7Pjzmk9Zgk+ZjTO7Ffuwz2t/Dw0OneL0ZOxXB4B1lW1+Q4S
p+AxOZ9S3Awg/OxWx/7a7LqqzJ4qSGVtpuZRvD0/Q+sY74RrsTs//rr/siPyanes
9BZr6DRyVmeRhXntJKiLqA0+k6AgKbdO5YaTzJmLHwzI8FBbdMwCxcN2S1voUdw7
IPi96JmIfdHJZUwXJswO4NOXk92uMPFyxJpJf3Ve4mhgis7AD8I4ba9uuWW+higu
peqkT9iJniI1hwGJY4zEgpN8LMoORE9Xkog0cMlOUPBvr4XIM1ir5Q/Dsjy9j7dB
Slxx4DR6bELAkKxg2n8J3Az/GVer0LhgKnuVTxmVc5tJpD09h85s11d+FNqNc97B
st+Wiu3fNCQnZc00TghlezfSjDjMXR7JG83KrTwSAWS8lNbyG2H50W/IK3avZ0SU
9EqMWUHAA9w14pxXOj7L3yxmjJShtwH7YgjnxtFj5h6TqmeRs8yRG2OpYxFDrBCp
d1dKAJoUcvaPzbzeddY1Xb5FnPvN8vd8BF56Ju710nXt+2BSjoNnY1NG2TeFZfm+
WhhdO1L0wUwlwUAZeZR2p2vGBbqs+Y8iPwlbSlMGB/rjuiR9N6Hqa4FE2rMPopHr
xTIrrqxxjdLcDV34G3DGjqdDjG3aflQZ/I+Vts/JZ9pucmLdt/F7sba419IQ4K1I
cKZcS9gJWqmbQ9Nm4RRUmVZ2yB0dl8yISnJt5jPA8aPZNh8s0j6UiJm2yoe/xs4I
Z0VRMhkP2pbvJOtGZzCZfBBaMrIOTPNe6/su4DAgPJuxw8cx8+T39lPA7OZHdJ8W
9tPvId/A1SFvXOKiakBbd01yMF1Y+ITRr8RPfeRG3nkKBi5JtwR1jrdo1lhIdFaF
HhP3wwSIK/Nvwgr7eYhLLocamcVHQcm36kfI85T0m3deHnY5nA/qLE5HbfrCzeEa
4AdForaVoDMNqf6fKcgQzZeuvivTxdqlSActw/tl/o1PZubs9526hwE9znBxr2EN
SWwcTq66huxLQEsF+wVzNpbKx+QOJ6DAg9DnjBcVHnC+ncp+K8phIMUbWlrUCuEO
QXMw316zSijNHBH+GNFlRQ0MXO/Wur+rDqhc2FP70dSwaU/VvoGIl7qqEZ7DSs4h
IsUnXrbbdavzddJj4Jje6qczhIlXd8rHNmMwZ92AI1swju/rU4zhkFlVsFhOkSs3
Gkhpr8uDFFj077KW2S5lrLZTcVqR/rip3Qh/XRrdCXzG1sYBXDQh2WzuAnloJsRs
5OxtRgRqql0keL8bqBa/jZjp1qa64sYyvfuIKcpJGzL3d6B9aF9fAAzFwFdLY9+C
35jSyQkK9tM20VIZ8m6xEIosc70btLHdrhUAYR/WotNmLRQg/afMbaMWNHiiemXq
Nx1lSOrY0ihcF7C3niP1qEgrOoIhujatj5ueJIYTIeIW6hrHBAh2VnW8jsRzAeYr
Q6wMgujk8TQFmP1qMMCxbCG+VwB6s8F3tCIRPk59bORKdJXfsaJy/fVJlbPcc4el
U2UKwagryjo4IX1gkazg2vlcAQzsH87dUjymd42STZE8mY8+VOK4UMKncHa/QnYR
xcYfH3exotVWHxTiyB4oC3ruhcQzDq/AaadqOft9fjiMuohr8n4DuetAOM3VZXAu
xsWGOFUmioGp/upHijZBdeUdGVWCsyyi5b/JF1h5XVEYrhSwxvFDbRB+D2GtjCCd
TVmsPAELH2wFSMrnA6cl5pq5JTPesFYAwXOp7MXypya7wRQM20aL/R5/iBA6DwKr
XgRtwuKDpXGA50+wvFgvMDLFqdBfOY5uekrCpNMhelSoHPexUcbllB3BfHuUvw4R
5la7yTY/5NssmIvh2Bzj9ED9+ym2Uu9A2DqAcMcYhh2VRVdcxezsuKstVn/d+gb7
qNlsiwVf6b9icqK7krrlSeC79k8S2P/7ZSC3i1AITxTTeHIfHepoGoIrGFEosvN6
q1AdNrLQtzNZCOKsGDhdFgt7uo1ZIyl1EpfM93Bd63sAXhdd/xs/OtV5LAHH7v5L
494QvEbgKKN1n7UpWbzgH1Nsyq1LFCPLvwm6B3omRvGC7/04DHbOUKsM6+z3f2zr
9PpCNeWPUKFGt+xyP7sfLBLblj1W5iCQwfQWv9hh+0hM8OUXC/JzVIAonlROtGOk
/L8PPW0emXdrn+EpxtWG4m0M6Hya9nTDoK8qomCxOEqWEAjArl6h6jZc607mMjfG
2k2dxrd+xpoXfCA1TahkeXWpjNuZw/68N9ipAZtASUlVaBl76P8KbxsQay4adfcT
k6hPrZZQ6LUleZx58MB+kNIIBDJxZcWpO6Kwqyl+6u5iZ1ryqTfAtmcDKRnTamdi
Walojir/SsfUtwaZVXyVLM2QK4/vvTeHhQmTmXw5F9Ocj5l9k2fQtuZOr7cIqT71
Xtb/XVowuNUilb4B9E1X+hNg7MPs0jh9xKn6E619N1khdULzreSaualzSP6OV333
sxPs7iWf0Wx+9ALTQBGYEb8lnIgYjoVy7ahzIpN+hFh6LfPBbepIez8dMg5C6eRC
IVdbELWP7ic6+iSgFOQNnJ+ZUMc9yxPqeg5sYS8RV11Z8Rgfi1owR8+48IrvDVyP
ghxdQPdJr7lZhKfAzxr6HkkPxc3p/BpG/PSQRecHQmGXT3c6j8fV0JQrauvCeAuI
Jh30gp+rsXeWge3Wurn6s5oZ1Dx3Bd8pihoH8k1kV2EPuaSEO2YdMJnpiYGxJtUT
LFHgkRqbynrU41ksuyd/Ch9RPRWqUDn4Q+KlMvHcjaWGCALDDlW/6GJnODROb6Ql
J+Oq23oZMd92c9xNxBjwwwjfKUghBKGjDlic4YGkjSBg/qz7EvpnNGut18s9h4jS
Y0+b2WgUbAfNBBSbKdosUInCyugFB9bLxAkS51cLcUJhNSA7/uHwGYrkWSGQO7vj
6aFs+P28yAQCSl1728S5VskvFJy+sGp+Pv4KkHO/fh7B4EVz5tVRWxSNA1x0o3sh
/ymxx+OvhL4fSrE2h51zri7J6tn1cH6MO+WsRkdLsA1ST28bbR51A9RRgDoxklfa
3of9iOwP0k8RpxaW25v0ZKEVhJWLOqy3n9/nFndJQ/SheoDerkZVWyrhFEvxvIcs
ysQhjNPRCwTJwiUHRDdaNN3zKtsK5rf7dm40NVIEXI8VSnS6sGFtiPlCZDewaZZJ
PnW7+95k7al7wY4qahHfYJpzwPoooqBrJUcVg1ii9gSx+0Cfqb+qjiFRhTccCaq0
5f5N87MncmR2rgQnv1ooqouRu1q/5+Rwgpcrp/QXbqlwy/g+FGl3IJo7/RGrhOtQ
G3RyLfXYm20T1QgTIVYFgdJS3/5SAZIz3jcaaRrVTAH/YgomcaFksmci5tRakxH3
dsDr/Qn1OjtMzHzqQ1CrQvOTSfL8n32LlmZNMNhsOiAyVLA624f1iFcpJiqEIOk1
b9c5cZb7/eqEI6zC8cPmVDRuYnQ4778X8OcCiz4glu0mD/j1AjrjZmeHubrGPyln
ecCa8NRWdQ5jm7ZZy3ejcm75bva6sGooloYo5Rhmm1tJ+0zmZ05FDTZlU24KhYt+
o6z9Cu7Aix31fbrO2j2DrKruF8ZaBKi/n7MukRy8xjP5phzh7Wl+Bpu9Wv1bgrct
5ImyMPUWWG10mwmNKvMSmUdIhZrwmC4F3FDJ6kq0ThD1g2tjT+n/A0ui545a0Fum
LzbOI+8SoxugNI1BwSPqbVJJ0DhzU7p+UpR5QHVVJWyZR2UohjkWQIrks+V5Sa8g
XUQLZGDyyBx62KqlPN1py6KgpTh2MXJR9jmxA8ZyuxsfmfCT1C1FJXgbq3KLgUke
u6u66gElcG51nlLzUjCA/yo+nC4U7jy+cZwTQFCXWem9UOwjUW3rRtDexBPYK6Ve
UXdwZFrIP/HISLaHg5aLRKletX9wKy93EJGugnl+JiztyVNyxTqIxyuFXAUr0lIW
UfhxbEqU79r/WucdGIcq39zf37+wEAo869/ysNKhSMfINaO9iVm/8HcsWUcOOgNv
XWcehcjo528Cz8iR3P27dc7frOlDngWqHBR1+k5OMgp+2xP4BFm/hmihh2j6BIhP
DGjEzYjCcOUy/1sRJIhj7Ma3DdYmmVcMyZjmdGsMIkAz1S01yoXlV3KkWeMLTlkg
gdbuaCYLG0LDpLq6zO96UY86UvreZ0jeSqzXTB7HKrUXKYTvV7ntRJUOBR3rqB2L
2wp1mWOE6RYbmMi19hQ36iQ7lCTHNcqCLU/kyAdXwrkZF9TzgDVtUucSNR0bpygK
wl72BVrYfRJXxAGauvrNfJwnWJfR/g6+g4qd7ehKpgJ0IwCoptc1yAE/vcuWbi6e
BQn68q/L8M285JPWHVzQ0KD5k9UKme7hG9am+kNXOc+8Kf/3IwreEcyBUeSuIm2s
zsDkoOpOUf2EAf1GxYUcmH3BTCGg0iOanrXo4tz+USXK4OXDx/6Kq5MXnQsBDh0F
3+O/PQF88zUyPaTgTetH8bigK6/zZop7zpftrK0Nn5uWThT1I2fVY1kbQUAgyrxM
4eMYtqFkLOUSBMgKUzxvuPLQ/5VRZuFiOkTRRDgdt1zhAJiSzq8cQG8RYYH4M7uY
ECn83L0kr5MOzU8ljeu/k0RtWmoPHgTRBjC+QL7npdThJr4JHo6mPk7V+hvP7/0U
Psp/zRUm/tV2mVVdoZQD7lK/IXOn2UxwMhIAD+pDpfOlSuzABP5vJLftSZJzbkG0
c5/4xAuKT78c+6u1dDqRsAhtHEHnzWNwvzU0LHRPxLub1hRBaHY8ePLWAl8nsPPK
v0tf/9WBdMF6kSfdii2QrykPF83yiQKMNLPJ+KUlF/I9IoayvKLrij9vTxoZtk7Q
x8zd1S8nD2anh0485zVr1gE4bf3l2A4LwCadG8M7URy6wGK4Wub2EsyOlAVqzT5n
63/521mI1ZOcEPpa9/8JPXbUQ3HUcqaacQtnqYkPuszPJHsek4mHrwWP6XTKiDcv
2Z5j5Sh01+Gv9bOO/LI9vDIVNEh8Pb5zTeuSR/wgT4ZaiNRPSt+3bfWpPo1mXxuo
bKdt7TOsOyPXA1vJYM0wHXB2J5ULYm0oBhARa7xu9pqb/yuFJkHK6i3FNzTKRvkV
0y09TJsrvEChGKxopCPou49l/Ch6FfVWeMJ2/ngjzwOKUBJufAharEyOzXL1nhHi
35G7fzmk+Bh9W6I8BCI+J9qZ1BLqmIGKTvK12WOXQL78FsRW98bI+HaoO7cJVb/A
8gTHPxwcak1OSU4V19kK3JYBmflmXljtM0TKiJssWhiB8QBCZsOt1/BdbCSYrChV
4jz4IIcd8+FvzbIh1AyYOHUgRx50EbpsnZSv1SKCnxwxc3IEr+rXgfh6pUZm4GD0
XjO8QYWlFx/m1oZ1AKu/ZXhDR2cw3m88Xgr+dH7+gFSRe3ZH8oh2AxR+8MzRZhGb
YwO6Dqnwy6ydA79lfMnc8n6MeEzhB0GLNDrv5Apk/7Kow0s3vxe1NXk5lo2Xu/aZ
koWTvgsVFgbTnfc2hY+U/UgxIZMtn3QoBCSLbB5Ot6I9nwde+YE4YfZK/yLdBoGh
tmTigUes7DOq6wzqeI+Dtek2SrsYhBrq+BOrixZtH/Bqr5BmzkFOyBafEycU8BRQ
kswUMi9AYBOKSNl6bemaqgfgq61fyJR6y3cG/pWgaXUZKeeMr7/JJlx6qsuAqNPY
Rs/VpEIMOSi1DREkfp2JcfGVhULK/4iolVZ6F5t+piZPHP/N1RcxfU40hPLEu4XO
I5+Yq35ZMMwl3jdlPkKem27DrUxt7uQ6UI10jL31zTneoCIQCri0wXpPW3FHA/rC
hwKxouwVEu5VD2kW24GF1ulwrUf2DU2aPpxHWKMuR4JisGNVzc61QPu4Vubh029A
M3Ljx3Ov/a8Vfq4b7Q8F+iznbd/xgjmHV254quZTDYppS0TTI7NDjA4N0n4464R9
aiIg9rwRHiokKhcI2ZuwtYPqGWT9q796EcPdN7Zzo92BEPHN2gRXiNN7R6UMBLMw
qiOEAt/WrAhSuRc997HlanpwdMHBl3XTn5ePRFzjHeq+uP8NxsX8w+jJPy6pcm1/
D25RC/i2Ei4lP7qm5TZufr4dxX84tVqRbRtqRIuLsT7qq4B2+sbE8Cta+686NHbo
9eMf7drozsTIhx98f8bezsRBZP9zgcUYX4Uu6x29Hx6UDOcNPZGtQSFvUkB2t7md
101fQ5JlbznAJbhswRx1NUTidpf6yI4RvpXl0k4GBACXwpgMNPwCfJ6i1UGEEEHE
6G1rjv9usSlmBSmQJZaFPhc4L9HSbd4/pfDAZaS2uSHI3h1F3fQZbBZEQdcApkKu
Gdyw4rMOWr41Kov+Hu43in9I03znmv4s3MdNo9cTxgkSVy5zfIp3PDi5Vp8Gd/G+
ufsVScztjMG8rZIm8zwhY4VKM3myR5fHMeqOX8BivfEhpItq7X++kVtuvZTzZoP1
RJsYhugW/4wlaP8MG65uZZpzXQCt8GKbL27ccR9mTPVY4DyJrx+CLhOSt06SXQjC
fD/Xd4M4C+B64ScrKSip+fLmxvB8jdiy3P8G3zSZ++Xx+FNkzsm9ROUJUsh9zBqa
Y8pDb/sTTEK+rgwlwKttL0CF+Xbm1Vvozaf1rbRDix/rHRBJjWelqlat+kf5xo3y
1e2zDjb1xiywTHiSRPF9Pi40EnmcZ7VRoqzsZg4GHT3rYvqSG5yMrPGQKJVoK3o7
F6jV0z3I27+2FTR1TG4xl5jvzOHCW1bs8AD2MMQQj+oEXGdLQabhR+LxlxZ/DFYa
zH8qfOWJ7bUjQ9ftxN8TN+MLBJL0pgKgIls3ZPrV4IXYI51dW8fHEYvpMZolf2gp
o29OpoNFYYCQxFjyAJ5dLWL3zabylyR9hUXF2Zg4VkHqgQgeYSef2bfQZHKKqQoc
evccREHdo9mngWVL+Qs0bKyZcPae1P2mzqQjTtHLanZJUT4BYBSRgiRsBQnvkEg3
6RHUXs6UuqQAFhH4GUX4Ty9nyV/jWTQT337jMC2ij7dHAKvV3yRkCDsRJI6+adBA
UIUOmb3HPLNSnAB5EznLSZqbOub9UVJ31IJ7tO3sya0VI/yVQBDImIVarBsKYM/o
6wl5egoJNGRgPQ/wa4f7vIn007UysND/B39t26QCYXVwFobsQLuqdYvM2mOWWcgM
+tWMzBNdeBT9iMHeIsRfzfIGC80lAKtP+L7vnFu/Wb3d/Y0H5+uxQY4HhopJ09t1
M5jcZrtALf6Lro3ooWxBTy5CUORWEKeSbfY0PlyfOjiAFYMN/ECrL8GT6LR/HXt1
3ckn4H3tO2iQYL1QsrFib0eFNIDJyLf2L/mQaidZWhY4ixyxfHVfBKzWImfuDVFo
vpHZ+h3tppFPhVpuW+khbtvDb2m+Lu067yeT31ZzxebzO+I2NF9jl4IXsg3jXdy7
qtFUXL/ZJHlfunEv2AhtDnRFKtmvfpG5iK58I933Nz4mFc7klHz/Tl5EletZ6GlD
fz2qHqjXlmcpFgKOlXSoMGc7oMy6ONYkEzAdd/Stf5WVCqqvp1/H9v6Uw9qZBsqC
FlcaUIyCwbe5tzFzOCuYUgd3jkGr8BByU7SFdwaRGZN5kegRA+OHYqoNvSnWOSUo
2uedvKk7Z4fEXCOtD7yOIuJ4hHffyiT/ZV5kPTOg0K/GVycBzSVDMwd12gRNTRWu
RAELknbAUiNmXLmLjt8LJ1p2xT9jp4SyD9TgkQH22pyoNdavfNvWg27zrSLT2rah
c8zmQD3HWuEayxmVt/e+Dp2QX6yqk81qYrj/AHq+yrU2P1+xa8OqfI7EVRytrTFu
sHG6KeiAN+FDL0+mnjjK8/xQ8bNld4ohWUHCYlqggBWnJiE76WOTpbPxD1TAoqCc
jBFg4dHTbsx7N/CGCpnlPHKfQ+B/08ZGczheUiFans6SKRZSZMxzGs2/5qiNluG0
+wYHWvP4IQ7W/nYTYo1uXPyAyN5+9+/xN9sWosCa89LCoPSnYFH599g4p7EgCQ1y
uI7qe5GSNwPfsVJhALBKbddtnWo/xfNUoLFRu29erD8xnh/k2C9vo1oAgNLMZ0DI
/cWdBHFqQ/0cKpOhao9RNcyitSVQC1gtKutaxb3tOntLY9CCOHRoqPrz+NXwnrUb
RKtsaSbXdCpSDCt1IQdDY09S9ft2d8zUvhyGCOAPIs0EW7YOL8Q+5SUay1Rlc9Eh
ub5vrPkwRsgjw/rgFgeIBmhbJSdVm8vHWLu6VbLIinrV1gNgiiuc1LNlSUIBvmgO
0JtiYzWdV03gYIn3slGPeGrrUzzimUxtp4IItcEYk46zCy+MCndGDZn60AXEpH+g
NSWDNWmEOPDO/87VXS2HXHfWqGX4cQ3i5TcG3EE5I1VHB3VToc3mMBEXkLBA0As9
qoRVG+9zMLERYQNhhjDoPr3rTt9nMrsiuCo85J3TZvscpANtcXH5sheBA1Ok9zAr
LNdGgH07fSfFXtrIzrp9fXZ6FWQlmb5s+5dv2Jonvo7kQn5cLExv+CmpXkNxwvbW
iJu8zbHhI+sj0u/p5LHEtt7Y8/CjGOuyMRTYcouD2rKGO7VDXYJi//L19uR7jXQ4
1pmwRti8Y/yTRnsJCEFdbO5vT7+BHbqspMdrvGZZtg9VnXry1Lr7wkLRxG7OsXtf
6kc9C4YAswaO2lyzhOTS0I7k6WB3AIWf6Zo/CVTP+7CqGsWGWJEBH5XkbN2SWnO8
blwK6Qc53zOewWnqunh7/ceVBGX3IhF2FqB7oP+NyYnnYhn5cFByoVoHpHCiZ94m
ff9gjLKfV4vWUTz3FySqcQ8itXe/fROrke1ykdRkrko7oYFceHA5C0YRre6k8GZy
H9P0ZdfQGJqho7E3k6r1JdxZszkFbcTG+NzsXYdsBFHts8tpPfz6FPrRZZElRKY3
Jpam0FTjliSRT1WaijF7Gldf1QhdA5zmwLvYC7YaIK6Zhy72D7ecPPfyCBMIuWh8
HMZzZaHW4YciifKNtd1czvcZ5Z63eOcJywJVhJVZ/m7C+9HiGHL4MkoywkNAUFpL
0VL46chOzoytoNOaqkrcCGHoBb30LMDRuGhwzR+EamBSzoXPAPG3PwIueq5N+MR+
7GPKyQFEMq/Dn1fT1KI4yqCo7WuMMAnwSR42LHH/9eE6x07f5yf4m4aULuEshj2w
2AQXZYQWYJY+hmfgqhf4xTVHqsxZknjz8sqeHkaxIksoyN8IjgzrfYhLcgqN5wFD
eAmgKQlWriRbrljQobSygiH5UG+KJsNaOK9niG0nZHH01ET3VPHIcvb/MAmTnlkx
907zdhG5ycU/36P04Axkb9NiA8j5/eiuN+1sgtHEUkYLOt9hJ24pnK5my5HGwOlr
AY2/bO5Mw1ENtE+C9Rjx4x/3UUNqWC7SkPi5OdAXVJ1Ox0/7QWdbGLFLLCWw71Jl
eQk5yCRLbS6o5FXsdkW5/MNQ7kBgVBEo2bV2BTy2F33u5hdGOWyHwl8egCN80a0P
nX91TFPsZsLlp2Zp1u7u3Xm0gupcVElJzTC45aqNkUXUh8SjW6rQVTmOJVla6q+u
N+4gvf9F7FZUGkGpQV1AxeazikLvtYsZSYpSLRHlm0CHPaNF4gX9I4TmbuOHJ8Lh
todo6U5rqDgJ1H+4HH+Hq2CORRisEU8/+wUtp1yGyvGQvUJs8G8/j3XPApOy12vD
kva5pkv6G3OVwpB7YddNNBDh9GaWzNMatwj8yKrrCWD82GcO7iZgMi5xbBoL+0Ds
5yNmEzaUUQ3KzuBfxMM/SCvjZ3iYdb1P2Qko2Zg79DRiAYIfKMZWolC6IfAxrePC
9BoLUTKPM9L+rn9p1yRFQ0peh86KU1XtG04gMaLPuAGaas64dQ0W2prVcopvPlV/
o2Lm1P3IjqWYHHNgnefsTOcDUsDsr6lawCkwcWmzU6PkK6AWj2t4KbCglPksVyY+
5o3q9csKnU/6fly+2L+5KpAuerKLM7bAa1sR2XLmdrETIX6YOj1W4havPGXKq5Kq
F4qaDuslMMB2F02vCCpMZuRj0fM92WjuO7sg7+gar4x2Ydjixp2+gZwgdGngg0mB
STE9rZSZT8bvMTwjlv2ddzvNEQDJPA383cNvRMnWdQh+AnCkuLUpfDSWOW44sY3o
yU6n4yLoXEzN0+7C9KkoMckRgFMyqjYKMPmlhsuKQ/uO60LgiW10ya7TTPpK1IX/
uV4PWBLjrrZfkcDBy8bl1L0bDQWgRzEXUkIY3h/J/JTrWZ0qpAtn/QNPVZyl0p/m
x50MRdjOJCOynVqgLpIA63CAnX7h6x+bmaZ+kFPSHHGnAERDh0pXxPUtL1Bg+9Fc
2WfgZwy3aSz4FOBJr/IvOVqEVJJYhxZc0cd/4cuSiBpV+rXfWIIiMZNHBAMF41dX
n+cUnk4982rVUmg5T4IIvBsfPfAQ3Wjekpa6kbnN/m1VK5bHakp4R7ECmq9m4oZH
s3edY1v88QsE8+o7mP7GuAmpQCVRppJyk3o1KMxoQl+41AkH8x0hPBCqZnjHZ8t/
PAG9RfnkfFqG9xVIeFrWfdXA2L4C9HOndDTjM20+QHX+ZLnBD6lxB3sHl8QXpTbo
AmbLE3mFfdKGKBhAopO/PjKlczEvLHbwTV0hA4gKdNV9L429TaNsphjra5+tKBO9
Ao06WyFB0yxsCKhnE2FgbAPJRmEsUs1m8hcGRO22QxDF82Kvlco6qnCmnuVIiRVe
6ZA//+VBmi2UxbztkAjqfaJ9VLoqyIaGSUZN6bTRtBkY8kp7CdShkQlhMwjvxhPh
BGlTrLmFa+IS5WLwHFpnbJYaeZ1PzWbqIYgPlrGiZKESWIEZdotd0m+371mQbSKF
CbeoKvrqm3oxePU2GHVN0smDBFaPzgf7oqzd1sXKsZ1TLjsHMDTYO4LQBeBumodB
/5GEWnq3zir4YgeHOfy2JGxP83dhtJ2QGWl7aWu1ff40gjYTn5BirF3/KMZ13WeP
aNKM2Z3DsOfVw6O3a5sM9Do3lMON2uo9ysul0ezCgBwexcyTffAYEUBHhQoF/TXv
ue5CRUGS6AJsVtOagstU0hvWHh7POSKtJ+Uv6de9frJPZtOGRCrdu0Dt25jv8nvp
ONzfiHsgeXyV2PdkVYpfNNNgftUAi/1XK5ATbSgVl12t9zQrtAMdHOo/nN4p5zNg
ygrPRjJ3pcrkVhyTZDBAECu/eohRfQ7pTXLaOjiOMlV6fRYARPFrITBMqsbbyO6P
w8bz15UZL6pd/yfAUlMIXRF84k8WkzjNtJPip6pG8fKGo3a9TyKEGkhsiMe053xX
c4zygcBM0BNzrttAhEe53r8N4rPy/RiqcXOR8xxq0CBp4wS8PFZwnAfwj3a9Ooh8
aUtbLPYuaTPO7AvKlcjzghW3akMsPRd3xhiXxTSaQ7cAq/NpLWCSzYGwVDPYL3Be
vOUGEU6N/ybhVu3IEOC/Ygabv+rh8AAu1zzRm+lsY0mMgV47BC3GIcp5Tq1v7PgH
/mA+a14xTsrl3s1+1C+72nFFJYcd3Y4o0MmkXfWYAXHMSNHiJgiXbIVRt1YsPK0t
u7QnSa54R6RkyQXwMrox7tz6tMzhoolmgWuSXfeILR2+x9SWdeGnli3edmyKl5fi
M9EOOTusWjhex0yVK1imCcxbUsxvnv3xpxlOFHuqz3W9kP8urrzaf4nOniw0gjM2
UcCUA8AVj4igtREVYFTPjiN7hdjsBsusKcV0TTakd3Ak2Mbo0sbFDGxajX9OFVBw
Xb/4NTiH1xxWRTsWueRrioImX/346kEuQxe1hnAoVZNBrLiESHh2xVDS3k7L9xwp
dBs4gTXHQ4bd40dAV7WNocxiaXFhlStxGAlSt5O9wsXBd0S5wlrjQ9VzLDSmfcS9
V2MZ5b6OEARnRWwiv+jwb/03mKqTWIbzp5Jdg5NmnBoE8RNJpaCiaVPmIdbJlkiI
3rpOPGn9vWv/vtn7Y8dgxcjWzTei8cXfQRb9N9I5J9nnPT0N15qC4uL5Avicenzi
54NEIdUN6YGko/MYsz/BuAPKKIkBSh4fWuQL8P07BHwDw0n2GR3ys4vs2jeS8oCD
tKJDWXo70H340QzfXURHFR5mTDXs8rX8ZPEktBQJWFlgELIgO7SlNTgz5vgrLLSV
mdg3F61v5Zo2JZqCyaKF7ZjNUgFuw5DG7o6Q6IM6sVlGu1JaBYc3vfwoDx6QdTLN
OwO9jLK0cLH0Ey8JM3CI2GYMAsU7vJcg2Ep460Ca3ontSAp66D8X9D8dwx3DNlhv
GbpwyLppYmdvBFr3EU8Vow7e+Oagrr289U90waohL3oavlyoapNWMlzy+4OUCP2R
3HyUNEFE/kGzJkUshXeTMvfNdhRQGj4UMvfd6Q1Vq5M81LPLG08trX9iN5RJsot0
+cnbo/vcs1z/hQL4vO8KEW8rvBHYoUDjQH6agg7/aoWiDrbEDUsbEY20jfUCsbGF
Bedl43uvtGImYg5ryRQqbavhB/BoReW/715m2hK+pil5wbCkAvN6YLMWyZgcJOSN
6zoeW8khV3imJ18gtn3dQv39NE70rVZ18hMXEN7vJgvDkx4tx1PUhiYsqSxDoxGd
NzzzHRYXQpT0L9GSEEtML2NGu0LdOfy1cwADWyrWr4F80D24VhmUY8cgpmjfkexe
DOrhgCrv/OaFPemv/Q0y3YtP5eGMqlkTv14TH1Isih6Hh8JdvCEIVz1F8HCkk4Mg
Kvz++QskyphbO4RnKIZqASzFOYWg8uqCrUYuE+j/X1A+oWRYu6w3AVg5d87Pap2y
HLewkMzV97TdfK6NoK/1pkrmJdloFE4SRPweilwB6J8bLwhLVeItQtX5goZsEJrh
we18EoYaGV6QYsv6ofpyPxxUHaLCC+8m9tIqauA5fqOHSb0ZrJNFFPeh4clv3A2W
J0Q8RcpQTvB6QAYpQ4bu7O6WUYP7NPoqRSeOAANwWrb4CPp0d+61w0ufrYFEV79E
nesdt7qH49e1Kf9lGA9aYbrB4lS5DK4rgvZFrPjYKHil36hP+Cw3ypfFNHmIsJJ2
thdg+aElm035M3Tzctok4P6W47jRHlbCFbwfUqaRzwuMK0aHyx2V2uzWTiWsjz3m
NBknVOcp/K45bQdFbOfoH7b7faN1JjDR8NVyE2oD0bgAUSBmbeIEPB6bURwMyTgL
a6vbDKGucMopKsFHDyZk+ryMQyBIb0V/HFJXSFiYspKFm87bnPYGXKkiR09acr+S
yRJZattxjP7lqvnAoa4FvCH4tdCaOtPT7oxHwCZd7SGNS3zml/9TwaMVLaNDyUSf
imM6vDEoGhZSQyD73d45qE4rjc4p8fvSmQKOz9WruhYEO/f2bYbiUuqzNwZEZUOM
mD/Pz3h8PcuViWx5WCaZ+1kmhemPz1RC3lr+yy1Qhy6iPQtkgdXRtXjA60HukEb6
DEOJwcUcqUpecmpMgOiKQV5KDWla0CYkLrGdcU9IDh5lwGmwOBTBE2ptpXzcJRBr
0F11ItUThvC43Ot+X5YncLwUkXWUK+yXuuU4syu05c3rUFvddkAyrZ1+gzX2KeYZ
g4Oj/fhuJ/wXGeKOvnqBPmEq79gGv9fyPX/4ePRZj4fubTD5XFdvdbxzKyndD+Oc
l/jMCpSI5OM4q8O4j2VnUigBuJq9zPMKhNCXkGisTF82/8PyAgEDPtprRVtK6Ofm
T2S6Bw0WZXo9Srjxt99pd8oLKmHn/wIO8cyBZ6PNk0GAN0DWRsT6tXmwffubH0rc
vgwiy1OZ+tnH/x5mRRj7ATa8mv7/kvrZeeQ75HGgs9LixB907f0p4LIQC/AoMuTJ
Be0p5UlBQIecDh7OzDQ43BhbsjisYVvPf+RrmqdukamK1VgfljycmoLRj3W56LJI
5vVyIZgAUKfQrSqxXszk0nucXQJcCt13iKl1csiXpRKVAf63BSVVE8+j9uMj2CxI
C748/A02vD4GQWohWZDoVP/Azw3BRDdcjRSVp/FCXjzcrcpER1+I6Q7+WZiLxdev
tF/urJifU2rFoTtN0yUUYcd3kMmb0J9n4EZijBhJDFbAAYeGXYCuEbJOsmJ7ypQY
F3oxD9OdvONfSqJvwi/8fQ7L0p4peZ0THRwRlZHWR6y/Ip0ssghG5jCt8tSiSxWL
gSL3Iv4yHlWMNjj+QOEa0KIHaNl8reR+YsvUY/ELia13cH4E6LPEayeh3aAHfdDO
tap4p8vI3mx8ClN9pNzlqkX+/egVcGdAq5GKTlIhU+h048BX6P13Jk34zVyyyum+
/zGZJIbfdYf6hFJv+AgJQBq3DKPUkzaSAdAIDIOIyKc+iQr3HLcgjb+ieV5ywcWQ
wYKIdRlzMPm15k37q4YXD59NKkN3rvc2zQdFf511FI0u1mXdEtCWBPTVlHCbEoU3
z0UK05dIRR88Lu/zYBwYZmp8HLUktlMxbfdYQzUB1DmJsPnbY09u5XHgn9Dqtzw/
ecctvRuizciDVWs3px7CyQZPbMqg94HdZCPB1dYhM2q1OqS5rZTKjTQeX/4uv9GP
AvqdeiuykQc4lG3jqKOaAhEkC14Z0T523YthXhpOGGq65M9yYKvi8wlJfeRcM6Kq
LShwX8pmj1hw/wNeLcQtPLmAoYcVqfpn9jbjScO2VmtU24lZ1jXDVzg4LKSMg2+L
glAb0qylBmqRkKw9loD5hi2lpf6qCsGDZAfni1OgJOO862IRtSPZXk0c9pr+XNZk
hNWhPXqs2nqRJLVBYRNclD1RXMFfJWA+Th9qyepNPk34BcIgErGGuIVLLgb5oG6J
0tj71EXK8eaZXi0qMFmv0ko3KHWwDVR8N1C5avqObuKg2P+jLRr/HFpA1ExUKusC
2DvBJ4FYICeSpa/kC982dV5QRjelADwTZgaUf7YsTRR3Jx8B5iIb2kjku0ota6vU
iBgxrCNgQ5cB8HLmBckpvOFq0Lac8VA87/BDr0zUEEt8wf2y1HkZmWYnw2pCIwMM
gp2uAQWStTXAgJLbLeuggPvTBpjBq12kkIpNVLgVuRlB+h6kw6jiISKBjA14loTM
exAkLzcdJqj3TC1YPbLkFPMIyU0R7vXofyGKue4ZnpQqClgcObmCHlN/KhhTIjfw
KDbM5U9viUJp0XWp+6UOMfuh3KV34n3gboWrehDPOVR7Y3PsVcCjHkAF1qpVSy0j
bDN7G8EvNSfTI1Cvj3uRlZ/dNrpgkI4FRquRzMed4HYgL9cYMBdDrTOY/OHFimpS
gH2anqpCtEbJd+9IleOw+kTDnOcK2/KgX5HTLMZC8Rd4yXZAdl6cZxSt7gWnT6nv
UvySA7QybSuGdpHbEl8QJQUz4j8bnPQBoxI8s/nUMOwDk9/uu0/ARejhZUopV974
CQEszpbWeOvcUMelesWnDcOipCXr881tG+OZzMTWH8woUT6FVmS1oD3uhUo/cZPY
fFSnDjsb5V3fv2hIrczgcHwkrvgnBIRlLb6DWoGr5joTy50qtM5hMuHwI0CIrgZS
tFZ4Z+RXCVnqxq4AeLOtI3hBulvJkr6WOvR/DvZFaFVWywb1QxrxGwIte7HwKBAU
vFbQxiOcAQrJc4MKZYMBKLB+XITbFRZyU6G8Ig43UcylJ3A4OThly1LIlOJocWSC
JNyXBJAQ+h6m6uaEvVRowi3Gnlpp+uG02mK1oqBbxsIRNnZKfmfJzbOJp6pgyATI
d8RWz6BlY7eW89M4BaymDkeHevyC74rmv0nn93zLFXO21kqWF3kOCP+1klR7dPbu
MNHkrTuglcc1BWGU9dcPY1iLzJiYyZyx9sCk6ReAiII8UYa0JgH3qIvf5Em12rYM
jhkJqljcbahmusbsN54lH5YVYw27K84Qw2E8w3gYjlJVb/wff8vdRuaSs3PU9Oht
UUMOTGhh4LG1uG29/ZYBMmvhGbjn8FWVHI6x+ZhDqyKPWQnVTg98WJ4ILH5yazJL
mWFLbJht3nV+2J/EgUn7mPdHqcN5NK5MLqg0yfGH/kUn75mXw6I8UW0Y6zBTbFG0
MXgyNLRxH41wCLptTrcwDXLRi6htYS43u4gK4it7V/1Dw0maLiMYnlYVixqzoET7
bFI2Tz3zTBJ6+vQLcl2ZOeeYeRffvQDj6njTB338u8cZXi/6svMUN3Ie/LEPrWWs
4vxkUNhM9GINGh6x/WjVCp9HN+TSiqJBuYnvCToshV/6I3CXCGZ6f8GDUce1qt6C
f3QVLFSkmwq6asUDLaw6+kcEolxeyR0LzFgzUuVpJQWvRehSgNLXLTwD1UrnwH4o
9uIeVHuM9TBSbU8Vre8KLoKZ1ZNemSK2ZkKXJFe0EwxRSGifB+lv030szw2T48YC
z3LA9ci5AyGh1uModQb6Zn8tl474IWztqx7Z2I46DUQq6CjLifOH3LRhtqFtFO9z
cRXEUSsJXdqyiOm6OiyDKBNLlW7xUmAayUfqlhoVQyQE8z5OO90cm+RYBx51X3uI
TxJak7iVTDkt7BdoDGBezDt3tsqKGX+s0JKPA3wIy7BKUogoUH87lOrKrICG781S
um5ITeEzH0C/HMtfTrsiqhnUWxc6N8oEMBUh8+mAPI0oMGenKYFBJ8B8TEOT+bR3
Y4looC6y0LHljuA2Oe2TD0XwDoN4moIxOcQ6r0sfdbyfJEDMs4rxD7PPD2NF1Hf0
v+6hgdyUlOtiotL8WSIiHC3VFkAV9rdpOHrTqNm/jlubIB6EwyFvP+FcMG30ggxd
sFSmfMw0uneTwNB+OeDw21UZ8i1faSRrwBAQxxBrInmTBiCWt/yG8ASGdiyp6bbU
kEVJ8Fzs2JSLl9eOemFTkdODxAdEgFm114hlDi4PSQ0Xcsi9Un7pKc7OiE7ra2HA
lNlqwLg7Cc3WUC4/Ivy0RfbtDmOBb+g3wSGFezJt9VlbvGtriPv84Gq8X60u/bv8
aQnam0+2CHKv3gyhZV3YhF08hA3qwZelOeFW72tr8W55oWM6bj1fyjqAPBymjFn8
jrBVVHdsin3cmQOMZ4AIpmQupvsC5i5AW05SPI10YNJqyNSTpdwIRhMppBrsjSa3
XG1v3rtmytL1Bg78J7KgA80nXiCvAmm2J9jEB04W3iuLcCdaqszLjFaVvaeEQMJs
9/kkyrPrPJd8apeIhxDnnUsVwnIQaQ7k8PJXZ9qldtMf5EaomfqJD0dNobDLI9qF
ganeXja4B9+21LjwqIhuFth6Y9j/p4SVHg6yfY+M9iBy2SBmpviZRCUikNe72/40
SKDT7JH/sE4w9jwZuklLQlliNxFlqqzEvtknZGZE7A7+OoyXCFj0+AATIW5aCZsN
Sorjxeq1a4YeWKAnQkLlWEz93ShRW7IXusaQhR/wK0aWNHcPEt5vRyZkiLGH4eXY
FUTbUQmBXlm2SNl6KrlmevHhvQN5OdnNQF/IoJi1lZ+d2rfBmrRRIGy5TmI5msz9
so5KykQ+NiYP6Zz7PYqs//y1xoByOFnQ7w7fPm2sIXUltIRc+hlZmCwE4tsvhMEb
z+RZ+W/fmGEY0+nonMs/Lk1mran7qDCATGzQPyhStrQx/1ySQkAYthZuyK1YRM5E
ghppJIPJwFqhSoG2GTjOFL6fafp8EJjPWVaBNcU2tHPRczL05rmK+4Sdgkbhe4Ef
xdUXts+4s5+6f4wOJ021EIBe7a9xhjdNt9vgupR9fygkpuW9IL/FwuxEPDsTrQrO
+gbiDV84nwcuqGrbFpPkb60zQXqBYKqKUTjz/urGAVS3FZgUY0q6yl6MeJhyc7yf
IKqbtEekv/fIl2WxoFgSuEdTneHCXV7ezjVSAwoaVgYpbsuLc1HnfzL1NQXFSfDj
qCzbMcI647GhhlXzqoata3Uu9Y2hl3IcorkDjgONC4Rzyurw11Dtrv5Gto+bYsUv
JPCdQZ/PbL+GNu4kDwy1l7GvH5p3gpJYwg+0yWL7kqj/t57hzc6IJvAEVmCcK7sU
bmCOcdOObxczby2+sIKGyRs+bUb1FCcFqHWI1/BYm37gOCd8Cq9AQtX9gmeaUe1W
6xBnFhYbykljxM4+u2sY0Sae7mthIZCGc7WuUur1iEKmZ4ox7AcsZpB/vv0iZXXR
6Nzl4hu+HS7EQVChTLs/KrFchpwJ30CQALaDEq8nhoewfun5C3VAeHW3iHqiPgpJ
88jz84x830pX+VJ/tD48vOsB9pNPpkpOJ2EbNcuhs2Db2FWRGLzsq8CeRMzEnY8G
gjrNyeyhc3u0gOpi8l/E1gBnJgIkLJB3Ny9XG+vcinob2qxXiDC2S9Eh/HCDzsbf
jpviPzxL4K82ST/u2c8NzYQV0V5NK7irXu4qnt5cuYSp/cV0DJsCzqAV+Ymm4v9r
RbQvhEvrHsY4zHf281gMQeO4si2y2f07Z3jY95EGJObTf18tkqdb9yd26IJ4eSzc
zQXcRMOsGyaMn7Zp8FN96lxO1VzJFVPM/v0N02z4cMSTr3b7Qyz6YZT0CJsaRWrl
Uf3SJyhV+ExU81oW2F+FeTorgvaC82jTmwSs2MieCIcHJQMgU+EKyakYOnSKchBs
NIzhBg9mO+o13vH2GS4mI3dockdZ8LdmKnVQ29bRsTt91XEgLTXFY355rhUDBCS4
9hHFD5KFj4IP6HtKPdXzOY9HxfskZrnGrehDpf4Lng7tqCKq8W/xpqZXZMF7nIEf
Q0qS1axdD7ZHVHc3pPAbzJCnZ8HC4XcBvDyN3PEXeEMDJ/tmnJlBtl7TWrXC5IeE
uGQUeN8XPZS77Eq3vE1XyGMg/+G0RxNRZRpEoqHoxKKl0J4JoTHXbZ4C0cs7wgLy
8SYs0KId9Iuu+9O7UD7rhM3+X5vh6AQxwTuPbK5pH8FdFK1MYc5nUcK1Tek9GBnY
CSFl79Q1cSU/D0MMQoaG2aYletpdKBkuvREzCo1wFYKbqbx1PhsMLarmGuFXW+xk
Ehk2QOVbT3cXmfS5SK4nOKW0vJUElc1ZiT2fN4/lA8V9EVlYGov4zyb9rVxUgZKZ
GrVajy7KivFIicwqat4wfeaVyeL6S5w/qZt5+KSmZVTrg5tcg/ngNzxp1AwfnCwR
z6qmo7rsXNCSgZuaE1XJTVs+IcoUQSgvMCz59miQ3+D916wl2UEoxlHq/RysX8l6
Q3qiyHLWlYUCtuPDACjdcbV8qUFoJcQDRg1N2kcPDQU20vVkE2ydFYQ74FTgMkCH
BRDMFr8Kw6muSZaByIyJ1GBvCn3ToFV8vkXGorXQMQaq3SZ/z/3WPONWnaxgMhwV
+F/R80At5hxCa2kC/SrkmdWqX127OSqe7KtjoWAdr2jxJVsgJ5H+6Ulw4Ilsto2x
ADKjFGjEwx61Z/NgmJ6H7Q8uvnx93kNGpOA1hAaDybC3Mh3reqE3NkTZOF8UYtpa
Ut38QfVtk9Gh3ge4GDEdV6gd9eV3dgrf3phVzVO5JzcUaYBRzpmEnc5OsfbISLnJ
OgTO44CB50kFrxK4sW/J8Na1SdtC6PuuRfmo0jwG8oU9OYou54BkDtiKalxF3wNi
PSmIQs8ZiaP31knCc1naYaVaCmBjd17Spp/tEuKKGwG7eAhkhGX+qfVqauM1VPif
48KY6MJnTmWeRfyh8GnZkRjpNXkGR04uyytw4Oe+BWtwvgzyCp8jyai2sx9AYP+S
qNoNpGunKZ7aINsnLIXWrhwovaAPIOYGVt0SDbJQqqAut7dXE6bCHXHj1soBe7bK
Sm5N+W6Q5BevHgpKw3ebo72ni8fxihu7hh2OQopojqMwPBH9BbrCxZjzUOQrazlJ
ES9VFgEkMWACteJ69lgwp8q0B9X72+O2jKxL4EpA9dqUqKElCN8dM43yNLd+FUUG
K4LC1bC0WDYkXBfBRa7rQ7f+yCm+DSCVDyndbho6FkM5B+TZbZbhaSIQtl1+B4BK
L2JWAtAQAnzK/flQnkob7MikLLYcZAehNsw5l6ZS7nMHQ146/z1LgWreabPKut7e
XVxHI5KN4OSlZ/cUySBIPTTe5G76ImwMzsfOrEH4LO4ksFir+YxnwYOMSWnlqFH9
bWNf17J1qlewv7FDWwS0WiQScwqB1p7C89vXVguuycr913XC5RA19yr5GYqFW6h0
DKP+5sBgJ33qjH+7Lmn8g0pCNEZawLQP3AflBuQvAQN/D+NYh6QUasBSQW1/R+4J
5GymxU6L+oU1SenOSWxQkfIz8O0ZTvSpGVB4pskxVf0Zs5sx334YQ2bb/s/nJhCt
SYgOVU5HDyDqIZ824bQklYDZNTnbqatWc7VWY4/SoClf8oJq/s8rj5mRK3HRyNbY
6Wg8vDGphXOyjSICgTKeT+j0wAkkjS227sJi2M/SonE14BeHnHKNJgQ5cozoCHa3
bUoILMbmu2M5KS8rkID9etQ62AacnlS4waYhglOByJYsPxI5fRIY15V8ulTcGXyI
fPbDcFWMk3UE5zS4UkmEi7f85POT5oNNLLE+wKGnobAsG48JcFKeNGT6pB0UUdPG
QWaemoB4MDmQMuOD9HB5hTzFodnvFf62+8x34LL8F84ReUuYWrRmr9OXHii7Xf+4
Z85PPb5JwahO1wXacj0AzuthqlVylryhRs4pzTWxdVyMHPyWVCtSlX0fv5o2eHW1
COXLYFzFMnhDHK6BqcrHRlIuR+jUws4HpsxV2OcAvbyWlJcvmtiiSkJqD9HucGUh
gx9jSlzADe8sRP09RdPryG5Kdke4BYgn5ocZvFlUwtktzGNP1175/QXvnrI5MTfQ
4SdNrNbmCR24xUovW8BLTIWv67rkgHOrmOt/o6WBZG+OBjfaB/5WW0qmCR8eGGDy
QIbOjr02GmGNBUWa35a9oFUt0SGqUapCZTF148QK5fexm3F2cmmocDfO6nzDDr7q
UtdWNQ4ftRgiYPRFW3nZyQL6+6kdeXbqRUIVM0krG/vw5OmZz0guCvyTUuNmp4jK
vRet05YfpjXBZn4/sQ+1Pga61TtnBrCBqPOgYGU5aZYuDUaOim5ESjb3Tqf1aQ5q
xgN3rjHCHyIV+iByYeC0+ljFU8gYhF5wGYsZFMy/LIRpts+2RJCuH+tCCaznPSXK
wWYIs/dzXUWhpkfSD4ElvydsZ74LZmQf03e0f2qfNJm1a0RaG1AS7VdwzFe5RCyJ
StR7oWcqJ0Pl46McWgia+js5dGXKAE8YhO6gXAq41qpeC/B2TyHIp8nwqU4gXFgO
p8e8TFlkGhJY/PM5sG/s9Uukstglngaz5HnTBE1Qlwk8XR/MIbhGtbSeQTCHSNeu
5zpJIthCm9SbF/8vtg7Lu2IZXyodt6TC1hMW7sZQeq/IgcNcqVXpxgP4vMA/2bWo
n+FIDTAeztW5v0oW2ekwdLJnJJpupSUHUn6Wnx2f5bDcjlu5+rr31HlGxUfYukZA
WGGEJLHkzdmc5HzpWX1wvCWfFRuFcEWlXeGDzK+1YKhm6SgOweP/Y86q5ArO0p62
w9g93fOWgsvDNWWOfrC56BybVmW0CkeZf7EoyP8812VFAC2NALlF7yuu6BNWZ7+Y
JwZlDteCS6JPAk1tsow8MEH3KhXYZypCncvIUL94gISdAdceo38FcQ4jrmamojCT
zdm8faBoJHyyyavXKjDiOuDLHFRnwAw25rMFL5JuYzFf+Vul/yPjMthxMTUBf6Y6
zeb5Sg/S+r3mWui8b7rR9CNuyxhfd6lh7OQCmvmB/qqdTCjiHK643PN9Ru8a8Ewx
2yWbard0rt4b+O1eU4/PAXn2nzecS8Eag3Y5sm3aADMeSsFlQ/P5p+MhPFmCMMDJ
hsQhgkQ9Q+N42LfKJ8w4mfT8bUFl7xK3AqjrN5EcmlBc5O+hNGkB7Kzlb79Zs3a7
x1uKCFtgHVWZGRFvdm0ZK/Bjjx8vuDrKXkklAv1aPGQplmrvKHhGGDjeNAM8C7ff
qh3+TZGoF3FVK7XqSbeXFoMQsd62UljCcOR1NhNhvFWbvN4gWDRF4VzvsTmlYDFX
4hix2oZ1PzFSvmrR6rpHKIQfqRPIyYgZpn5YeOswZidIqoSrJg51iK4ITO71sMvh
4DaBO9yxzuNsUY8Z+7rloNvn2fzEH1vEddAjktl4iuWJkbeL0YawcTxzaMQ4g1iq
XuYr/cx1IlwCPpyflcMpXD2G4qz1Rg991KAkaHGNToze8O2ZVAzHnVx6nVFSUVOG
5O+1ic6w34PWGeRbTJlXpefBYiLARscyLlwDLuQwklD5UbzWuc8ijDUPrqgB/hRK
XXmCa8wt/4RUJ0R+XPD3On2OfDXAX2OlSC7NZK4+rZ9r7JRVi74U7PM0qrtBhb/V
uqkzLj2HHB/mmxeJNg24VjSFaUcgf/Nm1o7/D84QFzfhJJ77rXL4x1SOPw0XPWw0
Qer86nm8v8T1lmohc6wiIQKKbSvj93dVCeRPRWTh7OZQzdMydOW2wfUauuw6/37I
d/7c91QKtlPt8GBz2MjGb4eTab/dhB4BDm/SHaKtEZPTD84iK15UHSsLzN3LtUA3
p5Lq3IMQX5K58FxSZ9gLmuvv5i0M27W9+bS9fFlNwCi44T+Nugh8j1hVa3TOvfPo
7b4OMSvqi3ut/mn8ITmNvyu5n3NkVKR1UbfQ5skLgIdRFotdJRgoQYLOCFUcABrj
LLclomX5u0BfIHGa6zXWol4e+0buIKnJgvM7IjWEtwlADGS6Pj2hHsVY7jcpWp+P
WMvAR3UHzHkpFE8T/7sYGQheeCtlKi1VfygjvWFEPZHcY3YfdUxPdkTwy4I72E07
vhYfI2dctPaj/5Zg2GNUujyI6wqYaqoz7sxSlTj/oA8yJbHBTQ6eEYRkILG3ZYfi
mJzoAqkO75RagxGJYBFqM9UFUDyNy+6TiQ00fMNkcFUAhEJ+N4NPQt3+AQmg1Kp9
Y9FbE+zm91icDFDtOgmrAfW0XH8b9QS971AMbmzJK1BYd/R66+X5XMuGyCWYGkTU
YUEuBD0GtSBvpe8KIKPM3iImSErBEBjEOUEtW2zKd3buPmxFYzpRl0MNcHDFZGxg
kPewp0Cp6Z0jwWAb1oHui7HdlxufjTKpwZBJzr/kjaxiFzl9iLZNOsHcTninDVWv
GawMesz36PAIFTzbzdSjFDdOxQT33jqBcOIBwUsPAGTQa0XWuJrC3g27OAahKi/F
fXSz0dsLODQ37DWBpcjhkLZnXf39oS5KFJXOpNd1z7221ume7g16wStm7nZ+LKl/
F+mAjfkFdEyJJ4zllbppOn+eeOcux5dLyoBhzo1Y/TJBUV9LAV/BuHzPLEaYjYVj
4H6QPdFq3qFywb6CPFXkM5vfmEUuxoyhByzQ7jYzBSqQod9Rs4kh2bDQM3B0BkQ5
26tvaGvj54006+4FD1GfTvZaYAzJ8X2kHOqYI/cuukULbVIA5xrjsg/PHhdLnZZH
Ny9pszS7h5GEtW2Csm19h+a54y7ELvbwD3p09pk/TbtesFJnMdebr7OTc0sWzbHA
PvkbOEYqprn1Hyro20yiGlcXOwqdRAo+97Hp5iffLeGDtZtE26z622TOQEieEF03
VkHen6YIVWGSUzqNFI5TXhbpwwm/IsYDUdfYEshibVcfMblRec4YozGh8M6gGhfB
6si0zIhuGpFgWPsosZ8B1eeAjoj/BMnIuCuvMK4r+6gs/oh7/eRcTOZjVJl/RS7K
F6TPEon7p/U7FUxMYEOFlIMgSwjrfiJntNloxQRM3HvfjXA/nCJmqqeFQjwQZ67d
NJk7f7E5lXB+GNoQsUPUG/SDGwxNCUnT1rfnw1ewPoIMiYmUQUiQo9MBIZ/hoW0k
A4TQTR4jeBYFZzNWB2z0cGgMlAmdzLp6ockNY4VJTdCraDOi6d7wcpmeUvXj0SzE
8WShy/SbRi3joYKPWAOqtSaPgYIjmuVXmYquSHwqodJsAYXLmsMpdOW2rIzp72Dl
l9tYWiM7dXwDxZjOjNVil+G4sqj3aLhSucIImcSKDWAvRfKem5SFCswprnZLa+rw
33O6bvdeIqjwn5dNZkwGly+KTbn9rhPW0r2Ku1VeUYe6i8YmqxQkO6xedmwCoMxt
+FSLXPBI9/XHvpF9GiCom35pWRTwBhe1ZSrGnaJM0dSAHfuLioG/hpLaFEnlTP/C
fRGoHk+flGQ52Jd0HRfQ+95kEMo4/cVEIP19t/Zs9DpkK0dzaPSejjZuLWYWN+Qm
Kygn5YLwjRgLNKOO/3gvXDk62pjEYXyz7neNhfgJna73TWasIrVwizOrmQhXjZ5O
13pVpOBtScAetWVsZZpoDiOoMB8RFuthHb3alee5dY1bWsZSH9Eh4GPpwLRNhtuU
T6EqQ2Xjnfxm6anddjjuZKog5z3vWkTbNLQtqTUuiIs16jC/TegiBVI3QZtzxzva
Kuz+2wqWmiveVu1yhYIMFbBWaSDBbKKfsZWC7ISIQWTiCuTpHCbSS/nnzBc1p+hY
+sTxD3W4lzlB0PpuKD4375nSi3i9S8EEOw6V5Ecevmqb0ehGETBOQA9Vjekfk0+z
X6Mw/r6N4qe2C6OfNT6bLGiQUwVA1VWQlsIvtq+Y3CImsWvxiYvmgymoDu1U4ul8
rsjiQljaq5QwciG2rOeVqMcTzePDNWJ47kegpCXFT4dN90V9F1kUKzm8TV9V0NEK
77nwzW7rEyXj8S7lLepyBqkJojx0dLLcJAs8z90GDvxZAgKvD0b3d/QVCzfaxGoV
SRgiy7fU050mCVx7SQ7sJjBBiP34Z2RriVAJZ0rj4clMWAVz49hojcwaim+gErjm
wznJQ4iTcI2Sji+g4PlMNoyR7K/2c5dxrnCTvn1AUbKeY2KXrUFOktAuPoMDWX2t
Cw+7yfnIwiy1L2+daV43ZSLCPgRgt1jXglBh17DjYw8VUXjuGAje4FpR5MG8SamQ
XhhQs9TtF3rHA8h8hevBBj4P3LpoWAd6YvJ0WCnHRZ6g2Si2nOp/zjuoysJEroq5
4xEn42shGNjiPlGNhnYILFdH4Gasu6X5YslBEvy65/HMoL/X2GASAlLHmYmJSkGP
tvSfj+Jm3zEP5iBaY5TUdzxY9GkrWvPJiNhFxTKfW5l6WxvIgDIjt1ackGcWKCjb
wAgf9iHq+Mjc77vSvhZJSwvE4/Z94BOhBH51zGGbEKju2/BfKVxUGXFxcTshYsh+
9dkk/u+mw5bh8w9jdd5ztGU/RwxhrOdVEV5wxQmqhTbxQUrlkxFfPt3TOLmYaYZG
+GHOGWEtEyr+d71n2eChoGVpFFtd5q0HhP7oKnKlIWTRsxujrPebPkqKERgDJiwb
VKndiVRafmII7pJx7LzQheH+WE2WxNOpQsf9j7GUOJKIlLHAMGfwddkJpw+3sqdK
FtXcSp+45Eqw3wAkkm8wy2k/CkSWd5eWiIckHV32jH7NJFW82BGhAZ3ARItyz1IJ
fnKGD4OVGezj8Qw8fduht8FYSfhcAFOWJ2L4F54WGMBp62yn+zXwwVAmi8LxzXgp
Qli92/in09wrq+xSOaWPSrv0r3mi6GolaNVkYedNdUQ2h7VFOuWynedAPuEoryjy
gPtTY14+MXKpHZezsIp9dVaOjcslcNIgYEl21iZ/qd73LnhJOUEt+VjrKrxThXim
CZb8tB09x68ERnajsQrEY4saZZ2A87CscxB6WHEOESW1NxMeb43SyQ31SrNO5lJZ
CtltdRFjD8gBVYxZmpQhjtioTQTjE4O0OwjF4NWvmNLkze5an9tQd9vaeB67b9+D
FxgsmZmGDAV+FDMd4E9qvEfvEFxnkWtQeMR0YqFGbQIN9N9Bm/Ku/dzlihc5phO3
Lj2MQpmXb3UhnqX051MCu2m0HN0aLma18dQYyAi0KxTQKNz8qS+unQiFJ1jLcU0Z
pXnYnVB9vw/oRlF9lIU6CPcTpzK0BN3HeJ38RwCMODCeh9wF98Con4MYxfKyHvkb
Re+7bEx1qS0IguLUlsd7/IV1/LB+RVbMfXZUIsjR3I/ReQpAtSrytFNH95wWv9ND
BLybejNoP2jCPxP/553p+E9O3V9tbJTjyDXTmfXJjK1Ur6wrbYSDfKNofgTnFRSN
MC43dOX/zQm6hCAh/eMWDwE27i1GxAZo3XKlvwHXxRBVtRiSjDdtIbjQPVuW/6HZ
15GZ2pfBiDUPK+HhMSCeYTaoAlYCGVshiCCybNAtICOsEdYYh2GrxIaXSbU2C7a3
8l9MIpd8TiNHHW3g22rf2VhaKHXfqQ6yufw4LPsI+6Kx7o9VYbcHo7GVhpiSsoxU
UHN8o1uRlQCD48lwGiS/i5zfWwDBCtszI+rzIK0X7pk2C72yE2mhZfEvmPf+nrxd
HRbviHXDOEwhNC5jsYsAEnKut0fJxakW2MLxe6KmnBaLRCsEMbinjaSDRJeXiMmz
LWihltJoZnra7w4kBPdzkjSFBTf9yYRqVukHo2wJfjbKzyK1KcFYEfJpDNBb87Aj
RnmsCXfflgJDq9WYQQUO3Bx0FMN/P3dai3QIOKpsA2cAj7n24YmH/IcSpSV4B+Q/
IxawHNzOPpSzmCHLSC6CGbFzGnhq+DH6/VzIoggKJO5u76kVJoT2SNb5CEHrFYNK
TdZ+oq3Iq2PtD2IJ4xSxmtwCS6miInoUXe/Rmk6aSet2G8SO/wZVwNJ+9zvpVHSK
mPrqHWBOHYhThmBF8PJ1EqeaoyGJYEFXu3t1/uk+jvkzsKqzm8GVUTzAbxAP70RI
dG+YW+47dW0OXKQWa4zN5zU7GyEKtRj3/+37qHhF3de3jDKbSCCmyrnbiJIcp9j3
KfEzRCT/Xa8x/xg/M38j/pfI2Aa8FhXbJIllA/3+qH4ptuMI5UJ+8rnALVxjBVz7
eKxERLcBW4Oc4Cgh5OmjdNjjQzOZlSZTljpfk5bN86djDcpQ3D1zmSj6osHWMdZ1
MhygW428903Hlyx4I+Ee4HR7GSClazr9avI8RzINY1Xy7ZAerFU2sgWEw8Uu024t
gKd8bbtE5Y1vegE1mduqLxl4k0acKzKGkNqxtnTs98/RlZCvs/RBcLtqCdxqXmM1
uj7NXoOLkEaOiwQQZEAC/X+lkgfIpFKLXosfhL51IIHqST7rt4p8UR6qC0bbYp+r
bntiFVH74wtfqz7TvXY0LZ7toD7Kt77536zU+0/ktNYnf2tN14OWGKrAxUMFwvZy
SUL0bfBvIfIND3XAjNpPKhC0RR8KoXjmEuYFcv1WwBvoPiyapiW1ZzpPtpfxekLW
Ahl/S87rsUrLf3tHe5j1u51tI4n5dCGxgJYTzJMXwru8zvVaL5RZSR+rZiGp8InX
D6Bfcfp8gmrDLR4xZQk4WVjGJBav9TTp4uh9VAVLb1GKQATmhKH689m4XPusZnhY
WJeTbRDxyVQrZRxY2JY/xrBjmbJNqYAMS+Mp2mten2nMtzlx+uEbtJuXaWlAqZs+
/K9kccb4VO56MHFkJ9nPR1TU4bNsuaR0e63xKri5U7yl8VkVAAYQfukSJqZwV5Mb
msLuLgvh0THBjqqDnFPiEv1i8QO4AZOG0qws88nKhWqBmoOWtMSpHFdNAGr690ia
r5+/CxkZEOKPXAN9DQ3/nrtM3+4jryLuUeMm93f0Bf8yEtgQGFpjMJZCPVqjFE5j
DYVpda5LRBlZ4ZvesxMwalWUZy+U5uDWssxz/fL8wh2hwe+LzH+wVklcEh5tpHaX
X6x3z3NF/8F3Ff0PvjR9mj6X3yQAmj+4VM2FzjC7s/RYyWDkqShvNgTFuXzy3Ahv
boxim1MIun2HcK7lNbMrV+ARV94UMnd1hVmZJSuhcpj0UCkrk85RvsBzaTRfI/s/
gcomH7NS2thk9B4Em18vuww4uxdfsiDoxB7DBUHulgoBeGrDrfwWyerbvvLhL1al
4PV9Ss/gEkKqY7m59EBg+KPeg3Zk7XACHtR7/egTC6kxrOKjQxM2xPNHW3QT8juz
wo3LVTl1/LEDqyVr8bUhLCAYJnoqkOH/tiHSNQ3zB8/Hq1pSlrZjQMmGluNdusel
kMmQccroM7WXY1+4tL7MfR0KUMkE4SHdhTh+fgHgxd+h/t9em6c0ZFe0EVPmIU7X
o73vmkI4mceirGXqx5sXEVc0V+leFi5jW/7i2+ai0kioykQ3aQ97PJhPptxg8wXq
Ep8PfiCRIQgnG8D/Ubr5c9gpTk3WS5WJMv+ytSiBFqqUvoXirKiL/8ygr79SHx4F
TYKIW3axkefn9zpylU6JHQyBISKBcBalVlZmv7YhD8J6VRHjmP6iCoP4PQ1wI8Oj
GPufSA3iRHRxSUkE/4WtD/MzT8wMPCax4hkq3lTr629HKMX4DlFA+MtVV6K/UzbO
jGx+1FZScpvVgE79STfhZy1yBCXa0plGgPjzt4asP4W2F46dkOdiShtbQ4N4w7jP
AH83mQGXOSKRtRB3fdxES49wQyz6ZkZ/uNA6L+7Ozuu4H2iC8VG83EKVRf78KrLK
UPYaSb1mSiDdZ3iPh3KltRA8n9fzs77Gcwp0xFBAj8+XnxfUjNWZzj8al7N8HZrW
wb/IarC0hhFP9VY4VJNlJURhNcEyq5+FjwGnq+arg0tXXXmpbrUnR+SjIFUBVvy0
04fF5OTmVYdrfg2biBA7xN42BFM370dkM9anKsuUr3Oi/El8c3h0I0ptCzdh2DBr
f5W45V7pQLLFOTs91ppRNNGgZ95cSRTKdAnC4s4h0yFjWx5lIoFc3HS+T8eR627m
L5YU6q7SQ9tTnryIMMGNNzvwcmRHzBWkDW2gaB8uQPFENGXJpSGzNvvSEpitzvDx
F8EXvTD8qVxL+sTUJOfTZqht5faKv8WuA+Cu+Us5/4CWOQlYbZxh8bU7MsvxKGyl
C3x7j9TYn6dHi3Iz0nCQzHz4Tn6SzTH5L94jVIH5scLmGyx8YBpBBwp/kg/bBdSu
IANGgOt7katFAo5pB39adUnUpu6KMCQF9JQdIUrz8+t81ew4ZF1Wr3boKGN21WrZ
yWNGG0hpMZZJgwMZcSLtu1KPEKyFUP/xOqjEFxISTj+d1X2gabR8n0H0PPHtV1tf
HTU4OSxVtqw/EiQ2tb7aGLqh/7VoC6ksuqDG+/Jnt7brsGOGYnaY+9A2bACXbgOc
6J54tvp5JXWxvq9xoiJSC1qgdyEchwf63bPejId6cz80i9f6vxuzLIx8fc2bFi9R
A/aINiSwr+h8ZIEjoAhoB2FM4OqDHCQ9FCX0w3iUKCzG90n0UdZf7wI7DEQvP0sF
nTrnLAUbLkL9L3tpKCzAjUNpx117g2HbpCVx/gvUWGnh/gjS2rMh7ZUT6To6fKT0
4U/kOXmnE1HrxN5P2enyQ6tAMh5IKVFgdpeH1PHNOMgrpyxEgBR1tpG690oHqPEp
HXz8xu2ImuTMAXe97rj7DMrvJCl/6ZQHACAVQDDCg76C0qU7d70Vo7WEe5sx6yZp
2dYO8lAVK3Gf0OcVvbR65UiMakxMqnd1z99doO0jaSs57EnF6Et0kBGQZb/0ZJb9
CPMXLWYWZqRk53+r5WM4SYVSLfYyYTf8PqfB4q2b5sAdLgLv0sQRhTKQ0L/kUM0+
NBgYMGBtcnXgzVSbVREekaXczAEtsJvBsf7GiiVgapGKV9Fh3qxfgiIX94Agh9zC
GjlNRd7k4B0cUE0VXusRKoJ7+/9qiC7NYVi+r70sZcgEfqphlJ9jMVOvjgUV9YdJ
9OG0Xo4qnbnuSdqaV8A7tJ6shywVSCFw9gP765TuFlV15qC6I3egwj7OVghWUKuG
ojJTjnSJTunhXAg7hGdvpDj82Qs95MvxDcl7jtSx0/3m9OTXdfSC56QlFaIr05Bu
HOo20bVzztgM9EWMOUYlGskkMyOidUGdfauuX5J67zU3cMGrg1nQWcgP1eTb2S8S
2DNlPufbSB2cbiqSle2pB4wq4i4yx0iJ64DRKuaVf72V9PXON5Ntbke1Illk6DEa
Lp6naCKRCuEgS0olh+Cf61ZF2gkr31B72voYqnSLbeHDlietyQnmBrKMya4nxtdt
X4+7tQHyit9taHJB8aCIhHPtH8mP9fOp8nm8kcm6PIiXfhDRQUR1vHGB+vEblmoi
BbYhGScVAWv1kEc7O07iTJpdTQe/DC57o+Y/hHEicq0stPJ6bgzKq5Ppe8J/mejA
aKzn5sY/gU9sxwIvbzeoXKJD5Bv67eoWT/+o7H9hMdJPzI0Wto+PSUnxyELmk5y2
5ysiMnz7igC/h5qcpuxekBL6mR7FEq4/LtlT2X/xnLyCHldrPKMX90frLKEYRIwn
syD3KEHbWT11X8FzJb91PqT+kM2DaBHcqEzm38L6jqQQ6LSJEHCYY5BWXTL/WFKi
l15VElcQMQXjPHcn3JrSKdTd8V0AzPOopJdYH2A4G6XfAbtP7Idyd92srz7Rc8TI
Jyw2LoR8qXjJNw931vtuGy2wlcMg/tVi5BD0XXjSSHY1DxJ4jFfGX/OOmYzed2/4
GcpmwOZgma7FV+xWJSEIYUl2jnZcWxsoGfGZbUQH2Lz5es6YphZQx409FbMbfiLy
6nJOYUevlc0PuVEhVy9zC2Yd+NSmI93vAVrqm/Mt4dsf9qtBxLctv7qMo/AO0MZm
rhjwraODYqm0lG0LksZKx/O/P1Jw6xWb7QBFmcBrCWvhBUbHgtMGgpyYPkRRCvc3
w5GK+dCkIhN+YfWKI4eswtgibKDYbGy7ubck2HGwnRLhN1HWCFAMDIDxlKbXpErR
CLfDHqmw7h2GQLTpnpBBHOq8M4MDjUB4WJA2GBvU5iT4PwRi2SdEbcksv8nkPSLx
PVyCBr0Uh30JAIk+3B1p8l6PDL47tGAkuqJrsf7S7EXQE+Son72a+4jqTgb+T/EL
Usk8BbcHNm+12E8wVB4dRH9NDxDgwQjlafi6lYAkIqv7PDo1IVg5YOxwxT3Arztv
7ANjWnh5mD8fjb1jBT/ksTy1RVSqcFul9YVAzjMukWzlZzj+tTlUJBkGZGfSqkh7
U10aQ1xuFkqxQlx45+gvcxH9DUdlVcKdeCkJjet2GBrc8ArmzQWfMezJbJQ9p6GN
CDGd/tyDVVoIWxk2tCD92U95Vf7/HwDnCVLwzxhje3ITVfG+4l62HoNfjfXVp99/
Ti7DtCaKosn9gjlfI8P3R/vslwHSz5j+YnpcRN+Dz3sEMlitLas5vIR5DcTSpHRn
S8cx2HQVCmlUOSBAWIUu8kV686KjKxEsjdRSQXPng6GXbGGkLmDyXIgMYYlBPaR2
vUWF6vKqW0Zjr3qADu3Ogvc09rFOj3REwzerLWnDiby6khP5n6bYT0pfZLUc+QRF
gMIHgymizuU+eMQTTf0WDIyKaGBGfn0Rq+YUjbCnwb/kAaP1yI0a9lbaVUpQPo1K
TaNptjWUY5CB2zSNUWLToIxybfk11l4O+YQTEqlNyOg7GTUbXZB6wgJIruwVa095
NOnFDzrNQOt3w6/h+EQBFJtiEkIlAE6Nu/4NBFLlYr9184sH05eQpYIP1eqNuvNV
FZ7w1uo1BamRPX8J7Gh/yR18l9NlIfnsQQ82Zl5DtMo8pRhZZpS0OWebxfeCHgC7
LuIhM/Y0lUOygdZNnBaS3flts+4+Cdnnbfes9nTI7rrD4FcHkp6F/MhOD+sr09RO
FXcSzx5Dl2ZkqCggu51r4vLxtStr2hXJtaXzSMI+wprzZcx3+f8WGDPvpFIa15Pc
c7ihDkHcOR85fNSEPRAkg6alJl2JrM+FvrTOcMmWayCp0rJgIBr89eYGAPEjaMlY
9EUBiD0WjLcS4UaORrRAgjpHJRbam51lrZTK/Kpf+tJMnPrkoeqd9ZIWqQxqjzTE
x0fp3Th/o7SyuvqK2XYTCiP/+KH3TXWzLKmdkUNN3b/zfe+TRatYR9gdNEfcCM3x
Vuvrs2/rQ97JgHk/ZmnYC0LImVr9KTNFu79SXxC5EUt5y1qb7HqDWwqchLDHIvuj
ijEGYMk/FaEiP8w1b2W4GN+hM5JV4hJrzUIaXqOeETqhisvbGK+cfO0rZ8Q/LmrW
x+c3fqtxuFDDD7vchzuQzx5xKHOVxQafTdM/ZZaHWoDQiAh1MBHUeiP34PUbXMzm
gBSvTqH5bwOmi0vk/TrhBa+7S/ZI50keEOlH0Zf34NIRj86838BS5lLUcqyngth+
bANBr5R2w2Qn2SZUbKsonOGmA6KTKAg5LBqHDIbsNaMbwvetMIsAFrwDw//qlQms
/7fcYys4/o0HAwg0ERYHPBdB2cNWgGHt4cs1r50S776nwt4szFEhy5g0pV0s1d/i
hb2F1qmZaGgpd7Cl7Z0HxDa3Ehd0XrltEyamFpyTtV/HfICvWNd/H7BEONH6KCXt
ugwcIeSyAhLV4X+kUFLGKKQWQjNMfcmZmn8gwREkveREPZRRXedV/IQrET75Nbrx
BUdpzdN7iEgyS3Dda6iF2BqWYxEhjMpiIIsEaJ3mqxoYymK6w9M48tqec3pVq8Pm
OwlMvXrDQZ6EM6ezuUMUWp+GYTiZxjQg6u76CbILVjlX0Kcrtj8dbt5Ouywj7cFQ
5WI2r4WwEFCFg+L6InCJJn8DtEjjUE2inW2RAuPP245YjeGNMuwi8m59JqVpR5CO
DXWlJdjKVnxr24VdwmZhRdBmL4g1Xnot4H55A7H49lG6ZKBB9ThyjitQzMncnkpi
zhuU3NFm0E80wdRKBFEJlM3CiR7JnwzIlgUCzNU+uOkvNDj77iQdLbC/ElKpTbQB
Vk9hN/UHEU2zPBd9lXk+qZh6iu7S/e3UtKnPzHXgFhZXanAahEvfOqDcBx2erqzS
mcMd0p4VhArr2oXBe3gnDeEjykqoJ5A0ZPQSrbTkxRKYkwnvNLmZoAD31AHNXTE4
rbqSrPCQY4CIzbUSFgksfY2/2wmcRoEBJwe+NNviOX71XIOVGzTBbrIkCQxTUr6m
pzYiPbh2HWsS63NTfFSjD0B9jg2HOIemNDf6KkpbmP8+/iB+S8xqprRX0/jB3yW1
sdN+tUqUws0UvklQ7vcVx0FckDJjl+Fhc29CXTNGjVDrZNqT+URFvU0kwXXxl7av
rKx4rh6eo2QR12fD4fsX3y4ySZy6oSf+v81PV1jHwc0l6hEKcrceWLRoqQmMmbS/
Q6ouRNDdeQbZibrJPK2R3WAk7pBdIj2HiYtcPqRxlsnsu0r1eZT03QAUWD/BgoUC
CgGxmkE8r0+yfAqv4E9hNbYIE5dMb+RFbL+AOYEdFyMkmILCl9vQ5KRvPPywSoc8
e1U8+ooCuOGfptmBfPoGLAG1yrfiCgoudTpq7GMPnKWQPp/mS3wgBbaJI3wwzzsZ
Jgwyc4/tepcja3ku+R3QKO2CsWkriIDKJvIFHraAUVibTkkAit71GK3B1t4ngUq5
GhMarb5XZvNfs/IJQpm/kdMuadEsSChdwpIoJY85u+iU0paoWhR1h6PNCIUK+QK/
mYNstJQ0mE4b4UP3qAl692nyz0nW4H4R9OrlcCSKRtuge8pGsafXV8qCi48BbboO
GSHyyRtm8BgeF0Sn31slbuIlN2QOI4U0Fb9DmGVsD1Bt/pX7pao4lV9I8lOwAUSm
IcWQugjAORiaTe+gI2Drxntcqy/GBAgb41fZuBzD0u2mKUSdmOaJPcMTc5K++vkS
p+1DnFC2UKX/Q/z4PB2+XGerDQFgcX7P63nGWykQHxN8H1DuttBD+E1St/NLa4vj
Z0LgZdwAQG/hQI7S/7dCllv+HFCIOlRBUsRAkTSxfrCUPFKCjNnSc/c20TpvQq7S
GAs3paVw/YEmanQnX3qHKUrw+D59TUp9ayf/fkwcJtRiaxiU7yGuJrQige/+Flvg
UvEwc0X3ui5z1PzRoTbEQJnuZaA2GOFWu151KMc6PMS5WTxcPYb2vnUIt06qT/AE
GDOnH1lo4jAgjAycFho+hgt8e89498ZpABGRxrurv5hPaM4A/EGR1kKschuAm/u7
Z3hNNhIruu2PHQU0T1Ou/2SdYq3yfePOUs0p3xFGmA9LI81b/unex9qDsTKS2wi2
1WvKS+UUenjgsgEr/7HjOh/2eRyV4/9PsV0u6dkig1UB+qiccBdXp6HMkh0bXsHS
0mHiCYsdea5nXj6aEFcX09Eyylzng4qKcOcW7HLvysTCrSYX+RADP0uGtMFj8k5G
98JC7tz/Q6O2mlAVRbdBkgtlqsMudjAj0zXKWW1c9RUCf0h2AftzVecJfthAZz/3
3jLrVVfeWtdrkUfz+hyMV0cBtHdjsQM4hk6l56JRlCemcOnKwzso+ZKFCn2DIx2l
373abt9XeE4mY4RDx+OdDqb2hQmplr1NH1d+E9Xt5JbW6ZrUyTPGUmxjVehcalAM
cwWbBGTExchzRrMnEXbNyLhUy5AgdkjABSXjcdGGmU13gzmoFh3oiKVOusPdVss+
dIm/Oj6RDA5v4GOQKSqknqBFSyLOdRsgPIhxgRKgNyj0bto40eCu85VGy7m7U0g5
IazfOb6/Jpab/4lTk2yLR57VYh0HI5G3pqvCYyWhOXP5aThU7KgMw6LMtdEW/hFf
Z2PJq3+9UcHDEJ5wy5lwWJlDDFdfzChtYQlEJtSHz9zoAV8d9PUB6y/BiSDCGg/2
VfyTpM1V03+OZ/mAXvX6fpDzovRgMh92MFcygut+tw1lK2wfxJ7nv/3o4fUQMYHO
JE75/3D+nrGSfMBmIWOjDdyrkGWe1aUab4NhfqNobhMVTx9BmihZ+JlVm61whoxL
VDJ9bh7nI+zUDEDSSYmfR2+9qtdgeFer4rrMMQljT2rI0ZPKvXBN/YSZs5wEUf0g
Qex1diVIUDP9ZtXDd4buhOmw0DNl58DAFMaEcG3AXm5JC70fakyy3iHQQM0m3SHt
QhvkXEiC1DIcmd9MUStzKfgFHrhtW4Co1BDx++NnEaosl9HWqH7hSLfc08HZxoW9
hCX/Gh9z6Dj6Hho1fgG4QA2jj8eJSEDPlE92CVSns93ucpzkWltRPz2JpOB7SUp9
XJZJ2MV8BSOo1dTMioTDNYcrYn1ERSnF1el0Cgxvya8lrhkup3jTnCirF4mV63+j
T4BfYJqg0ZXPcekxOBW6DUk8VtnR+jD49pXiPwa5VVsSthjWD0HO7KdvR4QEbwse
C8kuWTo44u8XE/uhRavalHKRLXJmhmmYaO282uo5qiTR65+MQuKMDwEKl2YafiLZ
q1oJEqkCIb/maz56T8fjJIhWWTgg4PfSQIICFxFRxVoRKFkRnm09cHwHYRExfRn2
L2VtrfkeAhpNuJnUolXYZsXu34qvXaiKzBje+6CnpHMEjXd/xAC64DogUa6lJXkt
WPAYwgcFIcbxlJ4xuF64SXa8ZUBBrw6AuAWvory6OF4HjdRyghTW5aH3LMFzRZuT
OKasaIn4Orz6mJmSuoHmZdnBAV89uKOdHJDFt6CIRC0y9HmHGhWe6IJPbxAV8H/I
lkHOueVaY9eAT6Tcg1XCGE3SKI1bXeOOPlkJUTohQwxYCU3/qYjYjk+aTIm2cchr
zIG+/jsSVh47a84/6HL23iDm0erDmpYldlBDSfIQNVjnimH0ljD3IrJoFL5rAmr6
NHZx9a1BtMA3O4KbbUw5uJPTaoTeSm/41V+k4/1/K079c5hXPPJ9tL9J4a5iVNnW
dD0YUJarvGahO9bSKVN0u8NGcZY3ckg2Z2cB1sGDdfunaSOdA5aPsEiwEfuJVqrL
hDr5P5caAvNJPl7gWBaR0f6vZfbMElEvaodhT6OfM0yc+HCa9EnotkGgFKt6p6m8
tVle2dokUnw/lLQqVg6HjADt6g6ls5+TpbcK6a97pzGaWmrXGylgSrWbhFSky1vA
mpC38m7gnJIsTkcXT8pTuk4JAUv6oWqpy1vw6njGRJkDWXrXvVoLrfqyXJZGRuz4
M9NgJE0aKN7KkQ11rlu8wH/GfDySrisWwDG+fDM4MlpEUblENk/I01SQ2SEQ0hqt
LdLK7UdKPPP+C4/4e5vkwl6JfdpwS27gIbl1vjLljWVkbR4NMP9/1ZwMtFkZtasH
dXkPXeNBfgmQs/pASdcuTkoJzwsN+tUdXTYG3VbEi7bRBR+LHw+Z82kn2IJrL3C4
31wG1pl50UfkAWYA2xQ3mx+vcHr5jkq5yVqUzn8sa2u3C/VZ/dA7VGtaFKVCOKog
aldenB9dZyiORL+wDqDIEvrtPcicFiFMIzlsqVWf0Q7NA6O+FmwYpzC62nE+G+Rs
kezCYqKyGDNo22/uyDUbo8BTsVAz0oJcCbxnlWTbDK2v9LbcLf9mBHTBTi2YJqfS
bVwSWZbNirBoAXC9Zb5YpLJ5dxC5wDfp8SwN9K5/k1J0TuK9qD8zNKVJQZa/gGaT
QrRCbbohG9r6tFUOmYAqREzb1lpBGpdW1apAkBbVfHFHoh98mxee7M1b1lswTayI
/uSFiUEfY6EZefuHQDYncs0pZwv22f66Zd7Jf2INlxAaGGHm6t/Fmf90S7iaEkE5
n/4H4bIxU8ahs/Bs3bhBNl0aJ7O15dP9l5kxzmkCXagn9m3Q9/bEJzVO08m10DrP
6gn7PIEPUb3II2pJ6SsDFlfXvVYzzVLbpejs9W0lI6z4RuJiOjT2+JjcQUtC5cKV
MAsj7rEOFbHzWK1XSxTFopYVJ33uETS7Oq1jSKt9A//YohI3ELl0OXsgzobLy5pP
ck/FTiVPlH+zMoravQ7n/8976MvAPk6i33KpLtkyhWC+93/HwZrjEen7hz8rysMd
BAti9IhQP7KfsUytbpYFepZOuqXGCzNWaueVEiq+TYc1MkPlrqhONGx/s7QYexeX
/rD5QzXQsfeSwofc4ipOxn3472/F27bfD7fqMddflq14LFysL6UbxHg3mEoUrb5B
MXbO0e+JZPHpL0rJAKjck6dZK90UU98mMPRgECLCLQG4Gf2ytZ86AmjxXSlNKIt3
diQpOd5oDdT/UJh4/IfYOjObIao6S5ElcT3qoMnPE8hvIWfsmx14iUpt8n5dui+l
Z6nv6IKPVT8bf3g+Q8Zy8wCHAILw6V/eJg60UawZE0diQcfwRJ1kZu/PgHiM3yOa
FsZSzSPkEi+XwCisg3+ertWCwWJSFx7vTC8ksb7frai/1Ft4v5jbFDCuXCFqco0y
k72dXqTSDnkL2BQTpFP9AG7jbeIsDgowOPzLT6owbCK9ttkqn3BtNYZZXXYkoLAw
w/rvd3vpWyttWfjxnylz0LaK53eSPfqLz/QotlrSbb34DJlfdsSmGgUBrV/vt4m/
KGoSSkOLrNaWMnrMqTDguH4YM+Z7XGdq3gT4wvTvZEu48yMXL1LXPDVG4Uvo8IqM
fT+HQnXioZiG048yJRolCOnd7fH+/zfVlC9AtxB42M+qYcwCgicV1HO2Nb3b9k8V
R4FB/kj+a4tjDG8LtCoDpG+PdVxFM5knXhh9MhDIimQUX0cFyktDnvmd0h7cNtIy
+0p8IxpageTyFtVKfuKfLjJOAI9oXvK7ZGh7lJ9CvhXHtc694egaTFUsJB33AbsD
4TXWIJ/0RZY4PBFrBq+vefrYVWhcO2EyiaEXh4E/9E5rAn/MOmxb93a5mqa/3kbO
ktRGMIT9r7TqCW1J1clQKPm1jzT63eYjDd+jSt6CBB+9NJPSdvW/E+QgE/A3C4zr
wDpYoA8H0Ft/eDsEHD2dWL6OsjjGE9JNgKyZkUHenyTK0w9KMXnjJKdoDNcZodpD
W2RsGtIgSbZLj1LFSol9xgKfrhmaV/5tormzjUjA8H1cuSYpaVYSLj7KB9xM6J2w
xf0l1aW6ywyvL0/1AQptdJlWRAeL/qLsgHsgtNCGYz4bEhiwquslJHheuRNDXCbg
n/uVnMlkkPR3MveeQ7xqwVrN24nYory8sPxVTKMxpfAzB6/IlV3uN5gj+JDE5tze
b/dCvxijBS3NkNSUE+P7evyLAzh6s+kHxqCc46Ejo2jbsVAkTniOqRY4CFhskAXZ
Iqd/qZlIBxntxDSh5Y40mdc1QBia4s/nC0n7Hh4jKEUrl0thr8YLSElNUNBiSH9j
JjTZIROvJ4u+Uc2uYRN6UTrAMtOgFpxAw7tvRJ4OHsp2gwzoj7qDDzwzwoNKGQTl
70ugk37pQSA2lfPNQPbaB8BqjWJZTNlJRXs/fg58HIqQs9TatCW4oJr7L7mYgliS
vS+0/WBP3CeoqOyZZRYATxSg3cFG5OmA1NripDNg9MEplaIQkvR1Z++kg6y7BpF1
LK3u6/UK3N9S4Q7X/+mIE/kG7KFyIDSr0uCu2bkpEcCWa+BAAuawSH3TFCqQlDLd
dhr75l9hqa8gmtjlkl6M+8wiOvz59ChMXXuwB2y/akhwJ7Pc+zXUBUHn0gE1fpUG
q3ziF0EoyBViboRJvRKq0OR4oRMbDceCTWg7xB/n4tj2G8IJrno4FMsoi24ldAzi
zVrRBKU7zhtvDeMIQXASJBDn6lIHyGDBmdox09yALGRm6JVBC+nVkqzSQ0PlhO77
fd01uFslmlOZWnO2Vhm8oGViHRNy0UlOc1Zle+3JY5Uz23MHDgkhCvJK2pKCLssC
Vol/EUORKb3d7pZfGNvA/VTjhmUpvTR4HzQJEy/7lPCeg27oOquimesp1x0oRgOK
j7Mo+B9UGcH6oOPtunO+6e9g2t18u/1cDYbPObLthtwuyQgSfQoDeKpUUnY9rGpf
dXJoi4Op9H/MOymerXgkDz7dB1L+haZYMnZm6tlFdZybC7Nk35LPlSeNr20RXKxx
oUsloAaRK42uzmr2fDBpe6zEJiMxsTW0sYDimgj8yZwjOkOccId3NmlPxrXojE8V
h7YkwXw6L5ILj2sq2EID1HOwC3s04ldGyaKt7C6RdNthl10Vv9ieRdWJA+D1IVP1
E0jAyIAy0w4LULMwrskJaB+1tbUeMhEqXJ2N0ut6CMByGasdi5F9j9gRg2NNWUrL
OpeuZX+5sgbM06hFNTD8i8mXSFicarGvSumbns9/YR6R8XA0V4CzppF+a/i5Po97
bKjQ0JLUsaokf/hQNtUViqrDT3n8TApmfL/HnbIau07V9yO6QakWYX1dUu5lysCw
7xhPHKkxlYvLPRglsdguWZ5bqTwwfvdKBXcEZrnFGDTmnzOrF1HZeuCr/7fKXq80
VQHn7x8ygpltqS123zFzg6A53OgMToP+7+cvpm2BctF5nb9+civLC7QiYAp0eeWG
AwUgHpSc8sYudhO8sGfXQv5cIqfqCfHTfzKlMpV92otLbPwH7iVisVyzmfbjppSn
PlH3n80YZpm2hFHf+RIqmk1Efd/ViUyVYWCxLUVCclj2kOW+cI01o+YQTgG/ZyJ7
OLX/1FlN12vTXdsOzf702E0lJn5EVCFcA2GZp7Yjcatq8c4bVzfMM7BngsTn29df
eRZRo5Z8Nulp9c6rIB+Rvexn3DtA1bv/bC0xBIRujNEtaH5sBSnwFZLSKrB8pWzk
YFpeNjXUcpvxEq8Hmo2ySYkJxjKJvsUzoynzz2kPmGNcLWK/xx0D4Zi3TKTr46SR
cm1UBtNDHl0C8NS6uJXHwy9Gtg8IB2+TTS89hakD3+2Qg3DMax2TtQzHesYL6qbV
BgV4Yg9/lhEA9FJXALIJEw83G+yYSsE2DvGFEZPanf8w/oeZ5D58IVwYYAUr3A6S
TKXZdMugYsH9+t3bRXgOS0JAeNc4Huk7EkFuU2udB5QhTIwYt6YhUoC75SkwkghN
swBJhefxsIkxJA4JAHbXh8H/zFiUPPGvGipfZEpLALdTZ9G9eKUqidjWDPOdb2qC
6NAIQzjhCXA8ICSYTnZq3Htil4cRake33jlXX3ZDIkdrA2+tn2z9FiMH0GqPzjaC
trOCkCP4NWhRYlJ+Y5c+z6qu83alKAgcxFe5V1e6QwdlgpJpFIkGukUQlpBbnd3t
xPi+dRONh+/rRQBOmDd5CCjhqNoPGxg1jJLz5XDXWWO/bJEIMgfKJCT6pVe/5e8U
HfTL4THJSjHx1GZozcEr7N/TGHztrxyD80tv4hTNXS9quiyPAEgpg1kJsdqWav8Y
Mh0Il2Xo/P5i/O00Gc0NpLx2GN9Z/9tzA07zkvw6fXAqyyWvMVMKswdZktEPolGD
NT+1soU8E2MjD22CGcGPGtcPyiTFh2u3z7o441hKT0STaKAWCyqMULC7eTTum7mx
crbRBx+QKdMPWOw7j2r2pasfJ7qccrzf/Zk8qNH69OZ4Mz7H/3UKtuv9nSXxOvYZ
kEr8hO990v+B4jNOCZrH3GLgxr/3lnkSgRh24Y8OPteXq+nCHt3v2h5pEJd5y386
8Srb7KGLK+y1OWRnE9187CKJ8wbDqbhupSHlNH0BLzix0iyc4MFVwPgVERiU5QXG
+Vr6UTWlmnHmhDveMHdsN4T1L3Q+mL4io28Pypn46sdhd2rYj3LHnEJ7i7ZD+N0o
4b7qjibztTJoqNlNcS/WNUecG2aWGcKEGReATKSfXG/Gn1tMBSymvoYCM0DANZkp
S0ZUboEnT7SZzrhYdwPNova8+CxjbKLYp6pgoYcp3H1XXGDVOxrKcdI5lkptFPiI
47067dWIXThoc8/SjnY6v3/Y4JDD+x+2sjbT7GPbmmLexn1hOYML3DbpSTq+0Tuj
v66xGnotDdPoMci65aTa/TxbC8iZOsznGdAZKSgNM3EjX9RJR11GQJVbYpLMDOxu
kGstP6PRH0J86q+8DbLVs9aDEo3EakKUI7ckdRjamqpA9vdEsACJF/yWkiTW7vPy
a4+GcwpLcHBINZXbJRVLQjuoqEmhy40nltew092Pdwv3pOAJr9njeHjG/eC/3SWb
/mu1Fo9M0m0xsIRWw7ZGeqUytcJKctC5ThqH3hhfzIBwKo8HWaTejP5GEfHiNjZE
tmZVasCC1CWMK3QI8+Bzanz2PyXvX0KhC0MVXZkGqksjkGuXm5SE0IGSFpJQLLym
FSbh/DUA/1wauLCeEqXejAWcR12ZjGS7fu0RnCHUsSFuIMGt+k1Wnn8jXh597P5q
l8BSsZldDCR0/aXi0pWidmqao0GFlNo+QkKPxaFF1gCcWlCvkTUA2IQxOM7XP3xs
dpTRq2UzFGhjY4DSc4dlCvWIrHDmqxh3y1ZHDrbH4AGaquI/Wnnw81sS66Tc5kWV
qztEcbtQFP9cFvFZGQOrd2zUQqeFjhXljQ1g5XaotHjF/27ATsqBPHtI8h/P6FqR
MpxjYZldyldkMs9x1MOv0dwrTMo68jPadVPpznCpRTSMD82pDhTyoMss/zrfYkJW
c4r3xIzf2ZtUpM+sw2T1MNLOi5v2OzgfZ7sidS1fDJ61d34jVitI+/pFy3tYuPFP
m1Hap9UXrhQmrorcIG8/nKVgM0L49/cvFe+DlDn25aEqaw5geBGb4U9hNGwkRnJX
yj7L2ZFnBPdhYZqQM8rPTHZo+KHMjNrsrkTZ5pOF4u3g3rmkQsEuKlRywU3R7e7C
Xwk3bGDDWsQ36wuefHc/cFeIiDAHc7st2Ar4g/IYs8kg5y9QMJ+Zo05i7mhbRgSg
AH885yIMDXsbarGvU1Ek7zFevkPhqWlA+qGhaevb2ZiSKy9bAqmO1HfV0rGJH2i0
eQ300LHhX9zm0k7Gdh4nYHOi7LZPok4FHHA3bYyeloy+GH+VOVV665sflmbkDTF0
7/boIQWGSZZ3dpveBMiA2OZD1rHNIvOdTKHH5gAX3/DGyXHK3tActVLC2hJMjJOE
P9bN3IEtdAK0cgQeSPxLpoFO94XcTWXvbIUWLQoO31Hh6yLz2G0AONpi1B6pZEmx
7IMeqxOXhRzTHlwzRtj4BuYKOMw3eHY20MPHoWKIbUzeDUVc4gXgXFp7Uub7OSQZ
+S2IcJP1cr9ocmu/i6Pi9jkkT+aY5iEcyB7d1FUCQqUYZcN2mAmBXgapIldmGOC+
+wAqlHTASinVdhtBczAWk3vqyv2eEmR5b1EAw+bX2KDqmspk2y9taKs18JEMNni5
kEX5HzL/0NotyeEItd4FMH09c3hUnRZFWa5jro+W0okR9bk9lHsOFOV5UxOq4Sva
x66UYjiot65babm8QjWqYiOUyncGLCjA67vBBTVXwsRtHS46ISQds8SvCsNpuFR3
+x34gHSCdwrwioJ5njz3BvUC3ysC2VNIcenA6V7A7IHSykflgRg87BMmha9W6eXS
Vemoph9ZkzjCC+d5oNNP0oE9tFZCayhizbcBIRhPpm3vSiXhdtV0858EsOy/P64W
yIGt1/KALFqt6DPglz/unB+VayOiksNnwn7mVelLv1vnJ+WZMbN2rJGDsl+wmBJf
/5XBA51da1TOvO3HhrzbPxPsEh7okhiAV1ThUHFmTpT2pc8+apHGIWcjEzwvsZ32
Usylv9ZSrYuyjw+tbCeWL8JhLMPEbpC09jG/3f4j4ZI1bH/fQAaok66wZBN6VgK4
HjqwKBsPxipy4X40rdbUsUS6mNr7e0y6jB1/d/8UvL9pi8EWL3wj5OBnl6uHcvii
ze4kvzORpU9A6vwazHQsiE3bAxfYS14mcl4NhqY5gVxhEgoFMQdvMKLQQc7wwiUc
tMZ7jdbD1TmTg+h+EJpyBRbqBGO/sS2Nz55i90ofzxsLrHUiDJntxnbJsqT9tgA5
sxHq4r6qcK8DhFdpE9Hki5CzKZFtlJSckttbeKv18iHtA+meB6Ztxhl5y1YDnk6Q
js8QyxmTcjN0m/0zT+Dfw4nTqEOi0nZxkqx1mVoptvLBuGPhWX0sIez3KL62ULSo
ImSFTJKJX4D70VEp2nEaCz+rAfcnOeEH8IQp5YsHKruIu1tjpXDjOV7TE41rtc0i
PKIo4Q8Ed2R3j4nBrdYqEurebhGRk2vNBw/n2L3BGr6zykbRh8kHvEbIVxTwfqrP
pAvd6nqBMq7X4SYZCzWr9qVQAU2GbIOfBmGUbf6f+Pf8MafT4xPTt9sYkMZDJ68F
DRGOGUUfJnfO/kPgehcEPZ4sjtyjCFttp8CSyPopVbPK8xqoXEBXdvMGsk+IE1Xx
TyLNZSEC230gyb7Ald732Hj0+rPtAuPt7lg7+TGGsF/hzmKfPkdfix9XB7/6y9fA
ESNVchi0flS3Z/GbUbVMboW4Uj8PbuqFoNvjnUKdUQYB9KXgJBfNVha60mG0LpkV
vbqttr44GM19MHPa4n0mOn74D9qRrqwWaOzsaywu/y7ujp5Qpryie7kb1pXDxbhx
RA6nd9k2cJGY4RpHmAx38KTVPawCh7GxRVWLgYtuuHNTecgvcewJ9T7FayrdZxxy
ORr3Xlqm6cPETc1l476T219AkmpPJfjNMhjAvKOQUe/StRqcDcaOcbxQqGW+Pr4o
7p1H2J4A2mjNlPbSkA6TJjaQBH5Djsj282wED/jWWcQpanasR3HvDyHtHSRaV+sM
jSj58nj8ctENcLe0DHNZlYkrYbow/b9G6kMxBe8BtNispTyLCEsJf+bge/c+eFhM
U31wepYGYQ8qmG8KogF8/b7z0hbMtJzCpl/Y3Fc4XEsICc/+EknibkgwC+xVx4+f
gCR+xGwG6uYxicZpGZkQYDiqY1zXPnyBSRfQIOqoawfRTNM7pS5IzhO06lpP5iZE
Ka+JR/21EEt09ovKWZUPmbuPrDDuwAyfvW2ACDfBEoeMO2+kYCcSpG/IEwURW/pH
gFw5iCHv4hcadsyYTIc2rnx80GMsvazX0/UKZjVJoWoH05D8/HlSDby+aBvNGnd9
iCcN6qgko0xa7vFez/sZgvNaHKk5P9OedAlJa5yk13YN9GyXnYd5tbgVzZ6YLllS
tomu01cGL3TOl1Pl+4wOPgLh0xPoN2m5rW/FWgsi+K1dJN+Qhhb9HoL8b1SVevLk
OWZGEb4YIkKisYcKVDdFzsoFRUjHfAAr5oHDKs+qCPLxNYtOvwWMlHSyjxYu452A
BvDisXqPM+2qs0sxqEt5pNgcJSzexx3NkEArG75SrCLCHQKueMUkQL34maLUajQ5
vB9c44GkerAJPyUOtKdaWPe7A2bs9JEvTSJQ2td+St4gOc6K9WctpE0pXDHK4Qe1
bphVx7xjXJFQ7gqEGIpz2SJXiD4cVtHnjaZ3qHXtmQG/0r9vGBbBepykOL8lB9e6
rfRD8TeQ3N1b3YMq8eBzemKniOxWQl+A9qXLJQ95qK/gRvdBnIRBQuTeCplxfJ7l
/Cd6QmJ2ELKVBO77ypuuhZZKg1oV6s+ds+QxAe5r4l/hs1U167Y9jf6dl3bBN2F7
3BgMvvlI6PhTxj40u3Vd90lHUjlO7zwdjgqwODxCRPJh4xr6N3d/rO7S1lNdTn03
Stg40p8gVHYYx3JwHYfYg5Gl444Xcay1DMvP5evX9rXnTHIgBNYktVTMYdD/UrhQ
BgaJp7m/KN7RXYDLv/MZ+ML4EFwHtM/D6erfZPI8ozblL9oxNlyR1BT8OxjjvGEP
oKVP3moM4oBQgwWVrdsSo6jCA/QW+VhFaS72PfB+fa7Ot02KF+f9awG3TRcV6UY6
Vxe54l6y5t5Bh83ByEXwVvvCbSy1PkkIPIJZdbxOIBxKfVJESmHRWCJxcGrl42hU
upaqXa7U7IEYMrRdTWv7UnMWXQpjkR+oby797j1q2oVYY4hdqqXBFhWyH1G1qQmq
WVxdZifoI2C++2/7tAUrhxOi8rGpwuVw8ZyGfXByRaeSa/tE4GqV2p2IqBeHJBzO
hiswogDDAjGpplJ6z4aRk+vA8XgUZ3SAYxMn4Z0Vt53+J20SvLSilHUheBjV/ayG
O7PTxssl52nS/D41B/ZZzVlm1nThUS3KDVLGEeAjwAa8axl7rLTJBtamvlvS2v65
I5MCK05qM93KBnQ4siFjLAngL2uLNlFuv902sAtxQztLzxWC0JH+vq0jrk+loGx8
/2uKYr4aMfFaxfFuyLXS6xORlBf2imUDaKrPq0uPziUuOo77uwtTjOdzalC7njUT
LSmYbCaUp+GM4nFU1nEg5/VZIS4yjsOFBCi4OxtaMQlILirZ71McL648i0pmN+nV
d/U6LtmpEVqyWPtKhLgHmg==
--pragma protect end_data_block
--pragma protect digest_block
jWiwzUS6exmMH6bLbUXjgKZ4YpY=
--pragma protect end_digest_block
--pragma protect end_protected
