-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Mw23qYZ4jPyE/Jv/n0gar+xYXe/+DIPBObLkUyCeblEkw+kusFVV/paDb6iSRkofJUM6jURSGtkY
PzE2WKB/myaZylbDXMVfQWnKJUsZbUlggNDO8LfP4BzukQNM8lIGQuLPl7m4hJ5akMeWAgcfhU1A
TXMlghrIFjy1BeuzjhLXHToEk+oYF7bJ/eZRu6+TfNDMcntzl8Y8JkNFG6NtjTSs3lbzN/MaQvwF
5Ow+btaDkjGitoLG4Yk8eXyzKRGQVaGdo1ObZlrDn9+yxPHuU2l1IjuxR/Iu2fHCMyv6JsC1BlVh
E7hbuDD/hIU5uBxSCvoiDR8UoYw0nd8oac6Ndw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 15488)
`protect data_block
adeDbsrGS3sdik4pwLqcPfvNlkHMCkel1BG/haxzgv5W4cleG72hC1n3dpHw+syrvZKmpyZrfRBu
KObwec+NJF2qgEMKN9r2JfY4p/osmXzKDGBZK9fnPAvkC7cg/a81plhigEjjx69XlYsYw8ejkLCV
WAaL2ZDdYuONnqppxmMhV1xwZLK7eELXf4GsqSdyQtBTVVXmzCWl346UcWVFb8brxIf1qDG9HqV2
bPv38Oplk63Rp/Sh1V7X4fvbczURAv9IGaDzHBpvGw2+/0hyYaSakVWJLecfTGYx4nfchp8vAnr7
JyQhEkDtlux4jQ3syE+tobABvDxO34gbPdz8HB8eSgcHuoFfHagEusaq2cebadmqcBviYOjqP/DQ
DMQy8xODuklmwUvTF+PSmEbsjXiRLCPztbziQovwROu2YbxNMybhKVM5Myl7JsZamKYn14fZxPJH
fC8ZqHYDVadtB8uwbAl86um1H11FTg1X7g9wCorWozaE3SesUZwjqvv9OV7cOYeKZjKF9EAgzSKp
myUSNH8Nei6Rn62CvyrRylcvkomTehDfxmgw7NZeyqZV5PwiZCcZE8dIz9aPJHkrNzXoE4BAvR/8
XHqekroo8bSm2O65oOpZI9at2bLm7Oa8WYEgwUF6cjkYXoSvNbU2Y0acF4uilc+B85WX1vzY3s4n
ZfY0Egygejrld4TtCPPYFlrozOLCzcTScogMX1pppsqsqH/taG09t28l6WHHwAhbFivSSQIgh7xd
xXYOb9dDmbISUKHRAkOd4d4IdsazzHVmNX2TH8Au/x308wwCHv49zo2UR/S0E3BOh5tsNPQEQJwh
YvL97P3Z2l4F6LuZgo2lqpc+l8m+Qcn2Jw75VJG++dFmh97+k5CixV+eXs+uamQ+/rACym3pE7Vk
4sfG5Tev9yHOPeIdfXH9j2+CtRn7Bz9iF1ic3LMIP+rZe3UvyCRLEBNRJEIdotYmfSziLAde6GMe
oLpdtdO5Z9BCUCASGzyMT8B2+qS/A9tJqj14jBSBGcLMUnZONueOcqvqJB7gCwJmcR760AUVxVEw
PFmQQiROSDkfm5/qyQay1J/carc0n+a/6qd/dm8gx/kJLYyNCdDHAFWbCc9CjBUZQkPOO3ZZbs+Z
jcgNmHVsSD/j/YuvkCi9IC37/pmRpPF9VhlfliVatbeI3ophOGcy/7r/mNkfwFuqsNzFzl7qRocF
Efz9F7SXyfGMtt0dgxke89mWQHtr8W8tRsgLOCxQBLrihpNgwZPlTjmbvFoRH0NA/QLLkcdv/xO0
yHocjBmZ8k/zXQEra9NKNlpJMcFAlfZcsUglAMzTh80E+h21s22Qb4oePxNBxksqrRYuNYp0ky2a
zcP86greKyDA9GdlTdWyhEDW9tTcJYFeqfxiGgTInbw3vG+uL0DJKiWB3GV+yua+m4c7wMCMIwna
gfyGX6gGIsbC1b8vUfvg+sM/D28EtlbZctzEMM1TRVNPQirxykRApfkJhYyp5jt9Skppkwp/8AIE
b84MDVIqlMt6Fluk6MtqKbDXtj0m+QKkGhGbTreNlcIqpvEFdvXJBMofWyXBKxSzyS81mJb2EXk6
lj1reOrCeFmhUyPbuP9qIBVarOFGAsIVd++OJiJ3rDrECBzbi8JOMGKVQY548HAEdwgrIhJTMdz8
oME84CtvW3myu/xi2oYGlFq78I/nWm9TaViF4WKCF9/J7x834zxIXO5RdBpoa7uuxny7cHOQPCcx
A18xrDMJur8fgacsDns4cdO2Zc5v/IKD21TlE/nPO+yev+txkuE9VJJe1WTD+wwR1k//MZGpEDL3
Y0f9swsl7G8ER1227AZB9WvPPnONa2iy718GgcOkk0WYgDJcqLxys9fCjq4mwhzGicPiXzzk72HM
zWIRv3LTfoo40KuRHwK+XY8vBDa2dtDhSJTIJzEPDfLMvCIGB/lHmtni/5bqTUbJrzlxnaD2qy1a
YIzGicM1zMv23br1m4oFw//TBTtY9GQr0FsIyZGUGAOoGc7Qk3RK8/GYwo2OfSELrKc/Cf1EvVcU
i/qPuNZSHGPRySxjdjy72/ThTamfcoglJaJosnSEw3Y5ziwHw+nyoWwFkgElfbJqyZAXUZiFpE5g
N9zt+vq6JWUr+D9euPoV/nZdnqhSYgr8NZzsrKMYQGD3GV2xH89Hg8fSzSEJZUlJTkCSjMRzld0r
yQPOirg+J9lPhw9ooOjsIY4A4JLPIE3n/nLethZEPB3SRo3Fbyz+v/GOq367GtP1zZAoUYxhq2M7
Nzkz4EyVBVNOy7njoJlcP+7aJRaXOoFsz3XDQkBSelNmillcD1gjDFMEOZa/MD2sCIqkIKTfuGG8
AtNa0XG2oe06bCo7sBs10zPPaloDWfcPNwBZjEVEAmmgi2l9+suds9VK++/f1NHNks4xwNTMylaj
zsLwOYMHfQ+dT8nAxUmDWRc3L3eWUUb6+PnlrgbvOaW0HngDNXCztgTVhaWVWnT3pQl8/yCe+hSV
OPeld7h/S56bR8l0pHhAMrJm9WlsmIsjp9H92ogM5VG6id+C9wD651esxxn7AQW/BPEVaja9E9zY
wBxPavoC5gs8WM1VECt6mWY55zy7/ECl2HLMoAU1Gu23fzNwbZZzcoNM5Ghje8FHVHk5E0m5Ux6h
qmBJGcb+SRrsgMlLxKlr51pwpNZ36wW4KonD0VyiH6YArw89VGtO953vCrwU24hvfG0Q6/oFaZxn
j8RYVgJmFg83OWl5Vbgqzr6GwVVGCskW+i6aNAbS4Y6ncm/2AzNPQXNu2KzBr/fQCQUvf1FmLvK/
8Dmd8jtll0yNqqk0ADi7L2rPdBO3MgZTC/9s5ZIVGHAl0LoZJwEk26HuiL4ovCOGEDzImLrkb9+A
XLZ2c83sZvL96R82woDYXDi40H7H9Wg1icpxjAMN51h7xvJEOuE4P/F2ocNyB7GCw/MLJn/z3MfX
9puGDbxrUdHZR8omEgJdmnKw+jzI5uCInJdLXFIzGEqSPgbJIYLlskHYcmjAK1RsT8EiJcnA+pAn
fTRADgNLLm9abGMze6Hf9Ll5e9X6y4VW+73ijbi/iqpev+zDDs0FvivkA/mNTupqalLJHEeEXuzT
S0yluqg07T53oOKKzc9zojEgFE467BtrRg2cVRjcDBAzaWk8jfbwm50ObunHxN3mytLVBBVwtrSE
Mv7HYnLFzx6nVzMm2biqc1XdpO5lZdyJHOmaz7WOCefHgqQZZ6ARKw7zl4Gq2ON04sggvHkmO7si
dOD3299P8SxEr03MF7T1YjDx07vdUG5nK7/nvExx1T33Bxcblig8UsVpkeUlWEAmQjf+UOUgtL6J
h7q69fU43RcRf6ZCEFtxezQpXPYWkwG9UDTrH95IAFIdZoIAMB6eIt1oLxnhCfjmQ6bnfov5rIBT
d+AvDkAkUf7quKXz+Qcdq/RGUCMr2XvJtkuzvwUbdfyZEjMFBFqtOGqxZCwpnPjw6r2AA2L33mMF
a5cmMsJCCEnmGd8cFon706ae9sLsDzoqTcs2BvPhqocLOR3poIRobbuPZiqA6Xvh0AH3kRS9MC2n
h1knTWd5TfnzcJFPhxvTQups7Its6bdJj8B+yFHyMfNtLkBzHNya3rr23KTgPI/6Qvy3Mn/MgNBc
XzxbDEZ52EpL67jrRi7ThG0Ii4TzVISIrHTWDp/AQUNYXPI5KoBNg1ZZK1o12azHVNkT822B6wl8
ACQFZqzzkMbheZ+DFgbmcLjiP7apYI64YzpweiCw2Hbc6jStG9GWk+DhFgYX5R3QuN8cDVIsnAAA
3Rrrf+WJa0z65ez7ItyIUCV99IJAolzMTeef6xRxmHfflbX1I7xpmNHrwEnwFBWsYdXAU97qVN/U
IRDrjqygbhBo+k8YMOTofUrzC7/QNxGNxFLupNeuqFXymU9RT8CWpEgGafgNceZcQv7aVrIKpK8A
KR9/v6ZCd9SwwAl/dCy5kDHRITHJRUmK0hgV8+x6CguylzpazBmu/ll7H1tMhAL5PEKLy4+Jhe0l
kmnxJpqxB3RAMvIHEteotQFm/2bACnnogRp2OgWxk7czQxk4NsJY3BWQmsst0ltg67ntGy67HS+3
n3tBNQiXUnrfby7FKXaXNjY46kgZj3iSENrRWBxB+g898Gb9ELD6s4dpQG7izZm46rQ9e+tYjvwH
RF3c8OtS1Gaf9Z3+IQznLM+yQXT0no6ynSoFBSRESEA0bNWjNhF+BVV3R3ni9AGzVT8XSibfPqNJ
uu0/PayxhoaGB8NF60SkkVo/CGOEowkHMiTqrAjKmt7FzU6dWHE2GYo72zJdvS+YBrJtiin43gCN
vyqKos6mKjNgtTqCcKPoBHzMIClDEk/PHrQNPU1e5c3G39C5LrpQ5JJoFfYS1egAioxpyCBz3qNc
5HtEeLuQlXRlhnryZfFTwz0Maj29hTpijPXYankLlqvsS0pzyKpQdLFk7a1nY8JyHr38OUP7itOa
bNalgRdiDZD1IENpCthYj+lJUV3Qx4MXc0z6ygb1SogbiU+tX97g65MlTdUtZo5gutKJUDqh2MX2
4B+xvEXbTd+C0y81lqTgo9TnRSg5gAbR9blkj4Ko6vMgvw/mbc5eRcWmVTl41I9MgEv2gSHlTF9i
nekbqHuprePuqmUnNEas31TuHkTwbbx3QbBLCeiJbUdXmjgsy8KRGl6Ze/gPxO5Z4289jZ0SCBA6
NNPakyMTflZCFEeEnUaBQuex4FDmzzEMeJrfs4coHRQcs6drO5BgmoDr8on09eWdEe/CKVQSyfLu
b+CKQX+Q74tuEDusw66+TYZnR6HMnza8kwwiAsIUNKmdAYZxWiAKZIPF1jYgG+t4sMcyri43krgA
l9S57/GJHTwUD1UZX2cXwtPnYfjWMG6r1dIeEdd2MPBkLaXU8aJVxUE2KA+lZAf58CxPICKyQaM6
arHjij30RiuMRUDrqO8Ym9kmAP/rxGGrFppjDEzbYH7OlkleNMuu+uiEoYkMpZo4hAjbQ7kzQyZM
59zW2/kD5akupYXapXcPDIfhRQIDqa8Q/UloT/igw7Zg331MAndbFlmy1ZO+eZZJFJFLFHrVJ2L2
1bUQCpm0HtOTuLgpTlsuTZqQYVXDIsuZx0nNHZZqZwlMFdEK4BfZF4AkTRtZAfUG2tk1ug2ODoKH
NQPNitLIEsBmoTx2RXBYs2HjSb0T/9s4dg9APfpQkqRG8aX6wqZ7Q098CUipz4cF0WJ580suUCSp
yQyL5VPO3qJ7A8W9WWs3W6D+kIJLFwewwVlEr3B9lDDNIH8jPOomQfW5YVyNthFvU451a2vTocQw
Y2Tn76KtLJ7rgqMwVKKA3dyoYzVntgf5RrA4a/iz74GtzMEm18fh8FTUEw9BK8R/n0of8ofuBbl/
Lh0MY6eN9PnX6DakboSR7yVJD3F5paPKoiHmH25glTTnsKt3nPKgtrgAYoneoOUqZufrGlo7W5oI
qdfV0yoKnkk8ZaFGBAMZcavDb5b7qJ0EKwofQxCdgX/YO1rTW2ltGyikgm574r3SyfYdcjIwM+f5
z8osjk91VXIzPM/ZVjA7eeouvB9kH5G1A7NjdZntTEBvu0zk9xLPOy9/Nxl1QXAtHIuk7irD4n5/
iQzdZDvKX+GLN939o1aqnY/wgnPYRCDMaU32vSUUJ8atKfByXdL/NuipPVXw/VOozsEXhSPM/n5s
WEfJCSJJJgwIwnN6WTlzu2Hmo6GdQ0K+pd022gpupp19mJfcNNLw+YueEwsc4HInWlAyNnQ0/U2M
7xzT0lsMSbZ/XZCzZSrfofa331P1n3zcoIIHDzG7Ck+14niiaQa3fKUI67lXnsNfKt7uJL2bYHRD
9zIt5C8qNxNqcZ+mzodimEbxAoarRkLcFkrvSl3jYhb6TcAhgFn7DqpDC8vzvMiJMGaPxZ1hWsPK
02azbDcZfGXKcQEB6UMCO2zw/KApoN5E1aBcq4KaDdwHeEQtu9oAcRHeuwn81cB/kwMKsKggZs+y
XJwCAWMH2Qns/SqU0UIIYGmnhyC8fU0U5Ji7mwABDSirhjIvwy14oG//wU51CZAiX1PrCfhPWCre
RW+rutsZvOGkJlX9/zCpNTUqxuOlII3wuEbdv7hbT4Nplj36KwGLfWBsp1VjZV9+aobiw/jdZZ/N
Qk8F3spBS9yWV0HTS3pZ3yqEDNxywdXYeexwDfAdDcFnAplzlV2lqh1Jk7lPr+Z9ER3uhYX/iyr3
8ZQd4cMlRckWwM2420SjnN20SoWPHiGlu/P9u6shJrJXHa9pRD3xtX7UkWLtrGM17Cwi9C95eETv
nclDqLnIMCOEH3WKy2JkY7Xh4w+vAqf+rJwwzzeFRB316yZP6huAVDEFif/UiJI0ESKfky8nc8j2
vzp3AQiuLfRBsnWGLmZ+vVNL3pkrjhFFKI6Dxk+uVFu8Iboj/dmUSa2tn/VDwzTTS1eA9A+Bjjic
M33x3Zz8uGbcf+NiDRemzYFiFEaTKpQSgQupDvrrbbImelhyjN0KV50rbUPXCTM42HV6e6vp+Dri
ADFrKQLDmzqgNQVSBTj95R+5+7U3xKSuYdbh/6pvdlXNcXy3VJ5+ByK6vRhIfMkstEbk0SEJrOta
ybgNuTrpfmk2Zvf1ITP6sdH1Z6pv3HZFqCGTYNWY9iEvNA5YaVIu65HuE18E65kb9qNDh/yjM553
PlkaHptsyyS5Y9xJk+x5CN8GAFmuSh8zqhzFoLQl04mzpUIqqmHwPXMqirs/SR9UcN6RD5RKUvsf
ugf4VtSWRegytobcRc4DBu8hkE3ccy+kAw5bWNiAmsplxWouCdJ/ng6A9l5RV+1hGfBWZDbNzJ3H
7wYaLZa3Om8XeVzvFxd79kPv1ilB7VFzj6IW5rhhJ6jV8tiEExVM2bs8IQbRdNu6p56R1QtCtxfF
BU+j7Xq8mupKfAwX4q3ZJnG1KQI58F4wRafQ0FhB5QQojug4mH1MaljKX7O65rznTa0UyWVBXXiT
u/SLAwhTcIKTCFsSJgNaAI6KkETdbd4M5XPR5Zyk1sFN80U0WYjp9JhIlHtPtb5XLz5hsXycZiXq
Z6L4Z4SooocA2djo9R3F0nwjj/0XJ2qN8ozYVwqxMCckPjRsig25v69L8wP02z+Lb6fsEOQCpDuk
gCQAhHie9mXdbtvLszwl9m3TRp+VIVEJj0raE0E1gwL5kO/IGjRWkH2Ypiozcb9GGiAINfeEAbvN
SL2N8CFEX4ezCHghueXoHLMfeKNZK6DMm0bhMHUUNUfFfxOOmEE+IDNGD2hNFISO9RqWBGpULvkq
MlenZztmsHN7qWT7AIsBP7csdQ3rjkbH/d53l8M/Sc+sck2KQyDqcmdvolUkZRqeKk15gZpfBvQl
4cjFVhhlcJVla6XMtEvKTvMqSi78MwrbYwLW41qIhkeCsE8+OUZV5H2pqQo6FumTSOx0d0lge5hj
pYssrjVaRF4r5Ypu8ncnmWuWQOmdN1NHc2JFA2TwxVMyUqeG/2mz2UGlkp4f2VuydYLnePBcPIfq
vgBo54G5Uz3cMBmfgBS2QpfRxg66XVwcDCbouOIFSfC7TLUxVOqPH+D+Ky9qaoB3GKzdPMYlg+B5
zPuC6H+k0sv/NS7hPdw6E63hzwlxmTL1NE5otgc08tcTcm5EAwubhqM7vzOpSrT4D/Bfq3xP7vdO
m95v0XeR1b1/B6lm5pr60RMV+rCzks0JsG0LOyu+VeWFWqWaXNoZEbNM47/apvJFXdr8G6K/fJH8
4TLjdIHnNo1Sux8Wf9wPIfWJNqYW4h2V5a/EAKO8miPl/TDQ9hDn/in0aKrKvbtJK2NckNVI3tum
jfAADwKWHObr3GNQD8Gd+82IUe8S/lNu7wvP/hOqHYFJ/qWMoom9NUliAeSdMUaFNWhRCpfOG6DD
3WtPR7SIa3S3Lk/XwJhyufTs/aCdRcviNeXkX/H2rf6P0bBK5F96rLmJadz1UBO/NTWeiko4WtFT
D/847d1xfHXQo1wYiOwpxeZxh7bp9KJVYlcKYdHO3cIINzmRzewa3+66kDrtG9lNqDPCRB99dTei
/Lst48tbN330Igt84ibNJfXbSrIPE+ReMs0xOWF9YsE5SI24Ny9dmLbAKwTKJb5nS9KgtcbiEwmf
0Ok7Y/xcrhDCCYXEPuyB1GB4gTev0CCGXMtaKrojPq9KaVD0KCM0oHGerMjF4lAAushpPz4fj7ZI
eMA9LKr0h3/30wUx/Im+2LNaaJltEUoJmzMS9FOAe/MJ06P5hlGwupjAo0/R7lbvrfiozIt09Wz3
59bOr9MbgEnHQhrCgBkDJEheGfpzE5qk74nqcc+GfDLiNTodBVzqyMNI4dalbNED3r2MLOPxdzk2
KCX9Oc9PiRUJ2mAGoHFoNIphZ59AMtOgf4oxseJ1XQfDRFb9zMtrZdHoFajBrR2VVOZOzfJpQHj7
26g824sEYeihFBbyGBNaOwp7N28iIaG1pi5gAi6SSQksuWCWexUDIV1j9jakNk6c9TQja1u8rzra
dlLKGPJI+VdQ1eTKi1pIEMukHvyYizNkEwFkqlw85IBl2WsfBBwUg9ZiesyNFV4qEBZA/pmlpaww
vRRpsn1pheEasnOyrRL3A28oTQVeGfF5cAmGjAYgIEORVNqs5IMG1YInTL3wpLEuUBIAknCLMy6F
/Y36K6iGYif8lXmgKKj/uqWQITyXT5kgaaTSjNmrXLpCI08uFkKZU2uIxb1WQa9LJuv1wpDB6/E8
nsGYPydZMS38Jn+G7zsweBeFYV/IP2mQebla2AXG+mSjr+TSEKl1zqrFNHQTVWTQP/UIxGBAKaWM
B6RS8+UJ8Q8NODU9q63Rga7gdR1sX+PnAmRBfpaV9MbrA6G/iICa32+zDrnFw7KMTp8oLTHr8c74
UDSjblcRwYFEILH1s2zdPA9K3ZNDbNhn9GnnWNGAMw8b6YKqB5TL8v14Q1Dprtf6FQVYycVlC6k8
gg0N54kmRB6+UPwZltWi9FIni1h873KpS4SPBaDtBVhDychOS/ZuSO8B8nYLurBuFjNhEmetWoqA
gW29/XZJ5TYTDJK6K7B8Rc1pmnBNbqlJnQl8n4G4KVSk67hRyilKbyoszIFWl57YSkeJbY4lULZb
mzN88Xr3uqORLfztoJxHEwWi7kivyQ7TxSTTn1lwIumWhzC57WjpKjpR3c2jctW3y90TnbaCIYn3
HMYo09LuvCgFPcV2UE6LsuG1YD9u14dfMkeThSCqIn2Q9mgwuMkuyofRDZAAFMWHQwistGdenais
fLbIWs0gJ4ZuFyqTJhPvZiKEOg2kDq102ePbc9MkqlEEHYrMLjCGQ00wJs6b4QEGcNjkKIJevo4u
tqaO8fmfeXZwXlZ7pagRd0xMQyhKLl+8kVycAUzBAnT/0G65lT4i5SsglYg5JPAuyqzD7a7yeraF
owxssiMtAUfT3jtw0KKsf8jSFzJFG8pMX380U8yczxJzYTIsNP7tyDF8dDVjk6f/ilGQjplvwThi
18RWvuxAcFhqCJ+ll8nA2ZJ2aoD8w3WrTxQIUrKQWk0yeSliNoDZlg7QXCJRCdjpclhQ3bVKGJhc
WBnQ0uQavF8djXMTfONDhMFtspUCYbJkhog7uYM5+IVq8g2GCCGcN0g68jW0KJ/uM0cq0X9SeSKl
GqnKh8SMYjfCeDamVdo/HN8E0zjLFcgZW5+rHtiWI2uZ4egk8pck7o6C90uW4exfd6zyM4whkhFe
wrHjNCsNem1lNBdzDuw+KWy6urac3I5ytw1wpqdHkiACKr6naoGcD87A6q0+z/eDb0iQJaHnLVXY
gt62yAQ1B+Z51+55QrXKBx+GciZVgsYE1heedGlIar+WLtrYA4XPQpscBZkssHk4kIP/KSbm6iIB
hxXLim0hFurubrsXDW4ajzy6EsWmavP1vWQ1c992Rj9fjCFdv2Ad+ZtKg649BV847mJtSiPTRwFr
pknh3V8scwfCrk0tMO1kCIA+8kv315GOs1dIpws/M2yqwLPZ/JUBpozU8BQia/u6OuQhI4lxwCdk
bmPAkBtOM8PN3NPRdK4aPFMWBLBHBtZcaWVODXLZqJL6qDDENdA3mMJqNWwi4hKxCLs5sglTV1wn
t0UXdFe966QwYMSjcTREJqYGRTVl/09xtCIQ3DTffvjlQmsErkMmUG3mx6u6kGW8hlBB3eponFI6
s4XFoWWzwZ0WDrbqhLrGbiC0jLik0m+OPTn6npqJPYj/yMoC5bdNcy7IxPYQR3Noff5dYFZ6hnz1
jTw2+J5DPWnqRjjo+cROX+EPBIS5TYrM/XRHn6jkFxD6V3J1XlMXwsD6Er2qTqDk6ChH/aGtQy2H
eHZaazqqd6oKjudrN/JAXSPNbM+Awqt7ku6yYQizsZFdIvm1TeLO1ibrNDowbSiTbo0ib5bnPLse
94pG9V8RL4feuEz1c302ZLTF5rIHexMkIzkB4lFh7Gzk6088hlZ99ZoH594scGCBE0SUxwgKA/pL
PfctmsYQRfeJ4OrxKQGWINQZ9ravc0X7E+51SwuiROVbAsdbYNDc1/hE3fWDx3bCQmRwgB7Xnasy
9WJayPlxKp+NaruDVW/o734CwJH/FqfWGOC6zt0nXemvzvlB+WxVHJ7LnVfOGoLT2bPSfHoiuKWj
GzVW3/cA2WovDX+C74ZbpIbF8St+HnDxu9K4H5okD/PlvquRjx/sECP1W5r5BEtvxQDTCalynlqJ
e/DrHw/Hm0KPXeUC9DsaZBKSwK+x3Ey7Q/fYA2y2rPoaTa0ls4171jtMs2eI2uzc1SYaNrZlk/+k
oLOZQ7Gmx6ZM5FuR8o4vyvQEQMmqvlt1hbbKYT3gpixxNG+qunW+Y718zfS49lifa0Mc6Z3LvE54
dQz0LZ+foBfxPgWvZepEkxevDEzJNmZFzR0JQ2aJmYuruRkmVU7GIvp3eIEFURPpOvAftJtQDlTs
BATlidMfOacUiyfS/6W8a4QAuoknPAArITENGLa1bP1A1Qz5oZeWkXiZi/KQa3qTsBXn12HSwBji
F9KnD07WCGc3Wuc5Ebm9ygsb48xTJBfFpniPwwx+4770o/ISp+PVkTfHtjTKL9jLO5f1gdnXjUqD
uvTgcRBtRUI13LHH698mPbwT4ut6JRInPEgAaZ9aFZS2HOTYfvxftrDp0nIADNZq9O1dvy788nc/
BIXyrZ/kM/Nv3YmDvRB6GonbQwZw6LJ+iuzybAiAyAMrz5PonrdhI2IKERw94hAzgPomKweBKKii
Q/aeVQCH4TzL8M1JXPpwPfB5rJt7gT+NQzhiK3vChXcb1CEwMJ96xUSyiW9QbbW5CmWH2OBG2+Ue
fF8bjNSaqR92waugf5zseWvKJcon/nukw7fKaGeM91P5n1RJSt8N9DEUog0/ytghqlKBYBU/XcvM
7Myr1i/fwdPH+pH9fW+B3J7iKkXu6hF9y6SWpg//qwfypRPar4p9H2FhivPIs2N59pV6G5C06O1h
DuNm3CtRn+ZC7yVNOfjFwF1OFRdNx5tqNchXtsHK4J9EngvDrt4XBBqH9Iom5+JC26FLGWZMSPmn
ro4kRvl9Vd4ZNyJTkhZOnu7JZuvLTDVdscrS7BHbGXwKPZAxGF28PQ+7DGjJFKj53WV6OgOQO1cw
ZDj+/BM8zC1+ZyeoU9WBau/k2xXsIBp/5DUmOKE9s9WcSZSRftRnxzKn2ELrQ9bfKU6kb7cO5RVX
9KHlAQU7K5kuI1OYmm7x1cefR/S2H6vE06ieRCKWzSe8grfjsFAo5sH1FE/JiZojyOY8mpVAFNnr
/t6I4jRxuYVTN2Ye/Qn50RnLIGNlxStgSJm2JQuLz8T8gd6DluJ5idnfvFITwWeQlBiUiSDRKwEi
iiI85vdvvS2vHQS513g2bHtTAHlmm7N25ENoCkvUgAbsO2wq/GnSg90Q9qgXeSpGd2Z8453YNjLm
OHHo5j/8ftZkVqloxVL+h9CPdzdqRDMKb2H/uGSzyWe5OhT1vs/h/mpcbL+aTrmoah0Y7H5nf5P9
8BnOhJQtnLI4K3h/SBnaZ2MjCxgbY6TlVYDnjZFCYrgdtzPkE9UB5Vg9YiWt37xi1ntN6EYlqp3g
r01t0qJZak/8Ix4NcC9Uj6+nl0PrZRLPhP1w+SCsXRlIwhUmTaYNF0VaecdtQkYLctTvLEYsahzD
T2AXcM/tNEeYIo/BnwniuONNF1R9lHwHfogKeByqqwUjituxX6rTekyV5CbdrPYu5WqDCkZUeZwO
+RivHoW3P4MY6clUn7Sm7rLrenwHQtc30D2QwEeHlIbu7yqjIW7VfvFD676743eERMhmOpy+l74Z
zUSzy/BuNpelGggdoZBNwqS43Y0kcPxBeWq4NqMv1pjXY1gyAD4HQ0po4x8zeUGuiJjr2lWIf83a
3F2oVMbmLdZDmKfcwFN37BILt0Z/EoR0stax8N5mnakzhKAm3IkedwLXYbpQ/sq+GRMVlDzP1ILE
EmuMtKVocMqwFctX5cyZrgvtD1gLCjEyvsouT1aShKF0eSvvQfcFMiAXgk36IHAi31oecQNKTlsJ
KBHbWQCInRxzfcdqDpgxQW6yM+WCs8nXWy71pbE7uErnMX9/2+/l4Cu0CfxiC8Nn/NNsHh37fiLu
1P9KZOX8XOe83byWermUxzpxS4BD9qkt3RpbfYuJ0g6PFdZWCWeWw5q4I3lL5Nmp6eiGQjRB0upd
WgqRiCpx9rBX0VRJtARsT2XOxrdZ2cneyKEOkZUXKZySoCDDoqsGoEa7TNUC9+IF/c2GDt+TmZpm
CGsPVSitvil3pu1fgTtBAeuKqQYBySK367fZ8IDZeLRHhDCP8exQtUsE4IQSBR+OZpZ/yYi1qYqw
BbfMN2FUkGlI3d28Rm/GwQlQDrgn3tYqa+/uIFx/CNcG+hG481h6FpPEIIz6URGoVbES0jQU3U3Z
A9RWJeD/6FjU1WKhjTh/IC3s6pcu4Im8jbl3ck5Ri8jG6lRr8W4XWgefAmwY4eTlk/FmT/5waQ2D
vnTmy1PMTSOhZuxmAgbZg0LjMrrcViq0kGMLw1LhZIGiQ0r/DTH7yW7M0R2aTSXVJAC18ykC9iEE
ND65wZXWDRKPEzkBm+NoFtVk5qyDpS0fGTUF5/AWnTd45hpVLaAPk4HMN/WOb75HpAK5p+H4dbY+
ORymoZA6UPWu7fTbRt0WdKiEIdBtpvPtOMX79vGQdLy+igtU1pa3Q3apMourXcpMiTk4vs/jf/4G
su9kGztWACtxp0wbhgTKYjudBMblo4+2ucfTpDJsqud9+liRZ4oyQwkjCz8PqGS6kBZ+ICV6ripY
6hz6ZuzdUlD5ehaB9XAKenoS6kadCVhp7OZ/hVJlbbCMBlXc+CtlnuS2f54pKyqrqlYIQFDgf0Fx
pja0P3T+DBkQ6/7OY1QJS7HAMme9kVKkBB7mMCe36+fidsxtxUVwJJ1srZ02mG94WtdvQOFMu4jk
Z/g06CTZAPXD2TTXeg3QsWaC9g/49mRCJL4/187DVmRlWgNNqGS9TXCd4ZpbNbpCLzUfSaw3siIi
KFeTS412wedWlEAW5bvP4fZS9u18XLxY+vjjGQzbOvWhVbzVcgE7p9v8N4yCw3ryD3UEjHYX6qed
znApcUMjtjpZgjz+Ux2YuzKWcbEAqdCZEGeojmRt6Ek/wFKEu2WgPzYx3xJj538QTBhdj/vMBWNJ
lmy18cF5K3oBDA4QjZ2Y+J29+YkcBL41Fd1kdoBLYdMV2AxY1kAPOZf3Ur3luno7PhqUXX+6lvHU
4rjOTuYx6n6WocjF1qsuB2g5maWI6CHZvtRGxzZf/Le7muY9Ue31AYJpxPbXEHys9u8d5FHaiCSR
dPrhwEQEXL1uR8Aw4+/rM/uUCdxl4Cn0xfrY/A69yd7nCWepBm+Jz4ARMZo12fRzQwWl71UwGyzH
OdclTZY0EF5iPh7AyeaEXad4Vt0f4M8YeIw6ZFJ1o3vDcZ6SRR5kAezompLFHiGYCLS1oqG2iZy4
Ev1zD+uHiVfz1pStRSiev3n93sv+GRQvoH1RHKA0iDHu6SjL7S/qz+U/WZ2ITlnegecaPn513H6V
JxRl0FFt4YS6nZzyygs8OKgHAEXcB+E/UjL7FeiYpESIm8AwA0tZj2mqTZEFke5TPh0yKt5k+xwL
hi/GyEcRCza90itTIw/KJy/99+4iRhIfRp1ul6F4XhVbRH7S/glNSTQ4gQWlZKuGi2cwvMhVHqPL
RcRGPELZCwvx28BCEPcVyzr/trUBr9Ppprx16kJ0jjgFi4um+YKFA8Oi0XDORMe47v8tLKi4qKaF
1fmUrMCYPx35XsmeeLH5qhvPuOUjDNRxR9VMsBuvfnv9ckCOxPyzzr/ytHlmgRD/dEfi4r/vBz1s
40grS4haP4WLIOgr3ZrlkS/ucwfnP9PsiZJ+ewAk0oqjDNxDqt1ghKJRGOnYrQl1jOMpGaCjumIa
ym9vL730hMikH3BEnBH4zBiFipdHXrbkhPV5UbF6LEkDx05sZLNJdWnLzdM327anD5akvUdUQ53B
dtk3L8sTQFdXb6STYNmU2huUR+o2ZsxjSJ+8EzJsuOJ5pUHU6FHT8x8YCNlTbaeoMwqCqLhEZICQ
vmOOVK3kyQJZ/8A0fYB1RAQigSzXacuzZ11sqkhBjCd/8yGdqoc8wdJPgPdVQeDFqq6mI1QbgPmt
dy4HoFS8Cfbxa8HuXcu0rHl57lRZveCtwwXW235SGGDjboZkNjc5hLQHrC47qDQCeZdzSbiooWcc
8lgt9tvf7CofpndGQLgWeU/Ir4FoHjbXbBk90u32gnHbDZZ6RB3EtH6WojBVK4AhNL8tpgMNsbwV
HnHALK/OgcWYn2Sfg3WKwKNpf8QDMRge8Pfjh18OEPVgKlk6/ISCITot3JGMaINLV/8i4NQX+QDd
ZySUk1ywrY0h6SSSU3lK611j6xGxGsCAzOrl++kcy63yvnEVfpsGUnuekCGAuJukxwLWCDMdvbOe
BIrU2Ho47+n4D8mu5scdg47u2dWPv5cOuq0veakxjMr3Nu8vp0DGfWHXtf5/A7+1+T+wYRszsv9/
x2J2BCNmoDkhnqKbrsc/1HNuvxlwPFC1DNkXTRYVqLumLuXt44MKjM7ELa2EyZr9I0xq1/v01qeD
zAYMv1423d8XJA5mzswIaJKs9qH8bardR2Cl3TBUeTs6S21Xa5Rd/RX96n9woECc23qG5G8W21bj
8j0cxwj9NNpoNaFDmhUvzMPtc7Av+gBDDqJS9tvGiEnq3g1rpR6pbwemDceNa7ekgejrbp8pwXHt
YFdyyHERsQYKZvcEVPB5z8ZcpUFSVuVgf8oxDYkgFPdHPSfPNX2dUYZeoYWnWI8PzI7onvpJVeMP
9JLF7PdNmlzAdQMgPW6FwSUPKwcs+akUHmB0B3yJl9rYnDYYeSq4m5VPnphJQeV/YneSodJ5PITw
SqP02H4TZ5vfQUf/rPuCFgzhjmX/fFtX2e+xu2M6+3tAk3n0Pr2B+j82oVqYdeJmlKarBEKqd62a
j3dk4QsZWeAIOhYnXXi/2UosRrlLZV4CM1OaSLHkkXYgCXut2RE2Mt0eUg6zL7vgGVESSN23ByLd
OF4qakJUzQehutt+SI/eoF4HqwvXFrGiNceBTfQZbmP7kiHxSwueIqks0WOk8nUICyszxjVgweQJ
a3i72gTg3AN91AHDgiqEiY3BRES9Jn2JixDdcFlYHLkcBHhtjkqtX+YVBy/b3mW4L4ybNELtqaV+
1afWCSVfmLMbK5KtSVE3MQOpSO1GPlksJ24vr6u97Cd/eTz5HJXQVNPICC55ETqsQgP084V25i3K
NoUKBkLacfCVFXPNbdQ63M3QYfVURR/O7bcqhTfDRPE3c8PKETCLjjuCk4eKugMacdr5jKuHFeFR
q07vyhPQXv0RdgTWIFLEUmDaP2EHIKQhipFf5hTNBfvbnazmXV4IreWgafvRAF/rGUuN1+x/m61R
FMk3XmsA89Sx4nSq+UPLisd1AmRX1oA1pzCHkRDndUqenjOPMHImxNwEaB3xzgIxMWV0WpXZZpVU
OczFbkMxI/GekazOuxbco1tbgzArAWHFVsFvGd5MOHBrix56bh9OFlhPgmJMkzsTMifC42cWw8dD
ccZ+EGqnq2iisECAzbpkEraW2+9R1pAV43iO3FJMWjebFiqAOMYn8ScBFsmXks9QZ4uKjSAtB/Dn
mIscftniE4nygbJd6cVkpB44ItbuBaFb+gSBaF/OTpjVsWqWz5HuCcE87idoTtMBu/hCodxD26Zu
xERhezWci2A+U8aAK9fYRYhj/1eGgZJp/XemwmURo9o4KgiQpfZfVmMwA9yiZ+zX0kNM4HIts6qb
uPvQeIudkZch0xocVp5f7egHQNk/wzWG8+Qm+qKr/hNvI4S7EaHU+C3D3oCKoYtOHr8Osbn3cXBT
32MB5avwhyhomH2hVOv3mG9VUsC95llYPMDTMIcZu2Oke05OnFUnNC8uILzrWda0gKuC8FAiMkw5
yvA4Jz+K5w3gNXYqOdFUbkxqRU5xJgWirNSUIIiotWUTH5RltsR6c/O1hSavp3Ai2ovLeOHBCiP6
5+gS1QpA8bVPhtPPm8c301zmKHwn7rWFyR99B/lYH2Ss4Qw2ijFAMALxwAmmQXpUD+a6t+4Pb6hF
7IoDtibzRwM02lT5GIK1T+1YeQz2AUIPg7dNMrgt9c4IRkZ0Jqbza/Ko6uGY5ap+C5Bq+dv/ozcV
/ST6kc0n/oh/SsUsL0sJHHjlnIhlLH+tEH7T6k7bOJxt4AskpdXa2IvcGKJyyEcM6aeh2oqqz5SM
MmBDvEPot4j/P+7T+QWZOQIVUKXNtv8ibSubkcxfX2ZiFOvDTVv+EkZK3+5BsqmFIxySwMjl6XBr
yBwy6Pu6aVLu8oV503aP5co8fTqIV87zU3zmLzZzwdPgmd7Qj2grylJpnSzqTnOLfqxZv00Z55FL
QFWO8H+cEXiyt3UkuL4rxBGGDSBBBuGO+ey+nEKeBe49GPmLtCCh8RHznkggBm8/Ds76EPBWZiKx
wlGPnDJokxVBWFjl+jt1/x29XT9HXpqBMoqtUHYkg9kwvMwp7iyRN93y4WfnzTe1byxBsB/phTtn
0Tv46/MA9wAAMmSZIfUjFT3nWY5P3VNugaAA0+VBWK1inrUeMTXFRVPHZXD1vON9E7pnAYHUQd0E
ZoU1jt1hpdFlKXftvn6hiGsvgc8d5J75CbtJ1hCVsJULFFFDZladNBTJTPeLeM4KPkZk30JJQruA
1qVX/ICsoajavhPkJ10Wh7TJGWGQwnbx2XiOL3Tg/7iqBsVxIszvbkwzhRJPODL19c5RonfVxHAR
st35N0jkFJxBcJiQ+Ok+W8PmGQMozVO+4FBsNRMN230FtkRT9oUTvpsbrggApzbIaHBB+tFrajb9
XhcerwtEPuPdwzXCLIZebRkWvLvqLba3oystviOq53fOw+7HWebV34HP4eTNKm0vna13gNZLa3oU
yT6Z8upCYawcNzB+qwj+LKrL4uQSe3wLT+F6dcOPCvyPw0cHVwgNxo1Woj3/TLjOfZZcWtuT7b7C
beXn34EP80gjQ3RWXd5pxrZavPf2I9H+KrwMuOqnKKtho8BmNmBBXcFPcai6RM/sDYy/p1XcpxT6
RG/emy/b0zW62u9iFbycEdBRCjCcWqLTQlVYJh3MXV5OfmkILpged0J6q+Ht6dF6yFZd8E/W899E
I6dbxyhc2h8W7yAZh/yicybT6LFVT3+jSnIYNX91nxxzkCPOT+W6YlYQMnhQCYYZFjD19D1j8uQt
rVw81VL73c7WOtnHfKp8HeSzML6Y15W7wWHBulu+Vmx+uHLW+XmEJ/Mtw+aK/R/7hMeuz6JAgKiA
nhlMEAR6QMIBxSybmjLkajsIoDFq5s8iD6UY1BxnskZIjxzVCMno77xvCm0y0Q/v9iTg7S2GdxVe
KHMZndvgkDPmi3rJXf0cO6eaG73KBcU3xeDA4Hchglgg9GRjTU2L30oDFF6L19EV36bYgTpuqf7Q
NNYYmIgd3u7V4hF6n/itNx9CjmP1QlYkI7iA4r0HrPpueCfV2NhymIBmwpkyjw6WH7mKxOgW2Jje
H9rXgUkt7qTWWYYGoS8UTHn1xxLMSS3j/p/2Sy36wICotst+JJWyz33lwVdQfjjNDQv3iejwyCf3
fO6EQGhYy0ChMuGf/vEKkmfiuJfZbuGoCcasK8L9Avj+EO4GvS1+UdfBUyEWc9MohENkCpis2vnv
gTfHHMwfCowKfpeSmWzgXl9iFpLXPtbN61AyTY1RU7emnHtFlM15JF9vXcPfGhQGpFL2HAt0WIAk
JoITWBcBbdA1O5IqIaxFbT3aJmG/k8Hjj/VD2Gps6UK753HUkbwpEyRm5kY6ff6V9qsnCFmHnxaz
Y+kvA0+p5xEgjXuqlHACTWmbV5/ZElkpfcB0phsM5tc4StqTKdCmk3lJpuxMPm+NwK5KpRh+bLgA
UH1PCaFRtWMf+3cOjNOztms3SonPforoZnMuz9pGf6kozcq6Ybfr2sqLvccqSd8jey1BFOj0Wczp
dPfQcyYXKV4F088pacikwifXIAVK8OR8m84Al+euqwSlHBIiuFzW5XHRzEGTgYvgNBM4aE+s1UoX
MfWafopFnrAZACLfhL+A+FHQ6lQTHIBTaRxNWLwlb9qUfDeE1X7LhxCJYEy7RzdL3fePJ/AlDUlZ
m+duTQeB09docUQXaM+GIEdfXyQh/rLHvIF0BzWNNgXKqDx0q/uv5GMO5rmdtfHghLJkDxywPPFH
hPzedmwJB5hOxHlN/aubLQeB4qAh+B7Ve94ufdmygIOFUuL967/y3knJAWbE/q9W6KyBmN8eJkm1
n7wIOqxy7yJY90r+gKBz7/8yWxNGoDJppYXfCE8h8c6G56K+DjNuM69b+gTK9JC4a+rxlo3QwR3u
UG7/Lvc2BI+HOUuKOhoZRdHMu3sbniXkRST6oS37OkDLouPTrc0lAsUN2CNUeYOntt6DZZbVlnS1
gliQAzkMzjjiBpyU3uoxFf2r6/DbuQ7wUoGHiLDDW6LVjzM+7vPigPbRdEythBddefz/JKA5Ab4F
VeAPbKEioZJVWH4XDwAfjuT701Ah2TfHuRYeIUgWNSkAxw1+0MWcwSeHZvocxS/SNylxu2zCIeQ7
J7FZ8EKfnr6rsG2Y7P1B6RwCjAVzJQJLXSp1tl4tbZEWOZ2wREqcGdba5r8h3pyuCNUSHyECNnKp
2FMlDz58ye+9uAuq/39u/9e4ytf18Lp3bZaiAQFOje+dlHoBTPyyBOzkxxsJsKjBZEOEe9SfTpvN
e6JlZSTUCR7Mjqmx9pTzMfnG7YfFBbsLx3LdT4MR+qbUN14SZjyq8lDV0wcrW9WjF+Iow6VIwVUV
YVivixwE3edeM5RZlowSZuhK9EXmJJXUAME5e+Us+KC+J1nhV1X6UXOIvHbC6Wbiunl12lTd+tPy
3Yb/GKfuZCOKZPpDwUiOAj74HRfc52FKPlbioVtyKI9cZZfT+ZcYzxHUJR57pgTV8S9XLZUdQLB5
YwGigyaC3K41onYZol6xIhi/I6JxwWS68YiJF3/Jim3x3/eZozKb+GujDD7V6zsx5zDtmqM5U+pC
Ylw7NUjjpZG00e9Q8JZ5Or/8Qxxti/89CVqCseM8BFj8dhSoVvH+WRco6Jrmmw6D3RyZIaahSTBM
3q5ne5PekZKHyTbY516+B+deBYpPknPIYAZEwvvDiubfUsuEMFuyX6ijHktO1g3jmbbNsM6oK0NZ
0b7uap1DAJCrQjjaWAzg/PMl+ee06hfWCXGz+UZ36F5iQ6Rhcpb3r/X/doYwcW0zYGc2wdazbjTt
WsgltLe10RMXjzrRXFLeVDTBoM1jksrpCFwCukfOuyssb1e6mB68o8O2AgLOFQtCLaTdt0mJcuDc
46ujbRW5x7wECZdKOOMUF7fXMoH1xwBgIHukcPyVoY9bI98+bEIlRbVd/MV+KGuEbHzaXV9s/cRG
WakxiMrarpHBUH7IIiA4YZscK+39P6n90KDqDiuxfICZAswyX6zXgrQDK/3u1+l4QDQWWmenr+D0
9lgSU9BODavKP+FXvaaOzKMQfR08rCPpQto3eHeAHcBGASKQjh8EU4sQYkc31MQMbr4fNPp2Y/B/
z8CaYOdA+FKsbWnmxfkmQAX381no+PRZsmhvpxTQy4xqotiNrAQMAJnJ5FtlhcLZnLh0gxlTZwwK
w9+e9ZDeVXWh3shGu9AKNk4/RkKGGIZxsTZbvSdIUm6nST/Gfj/ptiwtXvjAhT+XZI0Fj9HY4c86
KzPkoNCZLs0n0aLEFjsn2S3u60cSdQ8hwMG1tMiuwAR6B401Z1edkHIUW70fafWYi+duI2UoS3y0
Pdq8Lo7CPN0L86WFuKXgbp0j8m90+XBnX8mlnAfKV8w/+Dgn4OoDp7JMHJqk9BI6ogV5shHS7joP
YXCg6ptpkYTFMCl+6K5vi1YVqXgj7Dy2S55/IxA84a4Oj0tPNWFiegtSlOIvawuoQwKVccLv2N/G
yXqU4V2WzkXdhEUzuXAatU6tgNhCZx3PRytVJFyAFElwn+V9B2kH+lwzR5o2TxJT6pY4SmpKM42W
kEn6UGwF5aIDsvfzm9pGkvfXcjfwoAOl0mVS4ENOxHstdBKxd1iiktE=
`protect end_protected
