-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Z+gpFlV/MwDPKXbTJBuKTdyoQGpr1b33TfR5k93nsjAaIwAWcsmi5txHL/vDc5Qw
OF6ejVWlnILh1OhXozKuoZdjagyyLorTNOp/p7aOLqR28tPQvXHrOTgZAnkvw3PV
g5bFXcR3xtA/3aJHCo0N7cE7uT19uZqq46zv7403L7w=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 15488)
`protect data_block
VOLyGkHxehv6NhT7Y+BY+LjJEdOt79LBo84UP0AmtJBcR+H6vRIit6eTTM8QEmkL
GoV3lSqkCKqo+2mHUDjqZCy5UbkoZRtxCQo/hNfvTEzlaX6ZHXPCfmn+aUQkL0+r
Q9nrmd4bEmWVMaZMaDNpEZUQo6URNo5iYpYMKTzOTRooLO6SxvGRgEaTgmCYaOx2
ls+Z3Fri03zgr5IM+bx6LkqbQwYGy7jSUbiBw4s9aZb1bX281ievza6buQzVC76j
wORIxkNyFOHAChwyyrixFEzuaE0A+Q2HUiulJRyH8sP+bSVV440Cbafcm6mm1OdM
0VAtN/xwdELuAk/Lak2UfuJR2JKK3vqOWmGLFaq2wn1S3dn6cIzaOnC0UqnIdnFV
xyjZ1MMUMpp8C5UzgdhcnPPB1fiQoooh3+Ll55Bo9Fd5hNl+BVIlUVC91l6O3q+Q
o2HCp/HiXGdmHsnivNxH9cNMHpqxVlhCs6RcQjUwfnHQe6ma0HyHzbINKGiNt5Cj
7oHSR6qli3uQgkpOxBDhWbKMCpOCTBvpU8nz5lUT8ObZrwe7FHUun2CAnKEJmHXw
PvZbfhC123xFXwjJig9APWvq+hMAT3pweYJuGjXn+l4eAG6/9+3ApZyZEvxhnepv
YpBpKu+Y/hmMeu9voJwDfAuR4VwJoJiEr1Oh05a4jF8xzHVpmCKAOEUrpZ6KSrzN
y97PVIGNbN0y5cw5g9G+OA/xDNawOXMuoNWtZ/iNipyEEiaEMluADTXRxUk2JLTM
/kTp4O3BXhO1kbG5DGELE2sL/B4RjhEkzjIKLjk9k0KKTjcDs5BY95ZIEN/dcVO4
HW2bE1fldjce74BQVrf8j05KmYgbDTZ+NSBblTOnD3nIZg8cM8Wt6AoK9djlVeay
uUXX7wpWbhoTLe/ebpHVvBSTd5VCNVNEZjyEsmPgOz5ZxK/YB8PFC7Atkxx9rOmz
YOkDJlzG17yZyKeALZCS87SXtmEpypz6rQueCVnLUskC80ET37mRc5mueILh53qe
BBKt83nydS8MqfezZK84dHFJJBDLXo2pRLDaE49YRyuSHXwN1cj2A9/c3MYk4M+Y
/EX/3H/r1omvTyRECUJVTZDpyZC+ss095xN0JrwKR4PmM67GqHdNFKkvouG0DajA
ms6RkGucxA/hgCPOaoz/KEUJKKNdP8lrcJ+XWuMHLkAulZseCR0U0WPs6FXbUJKR
4i/KuB6G/pActDTFvRAOOcEVdtLfur0ZLLALsPOWZJ74wEsK9rvCyEYmHGVY3mf2
V/EzRoxz1VFiROJDFjcbUnHwLAPyHLST807FxZeuX14erwWK8zqMWfEWerTzR2uY
HRz9KE0I+2XjTux4ebVhUtoxbpxXmGbUk8RKxr7GJgzMIXOvPZIUyqekc61d3q0e
VUIys5XeE5PwMplAudksis5dibn3K2jKoaKF5xZgqM9gUoVfcSKfwlg1Rq+/QrY2
nUPekPPKnpGtrOLNGNQhZUwISANRRJVPqQyG73oxdE8sWmtm5XZlQjTD6URDNcGA
YTG0wqT5wUjhMKJZdMitZqlzf8lBh5pIXQ7ThQhp7Jo8Viq4syDzr5X+24IFqT5G
rlrJdOKyJm5Xh4DnQZZ0tMtdpCHNIqgm5ZTLuY0636t1qHmaqluDaIrdjBVsAIVe
RadHhRAWkvniPoBWt+pwJX+bcgfg67FCZi08dPEV+tw6DK6oTAM1zizhH9f42Kx4
ByDJunCmjqQb8EXHM+Rfb3WDT3ZG4BoLDXqQVvEn85PqTHL8gAG/CrreLbsGkSAC
F4R8L+1Z8Rc70ovewvSqPvhzXXVhOAgjC+jePN+LafZDezk79dVc+1ZiZqH0v8sV
pITLUV6shYD/gYbVx5GcITiQnqkVV+pwBbsnUjgAUV3uEieOsDMwi0ao1kOqukuB
LskBkQYTAcQDr46gkGy9i24+NYe2+rf0rgklf00N7p36Mtpa3bBMBLtNggnn4E0c
r++j6DOaE4BmfMRBkIL+XPssDAlf5ssoe/iHfrxLMjuHPx+IiBGfz1JCOjODIke/
Q609Hw1/54ApCgro7LKf4RUXm9VIlv4f3gd0jYqYBrLgXaRacXKPD0lVEnsGV8kN
Z+MZ693PUVd8SAHaJzuKvkH2jq89M8ogwnoIziL0cA3hpmGlJB5GuNapi8dI4Pjm
WX8m3NYey/2OVHib100Ge+oQpLVU8ql5BYmw7L2l9AL46q6ZukaYrhwJZch/shEP
lXqWjxiqwBA8egf2RxtkAoNCdlSQULKb7L+9A9dSCsK1R8rgtTQdLsFKMRNvkUsD
Lgj57d6w0w+IJoNWfNwkfGBm1C12i67REIt60llUNZuqyTWYyc7+WNv9yym77HiD
espKc5GxoguWsb9E0O/egvcyj1etGkH2tRWos2gaknWRVp4gdYb/ziCXxrGyiGW4
0e4MGUdjq+6HQXNZrGpPkJ4v2EmPWgwXz9UAk7IClqB8mmv2L9HigJ3MFGLWaorc
9FWhPo472X2sGP1YcjCqBtwTSK83TFcIY8qMGbsrAXLUaoAYtuZ874wGU3ZSi1bj
GvrpmrlUM2c3uLWKdcqkpCAZs9xn0RMGBTJZ3nM64Ew1Td/foaYHGvfLkTF1Meom
aTGo3ow2gTgsDX9ogaHSzKENNZu44lrRWQPoAHilLglR1kpvQoniRbHzWEx5mhf/
ByeEk7jSh2BOl6+hxJArxutFOmwXT6Y3dWmSoo+HQC7ruYyYVNkNCWXUU4XLLX5S
6RswlpZdmvehe6vtXDyq/bnCnHLqXeTlQmxWzBrdnbPyvzwbWRQ98yDvYsNJR1mK
7i8h9n7JVeGRK+tikQ2rpl3kX81VT9+Gn3+FtKR1SVam5RaryUFaHuvKt7M1QAkx
2j/yUtVWR4Ea+Cxc1VeWAvdhNSCn5twszkkOrKaHhtnynAwiqRKRI3PMPg1Z7WOi
I2CQMo5BSIn8iL8OfN9MLNUcvIi2Y3vCYlApiO6vak/ZSTPfBaDVe4cwax1kffiQ
tXu5BQcGiKKkYmiFdUhnAR8qvvpqigS2fOb+1ifoJJUVRg5+c/xbsrSzZGjG6lH8
AyZ74kZbcbMldD4g4tygXQg43mPV9y1gRWzQ4LHWuzHuiN3TelFJq4zDjV1ywOcw
vTIT0dEK9fz4sMn2WUBU1JiMG/80FLZAkxr65Ni7zLWmw5VoSGUAk5sz/bZiN9WF
z04oT+DWfQkk8uMu1tA7QEKDcWaF5ccHoCea2UKC0fJV+xpGcL7sFGndPx/QCWFB
6w+mUYBw/FxDGVpcKJuHKRFNuDgrQchCGuqSDuBukT30SndFDSAsxCFdRC90nlKg
POTgCm8XOVHFO2HNrBZxRVeELXOgCCv91fvSEaxkE51bWZyrsN/XUPbewZLiNKJe
tLwkIf0zBewbUT+Oxrgzl+MI+gbkNn4lfufJBinz7/by3gY4VcOgCwk47PxMqlC1
S57vlP3owJUmRGKAwNjeSFwVn5fpvd2U4jPhE95DKzu02t7eV6bd+LFunRKTzXqY
tDNDUIKyv1uh60YQA9hGzQqRA9NqB03XwpJNFdonbaof4+f7Lqct9xnrh34V4u3p
ba/V8usEd77oWS8Aa7KQd3wIKU5kal/Fq6kVi6PGZPSyAGq72+6MKBDfxKOBJHFy
jTKPRlmcrqJrtPKeX+28OBJMwwXFFgLAMsY9+niqPynrh9mrvDIGpIOKXioDjCKi
m6qV/xxbTs9kiWKTw1YON1YMtnDRa5PPNZZe0qbXMXvatnztUfOw46gp7+BL3Khn
HWmXCpZE5qV/GFmTF84ktJOSfmqvbqNaB5NHUubCY3W6Wjgi7jKUmRfc4bXh1/Pe
5ZgKDwJHvtVmWk6yaYNlfiN3crCq4q8ctFywtpoo3+ni7nLsQBmOO9Q2sf2umfcU
Zxi7JQYOLcuI9UJikB6GTc68CrpwcmiznxQnYjec2PYm1yVd3ppjOXbcYjhqQ5Dq
NeF84E6yi84cJGcFCgrEUqn3OhAz0tHa7DedjQqOs+P0Vxs1bwLEk0ddH8UQITeF
x/VSfZpW3Vk7gFX6MVogXCUAJzJJ2QOu4Ua2Y2hlnG8L1i3/QoleD6PhXoQpwLvg
kuN4QndBMF+K63+Hr4L9kr/O6tasOY2qHMXpnfYDpDyqwh1nBQevyiyFNYdTZouO
oy9hH7sPm+USxD4tpFxu3KswoB29pts0f9Zpabi9RRk1maZiAfPRrNfhmU7zVTAN
AH6yFWEIh09x2C/4tJvFOA6trpSf9IlrBiDPt/TCHRpLeuhIvXcPfLaGidRkZ4x6
ieMD+B1aB60m0TGykm+caWrGfqrHhJNZ4geQeRAyUTReHZ8D84k4iyK66wdAWy21
3vfVmyX3Yi4KBwW/r2e0cYbHYIvzDARDa0B06u95OHrg1ydxGtxQ9MdK24XSzMgH
HrH9e/SnG25eeZiNH/ELV/O6B2w81o8m11a7cyc8X+CbVUtZhjHsWmnbg5z5SnCl
WmtTduSXpB3ko9lN2tIS7D9uFLwDvw741FZZH2m84HZhmhK48JA1kjmA2CCxcJ+l
epTqy3vb5EiHietNHwTqjtaHLQfmionfM+BKJqjYEuYkZqG1teRe9S7terxbndav
PTIgS70HVoPgy37EWgKKQ7qQK9T/Z2Q93nuJDmlhWSp2W7tG5njFJayHm7Nkch/Q
GNibK1BIwu60XkpZ78IaWrjskOO9Ennwt/P0rftppUUMQTj0WNX2DWlUZ63PQPX+
QiuNU+iHPmy9VIlxiHqxJJNxbXf0aoaS0JAvZO6aDChH39rHZsb0Pb12s37kz8ic
Y3v36IIiKnJhNcOEntDg3fz7omQeWaflsbsizRnOknNaCFefwcUCkIStg0L4KrPe
PIlNoBoSbVnyne0mIrJRYo1uYCssL3tpbxw+VYh1wOHXDeHlSIct1x2F0nctW46Y
/vk4H2j8OxRCErSwHRQ0cbt4cYPSTsFpnwWzTqnwfFfnsKC/2rRynmWIvkF7J2SM
1eOEw5NQayyaPjDY0N1PfOWj+UAtwPehgYupU0LqLQ4SyRSKrkhIFO1k1zyJZsVE
ztb3uV49NZXTWL4ibo8hpwneiiksUl37eQcCyekAd97wELg95IW8+joeHahn+eek
tJlA0IEwLNY4XquL2F6VlOeChNXYbCS07St0l/mtTMCRXlsWa8SU4ySuVVUzm3ow
FjTM1sO4/5VzHFa2JmebbUHifchQMLeOlyoL71tP4jEHvQsg6zbN3eLxoei6ndls
miPRZi2ndbqqZYsVVTsiXxyPYkmymCwOdgpoMVAapL+yFtOl6jtB0PtIk/8Mirth
zVK98Ae2+mlie55tJg9tWQe932goaVLI+m9t8lnIy3C97cpPS8wJUCR1Fqb2lLUK
7QZXg61sSibbqgpzIlkJNimUUr9cu1D75heKDDBkgshJ5FlHrTNQkvja6lOOuMoL
T7opUNYj8NwvfQ7C300qtQb3J7u5KmjIZCjv1JU+g4OGesG5qD8PPRuxj/o97C1I
qWptX80bsMsM0/W/10uNZPsNkdBGznbx3gM45uPHoDC28xdvTR+Nxzye18NxSdK9
+CfJMBn9D0ne/2JEUxdIU7P4iFaZ0PrD9phn/udC884P8I4klOlTkpGE54/yWalu
msyEHEXO7LNJShPDEJzApULlufpGPONUElbsIrUKDw6KCF2+r+kGraLj+lxH513R
P06rPl2Bo5UKPkSYoMtdHLaGNYV3LMzHC29dYlQvSwnP5Ndc1er8fM1qctjm69vw
KC0/QsDFDV1H/lHpsfg+/k8a5j+prZFjtqhholnjGD7qOzXbe0Nvk87AdsEjaZis
peCPRK0flcSuTGSH3HZ1AXrWEqg7CxArSCc0hYjZ4NimNZG6fq08B9RhFr55b4xS
xCiGy4JeGY8sDWh3lszoFQSXMg5XsbpHBauCHuX7y6+Vn2t1ahWSeVM4UWsiYWqH
aJ7DgjgOAnxu6iFFjJVWL0HUbXt8F3yz3DXG7iQOdMVcclgSB6NMs3wy6XbtKUsD
giStBmmbaqtOI2MmhcyZ0GJoEsKKs8UD4uRVUy1MvWqyuv0dRkXSc2UD0rKJhQbX
dFzNFgrTjB4HvUVLva7dSQ30dZJLxI8TMNVnOtvRbMOrhuvvt1wtEvjVTcwV4McL
uAwi/tDn2m/waT5BfTkmnQq7XFcpOTCh2B9qGhmcg+JzI7Ilq+8SDoQYDta427Df
Ggp8uEVzAZj6PneWa8ZElORb5laf0x1mDvVzD294MzBlgtpFsqKNzMfYhuEu/wy3
/Yr6wZyRE97VBlag/Rdas/mG9uqskiJN3skW+0dLwUNqEhPGEHSKF3eVMOgrZBiJ
DHUhVeULvUqjksYydLhAl52EycCVf1JgXBHjXA4X7Aq70mbIGNnaxh2PJ/a4A1PM
sizDgHdj129RIu4L1pB/ehWHbwcjQXqllhaT1LPLGOPl+3T17tpN/xC562FkXFGL
WvffimlLFsq59SkdgY1qrxDP0SbLE0TFq+CY1EtRyAAU9eLwv2ErhBKRTMikBWdQ
HgsCtGJa+iNdrhYUl5v1v6CvKRIV9jjR60Mn9fcaWPwp6xajSz0+nJcDxP9Fkytn
Op47/i/1r3BbrS9+gwodq/mm7h/LMw7UTe4q1OU9/S23LLsZ5jmhS1pGXwFNnNlZ
O2fjSfjRkJBNgv7bhxpvz9+iaYfmsIvTXD242SH3rYU/2uokd1If2HwME5d3yktB
rrMNh6PE30iqVTXlLY9jY/xvvrxXDHMGM7WbK8Zxw0Q5LezF4BPNjz1wg5ui2LF0
96DeIt3muVby0YxMKWmWPOWQ/ODCXcfYcOhmr8caSfclQyuRYmJeejHWZzdH1nxz
SaiCFJeScVcuvjDA8gRN/sd8S7Se/0tH9VDYcNmxBnEUXX+5dC4hBpHa9uBYPq7u
H1BIoWR55a/QzoejHQ/NsYVXpfzl3tc/xXo1Q4G6ug90dIfBapEU7Kq05iE+BKUs
XuS8yEWJ4IQ0+bUH2tGUqwCIsLjumYzBs170EljAriV3q1c7kXBB0mm0UNc8VSXU
ZmWlIeujVGiSZXb//pgalBGyKyZAMir8TQT2PIs796M+lsj1GwjIeSxhdFmztutY
wXDJiKgp8uRwTO8xpk3SLX+Y3pwBqJlPsy69VSy/S906E90BeHLuTdMNk3Qagy3b
WM9DLgN6ehduZeaRG1gfrEJwnCQPsUYjVVpdtHI0YdtZKdHDeyJ8aUA/gT0/1fYh
VRjMlsw17WCM/3NU2GYCjzzjIA05Rj8xbKtlovuvfugSubwWYWOCZRp8m7oadTOn
3+nSkUCjIoMhBSIEbsYcsMkRnKjjGCMYwFrdEbKUd4dzXiVTkN+eLROXEr6X7Ag1
iX4kKTkIdgW7SGCJ9gdbSKlAuamdfHKm9bYLRSrDu+ilzvV7coptZBUz7yLqiki9
+sIFBoDeF+ku1pLZBsS40D5WfUvy8Ebp3JNRErYWnLPyDlazPNFwMiSdhZQbHzEE
Z6Jf4bMTn1wizbfhr0uFkvdPmwObmNB74JcSwZI7eMovUwWi0iaqaIasqt7XxcQN
51EuUItRC3SPobbTUBgJgqFhwElF3UM8ZnZO+6ZPgamnJYiBZzMTTXI7wT1I8uMF
wowbg4lhFmq9Ydqf7Arj1/dK1tfWSS1bIkcth2VVLvqlujjKgwq4f5oTUxNNrJP5
9DM0MLQv+SjHEtf/mXk2jWwNvW5Ku1m/JzesbLgqLaKwTlDj7qUI324AZEKP7wWI
6PlUuIFcxY7c0WYWqOBu19qaY7eiALGwVy48aFdszB1ObhbQv5NBuqEPFh03E02t
NFO0Fa/4UsXqx0RCdPeqjyqhaQdOllVvvFAH5yRvQEv93omrRLu8NQ7E5Patb1pC
BfAcC9ScmXQceaqWOm+oLIQ4qXTPzlO2mQUana0VEXjoBjLrl8PW4qkJpivjEGAa
7jmXsKYJGd9KUsH6RSLNSRtjW9tY9jWz8URsy1/H47RQnhExAcjGXZ3ON2HX9K7j
pPqumYEYRoQzh4E5DlpZ19Bg4mHPav0ZZZkkZsttqhu85Lq2ypk3YnYLfklqvK0j
G7ID22gYIuuYp4h0CV7ZjVpPa35f/AGwXyJTbuqWYnybHWy8OLJe/SObqaDOqkui
0YsXzm1mgWkXPXtGyWPcl58eoLxk/Gf+f92TaOBt47tdVqtypE/zYm3jKlepRnHZ
5BTUzmG9MnSwN+8Efir6ZQMOY0VqWg5KjJSIBcOrZRM62F6ji4bIEYR83wDZDMc+
3gQBqLj7zbpQF1T0sVoPTJQihVJ+l6qK73AycqsKJTgvwPSB9W+EEvvEDhbtoqs2
WNwgjPijBvpsW8ik/j8Q2thQmpEPAhIat3rMfyG7KC0HcrYww7ngiY/0mGr4pKAp
UXAftjLyg8EyvE1GeV0GfA+kSe1QQa5H+LGuY+rWlqlETGAe/0EAmoM2dzPB1ag/
3KfafIVmNSwCyx/BZQOWqbXwCgf1XPKC87nTAALw2AT7vSpvadU+KJELmA4SSr2C
BUUBF8ocUbA9exnB+MYA54OHpHihGA3IcgveyMNQuAC6iJBOquKkyfFVsa49jdzg
JFlvB93CzwVt5NuV8L9aqlhubQtBBM+EmQslDDlj+i0neqRkPq8PVpDRBF0u8s9A
c3dKppRCmlQP9PVhnivJGPwMYeZND5kRz3c9tS7hb/A3Hkb/gIVlF55pnfrGTLv6
vJz9sddFG7S7pR5ILPof+CEC7XhSTHVWj1QaOg4Ra1VI+tcfRYG/7hHsxH5fGQdg
ipaaSJd9Ybif4esdIpazeFmLDzB3jYEep0jCgZMoAAnXo3Aj0WaQ06LZAi8bTg+V
CbU4Bwv7CNMZpI4IEvbXifbJ6JAK4k4eTeUi0NHxMAKYM2sARu1aT7p7MsXPgimi
en51dilLi2r0k8tM+tQ3OYbjxwtAeK4kCkTj0knlmukvML88FOMMSlnngGWlEVF0
7iJlnCH2aOcjHwcJdIiol7XD00kJMncwk+09UGjy95yxRyrOXKkLXBusLaw2RTGO
teVeaghoAmBktOutzt/Tz+BGnfEwQO5k4xgGy4PnghqDAevGDhyTRM7Tu0a4Qlg6
HU80iu4aAT8UUAMzlTbp9ntwQxSyvaGHwzvgRQA4OTLZh3ZDxnPE1WZ4b4I3HUKq
xdJOCEJJpvSHAZbjMP+2wf1bm21NR+k4lPjebIv+Xfqw28Qi1D8O9TnKlE2D6uTb
aWDEy1jkB6SGl8tKNwuIf3n4Qq7on+qXsPLSbh1GrLw3yMn5JcazqAU/lbH1N3Yj
nPXik/RzLk3bLGnA4JR3wBLaF8OQ4NID7lzrSq3s0efiKmKZNso33NW0kwkP2EHD
Df2HgO78oi/9ZcIDLSYeNzxLAp/AGOpR8eKrc5PKIYVut2zP/NHhnMeS8BD59FrG
ikJxN6VLqcYJ4OG4l8igv7JjCVSp4eor2zExmaaD3mNP9Uig4Xnsj8KZReHacEBA
vu7G2H7o4wNMwnbkWg0gSgR1huEtroREbnPez/glCYioG5C6OVirSufMsNEXOqgE
r9nXwbOJVFVG+M+pkYCSkRUaQL9H1GUGf7j+Yv0jFgOAG7t5nyLwtgbBOrpiukhR
D70iVOtSz8eFroaQh4Mwi24HCT2hpm0hDP/KgPE2xN10hL/m+aFUPjWCONoFz/9b
B9H1WZmGYfBHi6DWn+tmSHiHaeh6MyFTpQJ9j0bHgowIZlcIN3FDYQezT8HLoKwz
+NfktzEGK2z/l7zIMAmgVf9GXQkiRZ1oIITaPhQJdQm+sBAmE78XOL0xYK0Hc9i5
KoKXU9zwhxI+rxgQNR4E8gNOD3dWkPn5825GWxoC4Iooz90VtjbPSAZhqeAMcPsr
L8fQmhUrSdtD+7+Nx88s3oFMTd2AsrwOzejFwL+CWju0P7B2NvxnJTVNX+PMGrWH
yB3gWsS5Ucqac+F2lfYmG1KlP8w2jQoY0V73AR1fjvHjWp8Hxyp45hlo9rDi6wGu
LzP4KARkLZQcwEQfLjmBxdej8yZ0eUiPIMfcj+So0vhC+QhDed1HCkVS7dLWo8NG
m6dJnzyHe4evPaGCXmeKdTzI9a/WKx53ep/W12xz8PD4M+oJWAdOQ1mL2BPr9gux
3RyvCwe2xCTmvgW7uqLCktdYcduiAzXs8Rl6tnGqrGlq+QeIObB+bp8lqBuxGDF6
XhdmpKZcAc3hIihjKXmP3kVLOeOHu3x40XVhCt7Y9yj5D0XDOBgha50YDphNXdo6
XFLqdKoANzdStzWwRLJQhStLrfHcRElWsN7GKGK+cwxKCQGcB09VFUWMQKrcxGE6
hUFg2+/cu0E/nTv3L96hs0mD9h+jOCrxghkbe6jm27RWuDxYgoFACmpTKIKQP9cg
zKa18uPHo0KxRy1vWzrTPD5lEAlR0bApCoS3IsOOZN8v76XPm8pFMc6Ptz0qL956
85mrAtotzPXh7plzqeYGnY3m9WPB79xkb62LRj1XdXpNLLACIvlR88W7FDgi3ggU
FFQb+0aOd99OwCgVHdkTadCSmL6hjD0XaebKwEYC8mHN03wwYKs0uHOaV1TtSkKj
WK2vWytl2TOKOBVVvvCDdeCIDo3kMVU7ekHuXAZSIGBc58MCurW2i4igwF5hrzSw
EcIkz5TUBb5Iu84CIwsajI3EuEd2pE9rvvGkwZUCHYPcfrhd0m3i2zyaYD2Hq03P
VSQ+s1Bu1XMSfqM/Jxnf8bg3d/aXFl1sdZG145BGH4OghTLPQJBKTu5dQbtL+48/
3RAdwAWpg9ZDRnLp1o/7lSYZnLlKFOzxfLdloVdIpdPWg1/gw4Kw9idNV/4IpzO3
GfVXZSmv6MyK1OFAqOykjKOTCfL/cU2EplG39plE8kbGIF5/ughf4co0IWkLKplU
8KYBv/Hc7hMK+VLZBReT2mW/Uu2Ih8KDXNp8MQaG2wG7cyZGL4gIDn5w4RbeW/WT
QEBnvHVqCClxeIyN1DXxiYG6TBcPFPCnsv/XyXf6lvle01XlM6F8RNMwJoDTgP6m
cK2TL9xbBbsSnu8o0kLyspgQVSa2JPONM/k+emKhAOzVkIwmf8SKFm8GRzglkFsE
W2xOemsxZmhrgcs9WKSo8yzyGEbBfbN3waVCa53uUaIwBbx94eh8shhftcE6ETKX
cwhLcyRfba/Tec6VdQtTN51ekn1CJ3iF5/2xhhe5ry6ZJm3X2MDZzDYdw1vvnGul
FmhJtxjVUy6aTf5G8FFKfdEnwNzFeDghxNiM00rBGWI6iCztRc5bTpKikSs2957F
9Gly43z3Fr0Z8a4l7WMf9RJ3TUc/KH17tfnS5IHtdfoHPxvz4IJGK80XAfxRt49a
6vCh4Ktikd5tnECBOnVGAE1Jhl7wYQfa1WRTwN1VCO9vtKyggI6CP0HyhGTBIzSu
G3lGR8Tc8cIPiI+xdifGf1L+Dyn+CkhixfN74XUu5DDw2MFKaHaYMaP1Uxu/LprL
THVDoH4Ma1r+afr5Ju1y0MCf9D+T4H2uh4//Yi3d56mZqgocF4DfKvdPA+nfSeuJ
IZojxI2FxxyAPZo0gEU45cHFU+C6iAOqVBnXdEKyRi/z3kcNdWoNtQqUCGJfuINK
GxL+kaoqQhuCgAnfVnzZ2Z3oDhBxd8eQFXPM2EYZNdApOFbpo8Dk72UJaWvCMuMH
fJhJoOSKzx01Q/T1HG1ea5g6YldkoZ2JQbEi+2wu/er1fEIjQ2FwRNDPv2/0Dxn0
hzC+Wxkk9rCifOipY0aSquBAnjzngbMK/HPFQJjp55NblDkimYfGl+p0uY3oFlVk
W4+VKeaDlC5Z9QULALsgdGLGa5v+EsI0xYrVRARfLkRhcqY2FgYSXX4V87FNnGtd
+olnguk+Gfxz40bk4jZEPcicd+EiXs5Dzp8STg0kFOz8++Ea6xpqSFIhAAU/oPhW
sKFDRj3YSNTVp8NYWnyB556frEfQKW2R+zcMHrkiGqDJeFL7JKPuPvZiTGAIfC+C
Q9DfVDz/nnWMTwmVQn+Zu8nY10Bs7IPmDP3oHSDiy0H4G2v4FpxPYxDoA4zIj79L
+I8o5EebrLkgRRKFnaUyzQUqArqvXEl+e4LhxtjuLjvn6nv41TcmLD8yU6SALA2X
2M5kTwqsWue/hdZyuv+mKwpppqCp5wbp9NLwApS4eAL8nrYrUHn60I20U3GVpE6s
omefJT2o3KdKjOUphALLK1g9UJidlGfAJsJUzrO0MRyqHCU4Dk9E+C+obY3L4Z99
uNh44pfueX47J41lfT5fayFCPKH3CZLoi8AioV0+tgl7rAK2tohOPCTO1ZG/ra7d
FmDq64pxjQ5pcKvFi8Qex1Po+4Mons8oPg12cJaoCKCEHiwzAb935GtE2xYNh3pi
l2yjO/jZjW+ER2mKZ8ac83Yy3A/BQHHvPhTrVnmFLDhaAaibYITOnr32TwXrbmGC
eRZ/HX+MS6zaujrXFoTf9AnXLBCv0VYAARQL1Ctt1BnnAnM9c0nGS/5gAUfoSyL2
jhE7omf2Fw1sqKTA9V7alJvIqwqqPawmXPrgO0NUImVSf1rhtA3+virGPHxZBXMW
B5iERavAqDk1Ysa/iXAm6W1BGLQcLo1YpWzNVmrt/kiTFsZQjdHM4MCeU8c3k6Ee
eKx4lFmrRVN0eY7Xx/dBVwoQ+YTmOYYp2GIQzc8yqK3WfZcxnyxrLamD6ffoqVcR
V2sIjWYTQeoFCCM6wFJWYZI1dCHEDguO7Hx/kuC9zBDUD9wHwQe/y2bSYsB9ihkJ
k/RzVZpMQmWV83Ca2Q6ac5QqiisLVDXfTNbaJ4suAboqRXu0H6y/uoSVY8otfXaV
Px9DfbelSxKQ8kvv737qJpI574hVUOdTUgRq4iyAUX5gtW6RyuVRMMLOWlCzPvOm
FsJjqrjmbh8oMdV6gbYUBcBOWlRPTRptu3zZZEPRcV+pVP1I2OhNRBEXOPapD0Tq
0oMZeap2zWbHFqUkaArr+h5N1t08GJnHaJiP9Z3GZBfftBx1qZck64gNakkqwY+y
RTZqweZZYhVp46Y1Z3tUv2FcQ1Fs7Stl9U5m9HY4WEHaagXDnSgkBoL7Qb3vsGjM
l4J7kP+pXDn34b3T6kcP5caAARgGsRi0/E0xrMbiLwnx0lPjyZ9JVBFceZa9MJeY
aYdbQPPuRUDCrzBQ7wBm0lGWcxNh6qf9hELeWwJLBUsORgdchjaO4CfDPk76adKl
o6kEQvK1ELEujPv1K0EWQNIGkhS70AMIhVqzeWQdtr/6a0bjnoxfXYt72XPtG1px
c9GRvJqZw8APe5F80nVBFTkPlOEJYMe+x2wArV8CmahlRmbWqVUogSq0YXfVY2qR
mwkTSTzMtCCKmIijRwoWlZii0tKWPQbylF9jVm6wgW3siVWmcpHBDZ83SC5DINL5
GBhtGiFvngc1tQb/gBc3YKb9C/isM746QWGAG8q689MkDoOB+kGPzRo2+XL2oDGq
mAsHCZ0XD4G9rJh8JGewwYlwGizsN2yucxZSBn3tnk7+J+WnrwviWA1hs6a7c97Y
HyYZ1c1QAIItA2vEC5o/fPJHA+cN5idD0VRsbxSuj1pTl1jKDz6CaNMN9VgSDKxx
grHWgifVFYVOl8gBd1m0f78aPM7/j3Ps18GdXiqFvtnWDZ6w+GWYyAnF8UBMAago
9O4mxsiYMrUxI7w7+viS1DRT2Hl512WMkpEkYqjrN3ulNZbSdIMPSJTpJlnQ/Yjz
3RQqyraIOnTl2JWRy4MnnKZqNUtSCbV7cN66SQbkojZz3bAHk/cEC7RAAP8BT1Va
GnVSSHcMbeSwFcTDsTi8W1Qe54e9hBBhCeC9ZiMwzZPeXaRnRwDLPHRSxH3mkEfP
bJtKzibgtaR4xvLphGSU6EklFZgsuR3A8/7d0nLg3UEeZtK0A4RA1ha/LCOWeXyv
LSoxOYc3bJz/AhdTXmBHts4mtOlj3jFct2SV/bMXLt97xFW0VCnRmHU7ve4iFgsB
wcTe+mkFnlAm5NIULdM/vH0+odkx0YlvGjk5AlkoBfV4Ko1Qsa7otTX+EV0k9wLP
51DECLG23tkBJqXV4ocQ099s530hUsJrVZ3xKD1XWJMSe4mKbvlLf1WaGPSPySu3
xla9jfiWMDrkAx2XBIgdRSvfT328peu3vmTch7JL5fJZNdG09Xz1DuY9SbZ3skMV
pyqnt6izhkNLOEOL3Gp1i5oL1FscxHeMEZrOmzWU+lOsMnH3AwKQJTH+2fYnmSn7
/Msh/oopcId93OVtpINGkIv5aPRCExmH1p6Qz4gjvyeQuu+iZZsR2F/PV+gXQgzC
uTKjzAMyFCIoOWJhu0E6tXrst1MYwbObjcY3spHDQSbpfqc3JTP0RsPQbrgFYofG
N93TwOMUnkijh6Goqjy2k7V00EnTLOGub51sHkFWBRE6lQRddNDTrMBEqWvBYlqK
D/uI7tv5QLMWoEaKQx9t53S9cHcv7zCL5O7S5tTcw1noZBIKINbfFu8PEm3A5Lpp
uutKAPhjAYi6UyXmYosutO1ApF1j5zkF5FvZ6lo+5cnpi8+OvqNY3Qr9AoLB8Ayb
usIiphhyswRjO/lnmYjp6gOPqoVtArz+GE9/cDMVhPhf91fbWddkBWGpFK3SbNjJ
CfhWMRjm8IpmB2PsPvsqqSMOMFL5vaVlCkXZqdFb02L6hOQnmYbPIirlzEwuYUX2
q6UtB3+Pz9eakc41wdyaIm+3zD1haf6nZSLiddf0oxjL8l2LOFVFQdQV/gSZQb8H
aHtSeOPaYXE9lgjytoKcdu1nkzsNkhFwp0DSktPaOtRD9EAlvloQKiBx8MVJ60el
svW3n4fLs57XMUVJ4On3TMJFaCxksXCubpYCxvMqFB8+7GjhRhrsfuewy+9CUNZa
Hl+5In6X/F4IVT2F8wzK9e0yu3cDo3cgpJjoaY0ld0FoeuY5Ds28Ws07cCa8+bJz
Xdc/XIy/45yqG+ZJsgB9MSfFX4u/3szva2PGvMjILkEDMrQSVx7mAHQwXPlLbJP+
4Q17o5K3oxCwUqK4w8ZFRoVSoQpq3wq7g75OMw0C8gRsjbg1rgiKA89RG3DBD/yG
+A5ZFk8NJds/xB2dG47YFH67nungwjazPHs1Z1BurjBnLBHpNPUpn7Kd8BoDPR8T
Go6QAdTIa0fnLwLQnlksbBkzjC0uL8clxggFaRyvEaXKFbYuaCZANQCL2s77s0d9
E6Y+kvvPJjsvpRzDStk0iV5fEqkq6YLyz8tGlip4Vt83J10AK0/Rw8sCTIcqTfcF
d56MU5Gj/jGvBYUzKe7OHQvjVHv3b3FAUKtJG/zTAiGoI5lf3QZy8mUfWojRcqcu
bmiJsK32uqCzdPkb+HCisisMzg0H5pVsZAsJak+SuQ3+HcXoZxEmUG6kiNXYzbzd
b3H0GnxhjXTXelG/ELjrzhsQ54EIlCiaq8TmvMskef3K6omkaddL65HewxTojNc9
9QWRkL98Xec+UhSthsbbnDXvuBN/I/3aN0XZfXgihiIvMQZvXbGHGGtVFMwBP72X
fS1XzIsNzRuj8s+oPUHWEPzIEKbk+ZYeh70AlTMuhPeRZKwlJ+OWIP9zDWZ1VU9X
Zs165XXUVhTWUkE6iwtZ2afylyIRYQyjxZMyGdqfACxqYpWYGIdOMZlI9Mmb1CjG
6Be27lHB/oQH+H7Yr1io6cAzVw43mvhLeFWZSZukVYk7wnzxTTU8gpOPKkGaf8Qg
HwX6xyLLHp2Rzo8LP03ISxgxZ+TSGlOi5SMFEYSgSD09fnW2IitcJxf7od6HfM+f
UFtrmadKiTbl9EJjFLLKcSkQUSK7OSh3HhKeg6U/rzeLbjrcC/pzPddF5ppasv6R
VAtgTcXDVVK7sYA+LJBYiPy/2qtNfkp/ptXxseIiLf3WkNOmfdJ9y5BeEchDb4GO
41qA3DNvGu6uX/B4Xo28v4a74ZENrXLULysVwYhwGeGb76A4xR0R5NMrB+hw5J9B
YSZ6whi3RmziB6XzqfDVUoZRyzAkFPnhLCxUECq7Repcznk+vUGqWd816ue8SmlL
FgWRKsIPU26B0fn0YF1BU/85TFhIJGZcb+eJGPeXX9uujwKi9PSMoAznixGGLbsG
YzBU4t2TmwmTudXhE3x1gHrq9pX1rjYWfAaasjfdO1lCvudUZUhNjGqsQFkfXLaJ
8PxeK31bhhHPUTL/WUbIkk6msCUbctYWaKLvOX8lmYeFSFDEWUL2Y/RqTtGhu8Wh
kkWEInER1JXmojxBcpUi/c0GPlKbY9xfiqYXPLvtPRLGPUlsQ3J7ePp0ihprjNBM
VXXyUihJ43c+2CkcZ1Y6gfVN/YlaAZQqSzTQ7Qq5500FgNz07s2dYz9MvBWWv+sw
YQgrAORnvwVHLKvBv8DeooGvvwi2mNKNHm6+ZkVyaC7ZtZT6FcjwghxJEAXyzSNN
O+INwpxAv+Mkx/sbdwVE+61yfsmCDjshu5Ww9jKRcAimUE8g+LRODpuv1s9l/Zzq
RvGC6CueucXcES9vy1UbFwlIoHnT4zn6B1O1YSi2KCriNaf/wG2vH/KY4jwO56E7
IlRUsNWEYOvqPoH/pa+YXMaHHYTRQpLap1nsvY4Ac+7C5CGweVd1ZuzXOBDMDyby
lA+BH5PveUMQZ6ElNyfftsi9GxBBGk27vhz/vl9jL3PW594VFzWd05laFfm1SyMG
q+XCri2i0Bzdz6QIA34zDtg4OeZQgdJNK7RIn8ZlHO8bQQkNiXHTd7/kFji6Dw49
UsMzgtyRFrOslnIIMdaTsX6EShjtpmFPmPdc5YUcFpOcJd5CNF/dRU2RXposSz9j
1jbxAZ0bjAPpfxzzRqPXY86MAIC9i3vy8kdt+c5BTJE7n+QxRfpuCk5B0C32K8ry
e5E8pqo3AFT7j4LP57pzN2f7K0iAfmSToFp1fDeMjL5axCU+TGY8v7aPnM4eEFMl
BcXOGkMlTM4wB/rbcLdDotZGOdALhRxhLkt5zd5ngpnrNz5do7dHMo8jpVrLvNz2
i7aTlp1NWz8aObU4m4Z0OsmN8r4yTKRJHlHRqrOZEhJXe3X6l+D/XBuphYVi7k0+
QSmYUXtTCpSqGYVet00/umfcreZ46pO9q+/aXSnfYpWQCdu5Txq19AxIKpJXQhTT
6aHGaH7Fg/KQt6kNb/rOhaAeMhIlfNzEpeP6ZBBWYZRig2bx5+q6cBQmu5JhXnjM
nHMMPhvjLRtnqJ/LIwNbUeV5BpqH8r68DoNQL//amzPtv6P7507CO7i/YBK1sxg/
44ZBYGl9R2N6r7gBJTh2lMk8OIYB7iZY6LUiWXJAHCpzbJfrvLcRfaf3/okqnrSs
2yHmw7Hudg/Co1jgNu9la/aqSmRbirqgpc6nPPYxYSr5HF8ljPQr+9seVP+36FGF
kjjfe7DFnuNDfCK1t0r9WSt7ZsUUyt+eubfyqYupGn837yPJESgLumChsjg/4F6e
o8DFkFDiNkxV/Agmce53IYt/c9rwx9rFIua4s54LoyOz4+8PsI5ls9uOrplu6ZQS
U/u0XL0aYnUX02bwNkjsxq4HRFNaENISZsFvNI2zagruTBjH9xF9RQG7VjP7hQcx
8zZa4ZHXRaCRWIulLoRtD/Stva3S4BLbz3Ca0Rm5Vy4y5Bml1gZezjJRmCygYe+t
mmJ6bDjiY5HNd1rEks2DgYiRsPPsn0FrCp2X2qsIIm4Uz4u2nxyIhhwLjyFK0B38
hZkP0UDtgoNDJK2eMHpPk7FNJZ9M+ev/IO8oJaHofhMVF6DInI0gSGVijB3dTx/Z
uQBbJPIm+3jco0M6MBnwdCgKz+8YYZdCH1nFvcaJXx7mIwmQzCXeaRnCbf1aGMoM
vwUmZY4/e9bgCMpsD+FDhgFDYMqtzI1imFUV3S26wamODfCr9YL4MN4323K0Iyt/
GRsjDBk2YxL5MUYUBuVZTBjAbsyflM4o5+P4BK0veWh2v8EZx+DHFXzeC+xkJFbh
ud8ADLiq6b+u0BhxwZrUqAFFvgJ7Kx+gRsNAwlWZ3vohwn/DwzIMHoQdQAWoLz7l
i+FKCCqz2UOEMrOFCXTE1afsfon3Gw2l8YRUXOi5Aoj3cf5sBHc7jF0xvzHKtd2n
Nllt8vzgl5pKj4pKJTt4N+dTtn0RRxBJgnAuzr6/1SxhujVJoSHBSXe4uJ9Y4g8i
GVX+dGJoN2rZQ+6lIIeX5VfYvPCzWrWnN56lJX5yDNW5lGFR7s5bY2pmj4Xzkeqr
Ef7KcBoCK0LRZ02bxvUrUmp1PfrpSihGBb3/C5Y9IQr2HIs3PYZ2GLlHfcBPbxza
mt16wQ77vtS5CI+ydjNeUm9oI2NeWtsvqTVO/UGndx9GjaHUCYpev9+EJ7wCjB8i
C3DINmSIvqCyCTCvuj6jGP2fSBL92A5DK/U/FTDicZWOUKQQ2CJQkfHsQ7gNzAee
Q9vWn7w3975LlPlVWmQ9VlIHabV4SMZ1B4+WOetIb/LYR08H0enUpi2pY1dUmdNT
rt/Va6Afhyn1+sh+xDr7iY1jWT/Xt6mlOH3ZdaAs+Vk2C90ePkWCS4EclCxo9T3t
44CnbI7hklTeEfqB4mIqTqOWvKzEZwQu74u0JeBnIkgn2atAXmlaGPT/RJlCpCts
FYnmyMPbzRZvgkZwW/P5RIbuXY5UNhAvYL988S5ZsvGTMwMXWBQbw6SlXW/Bm9nZ
lb+Y3Gn0Fca3rhBCF4reHMuLwiMJYx5NtVyb3sN5zjq3kRZ9pwgBPZ2OuQGj3Aqd
HnC50ASSt6n5VW2CPJmlv1HV5srO3GBybumKQq1IjnrDbJLXf6Np9A1QvkEaLp4h
k0Oemo7foT93wLY/DCsXcuVDPU0xKYMJoOjUPRjYjaUycq/HsIll9iuCExp4gOgd
lL8ZW9QCzxvN1BmdUML7+puUfsY0AZ2+JyinFCkSfApQTCVva6w9122zqv6ITo1h
FQk8nF4Tf/mFhlShtvgmAw4H2W5+Zvk8sN17xnfPbZIzyqHOH+mF61QOGf5tgwBG
L7QbxQBigGgsdJLZwOnpHLN9xT+AkqcGruyaCikk2qEhOtlVkdhJftVpsb8JMnBC
GazcjIQFQO1l5+yzx/pk74vRQz2DmwfbASGW2OPw5KAbmgqS2GHqaBp6fz9FD3mn
N353VhnyxW7MUfVZenwN7KM383/FWxXuVbBnHOGAZHneJo5or4QinHGokuQ375oh
GSYAHpwTb1P5GCL0jl4j8v2/3tMFsnkTlCKxYC1G5s0MiZG/gCutDrghSJ9wQw3g
OCVncc4WtXfc36GOrsFeynyJNWxNcTed8CGD5G3Pi7mc7UnFTQre2FwxeSXLN5x3
wCoZBJfRH29WbpuQvRpKbWRC+ll4alNGwcULPVtjvPF7kU0Iz1CEVdblP5jjYcg8
9LBhBSZI4xacWZ55OB93Zjf/6QSkuJe596yjCTHQ+IrobZPtO3LmFU02U84fSueb
Zi5vY1K0N1DkxddljluT2R4m3/Dcnjaxq9gNot+8W4tx/mklEsPchbtBM14Wa50I
z/W6f0xsFshK+G1bpS176zz4zPj4eXDGm3s/4dPSMcxncFFQIpBEP7Sh1weku8oE
87tqflEwGP6WnuWIF2W2eshSLNeNSVxYrVcz1Y63EyqE+KboSA5RcCHJlfGnbykh
KUvuuy84GLvmRN5bMqI58UJztDQPjahelv38VW0ub3rmVIEyXyJ3yhyUmXyHTB3H
Gndp2Q54PZsROwb5KcPQYPlofMGhybwiUDSZ6xV7W47Es6/yA1p93nHfDDj1fwKI
iRUHrCAm1HN8AQE19mn+1YT0OiV3INBR1/r2MzTFWECSWGknK3acSWOoaWwqrVZj
5bhFh1Bq9zRMvgn/ZJKlFgy5EVrc2cea2H52vGJcKBP9jidPb1kbJqRkrUwRukcv
dEtlE9dfMF6MNG+X/NtGrOaZcPSLLNlhO42RB0Fwu2Q8R+Fb5HgywGKY1BHoIhh1
KYGT4d3A59dm5UfNmLy7PYbn4TigV+iaNMqH0e+XWQxgYumgp6XuKKAnI6HeqyM+
0KI613dPpzCsHisFjyz1ufFjokvFB/UQHUy2ckZ11HPoWONo5UjZ+SpBdc7PCpEz
h+2ydlH3lToySvIpCNGGWuPe5aypX7unizn6cyU5WBtiYEs3eBHnpuACKMmuBS13
+xJen/MwEuvcN9plpl1Ym1vTgqxpAmz7G/BlLOixhNRUqpTRoIN8b73HhK9kfiVA
T3cg8K/0W8YpFYJJVhA5regXIsjavS8ynEN60DSjMEPnmSmNXr/LOwbj9AAwyI2l
E6DXIqVVW5ZSzlG3wFrv9wOZFGM9iTgLTk9p0TIyPuTJmPGU0sg2Rd9o+GoZqo14
kRj/NjdzacrgcozVBEcwNiJaF1laBOP3nbUMwfWQM8joaR704HlSL+XJXs5eJ10w
T8xfPj1F348moSHsqY0+4CeG/TS4s3JyNy0jFWAQks8AUMvUJHKSFG7un8LyICCB
HZmhG2WB3RtyaHKdtW1+U9NmYXNSe4IKBirNwRcaMEpcofofEUaaMJyC9utTkU7d
7MLMmtl10QzeNhDIJXrxD+jkmd8R1ZUuVQtodMlPnMDTWvUnrl/W+ouYq6lmiOok
+7HSQRxnbX4O0LJ3H55kWehoxrCjnKQXcpSP/VWHNrBWAz3K/1GW177JjKAcYVKj
1rEyG+EV4TNxBJxHSy1p8JRxdOmjdXncFvtl+fsQ+gg=
`protect end_protected
