-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NzndjELVy0kVKEmIKCucqnmaGwGqKkVdL2tMuiwrwCyMQ8f28B7OTpmsPauXh+H7GBF1rjT5hQ3G
60nhYvRsGn8CpfcfIjEhUy+ai1IIvBZyaUF65ZcJKcIPgUJJnN+Ja5JOI9eipn+JREJ7ni3q5IAn
mrQ7jwP36I+fhQ67M70QFlOQtE2C+pSCnUwYBFMuanVh3XtYu707zzOmBfoHX/ICUJSMu9xLFPfC
90+s/t+M9MVtLQNXpsm6HDfYABPcOnifgB7x/aIinbMNWVYP8VzPqbX2B52g+H4/bMPFZK2PwQV7
ZftE3nMqD1laVYX/sp22lFYUp+WQS2GakXJvxA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9856)
`protect data_block
K7Tja2MV9r1zucsIBUlVdlvccpylLoOmvN5ONgrwMPKMHZVpX0b0VW9zBtDmv9ojAblu0qTr1A9F
X+AjISoKBc8EolKyaxGzNfkeT9GbzsXMiwdfQPSWmDIKrUhKQm5nNEqhM6o+M5FKdV1gnHV+dkZU
/Uf+6dqOFQfoWQ3J2Ow17tBFneAbuVrICv6WpNP1uFpwA8fTx42dJpX/BdE9WvqDdYSJTu8O7Rf7
T/8RzHmducNjerfHuSPFhgqD7iFiRb6joWW0IYe7ameEIFoLooNuRC9nPjWWcSL9UMWv0UXoRufI
4RMRPtL980lxxAM4bevtiV0o5keYoAE8B5M+UBZMmlMgPQvBm5V/b94/NFSxNrsIx+wcpJPKybee
uNgi6xRVbB170QqzJyw3+J3hESHTa2wCR3FyZl5s67vQAl5lap8YXEbAuNJL5r41aCh1wkValAPA
F0i9uBOWvtzsppZILhUUsZ/2K2PtEXIIhHKHKkLpVzFLTnG6RlgjMAY5L++y+AJh/Qi2tSIDVkNk
iB5DoaPqiWZi31rbDtGbO2q65T2YCUyn15JMx7bYQ/E23YMVsD2kZwx2oBZvGVYIi+4K7CVgNL7l
9s84E7wQkXtyA3fLOu7yxZUDr4P43wBevsEvembGCOaE3lcbtHibtRRBBR4mUuwdVpdHv4RV565F
WKjjxyLIQm3ZKwqUayj/L/l1dmAAm6uZOmuwgCpCr4KDWSwY1WB+kNya/NGFcUtu9jV6CRg09h+r
FnQViFK9/3ICQ9I+3/Ikb7OdLpOcJsWWEhubWX+0D2W4s8OpgbB9q0U42BXzH+ak64BkU+nT9j3J
ENUEXIIfuhAETz294uqg4+Ouw2JRzDKmWsqYJw7RWAM5G9tbS+iBpbYn9F41w9XnN/2+AXaw+9Cu
STkwaamW2VozFG1AUXi06OZmy/MBVIpIZV6cGwuh+bRnCXHvRangg0F3VmfUeDl6WmbT3PaJ8//d
yKulHlwb5VUKfbjiOvAXiO74Btwk7JK1IsXmq927zj4wf0tBYbyx9DiK99C2nWLy4UjI+An7A0tr
3s3tb4E/tShELBmVwzyrSs6QmcAEIr3boqZf5vg0imswC/OPCCVbhUlj4upLRg93U4NaAcr/DWgl
sV/fFNqEon4tNPUfBK4haTdB8jEsapLYchS+AS8SUNTDdsbe7RlVE39sHFe+QMJQmOvTEAlgw4gy
kR2fnctQQ34zbDxbo2m8ZQn5WLZTLHDBFUl1x7n616NyRoEsISUX1VSVn+yrZLBu4DE3J0nSBvP3
gOyUYcshuHcWpemGSCx8YGgK7jZXIfuM4ZBVTpamqeCWGxCQH/e+mjfahd1jdty3RB/gSfK9od3L
05Hto4Oe+mm4uJ7nqLN1NpBkmt4p4l3NiX5nuErjOGegCL4U9rlaMkcRGwGmaCITf1faOHcg1VT2
4smDcpRbPUI0zh0uo0lRXJMWTaC1WHyEAkb6jfgJy2ZZ9Vw0dlD9Mt+kFnBmIPNTJnZH+abYWHIk
QR9io2Bic5fxVNo8CAuAKnWAnxoSBRbY3tJ5G9YtT+HKb/xT0lMmUmTBigwyFmwNcC6OiL0Pl2cD
OEmQICHOf5/RqkBNAEaqhdpGW4plpvpOUXfqMDJpI6vISooq7ZBZ20FkqI0z/W6VgbDAU1GSUANN
7gTRZ5dci02PdAVJYfV7naOyM0zw0Zmwt+3pVdnh0mBilkSYz+pxydFcAioZ2MtFKtb+8yyiwO75
qoC2LjSPLh6CrLnarDPWZ7rPSgN1XqXcsMhM/aOhf1F7yGKNtiUC91CC3yEOguh55h2hIFaBTfEp
cbHGvSXch44FsXvHfqr7vFkYwwzaWP1/uWl2+KOI5FhXpJM4QmqZSzesTv4oeMxn4AOcDhRFZCvl
0u0UpkEyEAskeQU7LkvS6YqjTf8YljcGa0jV1LiUjh4dRdg7mU5XhBR3P5heX2HAcW0NKiSxiiMu
f99oMwRRfsy6YxiG+Xm0tS+9VV05imlmK82vRYKxrC/rTt/HLynizvIBlLCZPZc59cRDVOYgv393
uqGhAz1YeCpiz4yo4nwS4mPeB1iDkAjQ1JY5dIZUeJ4APpoQ5YR0rcPLkMO4PcVdlB+T7hAlYnZ7
kZt/masDGcBxupwHkM9l8rRZpQNuRfIF55oEQpPUsLRt8lGZJj8y+qTaieJ/54/4NaPFipVfLwVM
uGleCloBTwVIvAarszoPb7Xa1r88lDLQBCZHTbaxt/zyQiHNKahDnmc+fwbk4dH7SaipDQEHDtp4
FdtEYSoO+1vBD95nqZqx+YF+VlCqKUMUQE01pW5aSbZpcvb1rVKIDnG8AMJtSURNuD1Uyr3HxBWO
WzOZ3ek5nJIbo+6nnDDvBtuEEf9t0vfkMo6e2uRJ3UEkzfDtfXkxp0NedhZvzWg/TVaXG8MXyrEY
fIMuxZuCXje0pKl64om/kKdNgLa1FzU6r2upe2/YTLvNKW4P6fGnDZy3clCr4fE4ife6NwMVw/aR
N0TPi/3OkWkwqlprmSs6oY4JuCU5gci5s0zVPAy62e1xUN9bWD4/tGKW1dUKI+gJ+T5i0IpB50id
iKCiJ3oqgC3eaT8YmK+Z+bDRYBu5vZrLmTmirgPJ91zqDZNRhnxaCe5x/Q+IyDmnWOrQZbn54q2W
fKGn2IC2EfxTUAl9SBG4Fh6CsBtBpagyiWdmEJr5Z+q6bL5eFO8EcsrS+wS80qOnesXouOciboeG
ZpHYaymU+/GFQY3xPTcKDDtMAayAD7aJvGxKkpeOApFH4lS9S9AmT3YdZpetDCIYH0ErIIAOXAdo
ciZcZe6zF8zls40OwiGJlsonsfOdsZcL++c/ORpShIBK4jsQiSnUXlUC2T9owQ08/8I0nxERKZ6t
QfGroA5hpOhQtvEwdNSK4pbGHNW/NnSvblwZQLNZ8EexFma9SVPKIO9fqzcHjQLPSNKWFMYHu/4x
mGSjISGT+PgidN3rrig2uH6RNI24oz89X0PLmvQcr+WD+4e7+ti34bqFjsviJ+wtXYZUYtDI5mY8
etmEOwBnH52V3+A3/pBCDQoIqVK6Z8Z8plYF+L7mjswf1ied+KXm1bAvov5NfKvl9p5jQJdMovSm
4v8U5ArcLnid6UMFCcAxNCrE/AFvV3OJZXm5oajquDWxI1PruGmdUeloVryck4iT1DA+93f1Mm/d
Xe1BfDUCyQeSSxDv4knSqfKY3tRawmxS8WR+s3H1Hc1yJRj7iUQ1sci9Zk1FU3tDpyB9WkyFSQGg
WQFSUR7ycpGCejgq1M9pnKfnu0Td/UyXl+RFCuU8wQsb2Dwz7P8zxndplKBF1ebUc0tQVHrysLcX
6Q45ca/xK7xsOu3EegCPcgY1ONSrn6BNBQQO/0VAyYd2Ckv2UOKlwbXrmF5yIJiJbL3Nn5tyvB1s
n0Kl8AQDU+G480eP1yyD7ahhkXRxO/hrYNC2J+4ExtbOa8w+lLxGlwZHnqeWeYvwIBkrzrYIPBKA
sY17TOSIvPIYrEFkbHCSdc2qDHDTx9vuuzJUq9V7quhu81rPfWXQeuQDayIkRGDwstJXeooIEERp
xL6PQu+qhXCg0g0VuC0o3y/rlRTmzaP6Fa4vL/VdYuM1tM/Jr6m81HL1mqk3pv4ZW6h4i4szPCBz
yxXIOHLvoeKFtUJQinQ+e2JWWC8ZCc4yVAuesTk3hRQWr/e4SmOtiLJa4FxaF5UVikxNw7DwAix/
gZsg97+Jn6qE+T85cyJZBR18ydID0CQpunoJ1VKjdD/kFrNKtFcHdnKaaaOafGDO/qAaniQzrI1d
OErWGx1duO9pLMPpazX1YJG55fOTBq6wct5wWLtQVPax0Ay0m34j5sDuWqQwyWWSnIGnqrX4cSjY
4I9Oyzzg9H2xseVWJD0sbZ87VXIefSuFSC5x+75dyg1NvPtMb+JWVE73iZKkfvi0OC/0y8HfywAt
Uk8DgkAJ/KjAGiYWpivhL9KlwoVbfdqbnH34J57Vz908pC6q4SHGamRlUOsh0RZVhDQwv0d5W4/D
2+qwxUqWEk24NgxByHnAFQNbj0q6WU/S4pkwKBAbqscj7rEOOp1KM8K73UKscAJTC9oLOlYvvVkP
DX5d5xdYQ5peR9+WvXkuze5Y+yajkvKWnf2e1cTX2UqKHVVPPOODvgUmIz16Rg5+AH0EtWnmuPE1
wMGGXdMhy6LW5gz76/UwiU3ZZtng2O8vJvWW5Sxtk9Qdn/PDzAlaZ/FsFgydQ2ZebRGOorh2HYT6
J9yy2y5OLK3DwABMb6TC6rfUNMUd94JuvOXYOm0OT5oOl1DSUKIbgVbGRoIvbAigET1Ykty5yAU2
sYiR4cT01w4GXWFhmKOQG1v5FXuazzstY8WsUjrUvr7M/VRDihP/z+oOR5XlOSGGYa0FN5WCJs8Q
czGR6NuTTeIN7eCm3+FSLVakwKCpjhO71at4zjCjMcxPaQUr0vrUmnS/7+b//cY18u1BRuYTBnE0
KlrgmpducSQMahYNzltVDLIQFc2rNb/9pUpFKHr4THrqyBlAN2fHDDJ5su1zhY83voUgmRkAluHS
aYy2Mski4EBLuuGRGDHBekTafzi+gFIPaWh1oMVWlJPhM+BWNu9Yi3SORPAM9qKdiy0C8ihk4T9L
uqsjDTxlwGoNiJvXS1yTVuEClALYftM5jWAObL2Et7XLKmIK/LxtTOeaLtIGEp5D+3KApXCzixPh
GiAadFOC0t2BlIlW72SiByAv6tWxkbjf8E/zVxT8H0QDcmOHXa4N62sDcrbRg9mdPoQIfzyV/gFw
BtVXAs5lDbJj1AZYJsc9jybLeD8Vm5V+wHC9Xyx1KBaag5jCiQ+lI68V+f2HvbixrdnZdN8Hh93X
EmUxyWPMnRa1hZeacQTh7n80C85UAgvdxYIRrTo7eqC+TKUPJMaojEHxXDdU1xsuwU9UsVu4Ojkf
tLhNCTW6N25Nb7LcpmZQDPnWHppt/RQUHSUWl1jjDw7234T+263QTcur8oAAOTu4YYgc8cziQlF1
Szy8a7CNajSAe3r5JTkNwoMQ5o6gtDgJzvCcQrSS4KS3dw9rIRe+mn3MUGoAnVouvq37/W906fFp
kXpln6bU9PUOQ4Mgq64Usdloo/afFqAUo2/xTe5KPzHCP44FOEXWpd2aNP9uEV4c8LG9k29zzGSC
D/u6a2dVsS6tC4xWnIzzBgK+6hNZjezHN6eJLnxCZNFb/KvnS0b96gqMtBioiYDdD8BWEFWQg6Pe
BDVJpEmOFMZ9SyfJv9cbbrDikc0AtSlHz/Q/XpPMJgw3ggBh6ryQ3U2ndFeUD3CpkZzSWfnKnsqx
Rf7Cu5bJ0TW3toFaTWX9X5vJCRRfyB4gbmK9C8xBaNMtj3GvPOeVBZhq/GZQ8YNNZRuhoI7EueyU
yLTOvWp8w+GJClzcJWhOu9OIHaHvw2ysEmZg6Zh+IvaYxbb/tUJzjOxx2dH/LWSX9hlHsjwUTs9l
YziMIOtTTwvtJxpLTp8ALJNKUFOxilV6qR4+moQW2VJZa+mgQgLiXypIgNA0zZ3c0Ejo8nNwpm1L
/koN0RXhA7/+3T16tZ2akIUmBjTYgsShNqOq+nUN6hD2P5QPxzJIqusd9Z/PXaUBI9KQ38E04ZUT
Wr8BM1a0y7P92KJIcu6LehO2afFM23lM5anzuanxcAwO/y6x4IS3gRgk4Y1jU1q1rXRFr067PSWU
C8ILAbil3ac0M3bcHpP3ogKhIFH8gJP5Ztgb2HPSl2LFQY5WIlukaj2TTlZB6YlBQ+QkCyBJuUlx
StQ5ZDxoS/ZO6dFm05mgBDdvkPldrQKh+qnat3HRuxFJzafJqlwpd1AhnmZGPa8wdSKTNMmA2bkO
cYMVmhn4zNiU7IFd8i9qAJc42l0RNkO7d98NUoQHzE0b6K3dwvTMoVLT43y+V5H3rs38DSjhImYu
bEsXJu0zcHmJWtf+s2+iqn4tV6g7t7HUBInGsv7fiVXnbp6E1r300F7vtbXAMAsTOES1tQpO05nO
cdF8cRc5ItqrtSmbEN2Jwj86jGGCvyTr8g9TB4ph+w/T3HloPmzU8pX/C2tTTXitPyORQ6FM0yFw
Tw+QpSa2jR3O1sW2/VHk7Z+U63Gi6wUvHB/wrFB3IjkzzVbbQTxi+XX/Y+jX1gNkqyXzocS6I/N3
19TWrEb10Gv90izcz5nmTew/cB3P3+LoS1+CPvbueTN56+AJBdXBdL6BgOu0XYwoWdqI3Lo7Vhy0
b6zkTbfidYV5Qpu+v8+so9rNUeiAXUgDgIWqAbs3ZDUanE1LPw0CfLFcJXRhILb1eADEU6B4Q+eX
mXfvl+eDONgKiMtq3vR5lZ9wyrhGUTcK8ejIMcKXn40Y0iIS0oRVudc2E7ve7OdmYeR0EKYQqhKL
9MqLwhuQkUHukZ3nA97jjmp0Rkp6dDl9IEEtP8PONyv2gHXabAzZ6hbQt2rKPbtsOhyICPst/nCI
+XfdQBkx2YI6+3p2/WvTw1yKlMfNotYV9tfFRjv6fSgk8vkLWwea09a/kzD01nZZ8xdHy6hNwKP1
n3CcYN/EJr64b6Dv79EhZTnrnnWkT0n+f+jnqSkjT4vxZ+4/huA5LoH71i1ieIHgBX2Ic0/B8r3h
wSi1GqlLsR0R79MgNiFoEpdXiYlW3k1rHek2iDQwhM7PCYx7IeS0OTPeh6BZQM244jANl+WYaCPr
bGfzZGF4e93a3fVFBoKEH1x7Js6Dn54T+w4gvCGnpOVC+h1Kj9EYrxISJEZQTwRsiWqKallM+0QK
M9M4ZuGPG9YF7jwk5MLlKJcAaJAOnYMGStLzGO5QHXX9WLf7WkEXOk/qnk76Rqfwccu8vPHu4w8x
7Nks15MKONg7RNplyZo63vdwzfk6EbxIDCjAJwe24HI7TwwgI5W84B4ouMJKD8A3DVb83XmRcIpD
zkYGQl4ybqE8jdfyW5pOTkdcjpfdFxopwsyf3tZTMjQoRJGahtllcuNTPjwfuNgWkdLwJnsXJBXG
yYd01amu6cEhI2pjpzq5j4MRPStVTF4qFmSq8a8zyxLSCkBrt5Z/CGLPyFo21ws60w++XsbOLmjm
i8XI9G4lAw+16kg6Oy+JyqqCZP4Fp2hkU+V65oHrqr4SB6WqlH8NBarfDzwhl25D374y1gMR9aVu
uLiH6BM3AAi9jUFl9pECaGSGNb2jYJFr4948OAer7u9Ujx65BoxGPT+y+PJprM3Tvt2S3vJMfeEU
5fdnzXWm51FstUWd42Us+FZVm79Iz6vI6mcqTuNNFiDqvNLCYUOck82H5h/bRlf/qsxLM5iD1Xf4
1GTW//jg0cHMboIgsHWm1VBvZJecNiC5Hrlw92h8hFO6ZmA3+L6C9BNQRtBdODNeVhyi70HsBjGf
zK4Bgxxzw9n+VcljaVUrViGdvJLfdkCJsYh9S2vTk8JdlJEUEsVL8taPeNa7KnWMnMb25DJfPo4q
m0kbDnpUXQ5eRE0QLOagPYqesLf9/JLoUn9jyT41cVm55nd2jxKP5GNQ9OAIIAUM5CEVvKzrsHEW
DgWsIBMKLDM8l4isWFZEcHdSTqR82oy8RiWPN01g1NRf1WVgq0i+uE6dhZrrribJXuqnXELmKsBN
9VP+i2xP3aPhlc7KvVDrtll6Lc6ugR/tJ9FK7VmtYF6EgsGB6MJQmGXRuYvPyq+45QFpJUQmK/Xc
zjrMdP2ht+YloYeuJ8AbIdX7Xt1BNwUQHUxlLN1RYVdc8y2qfJOLdOjwLBVFaDepwXl5IjDdvkr+
6qISQP+DoHiKIKaymMue+tYfnj9OZg88UW5tcyxfznscqAhpIcEixk4ADvDISeZqebpFr+dfWPFF
ndrTukGeCv8F8502LUEh6r8sNb8ZHRvis6+OJCvecGZuk1uOAtpgim/ZwbgokAHtehoEFMMweV13
WdnbN3MyFiDcr1DYbP2cm0T84Vc1SwQJQKziRFku5ugXp8Mt8hGx7pkc6ikzLTFRYXMxCrVEFxz0
u2YaXJnOm+EoGTEqusBD5lMbh6E/0zczd6k0pqEpXdw3OWgMCD0TnigkXSya2tU/gDxX4FchWE9E
eJpBC58Tma7d5/B614afJiaOE+zwWZIyvUtZwlkY0bkhDjZSweuWXmZwjo8i7KAvKZbMoBk26ODi
DTOrjPX2fmGxWl8FgLCjbwXPIDOIw5LAU7h3aaqjWabzdo0FELzc+qJm4evVghE6tUO3/4CjJPrX
bAIMlgyjk1so+I0/hAbvK+q2gY6uuvQ+2CrPc3knjMnZ1/JnrhzhF2xnoqoxAkb+tQoXFB1YfQmu
4m3UDQkWiKYLDYjIUfhIGO3kRYZQZf5M8KdClveguxqrSMhiGv4NqinbJJJS2K7d3W5FAERxkx/K
ssRdbm+4czewyO0Mx0RTAeAc7nfUlJMkLIFuGDaA68B6kSFLmzrNBCcqz+u/t8GIF5djjD7IIBVf
Kvk74UO5XODQ6UKcsdMd4V0XxxTKjvnvE5Swm8mA06cbKhNWpzEDXecJtj52qXKOnsd0IEbwaRQe
UpsLmZfQ3COZG83thJUtYR+F7//i4aRmdrGogJ+QkvgC1A/2vvW9fYbyYSggIRAT0MbUqAYdGVFo
N6zCIQuGTWIAjJDHWTwxlH0QHZe9X6mEcoL/87BM5+cKZbpGcV7KaNvS12ua+EE8C+vuOyv9LCoZ
tyX3id06tAX2WpdmimDvSFyLCCsujSaeKn+FoaR+0f2dH8gPouvMI3a91QYcR1Jkguk021ner+Ps
tyA6v9b3GsgOWaTVWePqpHP9eZYHRQLTRfDNNvgdRiHtFnG1zd92UaTEyMhi44j/V6jo4s2MAKOM
xTLtQqxsHX/6fPPES8GEAkpIoncWqWsPU6MWOasTBWe4nKPor8kGYk91PSZGN+OzaB/0a47T9e+Y
uxG95YhvQokY7rNZwE2JKz4JiaoFGgSx1J/AHAmjojxJo2akHFLaftPAq/LTXxfRJNVsv37iKYrM
mVZv/Q19u1bAQBEBvK72n+zA9yyICfZLRvLIxtw/kKHBJTJnHAMq8DlZzx2uod+JtTynxwa1vhXm
eEFKrAybIJSVDkwTjUA8GK7WqbEpbqP3MlH9CrndUEC8tnMKXRtnyunC8Gt04Bfr5Ga9fwaPBz1n
IYzYXK0+ih84R57WWB6P/tfxdOJLj7Eofn/0QeM1Ae6/46UcZDqzlYGlXEcakEU+CiR821J2tYYM
dGfUWIn2T4H0isOxDGgPHCsLyWXAFf1azO2k8oUkfxN7Hx0HKI3FCIt3ICUUDiXn8lXgXduW0if7
7LfPpM5737qTnEjqJYW81dJsqSlCo8KAoCU82f9HeDNMcb2+jIZksKVScjeCc6PwZtsVsZGUcGC2
KnX8wEw0LZkHyXocEQxWS/9cjCFpLMO5GCCykwFrs/ot+0l1/RE5s/p8H64loSiItL4JP90X8lrJ
aVY5/kYrSAhCGlwo2BfHkHn32G6LkYhPmrEt+GZPk78R0caQnxTMP8EBy0Xti0rJyVo1IaCzR2J2
sf4bHvi+gWMppBJHMt3roAzdqC5D30tsTxb3lenzEPs0LL3t/Ei1PEThgtnDQj22WR1e/5I7M2ZI
8sOj7k96k8SAejVbcqW0zDQ4fmLEi/zCa4HrguZ/Mxo5XvWDLh8rZzkxWoHuy4OVcreq43Htvb20
I9akKobj7vu9ivo8Oly72tSO/3f7gHlMuN4zLA3DvaBTk/Aj0/gLdvhshsCmRZ0IdBz5IbOXTo7D
oMr9wb43xZJCTpDLH8sxHLllVqDBM2vDqOCBiIHsQDEKVSneFgBlu6buMusKCV/tQGZYdE6zMxdR
5a2u9j1Z8BMA5Phwwqs2jjdfjWiwL0+ljTz0+hFGg1jYTXa2ELm55NfzKQ+IJ8iOWlbFEncgGlrz
bpZEwYu64Jr5j8dmgDDkq7RXeHd5C4jMVQx3uIDyOH8urSRUh9v/ZGIAoLm1PVlJgSPIHxANOnN2
Z1kGO9Ln0gx6lM9sBjt6joxWJoENKJkudR86OEV6owqP634bf7rLwVu1lo9tG84b0igfqVmLQz1Q
F4b4iYXynwPrEQm0x3hxXxb97WVt4vkxpQF0LC6S4MPEO+jJA0ACA43KSRN5FMbos8MfaxqXf2KR
CBOesqu7gP1YEEn0OU49jN+ruCxi18hLYfblNqh4f0sJEnsExAOBQf04tknCUkAdHxLbnvX2NWJe
7mtv+DxtFgX2nH6LSyIbLoICVCvkNN/PTUBwiLbeK0aN9QYs14yuJ8qeW8WrEa1Id2/XXv9VjBX+
J5bPtO464m8K1EL+51yUdMyfDMJOKmOzF4IjgRZQ/HeyKjod8fre5I3Cd9eiZvQnCiT6/qPzc3/4
QrfyJoSUcLflU8l4t0YXoUpzasmb7ODZSuBxRKYZKVhyeOa0UR57Lp6MTZfYjwkK5L0tR/FU31B+
1XN07lYrpaGTWXDjCCx9t7Nz/PFd6H28XRKvDZ0wUTlF1JVIuGXqutBnFzYe/IH0JL1LhBN/dEd1
1uWmqT0+i7m0FWlEWWsLMJB0ECQotL4YUGSHaLi46NSZi+FjY77qbdslASKvFCV/PfMjXRnkvpmk
ASZit/5BDNqcZPC3cvhpdK3yLpvGa9bJ1pieNxn8x98E9Ii8VH18orECRy9UZcUae6LpkC3Hr9/y
w5ZOgrDsAcouFm/kZ2ZkKjCuv1lx+DEyWPyd7ncneFroijbavGwRkwq8lAqi/x3NttY+MqJ1bgmV
iAEcKs/l6FNJO/6YY9Tcu4D5zMeEhu+qDyVygosupTJmtw3YI2P9eugrZxcV7tyRI8AAtr9XMeKO
f9TeBhBMTyCmtOLuPC/TfQubm5HAzSjlgqH3VQ53ym0jJo62v0fB27X4zyKUBSXQOn1Z6oQtrAWq
Mwcc2I9CFnZqYF9qSOZB/0EBJG+lWG/YiCZ4zPxVWF1qyJs793/77xWPkBrLoK2h6uk7OdkbsrGh
FI39ZropttTKEsukGOSp1ibiFSuWMnL+KPNa8WDI0d8RSUrQILRjeBl8aYNs8zlVHt4DHOi0++tG
FRsWqOF0Wp54NnYaCBlRE5ls6okcxK3xzCWDrq/roMSeME1CvQt754XRC3ptpa4sbEqDiMEU7PaL
y4p590+qmq7/lJq7M4TcUKRAebEJ+An0a3nxny/QwOCyTENXk7QtX7ZN9V/XUI6GCpDy/3n+nCDG
0Qcy290dxNYi/y5QQHe/lfjGoDd/1Z9NrRWQ36f7SmcXwxbuGI+UksWpuNKusxVBlE+5qvhUl7HM
NYOt8dcvJsEmefu9NewV6X5mpFGMf4XvG2xxyGkbIipeb9wRt2EtD8+PSDkzWOy5Tvt/SgRSwHKl
887hA3H4u33d5P/1CXDWS5LXNj8u7zIVVT6o9PgW8lESeZhW2xA5jxugmL0Az7W+rwvV8WmXlnfI
SozkfCCQG3+3m0yGJpWhbS1e4bVDoi0EPTYITC9A2Ic4X7R6Joe0ZOjJWy5QA8lWHqcJY4yG86MP
bLxThZrp5ZZ7OhTRB/psTYkQqxavG9hFIXCHnWZkSIpnaa7xPAIYEQoKqxHWc1xoUGaxeSaBL6Yt
4I+SHXc6QgJbi+Cz78VzAKzmlHnO8eDACq2csB1Nk+LnXDdMb82FxqmebpS1QD4uLNhnKWymDIFj
2cRs2dPn3v4y8Ugl3Jx54vHT/jz8qieKySrr5BEm9EoqUES1WynQoMBy8oOrGXjTlir4Tw8AWueX
7fkhbGsywT+8lM2SzKzQm4dC2W4aMO9z5UiptJyYS3SG9LX7TB2GVmhziSopKHQcNoDmP/q0hFZ6
wBHYimFOM/sVveHdeu0OQ6SIZAj2jHLB0Xr2dfXVR5Ry2yJXh1F3R+jtcAeXqJmN4G01Hf+9EAtl
jC9uzug5E8zbkPHPIgYVtgRK6z7uP58oDU6iuv4d2u7yVmsTktesNjMwJX6NDTMMxJ+bUJdUxsQi
CVWVPQ6zMfnnw5qXMpVJeUs/uaPvyCyHC6FOmNtXD/fKq7OSRHEl9V6hPC7a5tWldSk7DSNx5NOi
BZamZDpdTn9tkYTva46uQ8hBFG8WIx2MDs8vYUSXnd9zzElZdbi4l1eQYMt54LCrjR3ZQmDn1cqf
8e8P1NkBFId4tMIjEPNoNZ845PbrxP300CGZyueLgSzkBYFOI67j5z94FvvyW7rRCKw6Zdkb1760
IQZLNdHxOtUwPxgS/nPSw02v16UYUrWBKG5KPvNXQZkeZgwlq4U+yQ/xFql5dwWQdYahbLu4TWnk
+VTSfUHN7W5ES0OP/OgP6D4Qo2lQVIpOB68JGy/uCxQVNfdn+AXNkd7vb+7nEurUe04VRJJtqAEp
lp5ZOLqM0jo5Hk/281lW8MwSfgJ+G7pcktOgf65Lps2A/xYq5xhkVApMk02DsMiVoEQKKE2DoG3W
tfaPSu7d04x1ghAThbcrA/3syRYqn5ZAKmKbIZo4xYugEXpDAVaxfIDe1o7j9P9ohxVOlNw2bIt2
NKfGM9NcArLzEXCCwk6OJFd/V670dDqxFT+sZEfj5OSLASi+GtSzig5f7yBaLlp8rdY6smQ0OPIa
/wluIsPfUsljGrpyX/czlfo3D2t6LN1KsnsqZvdQ+OCA/8Ix7yumyzR5sQz6ihaDgrtrtiZu2jw8
JBYt8mOJmibCgxhKlVXvs90yLKQar/KM/1QUFgjqc2Unyo6hgmC9zzn86hsZ527bxUn1Yiqlwg8X
BglKntNAKdjCvPv2PST9im7haM1G3t+KE3uEp6/NtyaezQgV26Z+ewhDspGhxPxZ+ZTtjXORxgkg
lvIT0rg8xP4bXXt6teVonKUDDPLXp7hLg4/8v7KR+ygV2qu2xp/NGEPBX0mlGo1E0tge29c/7iXT
TxMk/a9tmRmj9yP3GpVYM+Lp3C7hSNKTNVToRUlKxj52OxYZAIcz/lnvHEOLuhN6ZwL5Co7aMKDc
+dL2cMhP6WNCquxY1tOfyAiinLDdABzWDeZO/Z0KpISbSeOZMnqgpd/wbyDykUUP/UKy5hHVO9am
ylfOxZDbzee/Ty2kMIv6jolBQ24RpLnoUYj9TesZFIrEMJf7nQq2Cq/FbjOdzpTka4MjyoAWah28
4vUf3oaDhYY2n89UcE12w38+ew0OxBbC1R8VDi+pNWuapnpRpPdJR42Y+DWcsbUHlnF3sw==
`protect end_protected
