localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTY_CHK = {
  {32'h3eadb08f, 32'hbe6eab13} /* (31, 31, 31) {real, imag} */,
  {32'hbe8c81aa, 32'h3e41a2f8} /* (31, 31, 30) {real, imag} */,
  {32'h3af2d970, 32'hbcae82e6} /* (31, 31, 29) {real, imag} */,
  {32'h3d8aba9c, 32'h3d5dba23} /* (31, 31, 28) {real, imag} */,
  {32'hbd6ff125, 32'h3c9abe34} /* (31, 31, 27) {real, imag} */,
  {32'h3af629c0, 32'hbc497c9a} /* (31, 31, 26) {real, imag} */,
  {32'hbc9bfc9a, 32'hbcf6848a} /* (31, 31, 25) {real, imag} */,
  {32'h3d0a7628, 32'h3d3ee6ee} /* (31, 31, 24) {real, imag} */,
  {32'hbd14d280, 32'h3c9852e5} /* (31, 31, 23) {real, imag} */,
  {32'hbc96cedb, 32'hbd0fbaf3} /* (31, 31, 22) {real, imag} */,
  {32'hbd0cd3d0, 32'h3c76c7cd} /* (31, 31, 21) {real, imag} */,
  {32'h3d1f948c, 32'hbd12eb88} /* (31, 31, 20) {real, imag} */,
  {32'h3c9101b8, 32'h3c5684b1} /* (31, 31, 19) {real, imag} */,
  {32'h3cdf04c4, 32'hbab3c2c8} /* (31, 31, 18) {real, imag} */,
  {32'h3c83bb16, 32'hbc7b7f98} /* (31, 31, 17) {real, imag} */,
  {32'hbb233e80, 32'h00000000} /* (31, 31, 16) {real, imag} */,
  {32'h3c83bb16, 32'h3c7b7f98} /* (31, 31, 15) {real, imag} */,
  {32'h3cdf04c4, 32'h3ab3c2c8} /* (31, 31, 14) {real, imag} */,
  {32'h3c9101b8, 32'hbc5684b1} /* (31, 31, 13) {real, imag} */,
  {32'h3d1f948c, 32'h3d12eb88} /* (31, 31, 12) {real, imag} */,
  {32'hbd0cd3d0, 32'hbc76c7cd} /* (31, 31, 11) {real, imag} */,
  {32'hbc96cedb, 32'h3d0fbaf3} /* (31, 31, 10) {real, imag} */,
  {32'hbd14d280, 32'hbc9852e5} /* (31, 31, 9) {real, imag} */,
  {32'h3d0a7628, 32'hbd3ee6ee} /* (31, 31, 8) {real, imag} */,
  {32'hbc9bfc9a, 32'h3cf6848a} /* (31, 31, 7) {real, imag} */,
  {32'h3af629c0, 32'h3c497c9a} /* (31, 31, 6) {real, imag} */,
  {32'hbd6ff125, 32'hbc9abe34} /* (31, 31, 5) {real, imag} */,
  {32'h3d8aba9c, 32'hbd5dba23} /* (31, 31, 4) {real, imag} */,
  {32'h3af2d970, 32'h3cae82e6} /* (31, 31, 3) {real, imag} */,
  {32'hbe8c81aa, 32'hbe41a2f8} /* (31, 31, 2) {real, imag} */,
  {32'h3eadb08f, 32'h3e6eab13} /* (31, 31, 1) {real, imag} */,
  {32'h3e61b5c3, 32'h00000000} /* (31, 31, 0) {real, imag} */,
  {32'h3f06c004, 32'hbe8db278} /* (31, 30, 31) {real, imag} */,
  {32'hbee68306, 32'h3e8c601a} /* (31, 30, 30) {real, imag} */,
  {32'h3ca503bc, 32'hb96cf200} /* (31, 30, 29) {real, imag} */,
  {32'h3d60a8d2, 32'h3a848b00} /* (31, 30, 28) {real, imag} */,
  {32'hbd331a3b, 32'h3cb4e6eb} /* (31, 30, 27) {real, imag} */,
  {32'h3d298a0a, 32'hbadc6040} /* (31, 30, 26) {real, imag} */,
  {32'hbd0da2f1, 32'hbda17a32} /* (31, 30, 25) {real, imag} */,
  {32'h3d9fd303, 32'h3cfa05ce} /* (31, 30, 24) {real, imag} */,
  {32'hbb28fc40, 32'hbd80b69a} /* (31, 30, 23) {real, imag} */,
  {32'hbd7098d0, 32'hbab30bc0} /* (31, 30, 22) {real, imag} */,
  {32'hbd1ca92a, 32'hbb5135a4} /* (31, 30, 21) {real, imag} */,
  {32'h3b3b81e0, 32'hbca89e92} /* (31, 30, 20) {real, imag} */,
  {32'h3c18aed2, 32'h3b357140} /* (31, 30, 19) {real, imag} */,
  {32'h3d8c26ba, 32'hbc3db234} /* (31, 30, 18) {real, imag} */,
  {32'hbc90fae4, 32'hbbe51205} /* (31, 30, 17) {real, imag} */,
  {32'hbd1e14e9, 32'h00000000} /* (31, 30, 16) {real, imag} */,
  {32'hbc90fae4, 32'h3be51205} /* (31, 30, 15) {real, imag} */,
  {32'h3d8c26ba, 32'h3c3db234} /* (31, 30, 14) {real, imag} */,
  {32'h3c18aed2, 32'hbb357140} /* (31, 30, 13) {real, imag} */,
  {32'h3b3b81e0, 32'h3ca89e92} /* (31, 30, 12) {real, imag} */,
  {32'hbd1ca92a, 32'h3b5135a4} /* (31, 30, 11) {real, imag} */,
  {32'hbd7098d0, 32'h3ab30bc0} /* (31, 30, 10) {real, imag} */,
  {32'hbb28fc40, 32'h3d80b69a} /* (31, 30, 9) {real, imag} */,
  {32'h3d9fd303, 32'hbcfa05ce} /* (31, 30, 8) {real, imag} */,
  {32'hbd0da2f1, 32'h3da17a32} /* (31, 30, 7) {real, imag} */,
  {32'h3d298a0a, 32'h3adc6040} /* (31, 30, 6) {real, imag} */,
  {32'hbd331a3b, 32'hbcb4e6eb} /* (31, 30, 5) {real, imag} */,
  {32'h3d60a8d2, 32'hba848b00} /* (31, 30, 4) {real, imag} */,
  {32'h3ca503bc, 32'h396cf200} /* (31, 30, 3) {real, imag} */,
  {32'hbee68306, 32'hbe8c601a} /* (31, 30, 2) {real, imag} */,
  {32'h3f06c004, 32'h3e8db278} /* (31, 30, 1) {real, imag} */,
  {32'h3e3a5132, 32'h00000000} /* (31, 30, 0) {real, imag} */,
  {32'h3f1ba38e, 32'hbe207cd1} /* (31, 29, 31) {real, imag} */,
  {32'hbec2b284, 32'h3e7a9433} /* (31, 29, 30) {real, imag} */,
  {32'hbc5e4818, 32'h3d905a4f} /* (31, 29, 29) {real, imag} */,
  {32'h3dc1f415, 32'h3baaa560} /* (31, 29, 28) {real, imag} */,
  {32'hbd80f407, 32'h3c636fac} /* (31, 29, 27) {real, imag} */,
  {32'hbd821fcc, 32'hbca91dcc} /* (31, 29, 26) {real, imag} */,
  {32'h3c8d592e, 32'hbd0a6626} /* (31, 29, 25) {real, imag} */,
  {32'hbcf2439b, 32'h3cbf5be2} /* (31, 29, 24) {real, imag} */,
  {32'hbc475fa7, 32'h3dd6ceb8} /* (31, 29, 23) {real, imag} */,
  {32'h3d76be28, 32'hbd270a68} /* (31, 29, 22) {real, imag} */,
  {32'hbd52fb64, 32'hbcf4fea7} /* (31, 29, 21) {real, imag} */,
  {32'hbc9ac18a, 32'h3d2c1d84} /* (31, 29, 20) {real, imag} */,
  {32'hbac447c0, 32'hbdece47f} /* (31, 29, 19) {real, imag} */,
  {32'hbcb0ba27, 32'hbcfaf237} /* (31, 29, 18) {real, imag} */,
  {32'hbcba963a, 32'hbcad5670} /* (31, 29, 17) {real, imag} */,
  {32'h3d93ec56, 32'h00000000} /* (31, 29, 16) {real, imag} */,
  {32'hbcba963a, 32'h3cad5670} /* (31, 29, 15) {real, imag} */,
  {32'hbcb0ba27, 32'h3cfaf237} /* (31, 29, 14) {real, imag} */,
  {32'hbac447c0, 32'h3dece47f} /* (31, 29, 13) {real, imag} */,
  {32'hbc9ac18a, 32'hbd2c1d84} /* (31, 29, 12) {real, imag} */,
  {32'hbd52fb64, 32'h3cf4fea7} /* (31, 29, 11) {real, imag} */,
  {32'h3d76be28, 32'h3d270a68} /* (31, 29, 10) {real, imag} */,
  {32'hbc475fa7, 32'hbdd6ceb8} /* (31, 29, 9) {real, imag} */,
  {32'hbcf2439b, 32'hbcbf5be2} /* (31, 29, 8) {real, imag} */,
  {32'h3c8d592e, 32'h3d0a6626} /* (31, 29, 7) {real, imag} */,
  {32'hbd821fcc, 32'h3ca91dcc} /* (31, 29, 6) {real, imag} */,
  {32'hbd80f407, 32'hbc636fac} /* (31, 29, 5) {real, imag} */,
  {32'h3dc1f415, 32'hbbaaa560} /* (31, 29, 4) {real, imag} */,
  {32'hbc5e4818, 32'hbd905a4f} /* (31, 29, 3) {real, imag} */,
  {32'hbec2b284, 32'hbe7a9433} /* (31, 29, 2) {real, imag} */,
  {32'h3f1ba38e, 32'h3e207cd1} /* (31, 29, 1) {real, imag} */,
  {32'h3e389a35, 32'h00000000} /* (31, 29, 0) {real, imag} */,
  {32'h3f0b6094, 32'hbde882c6} /* (31, 28, 31) {real, imag} */,
  {32'hbe96625b, 32'h3db48b90} /* (31, 28, 30) {real, imag} */,
  {32'hbd237ab7, 32'hbbe41b3e} /* (31, 28, 29) {real, imag} */,
  {32'h3e1d85c8, 32'h3d7a02c5} /* (31, 28, 28) {real, imag} */,
  {32'hbd97176f, 32'hbcedfe16} /* (31, 28, 27) {real, imag} */,
  {32'hbc78ccc0, 32'h3d96b304} /* (31, 28, 26) {real, imag} */,
  {32'h3bde2dc4, 32'hbd878784} /* (31, 28, 25) {real, imag} */,
  {32'hbda60d7c, 32'h3dc8e82e} /* (31, 28, 24) {real, imag} */,
  {32'h3d21c1c9, 32'h3cb6de37} /* (31, 28, 23) {real, imag} */,
  {32'hbc3c8226, 32'hbc45ff2b} /* (31, 28, 22) {real, imag} */,
  {32'hbc78758f, 32'hbc94a35e} /* (31, 28, 21) {real, imag} */,
  {32'h3bf6a138, 32'hbcb7484a} /* (31, 28, 20) {real, imag} */,
  {32'hbc4c789f, 32'h3d0a334f} /* (31, 28, 19) {real, imag} */,
  {32'hbd2b79ca, 32'h3d5a84ef} /* (31, 28, 18) {real, imag} */,
  {32'h3d30f1f1, 32'hbbfa8b83} /* (31, 28, 17) {real, imag} */,
  {32'hbc075eae, 32'h00000000} /* (31, 28, 16) {real, imag} */,
  {32'h3d30f1f1, 32'h3bfa8b83} /* (31, 28, 15) {real, imag} */,
  {32'hbd2b79ca, 32'hbd5a84ef} /* (31, 28, 14) {real, imag} */,
  {32'hbc4c789f, 32'hbd0a334f} /* (31, 28, 13) {real, imag} */,
  {32'h3bf6a138, 32'h3cb7484a} /* (31, 28, 12) {real, imag} */,
  {32'hbc78758f, 32'h3c94a35e} /* (31, 28, 11) {real, imag} */,
  {32'hbc3c8226, 32'h3c45ff2b} /* (31, 28, 10) {real, imag} */,
  {32'h3d21c1c9, 32'hbcb6de37} /* (31, 28, 9) {real, imag} */,
  {32'hbda60d7c, 32'hbdc8e82e} /* (31, 28, 8) {real, imag} */,
  {32'h3bde2dc4, 32'h3d878784} /* (31, 28, 7) {real, imag} */,
  {32'hbc78ccc0, 32'hbd96b304} /* (31, 28, 6) {real, imag} */,
  {32'hbd97176f, 32'h3cedfe16} /* (31, 28, 5) {real, imag} */,
  {32'h3e1d85c8, 32'hbd7a02c5} /* (31, 28, 4) {real, imag} */,
  {32'hbd237ab7, 32'h3be41b3e} /* (31, 28, 3) {real, imag} */,
  {32'hbe96625b, 32'hbdb48b90} /* (31, 28, 2) {real, imag} */,
  {32'h3f0b6094, 32'h3de882c6} /* (31, 28, 1) {real, imag} */,
  {32'h3e8ddf70, 32'h00000000} /* (31, 28, 0) {real, imag} */,
  {32'h3ee36cba, 32'hbe0579e5} /* (31, 27, 31) {real, imag} */,
  {32'hbecc8cdc, 32'h3dffcad0} /* (31, 27, 30) {real, imag} */,
  {32'hbc89f400, 32'hbd1feb64} /* (31, 27, 29) {real, imag} */,
  {32'hbc46aa00, 32'h3d9e4b84} /* (31, 27, 28) {real, imag} */,
  {32'h3d17741e, 32'h3bf8dc70} /* (31, 27, 27) {real, imag} */,
  {32'h3d094c93, 32'hbca4344d} /* (31, 27, 26) {real, imag} */,
  {32'hbd21dfa4, 32'hbda19258} /* (31, 27, 25) {real, imag} */,
  {32'hbd92d7c7, 32'hbc8d0fcd} /* (31, 27, 24) {real, imag} */,
  {32'hba33c9e0, 32'h3d1f17a8} /* (31, 27, 23) {real, imag} */,
  {32'h3d0bf176, 32'hbd227b7e} /* (31, 27, 22) {real, imag} */,
  {32'hbd7c6ee2, 32'hb93a2a00} /* (31, 27, 21) {real, imag} */,
  {32'h3cdc435a, 32'h3c33fa6e} /* (31, 27, 20) {real, imag} */,
  {32'hbc00fde0, 32'h3d6e8688} /* (31, 27, 19) {real, imag} */,
  {32'hbc09948c, 32'h3dbfc806} /* (31, 27, 18) {real, imag} */,
  {32'h3c97a49e, 32'hbd6ceac4} /* (31, 27, 17) {real, imag} */,
  {32'h3d23ceaa, 32'h00000000} /* (31, 27, 16) {real, imag} */,
  {32'h3c97a49e, 32'h3d6ceac4} /* (31, 27, 15) {real, imag} */,
  {32'hbc09948c, 32'hbdbfc806} /* (31, 27, 14) {real, imag} */,
  {32'hbc00fde0, 32'hbd6e8688} /* (31, 27, 13) {real, imag} */,
  {32'h3cdc435a, 32'hbc33fa6e} /* (31, 27, 12) {real, imag} */,
  {32'hbd7c6ee2, 32'h393a2a00} /* (31, 27, 11) {real, imag} */,
  {32'h3d0bf176, 32'h3d227b7e} /* (31, 27, 10) {real, imag} */,
  {32'hba33c9e0, 32'hbd1f17a8} /* (31, 27, 9) {real, imag} */,
  {32'hbd92d7c7, 32'h3c8d0fcd} /* (31, 27, 8) {real, imag} */,
  {32'hbd21dfa4, 32'h3da19258} /* (31, 27, 7) {real, imag} */,
  {32'h3d094c93, 32'h3ca4344d} /* (31, 27, 6) {real, imag} */,
  {32'h3d17741e, 32'hbbf8dc70} /* (31, 27, 5) {real, imag} */,
  {32'hbc46aa00, 32'hbd9e4b84} /* (31, 27, 4) {real, imag} */,
  {32'hbc89f400, 32'h3d1feb64} /* (31, 27, 3) {real, imag} */,
  {32'hbecc8cdc, 32'hbdffcad0} /* (31, 27, 2) {real, imag} */,
  {32'h3ee36cba, 32'h3e0579e5} /* (31, 27, 1) {real, imag} */,
  {32'h3ecc18c6, 32'h00000000} /* (31, 27, 0) {real, imag} */,
  {32'h3f00b433, 32'hbe151bde} /* (31, 26, 31) {real, imag} */,
  {32'hbf03c0fb, 32'h3e65101a} /* (31, 26, 30) {real, imag} */,
  {32'h3c9ca018, 32'hbc549fd9} /* (31, 26, 29) {real, imag} */,
  {32'h3d0b4f3c, 32'h3ccebd44} /* (31, 26, 28) {real, imag} */,
  {32'h3d18adee, 32'h3ced3c44} /* (31, 26, 27) {real, imag} */,
  {32'hbc086763, 32'h3d153755} /* (31, 26, 26) {real, imag} */,
  {32'hbd461488, 32'hbdaa928a} /* (31, 26, 25) {real, imag} */,
  {32'hbba32dba, 32'h3d53c0e3} /* (31, 26, 24) {real, imag} */,
  {32'hbdb30c44, 32'hbd70a386} /* (31, 26, 23) {real, imag} */,
  {32'hbc95e595, 32'h3d14a8a3} /* (31, 26, 22) {real, imag} */,
  {32'h3d13b8fa, 32'h396c6200} /* (31, 26, 21) {real, imag} */,
  {32'h3cf13308, 32'h3d1b008c} /* (31, 26, 20) {real, imag} */,
  {32'hbcc2ca25, 32'hbdbfa7e6} /* (31, 26, 19) {real, imag} */,
  {32'hbcbe1388, 32'h3cf99d08} /* (31, 26, 18) {real, imag} */,
  {32'h3c52b2b4, 32'hbcc6f1aa} /* (31, 26, 17) {real, imag} */,
  {32'hbc78511b, 32'h00000000} /* (31, 26, 16) {real, imag} */,
  {32'h3c52b2b4, 32'h3cc6f1aa} /* (31, 26, 15) {real, imag} */,
  {32'hbcbe1388, 32'hbcf99d08} /* (31, 26, 14) {real, imag} */,
  {32'hbcc2ca25, 32'h3dbfa7e6} /* (31, 26, 13) {real, imag} */,
  {32'h3cf13308, 32'hbd1b008c} /* (31, 26, 12) {real, imag} */,
  {32'h3d13b8fa, 32'hb96c6200} /* (31, 26, 11) {real, imag} */,
  {32'hbc95e595, 32'hbd14a8a3} /* (31, 26, 10) {real, imag} */,
  {32'hbdb30c44, 32'h3d70a386} /* (31, 26, 9) {real, imag} */,
  {32'hbba32dba, 32'hbd53c0e3} /* (31, 26, 8) {real, imag} */,
  {32'hbd461488, 32'h3daa928a} /* (31, 26, 7) {real, imag} */,
  {32'hbc086763, 32'hbd153755} /* (31, 26, 6) {real, imag} */,
  {32'h3d18adee, 32'hbced3c44} /* (31, 26, 5) {real, imag} */,
  {32'h3d0b4f3c, 32'hbccebd44} /* (31, 26, 4) {real, imag} */,
  {32'h3c9ca018, 32'h3c549fd9} /* (31, 26, 3) {real, imag} */,
  {32'hbf03c0fb, 32'hbe65101a} /* (31, 26, 2) {real, imag} */,
  {32'h3f00b433, 32'h3e151bde} /* (31, 26, 1) {real, imag} */,
  {32'h3ec8d262, 32'h00000000} /* (31, 26, 0) {real, imag} */,
  {32'h3f12f89d, 32'hbc3b7963} /* (31, 25, 31) {real, imag} */,
  {32'hbf096ca3, 32'h3e8b3aea} /* (31, 25, 30) {real, imag} */,
  {32'hbd4691f8, 32'h3b2508e0} /* (31, 25, 29) {real, imag} */,
  {32'h3d5bea2d, 32'hbd3e147a} /* (31, 25, 28) {real, imag} */,
  {32'hbbde0b48, 32'h3ce48782} /* (31, 25, 27) {real, imag} */,
  {32'h3ab05340, 32'hbd27d4b6} /* (31, 25, 26) {real, imag} */,
  {32'h3d4db3ea, 32'hbd0331d6} /* (31, 25, 25) {real, imag} */,
  {32'hbd9a9203, 32'h3cb4e7b8} /* (31, 25, 24) {real, imag} */,
  {32'hb9045c00, 32'h3d23cc4e} /* (31, 25, 23) {real, imag} */,
  {32'h3bb70928, 32'hbc7add52} /* (31, 25, 22) {real, imag} */,
  {32'hbda98860, 32'hbc84e68f} /* (31, 25, 21) {real, imag} */,
  {32'h3dd318c0, 32'hbcafe4a8} /* (31, 25, 20) {real, imag} */,
  {32'h3d86d4b8, 32'hbc4049ba} /* (31, 25, 19) {real, imag} */,
  {32'h3ca6ea8d, 32'h3ca51a27} /* (31, 25, 18) {real, imag} */,
  {32'hbd061826, 32'h3d9a9658} /* (31, 25, 17) {real, imag} */,
  {32'hbbc1411c, 32'h00000000} /* (31, 25, 16) {real, imag} */,
  {32'hbd061826, 32'hbd9a9658} /* (31, 25, 15) {real, imag} */,
  {32'h3ca6ea8d, 32'hbca51a27} /* (31, 25, 14) {real, imag} */,
  {32'h3d86d4b8, 32'h3c4049ba} /* (31, 25, 13) {real, imag} */,
  {32'h3dd318c0, 32'h3cafe4a8} /* (31, 25, 12) {real, imag} */,
  {32'hbda98860, 32'h3c84e68f} /* (31, 25, 11) {real, imag} */,
  {32'h3bb70928, 32'h3c7add52} /* (31, 25, 10) {real, imag} */,
  {32'hb9045c00, 32'hbd23cc4e} /* (31, 25, 9) {real, imag} */,
  {32'hbd9a9203, 32'hbcb4e7b8} /* (31, 25, 8) {real, imag} */,
  {32'h3d4db3ea, 32'h3d0331d6} /* (31, 25, 7) {real, imag} */,
  {32'h3ab05340, 32'h3d27d4b6} /* (31, 25, 6) {real, imag} */,
  {32'hbbde0b48, 32'hbce48782} /* (31, 25, 5) {real, imag} */,
  {32'h3d5bea2d, 32'h3d3e147a} /* (31, 25, 4) {real, imag} */,
  {32'hbd4691f8, 32'hbb2508e0} /* (31, 25, 3) {real, imag} */,
  {32'hbf096ca3, 32'hbe8b3aea} /* (31, 25, 2) {real, imag} */,
  {32'h3f12f89d, 32'h3c3b7963} /* (31, 25, 1) {real, imag} */,
  {32'h3ec0d8a8, 32'h00000000} /* (31, 25, 0) {real, imag} */,
  {32'h3f06417a, 32'hbd5612a0} /* (31, 24, 31) {real, imag} */,
  {32'hbef531a6, 32'h3e6bde3f} /* (31, 24, 30) {real, imag} */,
  {32'h3c306070, 32'hbdb098ee} /* (31, 24, 29) {real, imag} */,
  {32'hbc971b70, 32'hbdc4d7c7} /* (31, 24, 28) {real, imag} */,
  {32'hbd610b0b, 32'hbcdf4cc0} /* (31, 24, 27) {real, imag} */,
  {32'hbd2ba0bc, 32'hbd8cfdb9} /* (31, 24, 26) {real, imag} */,
  {32'h3d0f8b63, 32'h3da1f0b6} /* (31, 24, 25) {real, imag} */,
  {32'hbe0211e6, 32'h3c2b627e} /* (31, 24, 24) {real, imag} */,
  {32'hbd39b813, 32'h3dc13436} /* (31, 24, 23) {real, imag} */,
  {32'hbc18cd5b, 32'hbd1886a5} /* (31, 24, 22) {real, imag} */,
  {32'hbc8c58d2, 32'h3be18df0} /* (31, 24, 21) {real, imag} */,
  {32'h3d5ba92d, 32'hbcbbbb4f} /* (31, 24, 20) {real, imag} */,
  {32'h3d559846, 32'h3ceaed6c} /* (31, 24, 19) {real, imag} */,
  {32'hbcde3f1b, 32'hbcceb6a3} /* (31, 24, 18) {real, imag} */,
  {32'h3c92f5dc, 32'h3d66e2d3} /* (31, 24, 17) {real, imag} */,
  {32'h3ce22b16, 32'h00000000} /* (31, 24, 16) {real, imag} */,
  {32'h3c92f5dc, 32'hbd66e2d3} /* (31, 24, 15) {real, imag} */,
  {32'hbcde3f1b, 32'h3cceb6a3} /* (31, 24, 14) {real, imag} */,
  {32'h3d559846, 32'hbceaed6c} /* (31, 24, 13) {real, imag} */,
  {32'h3d5ba92d, 32'h3cbbbb4f} /* (31, 24, 12) {real, imag} */,
  {32'hbc8c58d2, 32'hbbe18df0} /* (31, 24, 11) {real, imag} */,
  {32'hbc18cd5b, 32'h3d1886a5} /* (31, 24, 10) {real, imag} */,
  {32'hbd39b813, 32'hbdc13436} /* (31, 24, 9) {real, imag} */,
  {32'hbe0211e6, 32'hbc2b627e} /* (31, 24, 8) {real, imag} */,
  {32'h3d0f8b63, 32'hbda1f0b6} /* (31, 24, 7) {real, imag} */,
  {32'hbd2ba0bc, 32'h3d8cfdb9} /* (31, 24, 6) {real, imag} */,
  {32'hbd610b0b, 32'h3cdf4cc0} /* (31, 24, 5) {real, imag} */,
  {32'hbc971b70, 32'h3dc4d7c7} /* (31, 24, 4) {real, imag} */,
  {32'h3c306070, 32'h3db098ee} /* (31, 24, 3) {real, imag} */,
  {32'hbef531a6, 32'hbe6bde3f} /* (31, 24, 2) {real, imag} */,
  {32'h3f06417a, 32'h3d5612a0} /* (31, 24, 1) {real, imag} */,
  {32'h3f10df63, 32'h00000000} /* (31, 24, 0) {real, imag} */,
  {32'h3ef647d1, 32'hbc3006bd} /* (31, 23, 31) {real, imag} */,
  {32'hbeb673b1, 32'h3e3991ae} /* (31, 23, 30) {real, imag} */,
  {32'h3e068e10, 32'h3b2c2780} /* (31, 23, 29) {real, imag} */,
  {32'hbcbb6e2a, 32'hbcfa569e} /* (31, 23, 28) {real, imag} */,
  {32'hbdd53cb8, 32'h3cc0f2ba} /* (31, 23, 27) {real, imag} */,
  {32'hbd3e7b46, 32'h3d8585ba} /* (31, 23, 26) {real, imag} */,
  {32'hbd5b0809, 32'hbd553b1e} /* (31, 23, 25) {real, imag} */,
  {32'hbd8ac656, 32'h3d169bda} /* (31, 23, 24) {real, imag} */,
  {32'hbd40f13b, 32'h3c40f607} /* (31, 23, 23) {real, imag} */,
  {32'h3db73b90, 32'h3d072ef4} /* (31, 23, 22) {real, imag} */,
  {32'h3d849aec, 32'h3d07450f} /* (31, 23, 21) {real, imag} */,
  {32'hbcf3fde6, 32'h3caa1068} /* (31, 23, 20) {real, imag} */,
  {32'h3a9e3540, 32'h3d1f063d} /* (31, 23, 19) {real, imag} */,
  {32'h3d0ab34a, 32'h3c67aa24} /* (31, 23, 18) {real, imag} */,
  {32'h3d534148, 32'h3cc406f2} /* (31, 23, 17) {real, imag} */,
  {32'hbca5f832, 32'h00000000} /* (31, 23, 16) {real, imag} */,
  {32'h3d534148, 32'hbcc406f2} /* (31, 23, 15) {real, imag} */,
  {32'h3d0ab34a, 32'hbc67aa24} /* (31, 23, 14) {real, imag} */,
  {32'h3a9e3540, 32'hbd1f063d} /* (31, 23, 13) {real, imag} */,
  {32'hbcf3fde6, 32'hbcaa1068} /* (31, 23, 12) {real, imag} */,
  {32'h3d849aec, 32'hbd07450f} /* (31, 23, 11) {real, imag} */,
  {32'h3db73b90, 32'hbd072ef4} /* (31, 23, 10) {real, imag} */,
  {32'hbd40f13b, 32'hbc40f607} /* (31, 23, 9) {real, imag} */,
  {32'hbd8ac656, 32'hbd169bda} /* (31, 23, 8) {real, imag} */,
  {32'hbd5b0809, 32'h3d553b1e} /* (31, 23, 7) {real, imag} */,
  {32'hbd3e7b46, 32'hbd8585ba} /* (31, 23, 6) {real, imag} */,
  {32'hbdd53cb8, 32'hbcc0f2ba} /* (31, 23, 5) {real, imag} */,
  {32'hbcbb6e2a, 32'h3cfa569e} /* (31, 23, 4) {real, imag} */,
  {32'h3e068e10, 32'hbb2c2780} /* (31, 23, 3) {real, imag} */,
  {32'hbeb673b1, 32'hbe3991ae} /* (31, 23, 2) {real, imag} */,
  {32'h3ef647d1, 32'h3c3006bd} /* (31, 23, 1) {real, imag} */,
  {32'h3f20dac0, 32'h00000000} /* (31, 23, 0) {real, imag} */,
  {32'h3ea6460f, 32'h3df438b6} /* (31, 22, 31) {real, imag} */,
  {32'hbeb334dc, 32'h3e80e432} /* (31, 22, 30) {real, imag} */,
  {32'h3e68f4ce, 32'h3e18044d} /* (31, 22, 29) {real, imag} */,
  {32'h3d0aad9a, 32'hbd028878} /* (31, 22, 28) {real, imag} */,
  {32'hbe1b7fba, 32'h3d5bd2de} /* (31, 22, 27) {real, imag} */,
  {32'hbd87e79c, 32'h3cf0307b} /* (31, 22, 26) {real, imag} */,
  {32'h3da434da, 32'hbd96c9c0} /* (31, 22, 25) {real, imag} */,
  {32'hbd6c099f, 32'h3d57184d} /* (31, 22, 24) {real, imag} */,
  {32'h3ac49490, 32'h3cc88ded} /* (31, 22, 23) {real, imag} */,
  {32'hbcd13d1c, 32'h3a8f26d0} /* (31, 22, 22) {real, imag} */,
  {32'h3d13e204, 32'h3c9bacec} /* (31, 22, 21) {real, imag} */,
  {32'hbd90c03f, 32'hbc59bbaf} /* (31, 22, 20) {real, imag} */,
  {32'h3d43ed7c, 32'h3bb8d0d8} /* (31, 22, 19) {real, imag} */,
  {32'h3d321282, 32'hbd9f0994} /* (31, 22, 18) {real, imag} */,
  {32'h3d7cb2c3, 32'hbc978318} /* (31, 22, 17) {real, imag} */,
  {32'h3d3e859c, 32'h00000000} /* (31, 22, 16) {real, imag} */,
  {32'h3d7cb2c3, 32'h3c978318} /* (31, 22, 15) {real, imag} */,
  {32'h3d321282, 32'h3d9f0994} /* (31, 22, 14) {real, imag} */,
  {32'h3d43ed7c, 32'hbbb8d0d8} /* (31, 22, 13) {real, imag} */,
  {32'hbd90c03f, 32'h3c59bbaf} /* (31, 22, 12) {real, imag} */,
  {32'h3d13e204, 32'hbc9bacec} /* (31, 22, 11) {real, imag} */,
  {32'hbcd13d1c, 32'hba8f26d0} /* (31, 22, 10) {real, imag} */,
  {32'h3ac49490, 32'hbcc88ded} /* (31, 22, 9) {real, imag} */,
  {32'hbd6c099f, 32'hbd57184d} /* (31, 22, 8) {real, imag} */,
  {32'h3da434da, 32'h3d96c9c0} /* (31, 22, 7) {real, imag} */,
  {32'hbd87e79c, 32'hbcf0307b} /* (31, 22, 6) {real, imag} */,
  {32'hbe1b7fba, 32'hbd5bd2de} /* (31, 22, 5) {real, imag} */,
  {32'h3d0aad9a, 32'h3d028878} /* (31, 22, 4) {real, imag} */,
  {32'h3e68f4ce, 32'hbe18044d} /* (31, 22, 3) {real, imag} */,
  {32'hbeb334dc, 32'hbe80e432} /* (31, 22, 2) {real, imag} */,
  {32'h3ea6460f, 32'hbdf438b6} /* (31, 22, 1) {real, imag} */,
  {32'h3eed0004, 32'h00000000} /* (31, 22, 0) {real, imag} */,
  {32'h3b064600, 32'h3dcd1da6} /* (31, 21, 31) {real, imag} */,
  {32'hbe250786, 32'h3d154c93} /* (31, 21, 30) {real, imag} */,
  {32'h3ddd6a28, 32'h3d910ff2} /* (31, 21, 29) {real, imag} */,
  {32'hbdb55600, 32'hbd6c0395} /* (31, 21, 28) {real, imag} */,
  {32'hbd9781f8, 32'hbb4055c8} /* (31, 21, 27) {real, imag} */,
  {32'hbd6d730e, 32'hbc837aa3} /* (31, 21, 26) {real, imag} */,
  {32'hbcf02309, 32'h3cf5f784} /* (31, 21, 25) {real, imag} */,
  {32'h3d1a849a, 32'hbc66216c} /* (31, 21, 24) {real, imag} */,
  {32'hbda657f4, 32'h3d23c0ad} /* (31, 21, 23) {real, imag} */,
  {32'h3c7eadc3, 32'hbd12f304} /* (31, 21, 22) {real, imag} */,
  {32'h3be91dc8, 32'h3d0db374} /* (31, 21, 21) {real, imag} */,
  {32'hbd46b9ae, 32'hbbbd1b9c} /* (31, 21, 20) {real, imag} */,
  {32'hbd895178, 32'h3d324d58} /* (31, 21, 19) {real, imag} */,
  {32'h3bc65ec8, 32'h3c813829} /* (31, 21, 18) {real, imag} */,
  {32'h3ca57d30, 32'hbc5a6966} /* (31, 21, 17) {real, imag} */,
  {32'h3cf369b1, 32'h00000000} /* (31, 21, 16) {real, imag} */,
  {32'h3ca57d30, 32'h3c5a6966} /* (31, 21, 15) {real, imag} */,
  {32'h3bc65ec8, 32'hbc813829} /* (31, 21, 14) {real, imag} */,
  {32'hbd895178, 32'hbd324d58} /* (31, 21, 13) {real, imag} */,
  {32'hbd46b9ae, 32'h3bbd1b9c} /* (31, 21, 12) {real, imag} */,
  {32'h3be91dc8, 32'hbd0db374} /* (31, 21, 11) {real, imag} */,
  {32'h3c7eadc3, 32'h3d12f304} /* (31, 21, 10) {real, imag} */,
  {32'hbda657f4, 32'hbd23c0ad} /* (31, 21, 9) {real, imag} */,
  {32'h3d1a849a, 32'h3c66216c} /* (31, 21, 8) {real, imag} */,
  {32'hbcf02309, 32'hbcf5f784} /* (31, 21, 7) {real, imag} */,
  {32'hbd6d730e, 32'h3c837aa3} /* (31, 21, 6) {real, imag} */,
  {32'hbd9781f8, 32'h3b4055c8} /* (31, 21, 5) {real, imag} */,
  {32'hbdb55600, 32'h3d6c0395} /* (31, 21, 4) {real, imag} */,
  {32'h3ddd6a28, 32'hbd910ff2} /* (31, 21, 3) {real, imag} */,
  {32'hbe250786, 32'hbd154c93} /* (31, 21, 2) {real, imag} */,
  {32'h3b064600, 32'hbdcd1da6} /* (31, 21, 1) {real, imag} */,
  {32'h3e29b110, 32'h00000000} /* (31, 21, 0) {real, imag} */,
  {32'hbef7b100, 32'h3d8307fe} /* (31, 20, 31) {real, imag} */,
  {32'h3e2fa0e0, 32'hbe4c94ec} /* (31, 20, 30) {real, imag} */,
  {32'h3da985e1, 32'h3dbb88da} /* (31, 20, 29) {real, imag} */,
  {32'hbe30be2d, 32'h3d2f58c5} /* (31, 20, 28) {real, imag} */,
  {32'h3d828483, 32'h3c21c40c} /* (31, 20, 27) {real, imag} */,
  {32'hb8ea77c0, 32'hbda2feb8} /* (31, 20, 26) {real, imag} */,
  {32'h3d0babc8, 32'hbd2b65bf} /* (31, 20, 25) {real, imag} */,
  {32'h3adb53c0, 32'h3d1ea775} /* (31, 20, 24) {real, imag} */,
  {32'hbd1212b6, 32'h3d354348} /* (31, 20, 23) {real, imag} */,
  {32'h3cb4fc42, 32'hbd695d8c} /* (31, 20, 22) {real, imag} */,
  {32'hbd9a3e4e, 32'hbd4e9ebd} /* (31, 20, 21) {real, imag} */,
  {32'hbd9eedac, 32'hbc5690e8} /* (31, 20, 20) {real, imag} */,
  {32'h3cdceefe, 32'h3d9ed2e1} /* (31, 20, 19) {real, imag} */,
  {32'hbc0bb260, 32'hbbf44d30} /* (31, 20, 18) {real, imag} */,
  {32'hb9ee0c80, 32'h3d4f0855} /* (31, 20, 17) {real, imag} */,
  {32'hbc9f84a7, 32'h00000000} /* (31, 20, 16) {real, imag} */,
  {32'hb9ee0c80, 32'hbd4f0855} /* (31, 20, 15) {real, imag} */,
  {32'hbc0bb260, 32'h3bf44d30} /* (31, 20, 14) {real, imag} */,
  {32'h3cdceefe, 32'hbd9ed2e1} /* (31, 20, 13) {real, imag} */,
  {32'hbd9eedac, 32'h3c5690e8} /* (31, 20, 12) {real, imag} */,
  {32'hbd9a3e4e, 32'h3d4e9ebd} /* (31, 20, 11) {real, imag} */,
  {32'h3cb4fc42, 32'h3d695d8c} /* (31, 20, 10) {real, imag} */,
  {32'hbd1212b6, 32'hbd354348} /* (31, 20, 9) {real, imag} */,
  {32'h3adb53c0, 32'hbd1ea775} /* (31, 20, 8) {real, imag} */,
  {32'h3d0babc8, 32'h3d2b65bf} /* (31, 20, 7) {real, imag} */,
  {32'hb8ea77c0, 32'h3da2feb8} /* (31, 20, 6) {real, imag} */,
  {32'h3d828483, 32'hbc21c40c} /* (31, 20, 5) {real, imag} */,
  {32'hbe30be2d, 32'hbd2f58c5} /* (31, 20, 4) {real, imag} */,
  {32'h3da985e1, 32'hbdbb88da} /* (31, 20, 3) {real, imag} */,
  {32'h3e2fa0e0, 32'h3e4c94ec} /* (31, 20, 2) {real, imag} */,
  {32'hbef7b100, 32'hbd8307fe} /* (31, 20, 1) {real, imag} */,
  {32'hbeae5500, 32'h00000000} /* (31, 20, 0) {real, imag} */,
  {32'hbf4afe9a, 32'h3d1efef0} /* (31, 19, 31) {real, imag} */,
  {32'h3eb303e8, 32'hbe37f0c8} /* (31, 19, 30) {real, imag} */,
  {32'hbc2c4bc6, 32'h3d8c467a} /* (31, 19, 29) {real, imag} */,
  {32'hbe3e77db, 32'hbd85d5ee} /* (31, 19, 28) {real, imag} */,
  {32'h3dcdb140, 32'hbddbd229} /* (31, 19, 27) {real, imag} */,
  {32'h3c848964, 32'h3d6ad2b9} /* (31, 19, 26) {real, imag} */,
  {32'hbc94d3ae, 32'h3d766f9c} /* (31, 19, 25) {real, imag} */,
  {32'hbd35f6ba, 32'hbcb36c10} /* (31, 19, 24) {real, imag} */,
  {32'h3c080985, 32'h3cfcc8b0} /* (31, 19, 23) {real, imag} */,
  {32'hbd5c9120, 32'hbd966fc4} /* (31, 19, 22) {real, imag} */,
  {32'hbd5cd2f1, 32'h3cdc6ec1} /* (31, 19, 21) {real, imag} */,
  {32'h3d16d3dc, 32'hbdaf4f3d} /* (31, 19, 20) {real, imag} */,
  {32'hbcdf72ca, 32'hbd931579} /* (31, 19, 19) {real, imag} */,
  {32'hbc8781bb, 32'hbdd922b2} /* (31, 19, 18) {real, imag} */,
  {32'hbba33488, 32'h3cefc944} /* (31, 19, 17) {real, imag} */,
  {32'h3cbfe1d6, 32'h00000000} /* (31, 19, 16) {real, imag} */,
  {32'hbba33488, 32'hbcefc944} /* (31, 19, 15) {real, imag} */,
  {32'hbc8781bb, 32'h3dd922b2} /* (31, 19, 14) {real, imag} */,
  {32'hbcdf72ca, 32'h3d931579} /* (31, 19, 13) {real, imag} */,
  {32'h3d16d3dc, 32'h3daf4f3d} /* (31, 19, 12) {real, imag} */,
  {32'hbd5cd2f1, 32'hbcdc6ec1} /* (31, 19, 11) {real, imag} */,
  {32'hbd5c9120, 32'h3d966fc4} /* (31, 19, 10) {real, imag} */,
  {32'h3c080985, 32'hbcfcc8b0} /* (31, 19, 9) {real, imag} */,
  {32'hbd35f6ba, 32'h3cb36c10} /* (31, 19, 8) {real, imag} */,
  {32'hbc94d3ae, 32'hbd766f9c} /* (31, 19, 7) {real, imag} */,
  {32'h3c848964, 32'hbd6ad2b9} /* (31, 19, 6) {real, imag} */,
  {32'h3dcdb140, 32'h3ddbd229} /* (31, 19, 5) {real, imag} */,
  {32'hbe3e77db, 32'h3d85d5ee} /* (31, 19, 4) {real, imag} */,
  {32'hbc2c4bc6, 32'hbd8c467a} /* (31, 19, 3) {real, imag} */,
  {32'h3eb303e8, 32'h3e37f0c8} /* (31, 19, 2) {real, imag} */,
  {32'hbf4afe9a, 32'hbd1efef0} /* (31, 19, 1) {real, imag} */,
  {32'hbeeed135, 32'h00000000} /* (31, 19, 0) {real, imag} */,
  {32'hbf53a90a, 32'hbd2d3beb} /* (31, 18, 31) {real, imag} */,
  {32'h3ea03c6c, 32'hbe06c17a} /* (31, 18, 30) {real, imag} */,
  {32'hbd2b3bb6, 32'h3dbd2c4d} /* (31, 18, 29) {real, imag} */,
  {32'hbe8776ff, 32'h3ce9a8d5} /* (31, 18, 28) {real, imag} */,
  {32'h3e048b1f, 32'hbd61865e} /* (31, 18, 27) {real, imag} */,
  {32'h3ba99dec, 32'hbb011e40} /* (31, 18, 26) {real, imag} */,
  {32'h3c778805, 32'hbc2edf16} /* (31, 18, 25) {real, imag} */,
  {32'h3d4f3ce0, 32'h3c064c1c} /* (31, 18, 24) {real, imag} */,
  {32'h3b0b9bb8, 32'h3d44e70c} /* (31, 18, 23) {real, imag} */,
  {32'h3d0a8487, 32'hbcc0de60} /* (31, 18, 22) {real, imag} */,
  {32'h3be7ecac, 32'h3c9678f2} /* (31, 18, 21) {real, imag} */,
  {32'h3d6824eb, 32'h3c63dc8c} /* (31, 18, 20) {real, imag} */,
  {32'h3dbf60cd, 32'h3c122e40} /* (31, 18, 19) {real, imag} */,
  {32'hbb872e22, 32'hbc4bacfe} /* (31, 18, 18) {real, imag} */,
  {32'h3c328088, 32'h3cbcda76} /* (31, 18, 17) {real, imag} */,
  {32'h3c4313fb, 32'h00000000} /* (31, 18, 16) {real, imag} */,
  {32'h3c328088, 32'hbcbcda76} /* (31, 18, 15) {real, imag} */,
  {32'hbb872e22, 32'h3c4bacfe} /* (31, 18, 14) {real, imag} */,
  {32'h3dbf60cd, 32'hbc122e40} /* (31, 18, 13) {real, imag} */,
  {32'h3d6824eb, 32'hbc63dc8c} /* (31, 18, 12) {real, imag} */,
  {32'h3be7ecac, 32'hbc9678f2} /* (31, 18, 11) {real, imag} */,
  {32'h3d0a8487, 32'h3cc0de60} /* (31, 18, 10) {real, imag} */,
  {32'h3b0b9bb8, 32'hbd44e70c} /* (31, 18, 9) {real, imag} */,
  {32'h3d4f3ce0, 32'hbc064c1c} /* (31, 18, 8) {real, imag} */,
  {32'h3c778805, 32'h3c2edf16} /* (31, 18, 7) {real, imag} */,
  {32'h3ba99dec, 32'h3b011e40} /* (31, 18, 6) {real, imag} */,
  {32'h3e048b1f, 32'h3d61865e} /* (31, 18, 5) {real, imag} */,
  {32'hbe8776ff, 32'hbce9a8d5} /* (31, 18, 4) {real, imag} */,
  {32'hbd2b3bb6, 32'hbdbd2c4d} /* (31, 18, 3) {real, imag} */,
  {32'h3ea03c6c, 32'h3e06c17a} /* (31, 18, 2) {real, imag} */,
  {32'hbf53a90a, 32'h3d2d3beb} /* (31, 18, 1) {real, imag} */,
  {32'hbeb518bb, 32'h00000000} /* (31, 18, 0) {real, imag} */,
  {32'hbf532f85, 32'hbe176cf1} /* (31, 17, 31) {real, imag} */,
  {32'h3e81587c, 32'hbd7b08a0} /* (31, 17, 30) {real, imag} */,
  {32'hbd69a700, 32'h3be46aa8} /* (31, 17, 29) {real, imag} */,
  {32'hbe186532, 32'h3ab82828} /* (31, 17, 28) {real, imag} */,
  {32'h3dce08bb, 32'hbd3733fb} /* (31, 17, 27) {real, imag} */,
  {32'hbc36faf3, 32'hbd08cd2b} /* (31, 17, 26) {real, imag} */,
  {32'hbd722c02, 32'h3d6200cd} /* (31, 17, 25) {real, imag} */,
  {32'h3ce6f0c0, 32'hbd929768} /* (31, 17, 24) {real, imag} */,
  {32'h3c268e9e, 32'hbd462382} /* (31, 17, 23) {real, imag} */,
  {32'hbcbf4967, 32'h3d01ca11} /* (31, 17, 22) {real, imag} */,
  {32'h3d71d9ce, 32'hbd33d88f} /* (31, 17, 21) {real, imag} */,
  {32'hbd8fe250, 32'hbc745ab7} /* (31, 17, 20) {real, imag} */,
  {32'h3cdf2d32, 32'h3b82b338} /* (31, 17, 19) {real, imag} */,
  {32'h3d1d2ba2, 32'hbd71fb9d} /* (31, 17, 18) {real, imag} */,
  {32'h3bedc480, 32'h3b829f34} /* (31, 17, 17) {real, imag} */,
  {32'h3d58e79f, 32'h00000000} /* (31, 17, 16) {real, imag} */,
  {32'h3bedc480, 32'hbb829f34} /* (31, 17, 15) {real, imag} */,
  {32'h3d1d2ba2, 32'h3d71fb9d} /* (31, 17, 14) {real, imag} */,
  {32'h3cdf2d32, 32'hbb82b338} /* (31, 17, 13) {real, imag} */,
  {32'hbd8fe250, 32'h3c745ab7} /* (31, 17, 12) {real, imag} */,
  {32'h3d71d9ce, 32'h3d33d88f} /* (31, 17, 11) {real, imag} */,
  {32'hbcbf4967, 32'hbd01ca11} /* (31, 17, 10) {real, imag} */,
  {32'h3c268e9e, 32'h3d462382} /* (31, 17, 9) {real, imag} */,
  {32'h3ce6f0c0, 32'h3d929768} /* (31, 17, 8) {real, imag} */,
  {32'hbd722c02, 32'hbd6200cd} /* (31, 17, 7) {real, imag} */,
  {32'hbc36faf3, 32'h3d08cd2b} /* (31, 17, 6) {real, imag} */,
  {32'h3dce08bb, 32'h3d3733fb} /* (31, 17, 5) {real, imag} */,
  {32'hbe186532, 32'hbab82828} /* (31, 17, 4) {real, imag} */,
  {32'hbd69a700, 32'hbbe46aa8} /* (31, 17, 3) {real, imag} */,
  {32'h3e81587c, 32'h3d7b08a0} /* (31, 17, 2) {real, imag} */,
  {32'hbf532f85, 32'h3e176cf1} /* (31, 17, 1) {real, imag} */,
  {32'hbebf0c9a, 32'h00000000} /* (31, 17, 0) {real, imag} */,
  {32'hbf42bdd8, 32'hbe26ac52} /* (31, 16, 31) {real, imag} */,
  {32'h3ea17533, 32'hbde7971e} /* (31, 16, 30) {real, imag} */,
  {32'hbd603081, 32'h3d8cd869} /* (31, 16, 29) {real, imag} */,
  {32'hbe0bbbb5, 32'h3bbbe650} /* (31, 16, 28) {real, imag} */,
  {32'h3dd03b02, 32'h3bc2f800} /* (31, 16, 27) {real, imag} */,
  {32'hbd33c628, 32'h3cc79be1} /* (31, 16, 26) {real, imag} */,
  {32'hbd6106e4, 32'hbd763793} /* (31, 16, 25) {real, imag} */,
  {32'h3dc069ba, 32'hbd81eae8} /* (31, 16, 24) {real, imag} */,
  {32'hbd0885d4, 32'hbd1be1f0} /* (31, 16, 23) {real, imag} */,
  {32'hbca074f4, 32'h3b0d7f68} /* (31, 16, 22) {real, imag} */,
  {32'hbcb54d5a, 32'hbc4e14f7} /* (31, 16, 21) {real, imag} */,
  {32'hbd223446, 32'hbd2652b5} /* (31, 16, 20) {real, imag} */,
  {32'h3cd8baf6, 32'hbca1def6} /* (31, 16, 19) {real, imag} */,
  {32'h3c393810, 32'h3cf9e8f6} /* (31, 16, 18) {real, imag} */,
  {32'hbd2b38ab, 32'h3c844c1e} /* (31, 16, 17) {real, imag} */,
  {32'h3d03f96d, 32'h00000000} /* (31, 16, 16) {real, imag} */,
  {32'hbd2b38ab, 32'hbc844c1e} /* (31, 16, 15) {real, imag} */,
  {32'h3c393810, 32'hbcf9e8f6} /* (31, 16, 14) {real, imag} */,
  {32'h3cd8baf6, 32'h3ca1def6} /* (31, 16, 13) {real, imag} */,
  {32'hbd223446, 32'h3d2652b5} /* (31, 16, 12) {real, imag} */,
  {32'hbcb54d5a, 32'h3c4e14f7} /* (31, 16, 11) {real, imag} */,
  {32'hbca074f4, 32'hbb0d7f68} /* (31, 16, 10) {real, imag} */,
  {32'hbd0885d4, 32'h3d1be1f0} /* (31, 16, 9) {real, imag} */,
  {32'h3dc069ba, 32'h3d81eae8} /* (31, 16, 8) {real, imag} */,
  {32'hbd6106e4, 32'h3d763793} /* (31, 16, 7) {real, imag} */,
  {32'hbd33c628, 32'hbcc79be1} /* (31, 16, 6) {real, imag} */,
  {32'h3dd03b02, 32'hbbc2f800} /* (31, 16, 5) {real, imag} */,
  {32'hbe0bbbb5, 32'hbbbbe650} /* (31, 16, 4) {real, imag} */,
  {32'hbd603081, 32'hbd8cd869} /* (31, 16, 3) {real, imag} */,
  {32'h3ea17533, 32'h3de7971e} /* (31, 16, 2) {real, imag} */,
  {32'hbf42bdd8, 32'h3e26ac52} /* (31, 16, 1) {real, imag} */,
  {32'hbf023467, 32'h00000000} /* (31, 16, 0) {real, imag} */,
  {32'hbf2bbffb, 32'hbe0edc53} /* (31, 15, 31) {real, imag} */,
  {32'h3e91341c, 32'hbdd51164} /* (31, 15, 30) {real, imag} */,
  {32'hbd6c305c, 32'h3db07aac} /* (31, 15, 29) {real, imag} */,
  {32'hbd8e9a53, 32'h3c862a0e} /* (31, 15, 28) {real, imag} */,
  {32'h3dd8dff9, 32'h3d90fc28} /* (31, 15, 27) {real, imag} */,
  {32'h39a1db20, 32'hbc37dce0} /* (31, 15, 26) {real, imag} */,
  {32'h3c00f470, 32'hbd061df9} /* (31, 15, 25) {real, imag} */,
  {32'h3ce4dc04, 32'hbc96bb5e} /* (31, 15, 24) {real, imag} */,
  {32'h3ce949a1, 32'h3c9433b8} /* (31, 15, 23) {real, imag} */,
  {32'hbc8a4931, 32'hbd9fd9d6} /* (31, 15, 22) {real, imag} */,
  {32'h3b5c40e0, 32'hbcf359f6} /* (31, 15, 21) {real, imag} */,
  {32'h3da158a0, 32'h3c95425a} /* (31, 15, 20) {real, imag} */,
  {32'h3d7f82cd, 32'h3d3697c1} /* (31, 15, 19) {real, imag} */,
  {32'h3c68b04b, 32'h3ca889d6} /* (31, 15, 18) {real, imag} */,
  {32'h3d27d79a, 32'h3d0f53ae} /* (31, 15, 17) {real, imag} */,
  {32'h3ceee59a, 32'h00000000} /* (31, 15, 16) {real, imag} */,
  {32'h3d27d79a, 32'hbd0f53ae} /* (31, 15, 15) {real, imag} */,
  {32'h3c68b04b, 32'hbca889d6} /* (31, 15, 14) {real, imag} */,
  {32'h3d7f82cd, 32'hbd3697c1} /* (31, 15, 13) {real, imag} */,
  {32'h3da158a0, 32'hbc95425a} /* (31, 15, 12) {real, imag} */,
  {32'h3b5c40e0, 32'h3cf359f6} /* (31, 15, 11) {real, imag} */,
  {32'hbc8a4931, 32'h3d9fd9d6} /* (31, 15, 10) {real, imag} */,
  {32'h3ce949a1, 32'hbc9433b8} /* (31, 15, 9) {real, imag} */,
  {32'h3ce4dc04, 32'h3c96bb5e} /* (31, 15, 8) {real, imag} */,
  {32'h3c00f470, 32'h3d061df9} /* (31, 15, 7) {real, imag} */,
  {32'h39a1db20, 32'h3c37dce0} /* (31, 15, 6) {real, imag} */,
  {32'h3dd8dff9, 32'hbd90fc28} /* (31, 15, 5) {real, imag} */,
  {32'hbd8e9a53, 32'hbc862a0e} /* (31, 15, 4) {real, imag} */,
  {32'hbd6c305c, 32'hbdb07aac} /* (31, 15, 3) {real, imag} */,
  {32'h3e91341c, 32'h3dd51164} /* (31, 15, 2) {real, imag} */,
  {32'hbf2bbffb, 32'h3e0edc53} /* (31, 15, 1) {real, imag} */,
  {32'hbf1853e1, 32'h00000000} /* (31, 15, 0) {real, imag} */,
  {32'hbf092f0c, 32'hbddfca0a} /* (31, 14, 31) {real, imag} */,
  {32'h3ea5ae28, 32'h3c9d2ad4} /* (31, 14, 30) {real, imag} */,
  {32'hbc90b0a0, 32'h3d29819e} /* (31, 14, 29) {real, imag} */,
  {32'h3ca5f75c, 32'h3d6cf3f2} /* (31, 14, 28) {real, imag} */,
  {32'h3d751a55, 32'h3cc44e44} /* (31, 14, 27) {real, imag} */,
  {32'h3d1588a6, 32'hb91b3100} /* (31, 14, 26) {real, imag} */,
  {32'hbd2a3fad, 32'h3d83cfb3} /* (31, 14, 25) {real, imag} */,
  {32'h3d45febe, 32'hbd732423} /* (31, 14, 24) {real, imag} */,
  {32'hbbefb44c, 32'hbc787ab8} /* (31, 14, 23) {real, imag} */,
  {32'h3c5efb1c, 32'h3ce52e08} /* (31, 14, 22) {real, imag} */,
  {32'h3d829d2c, 32'h3c3d83c9} /* (31, 14, 21) {real, imag} */,
  {32'hbda2105e, 32'hbb848730} /* (31, 14, 20) {real, imag} */,
  {32'hbcdfa17c, 32'hbc562d8c} /* (31, 14, 19) {real, imag} */,
  {32'hbca598b8, 32'hbc651fb6} /* (31, 14, 18) {real, imag} */,
  {32'h3ba4ac0f, 32'h3c389bdc} /* (31, 14, 17) {real, imag} */,
  {32'h3bcc129a, 32'h00000000} /* (31, 14, 16) {real, imag} */,
  {32'h3ba4ac0f, 32'hbc389bdc} /* (31, 14, 15) {real, imag} */,
  {32'hbca598b8, 32'h3c651fb6} /* (31, 14, 14) {real, imag} */,
  {32'hbcdfa17c, 32'h3c562d8c} /* (31, 14, 13) {real, imag} */,
  {32'hbda2105e, 32'h3b848730} /* (31, 14, 12) {real, imag} */,
  {32'h3d829d2c, 32'hbc3d83c9} /* (31, 14, 11) {real, imag} */,
  {32'h3c5efb1c, 32'hbce52e08} /* (31, 14, 10) {real, imag} */,
  {32'hbbefb44c, 32'h3c787ab8} /* (31, 14, 9) {real, imag} */,
  {32'h3d45febe, 32'h3d732423} /* (31, 14, 8) {real, imag} */,
  {32'hbd2a3fad, 32'hbd83cfb3} /* (31, 14, 7) {real, imag} */,
  {32'h3d1588a6, 32'h391b3100} /* (31, 14, 6) {real, imag} */,
  {32'h3d751a55, 32'hbcc44e44} /* (31, 14, 5) {real, imag} */,
  {32'h3ca5f75c, 32'hbd6cf3f2} /* (31, 14, 4) {real, imag} */,
  {32'hbc90b0a0, 32'hbd29819e} /* (31, 14, 3) {real, imag} */,
  {32'h3ea5ae28, 32'hbc9d2ad4} /* (31, 14, 2) {real, imag} */,
  {32'hbf092f0c, 32'h3ddfca0a} /* (31, 14, 1) {real, imag} */,
  {32'hbf273b1e, 32'h00000000} /* (31, 14, 0) {real, imag} */,
  {32'hbf011068, 32'hbdc48184} /* (31, 13, 31) {real, imag} */,
  {32'h3ed5f904, 32'hbdb13f80} /* (31, 13, 30) {real, imag} */,
  {32'hbd5bfc5e, 32'h3d59dc28} /* (31, 13, 29) {real, imag} */,
  {32'hbdf03132, 32'h3d026dcc} /* (31, 13, 28) {real, imag} */,
  {32'h3d3960db, 32'h3b45e560} /* (31, 13, 27) {real, imag} */,
  {32'h3d45872c, 32'hbccaf876} /* (31, 13, 26) {real, imag} */,
  {32'h3d0e977b, 32'h3d5d8dac} /* (31, 13, 25) {real, imag} */,
  {32'h3c6a3732, 32'hbd316052} /* (31, 13, 24) {real, imag} */,
  {32'h3c01309b, 32'hbd68d9fc} /* (31, 13, 23) {real, imag} */,
  {32'h3d567610, 32'h3cb8f926} /* (31, 13, 22) {real, imag} */,
  {32'hbb067340, 32'h3d40f474} /* (31, 13, 21) {real, imag} */,
  {32'hbd932ec7, 32'hbce69c1b} /* (31, 13, 20) {real, imag} */,
  {32'h3cd7b438, 32'h3c82c8bc} /* (31, 13, 19) {real, imag} */,
  {32'h38aca300, 32'h3c1fc4ac} /* (31, 13, 18) {real, imag} */,
  {32'h3bb47050, 32'hbca8df44} /* (31, 13, 17) {real, imag} */,
  {32'hbd345879, 32'h00000000} /* (31, 13, 16) {real, imag} */,
  {32'h3bb47050, 32'h3ca8df44} /* (31, 13, 15) {real, imag} */,
  {32'h38aca300, 32'hbc1fc4ac} /* (31, 13, 14) {real, imag} */,
  {32'h3cd7b438, 32'hbc82c8bc} /* (31, 13, 13) {real, imag} */,
  {32'hbd932ec7, 32'h3ce69c1b} /* (31, 13, 12) {real, imag} */,
  {32'hbb067340, 32'hbd40f474} /* (31, 13, 11) {real, imag} */,
  {32'h3d567610, 32'hbcb8f926} /* (31, 13, 10) {real, imag} */,
  {32'h3c01309b, 32'h3d68d9fc} /* (31, 13, 9) {real, imag} */,
  {32'h3c6a3732, 32'h3d316052} /* (31, 13, 8) {real, imag} */,
  {32'h3d0e977b, 32'hbd5d8dac} /* (31, 13, 7) {real, imag} */,
  {32'h3d45872c, 32'h3ccaf876} /* (31, 13, 6) {real, imag} */,
  {32'h3d3960db, 32'hbb45e560} /* (31, 13, 5) {real, imag} */,
  {32'hbdf03132, 32'hbd026dcc} /* (31, 13, 4) {real, imag} */,
  {32'hbd5bfc5e, 32'hbd59dc28} /* (31, 13, 3) {real, imag} */,
  {32'h3ed5f904, 32'h3db13f80} /* (31, 13, 2) {real, imag} */,
  {32'hbf011068, 32'h3dc48184} /* (31, 13, 1) {real, imag} */,
  {32'hbf30a0d8, 32'h00000000} /* (31, 13, 0) {real, imag} */,
  {32'hbef64d92, 32'hb83e3000} /* (31, 12, 31) {real, imag} */,
  {32'h3ec075d0, 32'hbd938c41} /* (31, 12, 30) {real, imag} */,
  {32'hbd91c6b3, 32'h3d8c2a42} /* (31, 12, 29) {real, imag} */,
  {32'hbddece3e, 32'h3c4cc33d} /* (31, 12, 28) {real, imag} */,
  {32'h3ab21b30, 32'hbdba70e4} /* (31, 12, 27) {real, imag} */,
  {32'hba7ef8c8, 32'h3c76bc74} /* (31, 12, 26) {real, imag} */,
  {32'hbdc6af64, 32'h3d84b6c8} /* (31, 12, 25) {real, imag} */,
  {32'h3db2f17f, 32'hbbbad4c8} /* (31, 12, 24) {real, imag} */,
  {32'h3d2bdd5e, 32'hbd6dda90} /* (31, 12, 23) {real, imag} */,
  {32'h3befadca, 32'hbd370a74} /* (31, 12, 22) {real, imag} */,
  {32'hbd58fb71, 32'hbcb72c56} /* (31, 12, 21) {real, imag} */,
  {32'h3ab375a0, 32'hbb62bd22} /* (31, 12, 20) {real, imag} */,
  {32'h3c260ae4, 32'hbda32895} /* (31, 12, 19) {real, imag} */,
  {32'h3ddb4424, 32'hbc6ceb10} /* (31, 12, 18) {real, imag} */,
  {32'hbd158ed2, 32'hbc88f942} /* (31, 12, 17) {real, imag} */,
  {32'hbd31a466, 32'h00000000} /* (31, 12, 16) {real, imag} */,
  {32'hbd158ed2, 32'h3c88f942} /* (31, 12, 15) {real, imag} */,
  {32'h3ddb4424, 32'h3c6ceb10} /* (31, 12, 14) {real, imag} */,
  {32'h3c260ae4, 32'h3da32895} /* (31, 12, 13) {real, imag} */,
  {32'h3ab375a0, 32'h3b62bd22} /* (31, 12, 12) {real, imag} */,
  {32'hbd58fb71, 32'h3cb72c56} /* (31, 12, 11) {real, imag} */,
  {32'h3befadca, 32'h3d370a74} /* (31, 12, 10) {real, imag} */,
  {32'h3d2bdd5e, 32'h3d6dda90} /* (31, 12, 9) {real, imag} */,
  {32'h3db2f17f, 32'h3bbad4c8} /* (31, 12, 8) {real, imag} */,
  {32'hbdc6af64, 32'hbd84b6c8} /* (31, 12, 7) {real, imag} */,
  {32'hba7ef8c8, 32'hbc76bc74} /* (31, 12, 6) {real, imag} */,
  {32'h3ab21b30, 32'h3dba70e4} /* (31, 12, 5) {real, imag} */,
  {32'hbddece3e, 32'hbc4cc33d} /* (31, 12, 4) {real, imag} */,
  {32'hbd91c6b3, 32'hbd8c2a42} /* (31, 12, 3) {real, imag} */,
  {32'h3ec075d0, 32'h3d938c41} /* (31, 12, 2) {real, imag} */,
  {32'hbef64d92, 32'h383e3000} /* (31, 12, 1) {real, imag} */,
  {32'hbf28df90, 32'h00000000} /* (31, 12, 0) {real, imag} */,
  {32'hbe82e638, 32'h3ca48a98} /* (31, 11, 31) {real, imag} */,
  {32'h3e78da9a, 32'h3d0c08a1} /* (31, 11, 30) {real, imag} */,
  {32'hbd458fed, 32'hbca91446} /* (31, 11, 29) {real, imag} */,
  {32'h3d09f048, 32'h3d763eff} /* (31, 11, 28) {real, imag} */,
  {32'h3db8a14e, 32'hbd85574c} /* (31, 11, 27) {real, imag} */,
  {32'h3c04209a, 32'h3d51ccd4} /* (31, 11, 26) {real, imag} */,
  {32'hbd90824f, 32'hbafeb220} /* (31, 11, 25) {real, imag} */,
  {32'h3d73202a, 32'h3c1ad730} /* (31, 11, 24) {real, imag} */,
  {32'h3d8f3cd2, 32'hbd085fcf} /* (31, 11, 23) {real, imag} */,
  {32'h3ca27fdc, 32'h3d6118b4} /* (31, 11, 22) {real, imag} */,
  {32'h3dc7f3e0, 32'hbd5f9cee} /* (31, 11, 21) {real, imag} */,
  {32'hbdbf5ac1, 32'h3d10df72} /* (31, 11, 20) {real, imag} */,
  {32'hbd8192cc, 32'hbd255c5a} /* (31, 11, 19) {real, imag} */,
  {32'hbca7cb2a, 32'h3b319e58} /* (31, 11, 18) {real, imag} */,
  {32'hbb2ec194, 32'hbcadca19} /* (31, 11, 17) {real, imag} */,
  {32'h3d1ffa9c, 32'h00000000} /* (31, 11, 16) {real, imag} */,
  {32'hbb2ec194, 32'h3cadca19} /* (31, 11, 15) {real, imag} */,
  {32'hbca7cb2a, 32'hbb319e58} /* (31, 11, 14) {real, imag} */,
  {32'hbd8192cc, 32'h3d255c5a} /* (31, 11, 13) {real, imag} */,
  {32'hbdbf5ac1, 32'hbd10df72} /* (31, 11, 12) {real, imag} */,
  {32'h3dc7f3e0, 32'h3d5f9cee} /* (31, 11, 11) {real, imag} */,
  {32'h3ca27fdc, 32'hbd6118b4} /* (31, 11, 10) {real, imag} */,
  {32'h3d8f3cd2, 32'h3d085fcf} /* (31, 11, 9) {real, imag} */,
  {32'h3d73202a, 32'hbc1ad730} /* (31, 11, 8) {real, imag} */,
  {32'hbd90824f, 32'h3afeb220} /* (31, 11, 7) {real, imag} */,
  {32'h3c04209a, 32'hbd51ccd4} /* (31, 11, 6) {real, imag} */,
  {32'h3db8a14e, 32'h3d85574c} /* (31, 11, 5) {real, imag} */,
  {32'h3d09f048, 32'hbd763eff} /* (31, 11, 4) {real, imag} */,
  {32'hbd458fed, 32'h3ca91446} /* (31, 11, 3) {real, imag} */,
  {32'h3e78da9a, 32'hbd0c08a1} /* (31, 11, 2) {real, imag} */,
  {32'hbe82e638, 32'hbca48a98} /* (31, 11, 1) {real, imag} */,
  {32'hbea1e3c1, 32'h00000000} /* (31, 11, 0) {real, imag} */,
  {32'h3e9c28bd, 32'h3d3513fb} /* (31, 10, 31) {real, imag} */,
  {32'hbe27fb8b, 32'h3dec3bea} /* (31, 10, 30) {real, imag} */,
  {32'h3d4685e8, 32'hbdeeecde} /* (31, 10, 29) {real, imag} */,
  {32'h3dac3c32, 32'h3cb8537f} /* (31, 10, 28) {real, imag} */,
  {32'h3b9a9b50, 32'hbe0d3a9e} /* (31, 10, 27) {real, imag} */,
  {32'hbc8f6dba, 32'h3ce77efb} /* (31, 10, 26) {real, imag} */,
  {32'hbcf75c40, 32'hbdd95afc} /* (31, 10, 25) {real, imag} */,
  {32'h3c30bcd4, 32'h3d50cfd3} /* (31, 10, 24) {real, imag} */,
  {32'hbd72a842, 32'hbd72887e} /* (31, 10, 23) {real, imag} */,
  {32'hbd4f351a, 32'h3d527988} /* (31, 10, 22) {real, imag} */,
  {32'hbd636dc8, 32'hbd9f035d} /* (31, 10, 21) {real, imag} */,
  {32'hbd20d244, 32'h3c51dabb} /* (31, 10, 20) {real, imag} */,
  {32'hbd9660ec, 32'hbba17be8} /* (31, 10, 19) {real, imag} */,
  {32'h3e01fe72, 32'h3d3861e5} /* (31, 10, 18) {real, imag} */,
  {32'hbd3d46e3, 32'hbd5ee7de} /* (31, 10, 17) {real, imag} */,
  {32'h3be9d420, 32'h00000000} /* (31, 10, 16) {real, imag} */,
  {32'hbd3d46e3, 32'h3d5ee7de} /* (31, 10, 15) {real, imag} */,
  {32'h3e01fe72, 32'hbd3861e5} /* (31, 10, 14) {real, imag} */,
  {32'hbd9660ec, 32'h3ba17be8} /* (31, 10, 13) {real, imag} */,
  {32'hbd20d244, 32'hbc51dabb} /* (31, 10, 12) {real, imag} */,
  {32'hbd636dc8, 32'h3d9f035d} /* (31, 10, 11) {real, imag} */,
  {32'hbd4f351a, 32'hbd527988} /* (31, 10, 10) {real, imag} */,
  {32'hbd72a842, 32'h3d72887e} /* (31, 10, 9) {real, imag} */,
  {32'h3c30bcd4, 32'hbd50cfd3} /* (31, 10, 8) {real, imag} */,
  {32'hbcf75c40, 32'h3dd95afc} /* (31, 10, 7) {real, imag} */,
  {32'hbc8f6dba, 32'hbce77efb} /* (31, 10, 6) {real, imag} */,
  {32'h3b9a9b50, 32'h3e0d3a9e} /* (31, 10, 5) {real, imag} */,
  {32'h3dac3c32, 32'hbcb8537f} /* (31, 10, 4) {real, imag} */,
  {32'h3d4685e8, 32'h3deeecde} /* (31, 10, 3) {real, imag} */,
  {32'hbe27fb8b, 32'hbdec3bea} /* (31, 10, 2) {real, imag} */,
  {32'h3e9c28bd, 32'hbd3513fb} /* (31, 10, 1) {real, imag} */,
  {32'h3c6d1990, 32'h00000000} /* (31, 10, 0) {real, imag} */,
  {32'h3f17dab0, 32'h3a896b58} /* (31, 9, 31) {real, imag} */,
  {32'hbe94fea3, 32'h3e3faf52} /* (31, 9, 30) {real, imag} */,
  {32'h3ce3d4bc, 32'hbcdc95f8} /* (31, 9, 29) {real, imag} */,
  {32'h3dbd9902, 32'hbd53f8bb} /* (31, 9, 28) {real, imag} */,
  {32'hbd086dd5, 32'hbb744b30} /* (31, 9, 27) {real, imag} */,
  {32'hbcdf9fe4, 32'hbd9ff680} /* (31, 9, 26) {real, imag} */,
  {32'hbb643630, 32'hbdf37c49} /* (31, 9, 25) {real, imag} */,
  {32'h3b86b9c0, 32'hba493f60} /* (31, 9, 24) {real, imag} */,
  {32'hbc9f64b6, 32'h3d23ac3c} /* (31, 9, 23) {real, imag} */,
  {32'hbb2e6310, 32'h3c49daea} /* (31, 9, 22) {real, imag} */,
  {32'hbdc1af58, 32'h3bcc7540} /* (31, 9, 21) {real, imag} */,
  {32'hbd5a9bad, 32'h3d42e674} /* (31, 9, 20) {real, imag} */,
  {32'hbc5d5714, 32'hbd5a0603} /* (31, 9, 19) {real, imag} */,
  {32'hbd57b514, 32'hbcd05dd4} /* (31, 9, 18) {real, imag} */,
  {32'hbceb9c90, 32'h3d5479e3} /* (31, 9, 17) {real, imag} */,
  {32'h3d6d1ffb, 32'h00000000} /* (31, 9, 16) {real, imag} */,
  {32'hbceb9c90, 32'hbd5479e3} /* (31, 9, 15) {real, imag} */,
  {32'hbd57b514, 32'h3cd05dd4} /* (31, 9, 14) {real, imag} */,
  {32'hbc5d5714, 32'h3d5a0603} /* (31, 9, 13) {real, imag} */,
  {32'hbd5a9bad, 32'hbd42e674} /* (31, 9, 12) {real, imag} */,
  {32'hbdc1af58, 32'hbbcc7540} /* (31, 9, 11) {real, imag} */,
  {32'hbb2e6310, 32'hbc49daea} /* (31, 9, 10) {real, imag} */,
  {32'hbc9f64b6, 32'hbd23ac3c} /* (31, 9, 9) {real, imag} */,
  {32'h3b86b9c0, 32'h3a493f60} /* (31, 9, 8) {real, imag} */,
  {32'hbb643630, 32'h3df37c49} /* (31, 9, 7) {real, imag} */,
  {32'hbcdf9fe4, 32'h3d9ff680} /* (31, 9, 6) {real, imag} */,
  {32'hbd086dd5, 32'h3b744b30} /* (31, 9, 5) {real, imag} */,
  {32'h3dbd9902, 32'h3d53f8bb} /* (31, 9, 4) {real, imag} */,
  {32'h3ce3d4bc, 32'h3cdc95f8} /* (31, 9, 3) {real, imag} */,
  {32'hbe94fea3, 32'hbe3faf52} /* (31, 9, 2) {real, imag} */,
  {32'h3f17dab0, 32'hba896b58} /* (31, 9, 1) {real, imag} */,
  {32'h3e83d4e4, 32'h00000000} /* (31, 9, 0) {real, imag} */,
  {32'h3f2d3502, 32'hbd855a40} /* (31, 8, 31) {real, imag} */,
  {32'hbe884ace, 32'h3e06031d} /* (31, 8, 30) {real, imag} */,
  {32'hbdd83c42, 32'h3ced1920} /* (31, 8, 29) {real, imag} */,
  {32'h3e1f8efc, 32'hb89a3800} /* (31, 8, 28) {real, imag} */,
  {32'hbc1246e4, 32'h3d7d75ae} /* (31, 8, 27) {real, imag} */,
  {32'hbcbd5630, 32'hbd2ff72a} /* (31, 8, 26) {real, imag} */,
  {32'h3c9e8002, 32'hba757240} /* (31, 8, 25) {real, imag} */,
  {32'hbce99202, 32'h3b39f548} /* (31, 8, 24) {real, imag} */,
  {32'h3ca63d22, 32'hbb9850c0} /* (31, 8, 23) {real, imag} */,
  {32'h3c3c9e05, 32'hbbb43ac0} /* (31, 8, 22) {real, imag} */,
  {32'hbc19c995, 32'h3db1731f} /* (31, 8, 21) {real, imag} */,
  {32'h3ce2b162, 32'h3d13b075} /* (31, 8, 20) {real, imag} */,
  {32'hbd90598d, 32'hbd3308ea} /* (31, 8, 19) {real, imag} */,
  {32'h3ce06cc5, 32'hbc8a73d9} /* (31, 8, 18) {real, imag} */,
  {32'h3c8f1238, 32'h3d16d8c5} /* (31, 8, 17) {real, imag} */,
  {32'hbb801648, 32'h00000000} /* (31, 8, 16) {real, imag} */,
  {32'h3c8f1238, 32'hbd16d8c5} /* (31, 8, 15) {real, imag} */,
  {32'h3ce06cc5, 32'h3c8a73d9} /* (31, 8, 14) {real, imag} */,
  {32'hbd90598d, 32'h3d3308ea} /* (31, 8, 13) {real, imag} */,
  {32'h3ce2b162, 32'hbd13b075} /* (31, 8, 12) {real, imag} */,
  {32'hbc19c995, 32'hbdb1731f} /* (31, 8, 11) {real, imag} */,
  {32'h3c3c9e05, 32'h3bb43ac0} /* (31, 8, 10) {real, imag} */,
  {32'h3ca63d22, 32'h3b9850c0} /* (31, 8, 9) {real, imag} */,
  {32'hbce99202, 32'hbb39f548} /* (31, 8, 8) {real, imag} */,
  {32'h3c9e8002, 32'h3a757240} /* (31, 8, 7) {real, imag} */,
  {32'hbcbd5630, 32'h3d2ff72a} /* (31, 8, 6) {real, imag} */,
  {32'hbc1246e4, 32'hbd7d75ae} /* (31, 8, 5) {real, imag} */,
  {32'h3e1f8efc, 32'h389a3800} /* (31, 8, 4) {real, imag} */,
  {32'hbdd83c42, 32'hbced1920} /* (31, 8, 3) {real, imag} */,
  {32'hbe884ace, 32'hbe06031d} /* (31, 8, 2) {real, imag} */,
  {32'h3f2d3502, 32'h3d855a40} /* (31, 8, 1) {real, imag} */,
  {32'h3e6daba5, 32'h00000000} /* (31, 8, 0) {real, imag} */,
  {32'h3f314943, 32'h3cf8cc5a} /* (31, 7, 31) {real, imag} */,
  {32'hbe2f94ab, 32'h3e4f9568} /* (31, 7, 30) {real, imag} */,
  {32'hbdb5fde2, 32'hbdcf2a6b} /* (31, 7, 29) {real, imag} */,
  {32'h3e17e195, 32'hbd1d9934} /* (31, 7, 28) {real, imag} */,
  {32'hbd701eb7, 32'hbcdfb0ea} /* (31, 7, 27) {real, imag} */,
  {32'hbdaa79bd, 32'h3d4a3a8a} /* (31, 7, 26) {real, imag} */,
  {32'h3d5770ba, 32'hbd8e3a29} /* (31, 7, 25) {real, imag} */,
  {32'hbd9b8c49, 32'hbcd0377a} /* (31, 7, 24) {real, imag} */,
  {32'hbc9d2e8b, 32'hbd27216a} /* (31, 7, 23) {real, imag} */,
  {32'h3d9686c6, 32'hbc23364e} /* (31, 7, 22) {real, imag} */,
  {32'hbdd9e840, 32'h3d4f5f18} /* (31, 7, 21) {real, imag} */,
  {32'hbbeea6b8, 32'hbd477e28} /* (31, 7, 20) {real, imag} */,
  {32'h3d1658ec, 32'hbd3d141c} /* (31, 7, 19) {real, imag} */,
  {32'h3ce34c65, 32'h3d6ccdf4} /* (31, 7, 18) {real, imag} */,
  {32'hbbcb7b7c, 32'hbcb1c0ee} /* (31, 7, 17) {real, imag} */,
  {32'hbd30ea48, 32'h00000000} /* (31, 7, 16) {real, imag} */,
  {32'hbbcb7b7c, 32'h3cb1c0ee} /* (31, 7, 15) {real, imag} */,
  {32'h3ce34c65, 32'hbd6ccdf4} /* (31, 7, 14) {real, imag} */,
  {32'h3d1658ec, 32'h3d3d141c} /* (31, 7, 13) {real, imag} */,
  {32'hbbeea6b8, 32'h3d477e28} /* (31, 7, 12) {real, imag} */,
  {32'hbdd9e840, 32'hbd4f5f18} /* (31, 7, 11) {real, imag} */,
  {32'h3d9686c6, 32'h3c23364e} /* (31, 7, 10) {real, imag} */,
  {32'hbc9d2e8b, 32'h3d27216a} /* (31, 7, 9) {real, imag} */,
  {32'hbd9b8c49, 32'h3cd0377a} /* (31, 7, 8) {real, imag} */,
  {32'h3d5770ba, 32'h3d8e3a29} /* (31, 7, 7) {real, imag} */,
  {32'hbdaa79bd, 32'hbd4a3a8a} /* (31, 7, 6) {real, imag} */,
  {32'hbd701eb7, 32'h3cdfb0ea} /* (31, 7, 5) {real, imag} */,
  {32'h3e17e195, 32'h3d1d9934} /* (31, 7, 4) {real, imag} */,
  {32'hbdb5fde2, 32'h3dcf2a6b} /* (31, 7, 3) {real, imag} */,
  {32'hbe2f94ab, 32'hbe4f9568} /* (31, 7, 2) {real, imag} */,
  {32'h3f314943, 32'hbcf8cc5a} /* (31, 7, 1) {real, imag} */,
  {32'h3e66fc68, 32'h00000000} /* (31, 7, 0) {real, imag} */,
  {32'h3f2e86e3, 32'h3be283c0} /* (31, 6, 31) {real, imag} */,
  {32'hbe5185b1, 32'h3e9efc87} /* (31, 6, 30) {real, imag} */,
  {32'hbca72718, 32'hbc17c1e9} /* (31, 6, 29) {real, imag} */,
  {32'h3d9a43f9, 32'hbe1d38e0} /* (31, 6, 28) {real, imag} */,
  {32'hba10f6a0, 32'h3d49fbf2} /* (31, 6, 27) {real, imag} */,
  {32'h3a253370, 32'h3d0156ab} /* (31, 6, 26) {real, imag} */,
  {32'hbc8761f7, 32'h3d2f7a3d} /* (31, 6, 25) {real, imag} */,
  {32'hbc9aaec6, 32'hbd71de9b} /* (31, 6, 24) {real, imag} */,
  {32'h3cc3aa06, 32'h3cf06ccd} /* (31, 6, 23) {real, imag} */,
  {32'h3d534466, 32'hbdca02e2} /* (31, 6, 22) {real, imag} */,
  {32'hbd981455, 32'h3da2ab4d} /* (31, 6, 21) {real, imag} */,
  {32'hbccb9d2c, 32'h3ba1796c} /* (31, 6, 20) {real, imag} */,
  {32'hbd4af628, 32'hbd1758e3} /* (31, 6, 19) {real, imag} */,
  {32'hbd52300c, 32'h3d333400} /* (31, 6, 18) {real, imag} */,
  {32'hbd805340, 32'h3b4395ec} /* (31, 6, 17) {real, imag} */,
  {32'hbb4877d4, 32'h00000000} /* (31, 6, 16) {real, imag} */,
  {32'hbd805340, 32'hbb4395ec} /* (31, 6, 15) {real, imag} */,
  {32'hbd52300c, 32'hbd333400} /* (31, 6, 14) {real, imag} */,
  {32'hbd4af628, 32'h3d1758e3} /* (31, 6, 13) {real, imag} */,
  {32'hbccb9d2c, 32'hbba1796c} /* (31, 6, 12) {real, imag} */,
  {32'hbd981455, 32'hbda2ab4d} /* (31, 6, 11) {real, imag} */,
  {32'h3d534466, 32'h3dca02e2} /* (31, 6, 10) {real, imag} */,
  {32'h3cc3aa06, 32'hbcf06ccd} /* (31, 6, 9) {real, imag} */,
  {32'hbc9aaec6, 32'h3d71de9b} /* (31, 6, 8) {real, imag} */,
  {32'hbc8761f7, 32'hbd2f7a3d} /* (31, 6, 7) {real, imag} */,
  {32'h3a253370, 32'hbd0156ab} /* (31, 6, 6) {real, imag} */,
  {32'hba10f6a0, 32'hbd49fbf2} /* (31, 6, 5) {real, imag} */,
  {32'h3d9a43f9, 32'h3e1d38e0} /* (31, 6, 4) {real, imag} */,
  {32'hbca72718, 32'h3c17c1e9} /* (31, 6, 3) {real, imag} */,
  {32'hbe5185b1, 32'hbe9efc87} /* (31, 6, 2) {real, imag} */,
  {32'h3f2e86e3, 32'hbbe283c0} /* (31, 6, 1) {real, imag} */,
  {32'h3e547bab, 32'h00000000} /* (31, 6, 0) {real, imag} */,
  {32'h3f033409, 32'hbe940fde} /* (31, 5, 31) {real, imag} */,
  {32'hbd8da6e8, 32'h3ea0d2ac} /* (31, 5, 30) {real, imag} */,
  {32'hbd1e39dc, 32'hbc704bfa} /* (31, 5, 29) {real, imag} */,
  {32'hbda7b1d8, 32'hbdc2cdea} /* (31, 5, 28) {real, imag} */,
  {32'hbd580b96, 32'h3cecc8c2} /* (31, 5, 27) {real, imag} */,
  {32'hbc843058, 32'h3d5d9540} /* (31, 5, 26) {real, imag} */,
  {32'hbb693a98, 32'h3d0438ec} /* (31, 5, 25) {real, imag} */,
  {32'h3cd51b0b, 32'hbd544fa6} /* (31, 5, 24) {real, imag} */,
  {32'h3d4f54b4, 32'h3ccded5b} /* (31, 5, 23) {real, imag} */,
  {32'h3d03cb56, 32'hbd3e0972} /* (31, 5, 22) {real, imag} */,
  {32'h3bbbb8c4, 32'h3d071d18} /* (31, 5, 21) {real, imag} */,
  {32'hbdc8a0b0, 32'hbd367158} /* (31, 5, 20) {real, imag} */,
  {32'hbe11f55c, 32'hbc08ee46} /* (31, 5, 19) {real, imag} */,
  {32'hbd6f1f65, 32'h3d03678c} /* (31, 5, 18) {real, imag} */,
  {32'hbc575e90, 32'hbb53ddc8} /* (31, 5, 17) {real, imag} */,
  {32'h39c81140, 32'h00000000} /* (31, 5, 16) {real, imag} */,
  {32'hbc575e90, 32'h3b53ddc8} /* (31, 5, 15) {real, imag} */,
  {32'hbd6f1f65, 32'hbd03678c} /* (31, 5, 14) {real, imag} */,
  {32'hbe11f55c, 32'h3c08ee46} /* (31, 5, 13) {real, imag} */,
  {32'hbdc8a0b0, 32'h3d367158} /* (31, 5, 12) {real, imag} */,
  {32'h3bbbb8c4, 32'hbd071d18} /* (31, 5, 11) {real, imag} */,
  {32'h3d03cb56, 32'h3d3e0972} /* (31, 5, 10) {real, imag} */,
  {32'h3d4f54b4, 32'hbccded5b} /* (31, 5, 9) {real, imag} */,
  {32'h3cd51b0b, 32'h3d544fa6} /* (31, 5, 8) {real, imag} */,
  {32'hbb693a98, 32'hbd0438ec} /* (31, 5, 7) {real, imag} */,
  {32'hbc843058, 32'hbd5d9540} /* (31, 5, 6) {real, imag} */,
  {32'hbd580b96, 32'hbcecc8c2} /* (31, 5, 5) {real, imag} */,
  {32'hbda7b1d8, 32'h3dc2cdea} /* (31, 5, 4) {real, imag} */,
  {32'hbd1e39dc, 32'h3c704bfa} /* (31, 5, 3) {real, imag} */,
  {32'hbd8da6e8, 32'hbea0d2ac} /* (31, 5, 2) {real, imag} */,
  {32'h3f033409, 32'h3e940fde} /* (31, 5, 1) {real, imag} */,
  {32'h3e33b76b, 32'h00000000} /* (31, 5, 0) {real, imag} */,
  {32'h3eb779fe, 32'hbebad384} /* (31, 4, 31) {real, imag} */,
  {32'h3d853443, 32'h3eb082e0} /* (31, 4, 30) {real, imag} */,
  {32'hbd8091c8, 32'h3c5d027f} /* (31, 4, 29) {real, imag} */,
  {32'hbd143cb6, 32'h3d4f4477} /* (31, 4, 28) {real, imag} */,
  {32'h3d3ee722, 32'h3dab729c} /* (31, 4, 27) {real, imag} */,
  {32'h3c0206fc, 32'h3d04cfab} /* (31, 4, 26) {real, imag} */,
  {32'h3d8ccf44, 32'hbdb12a30} /* (31, 4, 25) {real, imag} */,
  {32'h3d812788, 32'h3d6e7827} /* (31, 4, 24) {real, imag} */,
  {32'hbd2a4363, 32'h3ca34481} /* (31, 4, 23) {real, imag} */,
  {32'hbc34a8b6, 32'hbc18d6f5} /* (31, 4, 22) {real, imag} */,
  {32'hbcfd9a5a, 32'hbcf3da20} /* (31, 4, 21) {real, imag} */,
  {32'hbce60da6, 32'hbb23e6b0} /* (31, 4, 20) {real, imag} */,
  {32'h3cca41b0, 32'hbd236add} /* (31, 4, 19) {real, imag} */,
  {32'hbb1d0b28, 32'h3d660c27} /* (31, 4, 18) {real, imag} */,
  {32'h3be1ced0, 32'h3c93c1ec} /* (31, 4, 17) {real, imag} */,
  {32'h3cea2393, 32'h00000000} /* (31, 4, 16) {real, imag} */,
  {32'h3be1ced0, 32'hbc93c1ec} /* (31, 4, 15) {real, imag} */,
  {32'hbb1d0b28, 32'hbd660c27} /* (31, 4, 14) {real, imag} */,
  {32'h3cca41b0, 32'h3d236add} /* (31, 4, 13) {real, imag} */,
  {32'hbce60da6, 32'h3b23e6b0} /* (31, 4, 12) {real, imag} */,
  {32'hbcfd9a5a, 32'h3cf3da20} /* (31, 4, 11) {real, imag} */,
  {32'hbc34a8b6, 32'h3c18d6f5} /* (31, 4, 10) {real, imag} */,
  {32'hbd2a4363, 32'hbca34481} /* (31, 4, 9) {real, imag} */,
  {32'h3d812788, 32'hbd6e7827} /* (31, 4, 8) {real, imag} */,
  {32'h3d8ccf44, 32'h3db12a30} /* (31, 4, 7) {real, imag} */,
  {32'h3c0206fc, 32'hbd04cfab} /* (31, 4, 6) {real, imag} */,
  {32'h3d3ee722, 32'hbdab729c} /* (31, 4, 5) {real, imag} */,
  {32'hbd143cb6, 32'hbd4f4477} /* (31, 4, 4) {real, imag} */,
  {32'hbd8091c8, 32'hbc5d027f} /* (31, 4, 3) {real, imag} */,
  {32'h3d853443, 32'hbeb082e0} /* (31, 4, 2) {real, imag} */,
  {32'h3eb779fe, 32'h3ebad384} /* (31, 4, 1) {real, imag} */,
  {32'h3c7f47a0, 32'h00000000} /* (31, 4, 0) {real, imag} */,
  {32'h3eb86f93, 32'hbf10bf40} /* (31, 3, 31) {real, imag} */,
  {32'h3d58eec0, 32'h3ea6e63d} /* (31, 3, 30) {real, imag} */,
  {32'hbc2d9784, 32'h3c9043ed} /* (31, 3, 29) {real, imag} */,
  {32'h3ca6af94, 32'h3d8d7cb2} /* (31, 3, 28) {real, imag} */,
  {32'hbc587db8, 32'h3d2bd870} /* (31, 3, 27) {real, imag} */,
  {32'hbd832888, 32'h3d467a26} /* (31, 3, 26) {real, imag} */,
  {32'hbd28b3f7, 32'hbd111e32} /* (31, 3, 25) {real, imag} */,
  {32'h3d440acc, 32'hbc71269c} /* (31, 3, 24) {real, imag} */,
  {32'hbd2c224a, 32'h3d77678c} /* (31, 3, 23) {real, imag} */,
  {32'hbca4ebc0, 32'hbc7fdaa2} /* (31, 3, 22) {real, imag} */,
  {32'h3b9c6678, 32'h3c88fc1f} /* (31, 3, 21) {real, imag} */,
  {32'hbd73a3f7, 32'h3d9a8422} /* (31, 3, 20) {real, imag} */,
  {32'hbd8b69fd, 32'hbbfc98b0} /* (31, 3, 19) {real, imag} */,
  {32'hbbb0ce3c, 32'hbc0e9cba} /* (31, 3, 18) {real, imag} */,
  {32'h3d04c3ae, 32'h3cfa3e64} /* (31, 3, 17) {real, imag} */,
  {32'hbcd9016e, 32'h00000000} /* (31, 3, 16) {real, imag} */,
  {32'h3d04c3ae, 32'hbcfa3e64} /* (31, 3, 15) {real, imag} */,
  {32'hbbb0ce3c, 32'h3c0e9cba} /* (31, 3, 14) {real, imag} */,
  {32'hbd8b69fd, 32'h3bfc98b0} /* (31, 3, 13) {real, imag} */,
  {32'hbd73a3f7, 32'hbd9a8422} /* (31, 3, 12) {real, imag} */,
  {32'h3b9c6678, 32'hbc88fc1f} /* (31, 3, 11) {real, imag} */,
  {32'hbca4ebc0, 32'h3c7fdaa2} /* (31, 3, 10) {real, imag} */,
  {32'hbd2c224a, 32'hbd77678c} /* (31, 3, 9) {real, imag} */,
  {32'h3d440acc, 32'h3c71269c} /* (31, 3, 8) {real, imag} */,
  {32'hbd28b3f7, 32'h3d111e32} /* (31, 3, 7) {real, imag} */,
  {32'hbd832888, 32'hbd467a26} /* (31, 3, 6) {real, imag} */,
  {32'hbc587db8, 32'hbd2bd870} /* (31, 3, 5) {real, imag} */,
  {32'h3ca6af94, 32'hbd8d7cb2} /* (31, 3, 4) {real, imag} */,
  {32'hbc2d9784, 32'hbc9043ed} /* (31, 3, 3) {real, imag} */,
  {32'h3d58eec0, 32'hbea6e63d} /* (31, 3, 2) {real, imag} */,
  {32'h3eb86f93, 32'h3f10bf40} /* (31, 3, 1) {real, imag} */,
  {32'h3cd2c748, 32'h00000000} /* (31, 3, 0) {real, imag} */,
  {32'h3e976384, 32'hbf0ceb74} /* (31, 2, 31) {real, imag} */,
  {32'h3d5aa314, 32'h3e644774} /* (31, 2, 30) {real, imag} */,
  {32'h3d3a3c74, 32'h3bb0d650} /* (31, 2, 29) {real, imag} */,
  {32'hbda5a013, 32'h3dce1b3c} /* (31, 2, 28) {real, imag} */,
  {32'hbd74df5d, 32'h3d303bba} /* (31, 2, 27) {real, imag} */,
  {32'hbd5aff7a, 32'hbd83f549} /* (31, 2, 26) {real, imag} */,
  {32'hbc939c06, 32'hbd9939d2} /* (31, 2, 25) {real, imag} */,
  {32'h39da6200, 32'hbc3f9d3d} /* (31, 2, 24) {real, imag} */,
  {32'hbd0279fd, 32'hba7d1140} /* (31, 2, 23) {real, imag} */,
  {32'h3c47c3f0, 32'h3d9b7d8b} /* (31, 2, 22) {real, imag} */,
  {32'h3c44f1e2, 32'hbcc9a0b2} /* (31, 2, 21) {real, imag} */,
  {32'h3da646fe, 32'h3c8c48ea} /* (31, 2, 20) {real, imag} */,
  {32'h3c7a2702, 32'hbc2262ac} /* (31, 2, 19) {real, imag} */,
  {32'h3c3c0e34, 32'h3b286990} /* (31, 2, 18) {real, imag} */,
  {32'hbd5c94fa, 32'hbc629b26} /* (31, 2, 17) {real, imag} */,
  {32'h3c969ebe, 32'h00000000} /* (31, 2, 16) {real, imag} */,
  {32'hbd5c94fa, 32'h3c629b26} /* (31, 2, 15) {real, imag} */,
  {32'h3c3c0e34, 32'hbb286990} /* (31, 2, 14) {real, imag} */,
  {32'h3c7a2702, 32'h3c2262ac} /* (31, 2, 13) {real, imag} */,
  {32'h3da646fe, 32'hbc8c48ea} /* (31, 2, 12) {real, imag} */,
  {32'h3c44f1e2, 32'h3cc9a0b2} /* (31, 2, 11) {real, imag} */,
  {32'h3c47c3f0, 32'hbd9b7d8b} /* (31, 2, 10) {real, imag} */,
  {32'hbd0279fd, 32'h3a7d1140} /* (31, 2, 9) {real, imag} */,
  {32'h39da6200, 32'h3c3f9d3d} /* (31, 2, 8) {real, imag} */,
  {32'hbc939c06, 32'h3d9939d2} /* (31, 2, 7) {real, imag} */,
  {32'hbd5aff7a, 32'h3d83f549} /* (31, 2, 6) {real, imag} */,
  {32'hbd74df5d, 32'hbd303bba} /* (31, 2, 5) {real, imag} */,
  {32'hbda5a013, 32'hbdce1b3c} /* (31, 2, 4) {real, imag} */,
  {32'h3d3a3c74, 32'hbbb0d650} /* (31, 2, 3) {real, imag} */,
  {32'h3d5aa314, 32'hbe644774} /* (31, 2, 2) {real, imag} */,
  {32'h3e976384, 32'h3f0ceb74} /* (31, 2, 1) {real, imag} */,
  {32'hbd8c2bbc, 32'h00000000} /* (31, 2, 0) {real, imag} */,
  {32'h3e43ede6, 32'hbefdeb9c} /* (31, 1, 31) {real, imag} */,
  {32'hbcbd7c78, 32'h3e4083a6} /* (31, 1, 30) {real, imag} */,
  {32'hbc18b13e, 32'h3dd2f07a} /* (31, 1, 29) {real, imag} */,
  {32'hbd9cd22a, 32'h3d2c0aff} /* (31, 1, 28) {real, imag} */,
  {32'h3c3d355c, 32'hbc37e025} /* (31, 1, 27) {real, imag} */,
  {32'hbd8049b3, 32'hba09cde0} /* (31, 1, 26) {real, imag} */,
  {32'hbade7520, 32'hbd9488d0} /* (31, 1, 25) {real, imag} */,
  {32'h3d8c3575, 32'h3bde2b80} /* (31, 1, 24) {real, imag} */,
  {32'hbd8ae470, 32'hbd163c86} /* (31, 1, 23) {real, imag} */,
  {32'hbd9032a7, 32'h3b9dc2f6} /* (31, 1, 22) {real, imag} */,
  {32'hbd39d714, 32'h3c9caa4e} /* (31, 1, 21) {real, imag} */,
  {32'h3d41d148, 32'hbc363e36} /* (31, 1, 20) {real, imag} */,
  {32'h3d27035e, 32'h3b035abc} /* (31, 1, 19) {real, imag} */,
  {32'h3c244143, 32'hbc0dc19d} /* (31, 1, 18) {real, imag} */,
  {32'h3c75773e, 32'h3d93f625} /* (31, 1, 17) {real, imag} */,
  {32'hbcae9903, 32'h00000000} /* (31, 1, 16) {real, imag} */,
  {32'h3c75773e, 32'hbd93f625} /* (31, 1, 15) {real, imag} */,
  {32'h3c244143, 32'h3c0dc19d} /* (31, 1, 14) {real, imag} */,
  {32'h3d27035e, 32'hbb035abc} /* (31, 1, 13) {real, imag} */,
  {32'h3d41d148, 32'h3c363e36} /* (31, 1, 12) {real, imag} */,
  {32'hbd39d714, 32'hbc9caa4e} /* (31, 1, 11) {real, imag} */,
  {32'hbd9032a7, 32'hbb9dc2f6} /* (31, 1, 10) {real, imag} */,
  {32'hbd8ae470, 32'h3d163c86} /* (31, 1, 9) {real, imag} */,
  {32'h3d8c3575, 32'hbbde2b80} /* (31, 1, 8) {real, imag} */,
  {32'hbade7520, 32'h3d9488d0} /* (31, 1, 7) {real, imag} */,
  {32'hbd8049b3, 32'h3a09cde0} /* (31, 1, 6) {real, imag} */,
  {32'h3c3d355c, 32'h3c37e025} /* (31, 1, 5) {real, imag} */,
  {32'hbd9cd22a, 32'hbd2c0aff} /* (31, 1, 4) {real, imag} */,
  {32'hbc18b13e, 32'hbdd2f07a} /* (31, 1, 3) {real, imag} */,
  {32'hbcbd7c78, 32'hbe4083a6} /* (31, 1, 2) {real, imag} */,
  {32'h3e43ede6, 32'h3efdeb9c} /* (31, 1, 1) {real, imag} */,
  {32'h3ce35728, 32'h00000000} /* (31, 1, 0) {real, imag} */,
  {32'h3e3dd736, 32'hbeb2f0e7} /* (31, 0, 31) {real, imag} */,
  {32'hbe0d5d50, 32'h3e740a7f} /* (31, 0, 30) {real, imag} */,
  {32'h3cd25d5e, 32'h3c656708} /* (31, 0, 29) {real, imag} */,
  {32'hbb745fc0, 32'h3ce884d8} /* (31, 0, 28) {real, imag} */,
  {32'h3b7caa70, 32'hbd4384ae} /* (31, 0, 27) {real, imag} */,
  {32'h3c110580, 32'h3c328b12} /* (31, 0, 26) {real, imag} */,
  {32'hbcc226a0, 32'hbce6f212} /* (31, 0, 25) {real, imag} */,
  {32'h3ccef778, 32'hb9c45180} /* (31, 0, 24) {real, imag} */,
  {32'hbcabcd3d, 32'h3cfc0f38} /* (31, 0, 23) {real, imag} */,
  {32'h3cc1d12a, 32'hbc52b8e6} /* (31, 0, 22) {real, imag} */,
  {32'hbbb17a90, 32'hbc98b946} /* (31, 0, 21) {real, imag} */,
  {32'hbcc1e548, 32'h3d11d5c3} /* (31, 0, 20) {real, imag} */,
  {32'hbd34dfe5, 32'hbcdf0776} /* (31, 0, 19) {real, imag} */,
  {32'h3cc255f6, 32'hbce8c622} /* (31, 0, 18) {real, imag} */,
  {32'h3c423924, 32'h3b22b2f4} /* (31, 0, 17) {real, imag} */,
  {32'hbce6bf08, 32'h00000000} /* (31, 0, 16) {real, imag} */,
  {32'h3c423924, 32'hbb22b2f4} /* (31, 0, 15) {real, imag} */,
  {32'h3cc255f6, 32'h3ce8c622} /* (31, 0, 14) {real, imag} */,
  {32'hbd34dfe5, 32'h3cdf0776} /* (31, 0, 13) {real, imag} */,
  {32'hbcc1e548, 32'hbd11d5c3} /* (31, 0, 12) {real, imag} */,
  {32'hbbb17a90, 32'h3c98b946} /* (31, 0, 11) {real, imag} */,
  {32'h3cc1d12a, 32'h3c52b8e6} /* (31, 0, 10) {real, imag} */,
  {32'hbcabcd3d, 32'hbcfc0f38} /* (31, 0, 9) {real, imag} */,
  {32'h3ccef778, 32'h39c45180} /* (31, 0, 8) {real, imag} */,
  {32'hbcc226a0, 32'h3ce6f212} /* (31, 0, 7) {real, imag} */,
  {32'h3c110580, 32'hbc328b12} /* (31, 0, 6) {real, imag} */,
  {32'h3b7caa70, 32'h3d4384ae} /* (31, 0, 5) {real, imag} */,
  {32'hbb745fc0, 32'hbce884d8} /* (31, 0, 4) {real, imag} */,
  {32'h3cd25d5e, 32'hbc656708} /* (31, 0, 3) {real, imag} */,
  {32'hbe0d5d50, 32'hbe740a7f} /* (31, 0, 2) {real, imag} */,
  {32'h3e3dd736, 32'h3eb2f0e7} /* (31, 0, 1) {real, imag} */,
  {32'h3d0bf0bc, 32'h00000000} /* (31, 0, 0) {real, imag} */,
  {32'h3f5624b8, 32'hbf0cac78} /* (30, 31, 31) {real, imag} */,
  {32'hbec0a9ae, 32'h3ed10372} /* (30, 31, 30) {real, imag} */,
  {32'hbcf5ab1c, 32'hbcfa3e90} /* (30, 31, 29) {real, imag} */,
  {32'h3dd4afe9, 32'h3d7de6f2} /* (30, 31, 28) {real, imag} */,
  {32'hbd994eff, 32'h3cdaa400} /* (30, 31, 27) {real, imag} */,
  {32'hbd4dab27, 32'hbd2f5398} /* (30, 31, 26) {real, imag} */,
  {32'hbc6f07bc, 32'h3d20410e} /* (30, 31, 25) {real, imag} */,
  {32'hbbf9e95c, 32'h3dcf2593} /* (30, 31, 24) {real, imag} */,
  {32'h3d9f4969, 32'h3c26b794} /* (30, 31, 23) {real, imag} */,
  {32'hbd3fed74, 32'hbd90c04b} /* (30, 31, 22) {real, imag} */,
  {32'hbbd36408, 32'h3c0e1ddc} /* (30, 31, 21) {real, imag} */,
  {32'hbbc19da9, 32'h3c101b4e} /* (30, 31, 20) {real, imag} */,
  {32'h3d32acb4, 32'h3bc75390} /* (30, 31, 19) {real, imag} */,
  {32'h3bdd3f42, 32'hbc930e86} /* (30, 31, 18) {real, imag} */,
  {32'hbbc4bd6c, 32'hbd957000} /* (30, 31, 17) {real, imag} */,
  {32'hbd2df4c2, 32'h00000000} /* (30, 31, 16) {real, imag} */,
  {32'hbbc4bd6c, 32'h3d957000} /* (30, 31, 15) {real, imag} */,
  {32'h3bdd3f42, 32'h3c930e86} /* (30, 31, 14) {real, imag} */,
  {32'h3d32acb4, 32'hbbc75390} /* (30, 31, 13) {real, imag} */,
  {32'hbbc19da9, 32'hbc101b4e} /* (30, 31, 12) {real, imag} */,
  {32'hbbd36408, 32'hbc0e1ddc} /* (30, 31, 11) {real, imag} */,
  {32'hbd3fed74, 32'h3d90c04b} /* (30, 31, 10) {real, imag} */,
  {32'h3d9f4969, 32'hbc26b794} /* (30, 31, 9) {real, imag} */,
  {32'hbbf9e95c, 32'hbdcf2593} /* (30, 31, 8) {real, imag} */,
  {32'hbc6f07bc, 32'hbd20410e} /* (30, 31, 7) {real, imag} */,
  {32'hbd4dab27, 32'h3d2f5398} /* (30, 31, 6) {real, imag} */,
  {32'hbd994eff, 32'hbcdaa400} /* (30, 31, 5) {real, imag} */,
  {32'h3dd4afe9, 32'hbd7de6f2} /* (30, 31, 4) {real, imag} */,
  {32'hbcf5ab1c, 32'h3cfa3e90} /* (30, 31, 3) {real, imag} */,
  {32'hbec0a9ae, 32'hbed10372} /* (30, 31, 2) {real, imag} */,
  {32'h3f5624b8, 32'h3f0cac78} /* (30, 31, 1) {real, imag} */,
  {32'h3ed265ae, 32'h00000000} /* (30, 31, 0) {real, imag} */,
  {32'h3fa64438, 32'hbf0eff1e} /* (30, 30, 31) {real, imag} */,
  {32'hbf314c4e, 32'h3f060756} /* (30, 30, 30) {real, imag} */,
  {32'h3ce543ea, 32'hbd663d78} /* (30, 30, 29) {real, imag} */,
  {32'h3e695a64, 32'h3db09ae0} /* (30, 30, 28) {real, imag} */,
  {32'hbe40ded8, 32'h3cb12f50} /* (30, 30, 27) {real, imag} */,
  {32'h3d8fe00c, 32'hbe1cced5} /* (30, 30, 26) {real, imag} */,
  {32'hbd0bedfa, 32'h3d8aa031} /* (30, 30, 25) {real, imag} */,
  {32'h3d222345, 32'h3db9f86c} /* (30, 30, 24) {real, imag} */,
  {32'h3d82747a, 32'h3d9d3a4c} /* (30, 30, 23) {real, imag} */,
  {32'hbd1319a8, 32'h3d361605} /* (30, 30, 22) {real, imag} */,
  {32'h3d001fc9, 32'h3d51cc5a} /* (30, 30, 21) {real, imag} */,
  {32'h3b8dd968, 32'h3d26b26e} /* (30, 30, 20) {real, imag} */,
  {32'hbd588896, 32'h3c1dfcb6} /* (30, 30, 19) {real, imag} */,
  {32'h3c4d23c8, 32'h3d08e225} /* (30, 30, 18) {real, imag} */,
  {32'hbb1186d8, 32'hbd6ca192} /* (30, 30, 17) {real, imag} */,
  {32'hbc2c6958, 32'h00000000} /* (30, 30, 16) {real, imag} */,
  {32'hbb1186d8, 32'h3d6ca192} /* (30, 30, 15) {real, imag} */,
  {32'h3c4d23c8, 32'hbd08e225} /* (30, 30, 14) {real, imag} */,
  {32'hbd588896, 32'hbc1dfcb6} /* (30, 30, 13) {real, imag} */,
  {32'h3b8dd968, 32'hbd26b26e} /* (30, 30, 12) {real, imag} */,
  {32'h3d001fc9, 32'hbd51cc5a} /* (30, 30, 11) {real, imag} */,
  {32'hbd1319a8, 32'hbd361605} /* (30, 30, 10) {real, imag} */,
  {32'h3d82747a, 32'hbd9d3a4c} /* (30, 30, 9) {real, imag} */,
  {32'h3d222345, 32'hbdb9f86c} /* (30, 30, 8) {real, imag} */,
  {32'hbd0bedfa, 32'hbd8aa031} /* (30, 30, 7) {real, imag} */,
  {32'h3d8fe00c, 32'h3e1cced5} /* (30, 30, 6) {real, imag} */,
  {32'hbe40ded8, 32'hbcb12f50} /* (30, 30, 5) {real, imag} */,
  {32'h3e695a64, 32'hbdb09ae0} /* (30, 30, 4) {real, imag} */,
  {32'h3ce543ea, 32'h3d663d78} /* (30, 30, 3) {real, imag} */,
  {32'hbf314c4e, 32'hbf060756} /* (30, 30, 2) {real, imag} */,
  {32'h3fa64438, 32'h3f0eff1e} /* (30, 30, 1) {real, imag} */,
  {32'h3f41eb6e, 32'h00000000} /* (30, 30, 0) {real, imag} */,
  {32'h3fb27294, 32'hbeab1f66} /* (30, 29, 31) {real, imag} */,
  {32'hbf4a9b09, 32'h3eca0e2c} /* (30, 29, 30) {real, imag} */,
  {32'h3c043560, 32'hbcf2ac4c} /* (30, 29, 29) {real, imag} */,
  {32'h3e1015e2, 32'hbcb29fc8} /* (30, 29, 28) {real, imag} */,
  {32'hbe5d6993, 32'hbcfc72a6} /* (30, 29, 27) {real, imag} */,
  {32'hbe01668f, 32'hbcc06f08} /* (30, 29, 26) {real, imag} */,
  {32'h3d829348, 32'hbd00b666} /* (30, 29, 25) {real, imag} */,
  {32'hbcd04004, 32'h3d892f58} /* (30, 29, 24) {real, imag} */,
  {32'h3caa0c06, 32'h3d26195c} /* (30, 29, 23) {real, imag} */,
  {32'hbcbad18d, 32'hbdae23e9} /* (30, 29, 22) {real, imag} */,
  {32'h3d756f21, 32'h3d69e3c2} /* (30, 29, 21) {real, imag} */,
  {32'h3d5a035c, 32'h3d648ca7} /* (30, 29, 20) {real, imag} */,
  {32'h3d8cc015, 32'h3b76adb0} /* (30, 29, 19) {real, imag} */,
  {32'hbbfdee6c, 32'h3d1578da} /* (30, 29, 18) {real, imag} */,
  {32'h3c8fdc81, 32'h3d698c0a} /* (30, 29, 17) {real, imag} */,
  {32'hbda9610a, 32'h00000000} /* (30, 29, 16) {real, imag} */,
  {32'h3c8fdc81, 32'hbd698c0a} /* (30, 29, 15) {real, imag} */,
  {32'hbbfdee6c, 32'hbd1578da} /* (30, 29, 14) {real, imag} */,
  {32'h3d8cc015, 32'hbb76adb0} /* (30, 29, 13) {real, imag} */,
  {32'h3d5a035c, 32'hbd648ca7} /* (30, 29, 12) {real, imag} */,
  {32'h3d756f21, 32'hbd69e3c2} /* (30, 29, 11) {real, imag} */,
  {32'hbcbad18d, 32'h3dae23e9} /* (30, 29, 10) {real, imag} */,
  {32'h3caa0c06, 32'hbd26195c} /* (30, 29, 9) {real, imag} */,
  {32'hbcd04004, 32'hbd892f58} /* (30, 29, 8) {real, imag} */,
  {32'h3d829348, 32'h3d00b666} /* (30, 29, 7) {real, imag} */,
  {32'hbe01668f, 32'h3cc06f08} /* (30, 29, 6) {real, imag} */,
  {32'hbe5d6993, 32'h3cfc72a6} /* (30, 29, 5) {real, imag} */,
  {32'h3e1015e2, 32'h3cb29fc8} /* (30, 29, 4) {real, imag} */,
  {32'h3c043560, 32'h3cf2ac4c} /* (30, 29, 3) {real, imag} */,
  {32'hbf4a9b09, 32'hbeca0e2c} /* (30, 29, 2) {real, imag} */,
  {32'h3fb27294, 32'h3eab1f66} /* (30, 29, 1) {real, imag} */,
  {32'h3f1dc60c, 32'h00000000} /* (30, 29, 0) {real, imag} */,
  {32'h3fb89d90, 32'hbe363c34} /* (30, 28, 31) {real, imag} */,
  {32'hbf4d50fb, 32'h3dbc00ac} /* (30, 28, 30) {real, imag} */,
  {32'hbe0bbb30, 32'hbda19154} /* (30, 28, 29) {real, imag} */,
  {32'h3e228b48, 32'hbd04b56a} /* (30, 28, 28) {real, imag} */,
  {32'hbe314d84, 32'hbcf79cc8} /* (30, 28, 27) {real, imag} */,
  {32'hbd71209a, 32'hbb63e038} /* (30, 28, 26) {real, imag} */,
  {32'hbe002bce, 32'hbd1162ba} /* (30, 28, 25) {real, imag} */,
  {32'hbd941b51, 32'h3dc36309} /* (30, 28, 24) {real, imag} */,
  {32'hbb603cac, 32'h3de5bfa6} /* (30, 28, 23) {real, imag} */,
  {32'h3d4149d1, 32'hbc216a77} /* (30, 28, 22) {real, imag} */,
  {32'h3dc5a306, 32'h3da23fb8} /* (30, 28, 21) {real, imag} */,
  {32'h3d92e1a8, 32'hbcbca943} /* (30, 28, 20) {real, imag} */,
  {32'h3d0d89a4, 32'h3c81b992} /* (30, 28, 19) {real, imag} */,
  {32'hbd8651f7, 32'hbc430ebc} /* (30, 28, 18) {real, imag} */,
  {32'h398a7500, 32'hbd8b06ac} /* (30, 28, 17) {real, imag} */,
  {32'h3d674c33, 32'h00000000} /* (30, 28, 16) {real, imag} */,
  {32'h398a7500, 32'h3d8b06ac} /* (30, 28, 15) {real, imag} */,
  {32'hbd8651f7, 32'h3c430ebc} /* (30, 28, 14) {real, imag} */,
  {32'h3d0d89a4, 32'hbc81b992} /* (30, 28, 13) {real, imag} */,
  {32'h3d92e1a8, 32'h3cbca943} /* (30, 28, 12) {real, imag} */,
  {32'h3dc5a306, 32'hbda23fb8} /* (30, 28, 11) {real, imag} */,
  {32'h3d4149d1, 32'h3c216a77} /* (30, 28, 10) {real, imag} */,
  {32'hbb603cac, 32'hbde5bfa6} /* (30, 28, 9) {real, imag} */,
  {32'hbd941b51, 32'hbdc36309} /* (30, 28, 8) {real, imag} */,
  {32'hbe002bce, 32'h3d1162ba} /* (30, 28, 7) {real, imag} */,
  {32'hbd71209a, 32'h3b63e038} /* (30, 28, 6) {real, imag} */,
  {32'hbe314d84, 32'h3cf79cc8} /* (30, 28, 5) {real, imag} */,
  {32'h3e228b48, 32'h3d04b56a} /* (30, 28, 4) {real, imag} */,
  {32'hbe0bbb30, 32'h3da19154} /* (30, 28, 3) {real, imag} */,
  {32'hbf4d50fb, 32'hbdbc00ac} /* (30, 28, 2) {real, imag} */,
  {32'h3fb89d90, 32'h3e363c34} /* (30, 28, 1) {real, imag} */,
  {32'h3f419a58, 32'h00000000} /* (30, 28, 0) {real, imag} */,
  {32'h3fb39a36, 32'hbde1cfb0} /* (30, 27, 31) {real, imag} */,
  {32'hbf746f7c, 32'h3e439905} /* (30, 27, 30) {real, imag} */,
  {32'hbc5faad4, 32'hbe408951} /* (30, 27, 29) {real, imag} */,
  {32'h3e1c5eb6, 32'h3dbfdb68} /* (30, 27, 28) {real, imag} */,
  {32'hbde7ba5e, 32'h3d733baa} /* (30, 27, 27) {real, imag} */,
  {32'h3d738a19, 32'hbe08b7ea} /* (30, 27, 26) {real, imag} */,
  {32'hbddde7a1, 32'hbe02871d} /* (30, 27, 25) {real, imag} */,
  {32'hbd1ad470, 32'h3d488a38} /* (30, 27, 24) {real, imag} */,
  {32'hbd82918e, 32'h3d921f76} /* (30, 27, 23) {real, imag} */,
  {32'h3d384c1e, 32'hbc0a4534} /* (30, 27, 22) {real, imag} */,
  {32'h3d4941a0, 32'h3d7a384d} /* (30, 27, 21) {real, imag} */,
  {32'hbddf6850, 32'hbd4f1772} /* (30, 27, 20) {real, imag} */,
  {32'hbd00e04a, 32'hbe036b8c} /* (30, 27, 19) {real, imag} */,
  {32'hbbd3e6f5, 32'h3d9e8bd0} /* (30, 27, 18) {real, imag} */,
  {32'hbcf13533, 32'hbd02d879} /* (30, 27, 17) {real, imag} */,
  {32'h3cb7ac4e, 32'h00000000} /* (30, 27, 16) {real, imag} */,
  {32'hbcf13533, 32'h3d02d879} /* (30, 27, 15) {real, imag} */,
  {32'hbbd3e6f5, 32'hbd9e8bd0} /* (30, 27, 14) {real, imag} */,
  {32'hbd00e04a, 32'h3e036b8c} /* (30, 27, 13) {real, imag} */,
  {32'hbddf6850, 32'h3d4f1772} /* (30, 27, 12) {real, imag} */,
  {32'h3d4941a0, 32'hbd7a384d} /* (30, 27, 11) {real, imag} */,
  {32'h3d384c1e, 32'h3c0a4534} /* (30, 27, 10) {real, imag} */,
  {32'hbd82918e, 32'hbd921f76} /* (30, 27, 9) {real, imag} */,
  {32'hbd1ad470, 32'hbd488a38} /* (30, 27, 8) {real, imag} */,
  {32'hbddde7a1, 32'h3e02871d} /* (30, 27, 7) {real, imag} */,
  {32'h3d738a19, 32'h3e08b7ea} /* (30, 27, 6) {real, imag} */,
  {32'hbde7ba5e, 32'hbd733baa} /* (30, 27, 5) {real, imag} */,
  {32'h3e1c5eb6, 32'hbdbfdb68} /* (30, 27, 4) {real, imag} */,
  {32'hbc5faad4, 32'h3e408951} /* (30, 27, 3) {real, imag} */,
  {32'hbf746f7c, 32'hbe439905} /* (30, 27, 2) {real, imag} */,
  {32'h3fb39a36, 32'h3de1cfb0} /* (30, 27, 1) {real, imag} */,
  {32'h3f761818, 32'h00000000} /* (30, 27, 0) {real, imag} */,
  {32'h3fbae5d8, 32'hbd9ac036} /* (30, 26, 31) {real, imag} */,
  {32'hbf5ece16, 32'h3eab95be} /* (30, 26, 30) {real, imag} */,
  {32'hbdbce90a, 32'hbde2032a} /* (30, 26, 29) {real, imag} */,
  {32'h3e2a57f5, 32'h3d4dae6f} /* (30, 26, 28) {real, imag} */,
  {32'hbdd5ac3a, 32'h3d7951de} /* (30, 26, 27) {real, imag} */,
  {32'hbd747ca9, 32'h3d2b8fce} /* (30, 26, 26) {real, imag} */,
  {32'hbd9bbb6c, 32'hbd889d38} /* (30, 26, 25) {real, imag} */,
  {32'hbda0ca5e, 32'h3d5b3ae5} /* (30, 26, 24) {real, imag} */,
  {32'hbb230f50, 32'hbdc3a7bd} /* (30, 26, 23) {real, imag} */,
  {32'h3c28c010, 32'hbcf55170} /* (30, 26, 22) {real, imag} */,
  {32'h3ca37152, 32'h3d4b48ba} /* (30, 26, 21) {real, imag} */,
  {32'h3db34b96, 32'h3d483664} /* (30, 26, 20) {real, imag} */,
  {32'h3c94fe73, 32'hbad495b0} /* (30, 26, 19) {real, imag} */,
  {32'h3cb2adaf, 32'hbb5490b0} /* (30, 26, 18) {real, imag} */,
  {32'hbd1b6602, 32'hbbeaac8c} /* (30, 26, 17) {real, imag} */,
  {32'hb940dd00, 32'h00000000} /* (30, 26, 16) {real, imag} */,
  {32'hbd1b6602, 32'h3beaac8c} /* (30, 26, 15) {real, imag} */,
  {32'h3cb2adaf, 32'h3b5490b0} /* (30, 26, 14) {real, imag} */,
  {32'h3c94fe73, 32'h3ad495b0} /* (30, 26, 13) {real, imag} */,
  {32'h3db34b96, 32'hbd483664} /* (30, 26, 12) {real, imag} */,
  {32'h3ca37152, 32'hbd4b48ba} /* (30, 26, 11) {real, imag} */,
  {32'h3c28c010, 32'h3cf55170} /* (30, 26, 10) {real, imag} */,
  {32'hbb230f50, 32'h3dc3a7bd} /* (30, 26, 9) {real, imag} */,
  {32'hbda0ca5e, 32'hbd5b3ae5} /* (30, 26, 8) {real, imag} */,
  {32'hbd9bbb6c, 32'h3d889d38} /* (30, 26, 7) {real, imag} */,
  {32'hbd747ca9, 32'hbd2b8fce} /* (30, 26, 6) {real, imag} */,
  {32'hbdd5ac3a, 32'hbd7951de} /* (30, 26, 5) {real, imag} */,
  {32'h3e2a57f5, 32'hbd4dae6f} /* (30, 26, 4) {real, imag} */,
  {32'hbdbce90a, 32'h3de2032a} /* (30, 26, 3) {real, imag} */,
  {32'hbf5ece16, 32'hbeab95be} /* (30, 26, 2) {real, imag} */,
  {32'h3fbae5d8, 32'h3d9ac036} /* (30, 26, 1) {real, imag} */,
  {32'h3f73b27c, 32'h00000000} /* (30, 26, 0) {real, imag} */,
  {32'h3fc5e649, 32'hbdb0a720} /* (30, 25, 31) {real, imag} */,
  {32'hbf8527fa, 32'h3e8c7e20} /* (30, 25, 30) {real, imag} */,
  {32'hbdd89c4c, 32'hbddea51a} /* (30, 25, 29) {real, imag} */,
  {32'h3d8aa9e4, 32'h3c1aec16} /* (30, 25, 28) {real, imag} */,
  {32'hbe15fb2d, 32'hbd277855} /* (30, 25, 27) {real, imag} */,
  {32'h3d48d6ac, 32'hbdabed6a} /* (30, 25, 26) {real, imag} */,
  {32'hbd3b676e, 32'hbdb7b7be} /* (30, 25, 25) {real, imag} */,
  {32'hbdb1a3e8, 32'h3cab049d} /* (30, 25, 24) {real, imag} */,
  {32'h3ab56398, 32'h3d51a807} /* (30, 25, 23) {real, imag} */,
  {32'hbda5914c, 32'hbbfda338} /* (30, 25, 22) {real, imag} */,
  {32'hbd861006, 32'h3df39d01} /* (30, 25, 21) {real, imag} */,
  {32'h3d8c88ac, 32'hbda2145b} /* (30, 25, 20) {real, imag} */,
  {32'h3d6bc3b0, 32'h3d714b68} /* (30, 25, 19) {real, imag} */,
  {32'h3cd67c1a, 32'hbc37adac} /* (30, 25, 18) {real, imag} */,
  {32'h3ce89787, 32'hbcbcc8aa} /* (30, 25, 17) {real, imag} */,
  {32'hbce9c721, 32'h00000000} /* (30, 25, 16) {real, imag} */,
  {32'h3ce89787, 32'h3cbcc8aa} /* (30, 25, 15) {real, imag} */,
  {32'h3cd67c1a, 32'h3c37adac} /* (30, 25, 14) {real, imag} */,
  {32'h3d6bc3b0, 32'hbd714b68} /* (30, 25, 13) {real, imag} */,
  {32'h3d8c88ac, 32'h3da2145b} /* (30, 25, 12) {real, imag} */,
  {32'hbd861006, 32'hbdf39d01} /* (30, 25, 11) {real, imag} */,
  {32'hbda5914c, 32'h3bfda338} /* (30, 25, 10) {real, imag} */,
  {32'h3ab56398, 32'hbd51a807} /* (30, 25, 9) {real, imag} */,
  {32'hbdb1a3e8, 32'hbcab049d} /* (30, 25, 8) {real, imag} */,
  {32'hbd3b676e, 32'h3db7b7be} /* (30, 25, 7) {real, imag} */,
  {32'h3d48d6ac, 32'h3dabed6a} /* (30, 25, 6) {real, imag} */,
  {32'hbe15fb2d, 32'h3d277855} /* (30, 25, 5) {real, imag} */,
  {32'h3d8aa9e4, 32'hbc1aec16} /* (30, 25, 4) {real, imag} */,
  {32'hbdd89c4c, 32'h3ddea51a} /* (30, 25, 3) {real, imag} */,
  {32'hbf8527fa, 32'hbe8c7e20} /* (30, 25, 2) {real, imag} */,
  {32'h3fc5e649, 32'h3db0a720} /* (30, 25, 1) {real, imag} */,
  {32'h3f618a60, 32'h00000000} /* (30, 25, 0) {real, imag} */,
  {32'h3fb710d6, 32'h3d446ea4} /* (30, 24, 31) {real, imag} */,
  {32'hbf57c692, 32'h3e985608} /* (30, 24, 30) {real, imag} */,
  {32'h3c22eaa0, 32'hbd6725aa} /* (30, 24, 29) {real, imag} */,
  {32'h3d993f12, 32'hbdd4d546} /* (30, 24, 28) {real, imag} */,
  {32'hbe4c97a6, 32'hbb392ad0} /* (30, 24, 27) {real, imag} */,
  {32'hbd9fc565, 32'h3c664f5c} /* (30, 24, 26) {real, imag} */,
  {32'hbdb61439, 32'hbdea34ec} /* (30, 24, 25) {real, imag} */,
  {32'hbe0fdbb3, 32'h3d2f3fc9} /* (30, 24, 24) {real, imag} */,
  {32'h3ca09de4, 32'h3e01fa1e} /* (30, 24, 23) {real, imag} */,
  {32'h3c882ab4, 32'hbe014db3} /* (30, 24, 22) {real, imag} */,
  {32'h3d0012ea, 32'hbcaa5da6} /* (30, 24, 21) {real, imag} */,
  {32'h3cbf88c2, 32'hbdc3be31} /* (30, 24, 20) {real, imag} */,
  {32'hbc673f44, 32'hbd1e1e57} /* (30, 24, 19) {real, imag} */,
  {32'hbcc47aac, 32'h3dd80608} /* (30, 24, 18) {real, imag} */,
  {32'h3c460b54, 32'h3d005377} /* (30, 24, 17) {real, imag} */,
  {32'hbd013bb8, 32'h00000000} /* (30, 24, 16) {real, imag} */,
  {32'h3c460b54, 32'hbd005377} /* (30, 24, 15) {real, imag} */,
  {32'hbcc47aac, 32'hbdd80608} /* (30, 24, 14) {real, imag} */,
  {32'hbc673f44, 32'h3d1e1e57} /* (30, 24, 13) {real, imag} */,
  {32'h3cbf88c2, 32'h3dc3be31} /* (30, 24, 12) {real, imag} */,
  {32'h3d0012ea, 32'h3caa5da6} /* (30, 24, 11) {real, imag} */,
  {32'h3c882ab4, 32'h3e014db3} /* (30, 24, 10) {real, imag} */,
  {32'h3ca09de4, 32'hbe01fa1e} /* (30, 24, 9) {real, imag} */,
  {32'hbe0fdbb3, 32'hbd2f3fc9} /* (30, 24, 8) {real, imag} */,
  {32'hbdb61439, 32'h3dea34ec} /* (30, 24, 7) {real, imag} */,
  {32'hbd9fc565, 32'hbc664f5c} /* (30, 24, 6) {real, imag} */,
  {32'hbe4c97a6, 32'h3b392ad0} /* (30, 24, 5) {real, imag} */,
  {32'h3d993f12, 32'h3dd4d546} /* (30, 24, 4) {real, imag} */,
  {32'h3c22eaa0, 32'h3d6725aa} /* (30, 24, 3) {real, imag} */,
  {32'hbf57c692, 32'hbe985608} /* (30, 24, 2) {real, imag} */,
  {32'h3fb710d6, 32'hbd446ea4} /* (30, 24, 1) {real, imag} */,
  {32'h3f7c3498, 32'h00000000} /* (30, 24, 0) {real, imag} */,
  {32'h3f9257fa, 32'h3d866420} /* (30, 23, 31) {real, imag} */,
  {32'hbf258a3f, 32'h3ea6be8b} /* (30, 23, 30) {real, imag} */,
  {32'h3e18d446, 32'h3d2536c8} /* (30, 23, 29) {real, imag} */,
  {32'h3dd78c41, 32'hbde43a0a} /* (30, 23, 28) {real, imag} */,
  {32'hbe1a834e, 32'h3cf91a6a} /* (30, 23, 27) {real, imag} */,
  {32'hbc98a3ef, 32'h3db598b9} /* (30, 23, 26) {real, imag} */,
  {32'hbc9a3ba0, 32'hbdd43521} /* (30, 23, 25) {real, imag} */,
  {32'h3c97a611, 32'h3d0314aa} /* (30, 23, 24) {real, imag} */,
  {32'h3a39bf50, 32'h3d92acbe} /* (30, 23, 23) {real, imag} */,
  {32'hbb9684d0, 32'hbd8507fc} /* (30, 23, 22) {real, imag} */,
  {32'h3be6fe28, 32'h3ce66186} /* (30, 23, 21) {real, imag} */,
  {32'hbd2f1a2b, 32'hbbab2040} /* (30, 23, 20) {real, imag} */,
  {32'h3d9374f0, 32'h3c83dc0b} /* (30, 23, 19) {real, imag} */,
  {32'h3d0efb21, 32'h3d65ed5c} /* (30, 23, 18) {real, imag} */,
  {32'h3d77a1ca, 32'hbcb1bf7e} /* (30, 23, 17) {real, imag} */,
  {32'h3cba36f0, 32'h00000000} /* (30, 23, 16) {real, imag} */,
  {32'h3d77a1ca, 32'h3cb1bf7e} /* (30, 23, 15) {real, imag} */,
  {32'h3d0efb21, 32'hbd65ed5c} /* (30, 23, 14) {real, imag} */,
  {32'h3d9374f0, 32'hbc83dc0b} /* (30, 23, 13) {real, imag} */,
  {32'hbd2f1a2b, 32'h3bab2040} /* (30, 23, 12) {real, imag} */,
  {32'h3be6fe28, 32'hbce66186} /* (30, 23, 11) {real, imag} */,
  {32'hbb9684d0, 32'h3d8507fc} /* (30, 23, 10) {real, imag} */,
  {32'h3a39bf50, 32'hbd92acbe} /* (30, 23, 9) {real, imag} */,
  {32'h3c97a611, 32'hbd0314aa} /* (30, 23, 8) {real, imag} */,
  {32'hbc9a3ba0, 32'h3dd43521} /* (30, 23, 7) {real, imag} */,
  {32'hbc98a3ef, 32'hbdb598b9} /* (30, 23, 6) {real, imag} */,
  {32'hbe1a834e, 32'hbcf91a6a} /* (30, 23, 5) {real, imag} */,
  {32'h3dd78c41, 32'h3de43a0a} /* (30, 23, 4) {real, imag} */,
  {32'h3e18d446, 32'hbd2536c8} /* (30, 23, 3) {real, imag} */,
  {32'hbf258a3f, 32'hbea6be8b} /* (30, 23, 2) {real, imag} */,
  {32'h3f9257fa, 32'hbd866420} /* (30, 23, 1) {real, imag} */,
  {32'h3f729179, 32'h00000000} /* (30, 23, 0) {real, imag} */,
  {32'h3f46ca20, 32'h3dc81025} /* (30, 22, 31) {real, imag} */,
  {32'hbf134e96, 32'h3eb16e46} /* (30, 22, 30) {real, imag} */,
  {32'h3e3854ce, 32'h3dc03046} /* (30, 22, 29) {real, imag} */,
  {32'hbc9b4efc, 32'hbe1104d4} /* (30, 22, 28) {real, imag} */,
  {32'hbe44ba58, 32'h3b37cdd0} /* (30, 22, 27) {real, imag} */,
  {32'hbd62e9f4, 32'h3cc61352} /* (30, 22, 26) {real, imag} */,
  {32'h3d047f7a, 32'hbd4cebb7} /* (30, 22, 25) {real, imag} */,
  {32'hbd8cd7f6, 32'h3d8c944b} /* (30, 22, 24) {real, imag} */,
  {32'h3c888ce0, 32'h3d420f1a} /* (30, 22, 23) {real, imag} */,
  {32'h3d898fbb, 32'h3d5145b8} /* (30, 22, 22) {real, imag} */,
  {32'hbd8da602, 32'h3d242264} /* (30, 22, 21) {real, imag} */,
  {32'hbd3f633e, 32'hbb1d9e00} /* (30, 22, 20) {real, imag} */,
  {32'h3d9ecb43, 32'hbd2033f7} /* (30, 22, 19) {real, imag} */,
  {32'h3d6e5540, 32'hbae4a260} /* (30, 22, 18) {real, imag} */,
  {32'hbd076580, 32'h3ae4daa0} /* (30, 22, 17) {real, imag} */,
  {32'h3d12a3d5, 32'h00000000} /* (30, 22, 16) {real, imag} */,
  {32'hbd076580, 32'hbae4daa0} /* (30, 22, 15) {real, imag} */,
  {32'h3d6e5540, 32'h3ae4a260} /* (30, 22, 14) {real, imag} */,
  {32'h3d9ecb43, 32'h3d2033f7} /* (30, 22, 13) {real, imag} */,
  {32'hbd3f633e, 32'h3b1d9e00} /* (30, 22, 12) {real, imag} */,
  {32'hbd8da602, 32'hbd242264} /* (30, 22, 11) {real, imag} */,
  {32'h3d898fbb, 32'hbd5145b8} /* (30, 22, 10) {real, imag} */,
  {32'h3c888ce0, 32'hbd420f1a} /* (30, 22, 9) {real, imag} */,
  {32'hbd8cd7f6, 32'hbd8c944b} /* (30, 22, 8) {real, imag} */,
  {32'h3d047f7a, 32'h3d4cebb7} /* (30, 22, 7) {real, imag} */,
  {32'hbd62e9f4, 32'hbcc61352} /* (30, 22, 6) {real, imag} */,
  {32'hbe44ba58, 32'hbb37cdd0} /* (30, 22, 5) {real, imag} */,
  {32'hbc9b4efc, 32'h3e1104d4} /* (30, 22, 4) {real, imag} */,
  {32'h3e3854ce, 32'hbdc03046} /* (30, 22, 3) {real, imag} */,
  {32'hbf134e96, 32'hbeb16e46} /* (30, 22, 2) {real, imag} */,
  {32'h3f46ca20, 32'hbdc81025} /* (30, 22, 1) {real, imag} */,
  {32'h3f26a97c, 32'h00000000} /* (30, 22, 0) {real, imag} */,
  {32'h3e2e56ca, 32'h3e4e35d1} /* (30, 21, 31) {real, imag} */,
  {32'hbe669951, 32'h3db00cc4} /* (30, 21, 30) {real, imag} */,
  {32'h3dd10698, 32'h3d9dff73} /* (30, 21, 29) {real, imag} */,
  {32'hbcd4b9ee, 32'h3d944c80} /* (30, 21, 28) {real, imag} */,
  {32'hbd27463c, 32'hbce2a9a5} /* (30, 21, 27) {real, imag} */,
  {32'hbd521d81, 32'hbd75c02a} /* (30, 21, 26) {real, imag} */,
  {32'h3d449380, 32'h3cad257a} /* (30, 21, 25) {real, imag} */,
  {32'hbd990c84, 32'hbc6c46e8} /* (30, 21, 24) {real, imag} */,
  {32'hbc92b018, 32'h3c7e8b2c} /* (30, 21, 23) {real, imag} */,
  {32'hb8a80f00, 32'h3d2a8ad4} /* (30, 21, 22) {real, imag} */,
  {32'h3d364742, 32'h3ceef334} /* (30, 21, 21) {real, imag} */,
  {32'hbd4b4b82, 32'h3c8fb3ef} /* (30, 21, 20) {real, imag} */,
  {32'hbdf8a22a, 32'h3b5a1a00} /* (30, 21, 19) {real, imag} */,
  {32'h3d52bee4, 32'hbd751837} /* (30, 21, 18) {real, imag} */,
  {32'h3d4a352b, 32'h3c625ae9} /* (30, 21, 17) {real, imag} */,
  {32'hbbdb2428, 32'h00000000} /* (30, 21, 16) {real, imag} */,
  {32'h3d4a352b, 32'hbc625ae9} /* (30, 21, 15) {real, imag} */,
  {32'h3d52bee4, 32'h3d751837} /* (30, 21, 14) {real, imag} */,
  {32'hbdf8a22a, 32'hbb5a1a00} /* (30, 21, 13) {real, imag} */,
  {32'hbd4b4b82, 32'hbc8fb3ef} /* (30, 21, 12) {real, imag} */,
  {32'h3d364742, 32'hbceef334} /* (30, 21, 11) {real, imag} */,
  {32'hb8a80f00, 32'hbd2a8ad4} /* (30, 21, 10) {real, imag} */,
  {32'hbc92b018, 32'hbc7e8b2c} /* (30, 21, 9) {real, imag} */,
  {32'hbd990c84, 32'h3c6c46e8} /* (30, 21, 8) {real, imag} */,
  {32'h3d449380, 32'hbcad257a} /* (30, 21, 7) {real, imag} */,
  {32'hbd521d81, 32'h3d75c02a} /* (30, 21, 6) {real, imag} */,
  {32'hbd27463c, 32'h3ce2a9a5} /* (30, 21, 5) {real, imag} */,
  {32'hbcd4b9ee, 32'hbd944c80} /* (30, 21, 4) {real, imag} */,
  {32'h3dd10698, 32'hbd9dff73} /* (30, 21, 3) {real, imag} */,
  {32'hbe669951, 32'hbdb00cc4} /* (30, 21, 2) {real, imag} */,
  {32'h3e2e56ca, 32'hbe4e35d1} /* (30, 21, 1) {real, imag} */,
  {32'h3d823e70, 32'h00000000} /* (30, 21, 0) {real, imag} */,
  {32'hbf5b8ec2, 32'h3e3d81c9} /* (30, 20, 31) {real, imag} */,
  {32'h3ee7172a, 32'hbe93b590} /* (30, 20, 30) {real, imag} */,
  {32'h3e10c410, 32'h3d7a9154} /* (30, 20, 29) {real, imag} */,
  {32'hbe1d33eb, 32'h3d5b51b6} /* (30, 20, 28) {real, imag} */,
  {32'h3da6cec2, 32'hbd02f519} /* (30, 20, 27) {real, imag} */,
  {32'h3d1ce81b, 32'hbcbfb8c3} /* (30, 20, 26) {real, imag} */,
  {32'hbcadc952, 32'hbd067b42} /* (30, 20, 25) {real, imag} */,
  {32'hbd871bb2, 32'h3da62900} /* (30, 20, 24) {real, imag} */,
  {32'hbdcb6b12, 32'hbcb125e7} /* (30, 20, 23) {real, imag} */,
  {32'h3c2627fa, 32'hbd45765c} /* (30, 20, 22) {real, imag} */,
  {32'hbd0f2124, 32'hbdc723ff} /* (30, 20, 21) {real, imag} */,
  {32'hbdf54bba, 32'hbc0f012a} /* (30, 20, 20) {real, imag} */,
  {32'h3d9d95eb, 32'h3d80f269} /* (30, 20, 19) {real, imag} */,
  {32'h3d9697aa, 32'h3c271274} /* (30, 20, 18) {real, imag} */,
  {32'h3cc79dfa, 32'hbc904c04} /* (30, 20, 17) {real, imag} */,
  {32'hbdda65de, 32'h00000000} /* (30, 20, 16) {real, imag} */,
  {32'h3cc79dfa, 32'h3c904c04} /* (30, 20, 15) {real, imag} */,
  {32'h3d9697aa, 32'hbc271274} /* (30, 20, 14) {real, imag} */,
  {32'h3d9d95eb, 32'hbd80f269} /* (30, 20, 13) {real, imag} */,
  {32'hbdf54bba, 32'h3c0f012a} /* (30, 20, 12) {real, imag} */,
  {32'hbd0f2124, 32'h3dc723ff} /* (30, 20, 11) {real, imag} */,
  {32'h3c2627fa, 32'h3d45765c} /* (30, 20, 10) {real, imag} */,
  {32'hbdcb6b12, 32'h3cb125e7} /* (30, 20, 9) {real, imag} */,
  {32'hbd871bb2, 32'hbda62900} /* (30, 20, 8) {real, imag} */,
  {32'hbcadc952, 32'h3d067b42} /* (30, 20, 7) {real, imag} */,
  {32'h3d1ce81b, 32'h3cbfb8c3} /* (30, 20, 6) {real, imag} */,
  {32'h3da6cec2, 32'h3d02f519} /* (30, 20, 5) {real, imag} */,
  {32'hbe1d33eb, 32'hbd5b51b6} /* (30, 20, 4) {real, imag} */,
  {32'h3e10c410, 32'hbd7a9154} /* (30, 20, 3) {real, imag} */,
  {32'h3ee7172a, 32'h3e93b590} /* (30, 20, 2) {real, imag} */,
  {32'hbf5b8ec2, 32'hbe3d81c9} /* (30, 20, 1) {real, imag} */,
  {32'hbf3c40d6, 32'h00000000} /* (30, 20, 0) {real, imag} */,
  {32'hbfb31b67, 32'h3df9681a} /* (30, 19, 31) {real, imag} */,
  {32'h3f2e924b, 32'hbeb1721a} /* (30, 19, 30) {real, imag} */,
  {32'h3db14b02, 32'h3df3715b} /* (30, 19, 29) {real, imag} */,
  {32'hbe842553, 32'h3d617159} /* (30, 19, 28) {real, imag} */,
  {32'h3e1746e8, 32'hbe2cd7fc} /* (30, 19, 27) {real, imag} */,
  {32'h3d70342c, 32'h3c8a834d} /* (30, 19, 26) {real, imag} */,
  {32'h3c1c50e8, 32'h3ce38c24} /* (30, 19, 25) {real, imag} */,
  {32'hbd1b1ed2, 32'hbd45e8a8} /* (30, 19, 24) {real, imag} */,
  {32'h3bf1291c, 32'h3cdb0bc9} /* (30, 19, 23) {real, imag} */,
  {32'hbd360614, 32'hbd08daf1} /* (30, 19, 22) {real, imag} */,
  {32'hbc5b34ec, 32'hbdf5ad48} /* (30, 19, 21) {real, imag} */,
  {32'h3b28a460, 32'hbdbedf88} /* (30, 19, 20) {real, imag} */,
  {32'h3dca9bc0, 32'h3d0f5f9f} /* (30, 19, 19) {real, imag} */,
  {32'hbb81a980, 32'hbd2fa3d9} /* (30, 19, 18) {real, imag} */,
  {32'hbc96d5eb, 32'h3cc034f6} /* (30, 19, 17) {real, imag} */,
  {32'hbce78ac3, 32'h00000000} /* (30, 19, 16) {real, imag} */,
  {32'hbc96d5eb, 32'hbcc034f6} /* (30, 19, 15) {real, imag} */,
  {32'hbb81a980, 32'h3d2fa3d9} /* (30, 19, 14) {real, imag} */,
  {32'h3dca9bc0, 32'hbd0f5f9f} /* (30, 19, 13) {real, imag} */,
  {32'h3b28a460, 32'h3dbedf88} /* (30, 19, 12) {real, imag} */,
  {32'hbc5b34ec, 32'h3df5ad48} /* (30, 19, 11) {real, imag} */,
  {32'hbd360614, 32'h3d08daf1} /* (30, 19, 10) {real, imag} */,
  {32'h3bf1291c, 32'hbcdb0bc9} /* (30, 19, 9) {real, imag} */,
  {32'hbd1b1ed2, 32'h3d45e8a8} /* (30, 19, 8) {real, imag} */,
  {32'h3c1c50e8, 32'hbce38c24} /* (30, 19, 7) {real, imag} */,
  {32'h3d70342c, 32'hbc8a834d} /* (30, 19, 6) {real, imag} */,
  {32'h3e1746e8, 32'h3e2cd7fc} /* (30, 19, 5) {real, imag} */,
  {32'hbe842553, 32'hbd617159} /* (30, 19, 4) {real, imag} */,
  {32'h3db14b02, 32'hbdf3715b} /* (30, 19, 3) {real, imag} */,
  {32'h3f2e924b, 32'h3eb1721a} /* (30, 19, 2) {real, imag} */,
  {32'hbfb31b67, 32'hbdf9681a} /* (30, 19, 1) {real, imag} */,
  {32'hbf7f735e, 32'h00000000} /* (30, 19, 0) {real, imag} */,
  {32'hbfcd0918, 32'hbcc611a0} /* (30, 18, 31) {real, imag} */,
  {32'h3f268f4d, 32'hbe5fc4aa} /* (30, 18, 30) {real, imag} */,
  {32'h3d16b73b, 32'h3e6a85d3} /* (30, 18, 29) {real, imag} */,
  {32'hbe877c7e, 32'h3da44c72} /* (30, 18, 28) {real, imag} */,
  {32'h3e4b0ac5, 32'hbe6e463b} /* (30, 18, 27) {real, imag} */,
  {32'h3c2ae650, 32'h3df3c866} /* (30, 18, 26) {real, imag} */,
  {32'hbd08bdf4, 32'h3dde1a0d} /* (30, 18, 25) {real, imag} */,
  {32'h3d70c3cf, 32'hbb7acf40} /* (30, 18, 24) {real, imag} */,
  {32'h3d2d25ec, 32'h3d8ecc4e} /* (30, 18, 23) {real, imag} */,
  {32'hbd180838, 32'hbcc1008e} /* (30, 18, 22) {real, imag} */,
  {32'h3d90ae03, 32'hbddd60fc} /* (30, 18, 21) {real, imag} */,
  {32'h3d7eba70, 32'h3d8e2a33} /* (30, 18, 20) {real, imag} */,
  {32'hbd13f78c, 32'h3c168f78} /* (30, 18, 19) {real, imag} */,
  {32'h3b480a1c, 32'hbc9d3f72} /* (30, 18, 18) {real, imag} */,
  {32'h3d65283f, 32'hbd1704a5} /* (30, 18, 17) {real, imag} */,
  {32'h3c25dbb8, 32'h00000000} /* (30, 18, 16) {real, imag} */,
  {32'h3d65283f, 32'h3d1704a5} /* (30, 18, 15) {real, imag} */,
  {32'h3b480a1c, 32'h3c9d3f72} /* (30, 18, 14) {real, imag} */,
  {32'hbd13f78c, 32'hbc168f78} /* (30, 18, 13) {real, imag} */,
  {32'h3d7eba70, 32'hbd8e2a33} /* (30, 18, 12) {real, imag} */,
  {32'h3d90ae03, 32'h3ddd60fc} /* (30, 18, 11) {real, imag} */,
  {32'hbd180838, 32'h3cc1008e} /* (30, 18, 10) {real, imag} */,
  {32'h3d2d25ec, 32'hbd8ecc4e} /* (30, 18, 9) {real, imag} */,
  {32'h3d70c3cf, 32'h3b7acf40} /* (30, 18, 8) {real, imag} */,
  {32'hbd08bdf4, 32'hbdde1a0d} /* (30, 18, 7) {real, imag} */,
  {32'h3c2ae650, 32'hbdf3c866} /* (30, 18, 6) {real, imag} */,
  {32'h3e4b0ac5, 32'h3e6e463b} /* (30, 18, 5) {real, imag} */,
  {32'hbe877c7e, 32'hbda44c72} /* (30, 18, 4) {real, imag} */,
  {32'h3d16b73b, 32'hbe6a85d3} /* (30, 18, 3) {real, imag} */,
  {32'h3f268f4d, 32'h3e5fc4aa} /* (30, 18, 2) {real, imag} */,
  {32'hbfcd0918, 32'h3cc611a0} /* (30, 18, 1) {real, imag} */,
  {32'hbf869ff3, 32'h00000000} /* (30, 18, 0) {real, imag} */,
  {32'hbfde3232, 32'h3d21dad4} /* (30, 17, 31) {real, imag} */,
  {32'h3f2433f7, 32'hbe41182a} /* (30, 17, 30) {real, imag} */,
  {32'h3b8c49d8, 32'h3e207550} /* (30, 17, 29) {real, imag} */,
  {32'hbe2397fc, 32'h3de3aa31} /* (30, 17, 28) {real, imag} */,
  {32'h3e5c3fb8, 32'hbdf3dda5} /* (30, 17, 27) {real, imag} */,
  {32'h3acf94e0, 32'h3d8c4e9f} /* (30, 17, 26) {real, imag} */,
  {32'hbd99e7a2, 32'h3d75cc54} /* (30, 17, 25) {real, imag} */,
  {32'h3d4bcbf9, 32'hbd3513dc} /* (30, 17, 24) {real, imag} */,
  {32'h3d1f263e, 32'h3ced9a66} /* (30, 17, 23) {real, imag} */,
  {32'hba1b74a0, 32'h3dcdcc3e} /* (30, 17, 22) {real, imag} */,
  {32'h3dc417fa, 32'hbe2881f3} /* (30, 17, 21) {real, imag} */,
  {32'hbc2f1092, 32'h3c4e033e} /* (30, 17, 20) {real, imag} */,
  {32'hbcb26fd3, 32'hbbbb3920} /* (30, 17, 19) {real, imag} */,
  {32'h3cbef18a, 32'hbd46ec59} /* (30, 17, 18) {real, imag} */,
  {32'h38c09300, 32'h3dc20126} /* (30, 17, 17) {real, imag} */,
  {32'hbceeb35a, 32'h00000000} /* (30, 17, 16) {real, imag} */,
  {32'h38c09300, 32'hbdc20126} /* (30, 17, 15) {real, imag} */,
  {32'h3cbef18a, 32'h3d46ec59} /* (30, 17, 14) {real, imag} */,
  {32'hbcb26fd3, 32'h3bbb3920} /* (30, 17, 13) {real, imag} */,
  {32'hbc2f1092, 32'hbc4e033e} /* (30, 17, 12) {real, imag} */,
  {32'h3dc417fa, 32'h3e2881f3} /* (30, 17, 11) {real, imag} */,
  {32'hba1b74a0, 32'hbdcdcc3e} /* (30, 17, 10) {real, imag} */,
  {32'h3d1f263e, 32'hbced9a66} /* (30, 17, 9) {real, imag} */,
  {32'h3d4bcbf9, 32'h3d3513dc} /* (30, 17, 8) {real, imag} */,
  {32'hbd99e7a2, 32'hbd75cc54} /* (30, 17, 7) {real, imag} */,
  {32'h3acf94e0, 32'hbd8c4e9f} /* (30, 17, 6) {real, imag} */,
  {32'h3e5c3fb8, 32'h3df3dda5} /* (30, 17, 5) {real, imag} */,
  {32'hbe2397fc, 32'hbde3aa31} /* (30, 17, 4) {real, imag} */,
  {32'h3b8c49d8, 32'hbe207550} /* (30, 17, 3) {real, imag} */,
  {32'h3f2433f7, 32'h3e41182a} /* (30, 17, 2) {real, imag} */,
  {32'hbfde3232, 32'hbd21dad4} /* (30, 17, 1) {real, imag} */,
  {32'hbf914448, 32'h00000000} /* (30, 17, 0) {real, imag} */,
  {32'hbfe254ff, 32'hbc8e7540} /* (30, 16, 31) {real, imag} */,
  {32'h3f4ccf9c, 32'hbdf2b916} /* (30, 16, 30) {real, imag} */,
  {32'hbc0c0844, 32'hbd81b163} /* (30, 16, 29) {real, imag} */,
  {32'hbe494726, 32'h3d8a0240} /* (30, 16, 28) {real, imag} */,
  {32'h3e873877, 32'h3deb9e58} /* (30, 16, 27) {real, imag} */,
  {32'h3d570dda, 32'h3c9297bc} /* (30, 16, 26) {real, imag} */,
  {32'hbc7d8658, 32'hbdcb0bfd} /* (30, 16, 25) {real, imag} */,
  {32'h3e072472, 32'hbdc9bdef} /* (30, 16, 24) {real, imag} */,
  {32'hb9ff6c40, 32'h3dd83773} /* (30, 16, 23) {real, imag} */,
  {32'h3c569112, 32'hbd740ec6} /* (30, 16, 22) {real, imag} */,
  {32'hbb44ba20, 32'hbdc995f4} /* (30, 16, 21) {real, imag} */,
  {32'hbda13814, 32'h3d37f743} /* (30, 16, 20) {real, imag} */,
  {32'h3c2a80c2, 32'h3d88b2c6} /* (30, 16, 19) {real, imag} */,
  {32'h3d7434be, 32'h3d070e62} /* (30, 16, 18) {real, imag} */,
  {32'h3d4467a0, 32'hbd5b38bd} /* (30, 16, 17) {real, imag} */,
  {32'hbd92c86a, 32'h00000000} /* (30, 16, 16) {real, imag} */,
  {32'h3d4467a0, 32'h3d5b38bd} /* (30, 16, 15) {real, imag} */,
  {32'h3d7434be, 32'hbd070e62} /* (30, 16, 14) {real, imag} */,
  {32'h3c2a80c2, 32'hbd88b2c6} /* (30, 16, 13) {real, imag} */,
  {32'hbda13814, 32'hbd37f743} /* (30, 16, 12) {real, imag} */,
  {32'hbb44ba20, 32'h3dc995f4} /* (30, 16, 11) {real, imag} */,
  {32'h3c569112, 32'h3d740ec6} /* (30, 16, 10) {real, imag} */,
  {32'hb9ff6c40, 32'hbdd83773} /* (30, 16, 9) {real, imag} */,
  {32'h3e072472, 32'h3dc9bdef} /* (30, 16, 8) {real, imag} */,
  {32'hbc7d8658, 32'h3dcb0bfd} /* (30, 16, 7) {real, imag} */,
  {32'h3d570dda, 32'hbc9297bc} /* (30, 16, 6) {real, imag} */,
  {32'h3e873877, 32'hbdeb9e58} /* (30, 16, 5) {real, imag} */,
  {32'hbe494726, 32'hbd8a0240} /* (30, 16, 4) {real, imag} */,
  {32'hbc0c0844, 32'h3d81b163} /* (30, 16, 3) {real, imag} */,
  {32'h3f4ccf9c, 32'h3df2b916} /* (30, 16, 2) {real, imag} */,
  {32'hbfe254ff, 32'h3c8e7540} /* (30, 16, 1) {real, imag} */,
  {32'hbfa148ab, 32'h00000000} /* (30, 16, 0) {real, imag} */,
  {32'hbfd0c1a2, 32'hbddcfd22} /* (30, 15, 31) {real, imag} */,
  {32'h3f544331, 32'hbe063d7a} /* (30, 15, 30) {real, imag} */,
  {32'hbce0cf0a, 32'h3dd71a41} /* (30, 15, 29) {real, imag} */,
  {32'hbd42198c, 32'h3d5e731a} /* (30, 15, 28) {real, imag} */,
  {32'h3e503f00, 32'h3bd93890} /* (30, 15, 27) {real, imag} */,
  {32'h3b8a6f08, 32'h3afd2a40} /* (30, 15, 26) {real, imag} */,
  {32'h3c2f26e0, 32'hbc4fcda0} /* (30, 15, 25) {real, imag} */,
  {32'hbcba756a, 32'hbe030193} /* (30, 15, 24) {real, imag} */,
  {32'h3c60a901, 32'h3c64d3b5} /* (30, 15, 23) {real, imag} */,
  {32'h3d18caca, 32'hbbffa408} /* (30, 15, 22) {real, imag} */,
  {32'h3cf128f8, 32'h3cff5178} /* (30, 15, 21) {real, imag} */,
  {32'h3cb8c23f, 32'hbcb91a2d} /* (30, 15, 20) {real, imag} */,
  {32'hbda186a3, 32'hbd59294d} /* (30, 15, 19) {real, imag} */,
  {32'h3c883cee, 32'hbbf1dc08} /* (30, 15, 18) {real, imag} */,
  {32'h3d67543c, 32'hbceb5a26} /* (30, 15, 17) {real, imag} */,
  {32'h3c2eba05, 32'h00000000} /* (30, 15, 16) {real, imag} */,
  {32'h3d67543c, 32'h3ceb5a26} /* (30, 15, 15) {real, imag} */,
  {32'h3c883cee, 32'h3bf1dc08} /* (30, 15, 14) {real, imag} */,
  {32'hbda186a3, 32'h3d59294d} /* (30, 15, 13) {real, imag} */,
  {32'h3cb8c23f, 32'h3cb91a2d} /* (30, 15, 12) {real, imag} */,
  {32'h3cf128f8, 32'hbcff5178} /* (30, 15, 11) {real, imag} */,
  {32'h3d18caca, 32'h3bffa408} /* (30, 15, 10) {real, imag} */,
  {32'h3c60a901, 32'hbc64d3b5} /* (30, 15, 9) {real, imag} */,
  {32'hbcba756a, 32'h3e030193} /* (30, 15, 8) {real, imag} */,
  {32'h3c2f26e0, 32'h3c4fcda0} /* (30, 15, 7) {real, imag} */,
  {32'h3b8a6f08, 32'hbafd2a40} /* (30, 15, 6) {real, imag} */,
  {32'h3e503f00, 32'hbbd93890} /* (30, 15, 5) {real, imag} */,
  {32'hbd42198c, 32'hbd5e731a} /* (30, 15, 4) {real, imag} */,
  {32'hbce0cf0a, 32'hbdd71a41} /* (30, 15, 3) {real, imag} */,
  {32'h3f544331, 32'h3e063d7a} /* (30, 15, 2) {real, imag} */,
  {32'hbfd0c1a2, 32'h3ddcfd22} /* (30, 15, 1) {real, imag} */,
  {32'hbfa9d3b8, 32'h00000000} /* (30, 15, 0) {real, imag} */,
  {32'hbfbba010, 32'hbcaaf020} /* (30, 14, 31) {real, imag} */,
  {32'h3f53babb, 32'hbe03b202} /* (30, 14, 30) {real, imag} */,
  {32'hbc3aa3bc, 32'h3e081961} /* (30, 14, 29) {real, imag} */,
  {32'hbdd47eba, 32'h3dc62e52} /* (30, 14, 28) {real, imag} */,
  {32'h3e2bf0d7, 32'h3d7b5194} /* (30, 14, 27) {real, imag} */,
  {32'h3deccb4c, 32'h3cfab60a} /* (30, 14, 26) {real, imag} */,
  {32'hbcbdf1ef, 32'h3db7334b} /* (30, 14, 25) {real, imag} */,
  {32'h3ce5ba52, 32'hbde920fe} /* (30, 14, 24) {real, imag} */,
  {32'h3c51d3cf, 32'hbbd50e08} /* (30, 14, 23) {real, imag} */,
  {32'h3ca48ace, 32'h3d7d8c2f} /* (30, 14, 22) {real, imag} */,
  {32'h3d192e5a, 32'h3d1c1d67} /* (30, 14, 21) {real, imag} */,
  {32'hbc46be46, 32'hbd3429aa} /* (30, 14, 20) {real, imag} */,
  {32'hbd89ecba, 32'h3d5cf488} /* (30, 14, 19) {real, imag} */,
  {32'hbc1f43e9, 32'hbdd36a26} /* (30, 14, 18) {real, imag} */,
  {32'hbd42763d, 32'h3cd4fe6e} /* (30, 14, 17) {real, imag} */,
  {32'h3d0aa920, 32'h00000000} /* (30, 14, 16) {real, imag} */,
  {32'hbd42763d, 32'hbcd4fe6e} /* (30, 14, 15) {real, imag} */,
  {32'hbc1f43e9, 32'h3dd36a26} /* (30, 14, 14) {real, imag} */,
  {32'hbd89ecba, 32'hbd5cf488} /* (30, 14, 13) {real, imag} */,
  {32'hbc46be46, 32'h3d3429aa} /* (30, 14, 12) {real, imag} */,
  {32'h3d192e5a, 32'hbd1c1d67} /* (30, 14, 11) {real, imag} */,
  {32'h3ca48ace, 32'hbd7d8c2f} /* (30, 14, 10) {real, imag} */,
  {32'h3c51d3cf, 32'h3bd50e08} /* (30, 14, 9) {real, imag} */,
  {32'h3ce5ba52, 32'h3de920fe} /* (30, 14, 8) {real, imag} */,
  {32'hbcbdf1ef, 32'hbdb7334b} /* (30, 14, 7) {real, imag} */,
  {32'h3deccb4c, 32'hbcfab60a} /* (30, 14, 6) {real, imag} */,
  {32'h3e2bf0d7, 32'hbd7b5194} /* (30, 14, 5) {real, imag} */,
  {32'hbdd47eba, 32'hbdc62e52} /* (30, 14, 4) {real, imag} */,
  {32'hbc3aa3bc, 32'hbe081961} /* (30, 14, 3) {real, imag} */,
  {32'h3f53babb, 32'h3e03b202} /* (30, 14, 2) {real, imag} */,
  {32'hbfbba010, 32'h3caaf020} /* (30, 14, 1) {real, imag} */,
  {32'hbfa2b867, 32'h00000000} /* (30, 14, 0) {real, imag} */,
  {32'hbfb040bb, 32'h3cce2ab8} /* (30, 13, 31) {real, imag} */,
  {32'h3f5e455d, 32'hbe3efae4} /* (30, 13, 30) {real, imag} */,
  {32'h3d0e74b0, 32'hbcb09a94} /* (30, 13, 29) {real, imag} */,
  {32'hbdbe7c3c, 32'h3e0b8a06} /* (30, 13, 28) {real, imag} */,
  {32'h3dd5e4c4, 32'h3d87e3b4} /* (30, 13, 27) {real, imag} */,
  {32'h3d9d38a0, 32'hbc7e29c6} /* (30, 13, 26) {real, imag} */,
  {32'hbe0ccef0, 32'h3dd35107} /* (30, 13, 25) {real, imag} */,
  {32'hbcfd540d, 32'hbd2b8c38} /* (30, 13, 24) {real, imag} */,
  {32'h3c2fd3a2, 32'h3d2e3798} /* (30, 13, 23) {real, imag} */,
  {32'h3d4d4efc, 32'hbc5d43e4} /* (30, 13, 22) {real, imag} */,
  {32'hbbaabf48, 32'hbdfaa8ae} /* (30, 13, 21) {real, imag} */,
  {32'hbda78ccf, 32'h3cad35e2} /* (30, 13, 20) {real, imag} */,
  {32'h3d26c3e0, 32'hbd40877d} /* (30, 13, 19) {real, imag} */,
  {32'hbc8b8a16, 32'hbd85cfba} /* (30, 13, 18) {real, imag} */,
  {32'h3d222560, 32'hba0d3830} /* (30, 13, 17) {real, imag} */,
  {32'h3d0a1228, 32'h00000000} /* (30, 13, 16) {real, imag} */,
  {32'h3d222560, 32'h3a0d3830} /* (30, 13, 15) {real, imag} */,
  {32'hbc8b8a16, 32'h3d85cfba} /* (30, 13, 14) {real, imag} */,
  {32'h3d26c3e0, 32'h3d40877d} /* (30, 13, 13) {real, imag} */,
  {32'hbda78ccf, 32'hbcad35e2} /* (30, 13, 12) {real, imag} */,
  {32'hbbaabf48, 32'h3dfaa8ae} /* (30, 13, 11) {real, imag} */,
  {32'h3d4d4efc, 32'h3c5d43e4} /* (30, 13, 10) {real, imag} */,
  {32'h3c2fd3a2, 32'hbd2e3798} /* (30, 13, 9) {real, imag} */,
  {32'hbcfd540d, 32'h3d2b8c38} /* (30, 13, 8) {real, imag} */,
  {32'hbe0ccef0, 32'hbdd35107} /* (30, 13, 7) {real, imag} */,
  {32'h3d9d38a0, 32'h3c7e29c6} /* (30, 13, 6) {real, imag} */,
  {32'h3dd5e4c4, 32'hbd87e3b4} /* (30, 13, 5) {real, imag} */,
  {32'hbdbe7c3c, 32'hbe0b8a06} /* (30, 13, 4) {real, imag} */,
  {32'h3d0e74b0, 32'h3cb09a94} /* (30, 13, 3) {real, imag} */,
  {32'h3f5e455d, 32'h3e3efae4} /* (30, 13, 2) {real, imag} */,
  {32'hbfb040bb, 32'hbcce2ab8} /* (30, 13, 1) {real, imag} */,
  {32'hbfb2da65, 32'h00000000} /* (30, 13, 0) {real, imag} */,
  {32'hbf9007fc, 32'h3d72f724} /* (30, 12, 31) {real, imag} */,
  {32'h3f3038e9, 32'hbe3a6e8b} /* (30, 12, 30) {real, imag} */,
  {32'hbcfa88cc, 32'hbdd23992} /* (30, 12, 29) {real, imag} */,
  {32'hbd5f65cc, 32'h3d79197e} /* (30, 12, 28) {real, imag} */,
  {32'h3de7b8aa, 32'hbde4eeb0} /* (30, 12, 27) {real, imag} */,
  {32'hbd933aca, 32'h3d2c4636} /* (30, 12, 26) {real, imag} */,
  {32'hbc5bd544, 32'h3db74c74} /* (30, 12, 25) {real, imag} */,
  {32'h3ca811a2, 32'h3c001750} /* (30, 12, 24) {real, imag} */,
  {32'hbd6b122d, 32'h3d079886} /* (30, 12, 23) {real, imag} */,
  {32'hbbc5aac4, 32'hbc5e92d0} /* (30, 12, 22) {real, imag} */,
  {32'hbc8b5040, 32'hbd0ec64a} /* (30, 12, 21) {real, imag} */,
  {32'hbccd8fb6, 32'hbd2a1f44} /* (30, 12, 20) {real, imag} */,
  {32'hbd297776, 32'h3c89ac7d} /* (30, 12, 19) {real, imag} */,
  {32'hbc86c0ff, 32'h3d2363a9} /* (30, 12, 18) {real, imag} */,
  {32'h3c73b488, 32'h3c9b02e6} /* (30, 12, 17) {real, imag} */,
  {32'hbc48e56c, 32'h00000000} /* (30, 12, 16) {real, imag} */,
  {32'h3c73b488, 32'hbc9b02e6} /* (30, 12, 15) {real, imag} */,
  {32'hbc86c0ff, 32'hbd2363a9} /* (30, 12, 14) {real, imag} */,
  {32'hbd297776, 32'hbc89ac7d} /* (30, 12, 13) {real, imag} */,
  {32'hbccd8fb6, 32'h3d2a1f44} /* (30, 12, 12) {real, imag} */,
  {32'hbc8b5040, 32'h3d0ec64a} /* (30, 12, 11) {real, imag} */,
  {32'hbbc5aac4, 32'h3c5e92d0} /* (30, 12, 10) {real, imag} */,
  {32'hbd6b122d, 32'hbd079886} /* (30, 12, 9) {real, imag} */,
  {32'h3ca811a2, 32'hbc001750} /* (30, 12, 8) {real, imag} */,
  {32'hbc5bd544, 32'hbdb74c74} /* (30, 12, 7) {real, imag} */,
  {32'hbd933aca, 32'hbd2c4636} /* (30, 12, 6) {real, imag} */,
  {32'h3de7b8aa, 32'h3de4eeb0} /* (30, 12, 5) {real, imag} */,
  {32'hbd5f65cc, 32'hbd79197e} /* (30, 12, 4) {real, imag} */,
  {32'hbcfa88cc, 32'h3dd23992} /* (30, 12, 3) {real, imag} */,
  {32'h3f3038e9, 32'h3e3a6e8b} /* (30, 12, 2) {real, imag} */,
  {32'hbf9007fc, 32'hbd72f724} /* (30, 12, 1) {real, imag} */,
  {32'hbf9092ab, 32'h00000000} /* (30, 12, 0) {real, imag} */,
  {32'hbf29331c, 32'h3d644dbc} /* (30, 11, 31) {real, imag} */,
  {32'h3efcb6ee, 32'hbcb218e0} /* (30, 11, 30) {real, imag} */,
  {32'hbe034400, 32'hbd37f904} /* (30, 11, 29) {real, imag} */,
  {32'hbbfd8798, 32'hbcf70113} /* (30, 11, 28) {real, imag} */,
  {32'h3dfa1728, 32'hbdabd694} /* (30, 11, 27) {real, imag} */,
  {32'h3d5a4779, 32'h3c4abe08} /* (30, 11, 26) {real, imag} */,
  {32'hbd28e22a, 32'h3d90a042} /* (30, 11, 25) {real, imag} */,
  {32'h3cd3ba32, 32'hbdfd453d} /* (30, 11, 24) {real, imag} */,
  {32'hbda2fd7e, 32'hbcfe092e} /* (30, 11, 23) {real, imag} */,
  {32'hbd5bb13a, 32'h3e715ff7} /* (30, 11, 22) {real, imag} */,
  {32'hbd74aa0e, 32'hbd0421fc} /* (30, 11, 21) {real, imag} */,
  {32'h3d54217a, 32'hbd7a34d0} /* (30, 11, 20) {real, imag} */,
  {32'hbdbb4aae, 32'hbdab3d68} /* (30, 11, 19) {real, imag} */,
  {32'h3c436dce, 32'h3ccc4e9e} /* (30, 11, 18) {real, imag} */,
  {32'h3d3f1791, 32'hbcc42174} /* (30, 11, 17) {real, imag} */,
  {32'h3d3e19b7, 32'h00000000} /* (30, 11, 16) {real, imag} */,
  {32'h3d3f1791, 32'h3cc42174} /* (30, 11, 15) {real, imag} */,
  {32'h3c436dce, 32'hbccc4e9e} /* (30, 11, 14) {real, imag} */,
  {32'hbdbb4aae, 32'h3dab3d68} /* (30, 11, 13) {real, imag} */,
  {32'h3d54217a, 32'h3d7a34d0} /* (30, 11, 12) {real, imag} */,
  {32'hbd74aa0e, 32'h3d0421fc} /* (30, 11, 11) {real, imag} */,
  {32'hbd5bb13a, 32'hbe715ff7} /* (30, 11, 10) {real, imag} */,
  {32'hbda2fd7e, 32'h3cfe092e} /* (30, 11, 9) {real, imag} */,
  {32'h3cd3ba32, 32'h3dfd453d} /* (30, 11, 8) {real, imag} */,
  {32'hbd28e22a, 32'hbd90a042} /* (30, 11, 7) {real, imag} */,
  {32'h3d5a4779, 32'hbc4abe08} /* (30, 11, 6) {real, imag} */,
  {32'h3dfa1728, 32'h3dabd694} /* (30, 11, 5) {real, imag} */,
  {32'hbbfd8798, 32'h3cf70113} /* (30, 11, 4) {real, imag} */,
  {32'hbe034400, 32'h3d37f904} /* (30, 11, 3) {real, imag} */,
  {32'h3efcb6ee, 32'h3cb218e0} /* (30, 11, 2) {real, imag} */,
  {32'hbf29331c, 32'hbd644dbc} /* (30, 11, 1) {real, imag} */,
  {32'hbf1504f0, 32'h00000000} /* (30, 11, 0) {real, imag} */,
  {32'h3ee51c20, 32'h3d10120e} /* (30, 10, 31) {real, imag} */,
  {32'hbe288678, 32'h3e527f03} /* (30, 10, 30) {real, imag} */,
  {32'hbdc2b0f0, 32'hbd949fb6} /* (30, 10, 29) {real, imag} */,
  {32'h3dfaf1d1, 32'hbc88936e} /* (30, 10, 28) {real, imag} */,
  {32'h3bc761b0, 32'hbdd87ee8} /* (30, 10, 27) {real, imag} */,
  {32'h3d03ec6e, 32'hba4d3ab0} /* (30, 10, 26) {real, imag} */,
  {32'hbd1a4d82, 32'hbd193ef1} /* (30, 10, 25) {real, imag} */,
  {32'hbd83f08e, 32'hbdcda19d} /* (30, 10, 24) {real, imag} */,
  {32'h3cea0932, 32'h3ca09cc4} /* (30, 10, 23) {real, imag} */,
  {32'h3bec47f0, 32'h3d87632c} /* (30, 10, 22) {real, imag} */,
  {32'hbcf36eb4, 32'hbcc83b48} /* (30, 10, 21) {real, imag} */,
  {32'hbd8fd4d8, 32'h3d90ef90} /* (30, 10, 20) {real, imag} */,
  {32'hbcdc0ceb, 32'h3bee8bb0} /* (30, 10, 19) {real, imag} */,
  {32'hbbf41880, 32'hbd75841b} /* (30, 10, 18) {real, imag} */,
  {32'h3c340076, 32'hbd3e9c3a} /* (30, 10, 17) {real, imag} */,
  {32'h3d33c78d, 32'h00000000} /* (30, 10, 16) {real, imag} */,
  {32'h3c340076, 32'h3d3e9c3a} /* (30, 10, 15) {real, imag} */,
  {32'hbbf41880, 32'h3d75841b} /* (30, 10, 14) {real, imag} */,
  {32'hbcdc0ceb, 32'hbbee8bb0} /* (30, 10, 13) {real, imag} */,
  {32'hbd8fd4d8, 32'hbd90ef90} /* (30, 10, 12) {real, imag} */,
  {32'hbcf36eb4, 32'h3cc83b48} /* (30, 10, 11) {real, imag} */,
  {32'h3bec47f0, 32'hbd87632c} /* (30, 10, 10) {real, imag} */,
  {32'h3cea0932, 32'hbca09cc4} /* (30, 10, 9) {real, imag} */,
  {32'hbd83f08e, 32'h3dcda19d} /* (30, 10, 8) {real, imag} */,
  {32'hbd1a4d82, 32'h3d193ef1} /* (30, 10, 7) {real, imag} */,
  {32'h3d03ec6e, 32'h3a4d3ab0} /* (30, 10, 6) {real, imag} */,
  {32'h3bc761b0, 32'h3dd87ee8} /* (30, 10, 5) {real, imag} */,
  {32'h3dfaf1d1, 32'h3c88936e} /* (30, 10, 4) {real, imag} */,
  {32'hbdc2b0f0, 32'h3d949fb6} /* (30, 10, 3) {real, imag} */,
  {32'hbe288678, 32'hbe527f03} /* (30, 10, 2) {real, imag} */,
  {32'h3ee51c20, 32'hbd10120e} /* (30, 10, 1) {real, imag} */,
  {32'h3e4559e5, 32'h00000000} /* (30, 10, 0) {real, imag} */,
  {32'h3f94f304, 32'hbde6d254} /* (30, 9, 31) {real, imag} */,
  {32'hbed314ae, 32'h3e847efd} /* (30, 9, 30) {real, imag} */,
  {32'hbc65ff80, 32'hbb1ecc78} /* (30, 9, 29) {real, imag} */,
  {32'h3d0641c6, 32'hbc0e7c44} /* (30, 9, 28) {real, imag} */,
  {32'hbca13700, 32'h3c91323a} /* (30, 9, 27) {real, imag} */,
  {32'hbd20d4f6, 32'hbc18dc20} /* (30, 9, 26) {real, imag} */,
  {32'h3cd72900, 32'hbc5efc68} /* (30, 9, 25) {real, imag} */,
  {32'hbd76422c, 32'h3db50f40} /* (30, 9, 24) {real, imag} */,
  {32'h3bc02f4e, 32'h3cec043e} /* (30, 9, 23) {real, imag} */,
  {32'hbdac8037, 32'hbcbbddce} /* (30, 9, 22) {real, imag} */,
  {32'hbc965ace, 32'h3d8d9cdc} /* (30, 9, 21) {real, imag} */,
  {32'hbc684ccc, 32'hbd150709} /* (30, 9, 20) {real, imag} */,
  {32'h3db9991c, 32'h3d841c23} /* (30, 9, 19) {real, imag} */,
  {32'h3d0fa6b5, 32'h3da32e1e} /* (30, 9, 18) {real, imag} */,
  {32'h3c222836, 32'h3d78ee35} /* (30, 9, 17) {real, imag} */,
  {32'hbdb99dc2, 32'h00000000} /* (30, 9, 16) {real, imag} */,
  {32'h3c222836, 32'hbd78ee35} /* (30, 9, 15) {real, imag} */,
  {32'h3d0fa6b5, 32'hbda32e1e} /* (30, 9, 14) {real, imag} */,
  {32'h3db9991c, 32'hbd841c23} /* (30, 9, 13) {real, imag} */,
  {32'hbc684ccc, 32'h3d150709} /* (30, 9, 12) {real, imag} */,
  {32'hbc965ace, 32'hbd8d9cdc} /* (30, 9, 11) {real, imag} */,
  {32'hbdac8037, 32'h3cbbddce} /* (30, 9, 10) {real, imag} */,
  {32'h3bc02f4e, 32'hbcec043e} /* (30, 9, 9) {real, imag} */,
  {32'hbd76422c, 32'hbdb50f40} /* (30, 9, 8) {real, imag} */,
  {32'h3cd72900, 32'h3c5efc68} /* (30, 9, 7) {real, imag} */,
  {32'hbd20d4f6, 32'h3c18dc20} /* (30, 9, 6) {real, imag} */,
  {32'hbca13700, 32'hbc91323a} /* (30, 9, 5) {real, imag} */,
  {32'h3d0641c6, 32'h3c0e7c44} /* (30, 9, 4) {real, imag} */,
  {32'hbc65ff80, 32'h3b1ecc78} /* (30, 9, 3) {real, imag} */,
  {32'hbed314ae, 32'hbe847efd} /* (30, 9, 2) {real, imag} */,
  {32'h3f94f304, 32'h3de6d254} /* (30, 9, 1) {real, imag} */,
  {32'h3f075467, 32'h00000000} /* (30, 9, 0) {real, imag} */,
  {32'h3fc2193a, 32'hbe9356a4} /* (30, 8, 31) {real, imag} */,
  {32'hbf01b462, 32'h3ebcf034} /* (30, 8, 30) {real, imag} */,
  {32'hbd94dac4, 32'hbcc194bb} /* (30, 8, 29) {real, imag} */,
  {32'h3e08962b, 32'h3cd9d550} /* (30, 8, 28) {real, imag} */,
  {32'hbe2ce2be, 32'h3d89e1e6} /* (30, 8, 27) {real, imag} */,
  {32'h3b31aca0, 32'hbd4d9325} /* (30, 8, 26) {real, imag} */,
  {32'hbccde51c, 32'hbcb85bb0} /* (30, 8, 25) {real, imag} */,
  {32'hbde4cdaa, 32'h3cf2cb46} /* (30, 8, 24) {real, imag} */,
  {32'h3c64ccac, 32'hbcbf0610} /* (30, 8, 23) {real, imag} */,
  {32'h3dc9b2e9, 32'h3c065f4c} /* (30, 8, 22) {real, imag} */,
  {32'hbaae5500, 32'h3dd1700c} /* (30, 8, 21) {real, imag} */,
  {32'h3db2cbce, 32'hbd0d68d6} /* (30, 8, 20) {real, imag} */,
  {32'hbd19a16a, 32'h3d3f74cd} /* (30, 8, 19) {real, imag} */,
  {32'hbd18f81f, 32'hbd0ba321} /* (30, 8, 18) {real, imag} */,
  {32'h3d9afaa8, 32'h3d6f1da1} /* (30, 8, 17) {real, imag} */,
  {32'hbdfb0862, 32'h00000000} /* (30, 8, 16) {real, imag} */,
  {32'h3d9afaa8, 32'hbd6f1da1} /* (30, 8, 15) {real, imag} */,
  {32'hbd18f81f, 32'h3d0ba321} /* (30, 8, 14) {real, imag} */,
  {32'hbd19a16a, 32'hbd3f74cd} /* (30, 8, 13) {real, imag} */,
  {32'h3db2cbce, 32'h3d0d68d6} /* (30, 8, 12) {real, imag} */,
  {32'hbaae5500, 32'hbdd1700c} /* (30, 8, 11) {real, imag} */,
  {32'h3dc9b2e9, 32'hbc065f4c} /* (30, 8, 10) {real, imag} */,
  {32'h3c64ccac, 32'h3cbf0610} /* (30, 8, 9) {real, imag} */,
  {32'hbde4cdaa, 32'hbcf2cb46} /* (30, 8, 8) {real, imag} */,
  {32'hbccde51c, 32'h3cb85bb0} /* (30, 8, 7) {real, imag} */,
  {32'h3b31aca0, 32'h3d4d9325} /* (30, 8, 6) {real, imag} */,
  {32'hbe2ce2be, 32'hbd89e1e6} /* (30, 8, 5) {real, imag} */,
  {32'h3e08962b, 32'hbcd9d550} /* (30, 8, 4) {real, imag} */,
  {32'hbd94dac4, 32'h3cc194bb} /* (30, 8, 3) {real, imag} */,
  {32'hbf01b462, 32'hbebcf034} /* (30, 8, 2) {real, imag} */,
  {32'h3fc2193a, 32'h3e9356a4} /* (30, 8, 1) {real, imag} */,
  {32'h3ee53d7c, 32'h00000000} /* (30, 8, 0) {real, imag} */,
  {32'h3fbf7809, 32'hbe360d46} /* (30, 7, 31) {real, imag} */,
  {32'hbef58014, 32'h3eeed588} /* (30, 7, 30) {real, imag} */,
  {32'hbdfb48c0, 32'h3d883798} /* (30, 7, 29) {real, imag} */,
  {32'h3e252b70, 32'hbcc2f151} /* (30, 7, 28) {real, imag} */,
  {32'hbe1940c5, 32'h3d9afd42} /* (30, 7, 27) {real, imag} */,
  {32'hbd38ea92, 32'h3ba059b0} /* (30, 7, 26) {real, imag} */,
  {32'h3da9c6bb, 32'hbb3d40c0} /* (30, 7, 25) {real, imag} */,
  {32'hbd9863ba, 32'h3ccece57} /* (30, 7, 24) {real, imag} */,
  {32'hbbcbcebe, 32'hbd34137f} /* (30, 7, 23) {real, imag} */,
  {32'h3d42ca34, 32'hbdbdd154} /* (30, 7, 22) {real, imag} */,
  {32'hbdc7025e, 32'hbcfa519c} /* (30, 7, 21) {real, imag} */,
  {32'hbd42aed8, 32'hbd2c110a} /* (30, 7, 20) {real, imag} */,
  {32'h3d1c2488, 32'h3b000438} /* (30, 7, 19) {real, imag} */,
  {32'hbd0bd38f, 32'h3d3b2b25} /* (30, 7, 18) {real, imag} */,
  {32'hbb58e758, 32'h3b8c01da} /* (30, 7, 17) {real, imag} */,
  {32'hbc1c7ed6, 32'h00000000} /* (30, 7, 16) {real, imag} */,
  {32'hbb58e758, 32'hbb8c01da} /* (30, 7, 15) {real, imag} */,
  {32'hbd0bd38f, 32'hbd3b2b25} /* (30, 7, 14) {real, imag} */,
  {32'h3d1c2488, 32'hbb000438} /* (30, 7, 13) {real, imag} */,
  {32'hbd42aed8, 32'h3d2c110a} /* (30, 7, 12) {real, imag} */,
  {32'hbdc7025e, 32'h3cfa519c} /* (30, 7, 11) {real, imag} */,
  {32'h3d42ca34, 32'h3dbdd154} /* (30, 7, 10) {real, imag} */,
  {32'hbbcbcebe, 32'h3d34137f} /* (30, 7, 9) {real, imag} */,
  {32'hbd9863ba, 32'hbccece57} /* (30, 7, 8) {real, imag} */,
  {32'h3da9c6bb, 32'h3b3d40c0} /* (30, 7, 7) {real, imag} */,
  {32'hbd38ea92, 32'hbba059b0} /* (30, 7, 6) {real, imag} */,
  {32'hbe1940c5, 32'hbd9afd42} /* (30, 7, 5) {real, imag} */,
  {32'h3e252b70, 32'h3cc2f151} /* (30, 7, 4) {real, imag} */,
  {32'hbdfb48c0, 32'hbd883798} /* (30, 7, 3) {real, imag} */,
  {32'hbef58014, 32'hbeeed588} /* (30, 7, 2) {real, imag} */,
  {32'h3fbf7809, 32'h3e360d46} /* (30, 7, 1) {real, imag} */,
  {32'h3f4361e0, 32'h00000000} /* (30, 7, 0) {real, imag} */,
  {32'h3fa76a60, 32'hbeb795fe} /* (30, 6, 31) {real, imag} */,
  {32'hbef1750c, 32'h3efaa71e} /* (30, 6, 30) {real, imag} */,
  {32'h3cffc7e6, 32'h39053d00} /* (30, 6, 29) {real, imag} */,
  {32'h3e19be17, 32'hbdcaec8c} /* (30, 6, 28) {real, imag} */,
  {32'hbde1595c, 32'h3d8698ed} /* (30, 6, 27) {real, imag} */,
  {32'hbe18fd6a, 32'h3d650ab8} /* (30, 6, 26) {real, imag} */,
  {32'hbc6610e2, 32'h3d1693d0} /* (30, 6, 25) {real, imag} */,
  {32'hbd078665, 32'h3de7fde8} /* (30, 6, 24) {real, imag} */,
  {32'hbd86e432, 32'hbd136cca} /* (30, 6, 23) {real, imag} */,
  {32'h3d804654, 32'hbe0e0eba} /* (30, 6, 22) {real, imag} */,
  {32'hbce4f97e, 32'h3e19e462} /* (30, 6, 21) {real, imag} */,
  {32'h3c3dd90c, 32'hbda71d06} /* (30, 6, 20) {real, imag} */,
  {32'h3d13ffe2, 32'hbcaa4a71} /* (30, 6, 19) {real, imag} */,
  {32'h3d1eba80, 32'hbd1f054b} /* (30, 6, 18) {real, imag} */,
  {32'h3bb82864, 32'h3c3aea26} /* (30, 6, 17) {real, imag} */,
  {32'hbdbc0852, 32'h00000000} /* (30, 6, 16) {real, imag} */,
  {32'h3bb82864, 32'hbc3aea26} /* (30, 6, 15) {real, imag} */,
  {32'h3d1eba80, 32'h3d1f054b} /* (30, 6, 14) {real, imag} */,
  {32'h3d13ffe2, 32'h3caa4a71} /* (30, 6, 13) {real, imag} */,
  {32'h3c3dd90c, 32'h3da71d06} /* (30, 6, 12) {real, imag} */,
  {32'hbce4f97e, 32'hbe19e462} /* (30, 6, 11) {real, imag} */,
  {32'h3d804654, 32'h3e0e0eba} /* (30, 6, 10) {real, imag} */,
  {32'hbd86e432, 32'h3d136cca} /* (30, 6, 9) {real, imag} */,
  {32'hbd078665, 32'hbde7fde8} /* (30, 6, 8) {real, imag} */,
  {32'hbc6610e2, 32'hbd1693d0} /* (30, 6, 7) {real, imag} */,
  {32'hbe18fd6a, 32'hbd650ab8} /* (30, 6, 6) {real, imag} */,
  {32'hbde1595c, 32'hbd8698ed} /* (30, 6, 5) {real, imag} */,
  {32'h3e19be17, 32'h3dcaec8c} /* (30, 6, 4) {real, imag} */,
  {32'h3cffc7e6, 32'hb9053d00} /* (30, 6, 3) {real, imag} */,
  {32'hbef1750c, 32'hbefaa71e} /* (30, 6, 2) {real, imag} */,
  {32'h3fa76a60, 32'h3eb795fe} /* (30, 6, 1) {real, imag} */,
  {32'h3f381878, 32'h00000000} /* (30, 6, 0) {real, imag} */,
  {32'h3f88925e, 32'hbf4a9406} /* (30, 5, 31) {real, imag} */,
  {32'hbdf35854, 32'h3f210e35} /* (30, 5, 30) {real, imag} */,
  {32'hbd078cab, 32'hbc856ab8} /* (30, 5, 29) {real, imag} */,
  {32'hbd8720ba, 32'h3cbd2f76} /* (30, 5, 28) {real, imag} */,
  {32'hbe0208e2, 32'h3c6e88be} /* (30, 5, 27) {real, imag} */,
  {32'hbd859582, 32'hbca3ba7c} /* (30, 5, 26) {real, imag} */,
  {32'h3c754640, 32'h3d3a37bb} /* (30, 5, 25) {real, imag} */,
  {32'h3d76a770, 32'h3dddb486} /* (30, 5, 24) {real, imag} */,
  {32'hbd4c383d, 32'hbc09a484} /* (30, 5, 23) {real, imag} */,
  {32'h3ca0f2cd, 32'h3bd1a368} /* (30, 5, 22) {real, imag} */,
  {32'hbcc1d797, 32'hbcec668a} /* (30, 5, 21) {real, imag} */,
  {32'hb981dc80, 32'hbd4ce0f2} /* (30, 5, 20) {real, imag} */,
  {32'hbd836052, 32'hbca26390} /* (30, 5, 19) {real, imag} */,
  {32'h3c0c363a, 32'h3c856cd2} /* (30, 5, 18) {real, imag} */,
  {32'h3c46e86a, 32'h3d7f898b} /* (30, 5, 17) {real, imag} */,
  {32'h3dc24ae2, 32'h00000000} /* (30, 5, 16) {real, imag} */,
  {32'h3c46e86a, 32'hbd7f898b} /* (30, 5, 15) {real, imag} */,
  {32'h3c0c363a, 32'hbc856cd2} /* (30, 5, 14) {real, imag} */,
  {32'hbd836052, 32'h3ca26390} /* (30, 5, 13) {real, imag} */,
  {32'hb981dc80, 32'h3d4ce0f2} /* (30, 5, 12) {real, imag} */,
  {32'hbcc1d797, 32'h3cec668a} /* (30, 5, 11) {real, imag} */,
  {32'h3ca0f2cd, 32'hbbd1a368} /* (30, 5, 10) {real, imag} */,
  {32'hbd4c383d, 32'h3c09a484} /* (30, 5, 9) {real, imag} */,
  {32'h3d76a770, 32'hbdddb486} /* (30, 5, 8) {real, imag} */,
  {32'h3c754640, 32'hbd3a37bb} /* (30, 5, 7) {real, imag} */,
  {32'hbd859582, 32'h3ca3ba7c} /* (30, 5, 6) {real, imag} */,
  {32'hbe0208e2, 32'hbc6e88be} /* (30, 5, 5) {real, imag} */,
  {32'hbd8720ba, 32'hbcbd2f76} /* (30, 5, 4) {real, imag} */,
  {32'hbd078cab, 32'h3c856ab8} /* (30, 5, 3) {real, imag} */,
  {32'hbdf35854, 32'hbf210e35} /* (30, 5, 2) {real, imag} */,
  {32'h3f88925e, 32'h3f4a9406} /* (30, 5, 1) {real, imag} */,
  {32'h3f34f976, 32'h00000000} /* (30, 5, 0) {real, imag} */,
  {32'h3f452738, 32'hbf877ed6} /* (30, 4, 31) {real, imag} */,
  {32'h3db44fe8, 32'h3f3c3232} /* (30, 4, 30) {real, imag} */,
  {32'hbe5716bc, 32'hbb02ec50} /* (30, 4, 29) {real, imag} */,
  {32'hbe23ec40, 32'h3ce38bdb} /* (30, 4, 28) {real, imag} */,
  {32'hbc9b97d0, 32'h3d1e941e} /* (30, 4, 27) {real, imag} */,
  {32'hbaca26f0, 32'h3d30b574} /* (30, 4, 26) {real, imag} */,
  {32'h3bca32d8, 32'hbd5aad3c} /* (30, 4, 25) {real, imag} */,
  {32'h3daba8ff, 32'h3c556e78} /* (30, 4, 24) {real, imag} */,
  {32'hbb987f1a, 32'hbc8ad09a} /* (30, 4, 23) {real, imag} */,
  {32'h3cf6ecd2, 32'hbb9e047e} /* (30, 4, 22) {real, imag} */,
  {32'hbc0af0fc, 32'hbd1b7564} /* (30, 4, 21) {real, imag} */,
  {32'h3d059c7f, 32'h3d4c551c} /* (30, 4, 20) {real, imag} */,
  {32'hbc8bdac1, 32'h3d01ae46} /* (30, 4, 19) {real, imag} */,
  {32'h3d5ddc7a, 32'h3dc5851c} /* (30, 4, 18) {real, imag} */,
  {32'hbd605db7, 32'h3d3ea624} /* (30, 4, 17) {real, imag} */,
  {32'h3b10a8f0, 32'h00000000} /* (30, 4, 16) {real, imag} */,
  {32'hbd605db7, 32'hbd3ea624} /* (30, 4, 15) {real, imag} */,
  {32'h3d5ddc7a, 32'hbdc5851c} /* (30, 4, 14) {real, imag} */,
  {32'hbc8bdac1, 32'hbd01ae46} /* (30, 4, 13) {real, imag} */,
  {32'h3d059c7f, 32'hbd4c551c} /* (30, 4, 12) {real, imag} */,
  {32'hbc0af0fc, 32'h3d1b7564} /* (30, 4, 11) {real, imag} */,
  {32'h3cf6ecd2, 32'h3b9e047e} /* (30, 4, 10) {real, imag} */,
  {32'hbb987f1a, 32'h3c8ad09a} /* (30, 4, 9) {real, imag} */,
  {32'h3daba8ff, 32'hbc556e78} /* (30, 4, 8) {real, imag} */,
  {32'h3bca32d8, 32'h3d5aad3c} /* (30, 4, 7) {real, imag} */,
  {32'hbaca26f0, 32'hbd30b574} /* (30, 4, 6) {real, imag} */,
  {32'hbc9b97d0, 32'hbd1e941e} /* (30, 4, 5) {real, imag} */,
  {32'hbe23ec40, 32'hbce38bdb} /* (30, 4, 4) {real, imag} */,
  {32'hbe5716bc, 32'h3b02ec50} /* (30, 4, 3) {real, imag} */,
  {32'h3db44fe8, 32'hbf3c3232} /* (30, 4, 2) {real, imag} */,
  {32'h3f452738, 32'h3f877ed6} /* (30, 4, 1) {real, imag} */,
  {32'h3f189924, 32'h00000000} /* (30, 4, 0) {real, imag} */,
  {32'h3f3a6dbb, 32'hbfa5d0ec} /* (30, 3, 31) {real, imag} */,
  {32'h3e2d18e4, 32'h3f2931a8} /* (30, 3, 30) {real, imag} */,
  {32'hbd8907d6, 32'h3d310f36} /* (30, 3, 29) {real, imag} */,
  {32'hbd9269a5, 32'h3e055439} /* (30, 3, 28) {real, imag} */,
  {32'hbdfa0e86, 32'h3de62f06} /* (30, 3, 27) {real, imag} */,
  {32'hbca9eb20, 32'hbdbb33c2} /* (30, 3, 26) {real, imag} */,
  {32'hbd11f527, 32'hbe084cb0} /* (30, 3, 25) {real, imag} */,
  {32'hbdbbf523, 32'h3e471738} /* (30, 3, 24) {real, imag} */,
  {32'hbd339005, 32'hbd044964} /* (30, 3, 23) {real, imag} */,
  {32'hbc285b8a, 32'h3d8ae64f} /* (30, 3, 22) {real, imag} */,
  {32'hbd5b8a75, 32'hbcf976fc} /* (30, 3, 21) {real, imag} */,
  {32'h3d896842, 32'hbc9593b2} /* (30, 3, 20) {real, imag} */,
  {32'hbcc7f34b, 32'hbd452b35} /* (30, 3, 19) {real, imag} */,
  {32'hbcb90ac9, 32'hbe0f9538} /* (30, 3, 18) {real, imag} */,
  {32'h3d890a11, 32'h3bdddde0} /* (30, 3, 17) {real, imag} */,
  {32'hbc6b246c, 32'h00000000} /* (30, 3, 16) {real, imag} */,
  {32'h3d890a11, 32'hbbdddde0} /* (30, 3, 15) {real, imag} */,
  {32'hbcb90ac9, 32'h3e0f9538} /* (30, 3, 14) {real, imag} */,
  {32'hbcc7f34b, 32'h3d452b35} /* (30, 3, 13) {real, imag} */,
  {32'h3d896842, 32'h3c9593b2} /* (30, 3, 12) {real, imag} */,
  {32'hbd5b8a75, 32'h3cf976fc} /* (30, 3, 11) {real, imag} */,
  {32'hbc285b8a, 32'hbd8ae64f} /* (30, 3, 10) {real, imag} */,
  {32'hbd339005, 32'h3d044964} /* (30, 3, 9) {real, imag} */,
  {32'hbdbbf523, 32'hbe471738} /* (30, 3, 8) {real, imag} */,
  {32'hbd11f527, 32'h3e084cb0} /* (30, 3, 7) {real, imag} */,
  {32'hbca9eb20, 32'h3dbb33c2} /* (30, 3, 6) {real, imag} */,
  {32'hbdfa0e86, 32'hbde62f06} /* (30, 3, 5) {real, imag} */,
  {32'hbd9269a5, 32'hbe055439} /* (30, 3, 4) {real, imag} */,
  {32'hbd8907d6, 32'hbd310f36} /* (30, 3, 3) {real, imag} */,
  {32'h3e2d18e4, 32'hbf2931a8} /* (30, 3, 2) {real, imag} */,
  {32'h3f3a6dbb, 32'h3fa5d0ec} /* (30, 3, 1) {real, imag} */,
  {32'h3efc264c, 32'h00000000} /* (30, 3, 0) {real, imag} */,
  {32'h3f1d0e60, 32'hbfa6db96} /* (30, 2, 31) {real, imag} */,
  {32'h3e48c590, 32'h3ef97a35} /* (30, 2, 30) {real, imag} */,
  {32'hbd67f341, 32'h3d0c1358} /* (30, 2, 29) {real, imag} */,
  {32'hbe2a5966, 32'h3e13965e} /* (30, 2, 28) {real, imag} */,
  {32'hbde3f9a0, 32'h3ccaf3b8} /* (30, 2, 27) {real, imag} */,
  {32'hbdc2d0ce, 32'hbdb58c7e} /* (30, 2, 26) {real, imag} */,
  {32'hbcaa141d, 32'hbdc968b5} /* (30, 2, 25) {real, imag} */,
  {32'h3ce418f6, 32'h3df168f4} /* (30, 2, 24) {real, imag} */,
  {32'hbc8e9cca, 32'hbbd0ed58} /* (30, 2, 23) {real, imag} */,
  {32'hbc030286, 32'h3db2ee22} /* (30, 2, 22) {real, imag} */,
  {32'hbb1eda00, 32'hbd5bacfc} /* (30, 2, 21) {real, imag} */,
  {32'h3d9bcd6e, 32'hbd21b156} /* (30, 2, 20) {real, imag} */,
  {32'hbd91e7c7, 32'h3c715302} /* (30, 2, 19) {real, imag} */,
  {32'hbd6493e2, 32'h3daaa72c} /* (30, 2, 18) {real, imag} */,
  {32'h3d24f242, 32'h3d0e39ca} /* (30, 2, 17) {real, imag} */,
  {32'h3d7c6fa4, 32'h00000000} /* (30, 2, 16) {real, imag} */,
  {32'h3d24f242, 32'hbd0e39ca} /* (30, 2, 15) {real, imag} */,
  {32'hbd6493e2, 32'hbdaaa72c} /* (30, 2, 14) {real, imag} */,
  {32'hbd91e7c7, 32'hbc715302} /* (30, 2, 13) {real, imag} */,
  {32'h3d9bcd6e, 32'h3d21b156} /* (30, 2, 12) {real, imag} */,
  {32'hbb1eda00, 32'h3d5bacfc} /* (30, 2, 11) {real, imag} */,
  {32'hbc030286, 32'hbdb2ee22} /* (30, 2, 10) {real, imag} */,
  {32'hbc8e9cca, 32'h3bd0ed58} /* (30, 2, 9) {real, imag} */,
  {32'h3ce418f6, 32'hbdf168f4} /* (30, 2, 8) {real, imag} */,
  {32'hbcaa141d, 32'h3dc968b5} /* (30, 2, 7) {real, imag} */,
  {32'hbdc2d0ce, 32'h3db58c7e} /* (30, 2, 6) {real, imag} */,
  {32'hbde3f9a0, 32'hbccaf3b8} /* (30, 2, 5) {real, imag} */,
  {32'hbe2a5966, 32'hbe13965e} /* (30, 2, 4) {real, imag} */,
  {32'hbd67f341, 32'hbd0c1358} /* (30, 2, 3) {real, imag} */,
  {32'h3e48c590, 32'hbef97a35} /* (30, 2, 2) {real, imag} */,
  {32'h3f1d0e60, 32'h3fa6db96} /* (30, 2, 1) {real, imag} */,
  {32'h3e9d9804, 32'h00000000} /* (30, 2, 0) {real, imag} */,
  {32'h3f001c50, 32'hbf91b9c6} /* (30, 1, 31) {real, imag} */,
  {32'h3e14636c, 32'h3f0bff6c} /* (30, 1, 30) {real, imag} */,
  {32'hbdb034ec, 32'h3d24e5c8} /* (30, 1, 29) {real, imag} */,
  {32'hbdc9c6b5, 32'h3e253b3a} /* (30, 1, 28) {real, imag} */,
  {32'hbdc0e6d1, 32'hbd85eb4a} /* (30, 1, 27) {real, imag} */,
  {32'hbdf6fedc, 32'hba167220} /* (30, 1, 26) {real, imag} */,
  {32'hbcd1642c, 32'hbe3a2a4a} /* (30, 1, 25) {real, imag} */,
  {32'h3c52b638, 32'h3deeaafd} /* (30, 1, 24) {real, imag} */,
  {32'h3d4e903f, 32'hbd0481ad} /* (30, 1, 23) {real, imag} */,
  {32'h3c6ddae2, 32'h3ca6d681} /* (30, 1, 22) {real, imag} */,
  {32'hbdac3bd4, 32'h3c4cdd64} /* (30, 1, 21) {real, imag} */,
  {32'hbbe32cf9, 32'h3d577852} /* (30, 1, 20) {real, imag} */,
  {32'h3db7920c, 32'hbdee1a55} /* (30, 1, 19) {real, imag} */,
  {32'h3cac354e, 32'h3d5ce5a1} /* (30, 1, 18) {real, imag} */,
  {32'hbbe386ac, 32'hbc4d98b4} /* (30, 1, 17) {real, imag} */,
  {32'hbcfc61b8, 32'h00000000} /* (30, 1, 16) {real, imag} */,
  {32'hbbe386ac, 32'h3c4d98b4} /* (30, 1, 15) {real, imag} */,
  {32'h3cac354e, 32'hbd5ce5a1} /* (30, 1, 14) {real, imag} */,
  {32'h3db7920c, 32'h3dee1a55} /* (30, 1, 13) {real, imag} */,
  {32'hbbe32cf9, 32'hbd577852} /* (30, 1, 12) {real, imag} */,
  {32'hbdac3bd4, 32'hbc4cdd64} /* (30, 1, 11) {real, imag} */,
  {32'h3c6ddae2, 32'hbca6d681} /* (30, 1, 10) {real, imag} */,
  {32'h3d4e903f, 32'h3d0481ad} /* (30, 1, 9) {real, imag} */,
  {32'h3c52b638, 32'hbdeeaafd} /* (30, 1, 8) {real, imag} */,
  {32'hbcd1642c, 32'h3e3a2a4a} /* (30, 1, 7) {real, imag} */,
  {32'hbdf6fedc, 32'h3a167220} /* (30, 1, 6) {real, imag} */,
  {32'hbdc0e6d1, 32'h3d85eb4a} /* (30, 1, 5) {real, imag} */,
  {32'hbdc9c6b5, 32'hbe253b3a} /* (30, 1, 4) {real, imag} */,
  {32'hbdb034ec, 32'hbd24e5c8} /* (30, 1, 3) {real, imag} */,
  {32'h3e14636c, 32'hbf0bff6c} /* (30, 1, 2) {real, imag} */,
  {32'h3f001c50, 32'h3f91b9c6} /* (30, 1, 1) {real, imag} */,
  {32'h3eb16c62, 32'h00000000} /* (30, 1, 0) {real, imag} */,
  {32'h3f07ae0e, 32'hbf57a7da} /* (30, 0, 31) {real, imag} */,
  {32'hbdde05a0, 32'h3efe4f10} /* (30, 0, 30) {real, imag} */,
  {32'hbcfe739c, 32'hbc80562c} /* (30, 0, 29) {real, imag} */,
  {32'hbc7d9ae8, 32'h3e345ee7} /* (30, 0, 28) {real, imag} */,
  {32'hbe0eb8b3, 32'hbdab2fbe} /* (30, 0, 27) {real, imag} */,
  {32'h3d84fc83, 32'hbca1c94e} /* (30, 0, 26) {real, imag} */,
  {32'hbc4114c8, 32'hbdcdb9bb} /* (30, 0, 25) {real, imag} */,
  {32'h3b297ba0, 32'h3d3182de} /* (30, 0, 24) {real, imag} */,
  {32'hbb5ff2a8, 32'hbb959cb0} /* (30, 0, 23) {real, imag} */,
  {32'hbc691bce, 32'hbd870e43} /* (30, 0, 22) {real, imag} */,
  {32'h3b2bef40, 32'h3b054fb0} /* (30, 0, 21) {real, imag} */,
  {32'hbd3a1ffb, 32'h3cbaefc2} /* (30, 0, 20) {real, imag} */,
  {32'hbc304c3e, 32'hbc4f82cc} /* (30, 0, 19) {real, imag} */,
  {32'hbd3e6790, 32'h3cb096e1} /* (30, 0, 18) {real, imag} */,
  {32'h3cb4ea84, 32'hbbc25290} /* (30, 0, 17) {real, imag} */,
  {32'h3c16074c, 32'h00000000} /* (30, 0, 16) {real, imag} */,
  {32'h3cb4ea84, 32'h3bc25290} /* (30, 0, 15) {real, imag} */,
  {32'hbd3e6790, 32'hbcb096e1} /* (30, 0, 14) {real, imag} */,
  {32'hbc304c3e, 32'h3c4f82cc} /* (30, 0, 13) {real, imag} */,
  {32'hbd3a1ffb, 32'hbcbaefc2} /* (30, 0, 12) {real, imag} */,
  {32'h3b2bef40, 32'hbb054fb0} /* (30, 0, 11) {real, imag} */,
  {32'hbc691bce, 32'h3d870e43} /* (30, 0, 10) {real, imag} */,
  {32'hbb5ff2a8, 32'h3b959cb0} /* (30, 0, 9) {real, imag} */,
  {32'h3b297ba0, 32'hbd3182de} /* (30, 0, 8) {real, imag} */,
  {32'hbc4114c8, 32'h3dcdb9bb} /* (30, 0, 7) {real, imag} */,
  {32'h3d84fc83, 32'h3ca1c94e} /* (30, 0, 6) {real, imag} */,
  {32'hbe0eb8b3, 32'h3dab2fbe} /* (30, 0, 5) {real, imag} */,
  {32'hbc7d9ae8, 32'hbe345ee7} /* (30, 0, 4) {real, imag} */,
  {32'hbcfe739c, 32'h3c80562c} /* (30, 0, 3) {real, imag} */,
  {32'hbdde05a0, 32'hbefe4f10} /* (30, 0, 2) {real, imag} */,
  {32'h3f07ae0e, 32'h3f57a7da} /* (30, 0, 1) {real, imag} */,
  {32'h3eb4e2a8, 32'h00000000} /* (30, 0, 0) {real, imag} */,
  {32'h3f633da2, 32'hbf0edabb} /* (29, 31, 31) {real, imag} */,
  {32'hbedda059, 32'h3efcd1bd} /* (29, 31, 30) {real, imag} */,
  {32'hbd1f1187, 32'hbd48b96c} /* (29, 31, 29) {real, imag} */,
  {32'h3dce8922, 32'h3d983d1f} /* (29, 31, 28) {real, imag} */,
  {32'hbe02820f, 32'h3d727082} /* (29, 31, 27) {real, imag} */,
  {32'hbd3e845c, 32'hbc5c906e} /* (29, 31, 26) {real, imag} */,
  {32'h3cc4cdff, 32'h3d1239f4} /* (29, 31, 25) {real, imag} */,
  {32'hbc539930, 32'h3d17e41a} /* (29, 31, 24) {real, imag} */,
  {32'hbc533b11, 32'hbbb7ef30} /* (29, 31, 23) {real, imag} */,
  {32'h3d8e89b6, 32'h3c33bf8e} /* (29, 31, 22) {real, imag} */,
  {32'h3c922c0a, 32'h3d32f2f3} /* (29, 31, 21) {real, imag} */,
  {32'h3af0ec38, 32'h3c89d654} /* (29, 31, 20) {real, imag} */,
  {32'hbbe06ed4, 32'hbd849464} /* (29, 31, 19) {real, imag} */,
  {32'hbd7d6f68, 32'hbd0aa69b} /* (29, 31, 18) {real, imag} */,
  {32'h3c995092, 32'h3d298370} /* (29, 31, 17) {real, imag} */,
  {32'hbccbbe10, 32'h00000000} /* (29, 31, 16) {real, imag} */,
  {32'h3c995092, 32'hbd298370} /* (29, 31, 15) {real, imag} */,
  {32'hbd7d6f68, 32'h3d0aa69b} /* (29, 31, 14) {real, imag} */,
  {32'hbbe06ed4, 32'h3d849464} /* (29, 31, 13) {real, imag} */,
  {32'h3af0ec38, 32'hbc89d654} /* (29, 31, 12) {real, imag} */,
  {32'h3c922c0a, 32'hbd32f2f3} /* (29, 31, 11) {real, imag} */,
  {32'h3d8e89b6, 32'hbc33bf8e} /* (29, 31, 10) {real, imag} */,
  {32'hbc533b11, 32'h3bb7ef30} /* (29, 31, 9) {real, imag} */,
  {32'hbc539930, 32'hbd17e41a} /* (29, 31, 8) {real, imag} */,
  {32'h3cc4cdff, 32'hbd1239f4} /* (29, 31, 7) {real, imag} */,
  {32'hbd3e845c, 32'h3c5c906e} /* (29, 31, 6) {real, imag} */,
  {32'hbe02820f, 32'hbd727082} /* (29, 31, 5) {real, imag} */,
  {32'h3dce8922, 32'hbd983d1f} /* (29, 31, 4) {real, imag} */,
  {32'hbd1f1187, 32'h3d48b96c} /* (29, 31, 3) {real, imag} */,
  {32'hbedda059, 32'hbefcd1bd} /* (29, 31, 2) {real, imag} */,
  {32'h3f633da2, 32'h3f0edabb} /* (29, 31, 1) {real, imag} */,
  {32'h3ed1a884, 32'h00000000} /* (29, 31, 0) {real, imag} */,
  {32'h3fb3033e, 32'hbedb3d88} /* (29, 30, 31) {real, imag} */,
  {32'hbf4c31f6, 32'h3ef868eb} /* (29, 30, 30) {real, imag} */,
  {32'hbd8609cd, 32'hbc022a70} /* (29, 30, 29) {real, imag} */,
  {32'h3e2d71d0, 32'h3debc1de} /* (29, 30, 28) {real, imag} */,
  {32'hbe301171, 32'h3e2a965e} /* (29, 30, 27) {real, imag} */,
  {32'hbd80d100, 32'hbd14cc8c} /* (29, 30, 26) {real, imag} */,
  {32'h3d758a93, 32'h3cb7dcb0} /* (29, 30, 25) {real, imag} */,
  {32'h3c06d10a, 32'h3dc25920} /* (29, 30, 24) {real, imag} */,
  {32'hbc3979e4, 32'h3ce18d41} /* (29, 30, 23) {real, imag} */,
  {32'h3d8d78e7, 32'hbdaf453f} /* (29, 30, 22) {real, imag} */,
  {32'h3d903195, 32'h3da01d23} /* (29, 30, 21) {real, imag} */,
  {32'h3bf1cc70, 32'h3deca77b} /* (29, 30, 20) {real, imag} */,
  {32'hbd160790, 32'h3da3006c} /* (29, 30, 19) {real, imag} */,
  {32'h3cfc7e2c, 32'h3beaa073} /* (29, 30, 18) {real, imag} */,
  {32'h3c3ae68e, 32'hbd0609ba} /* (29, 30, 17) {real, imag} */,
  {32'hbd339573, 32'h00000000} /* (29, 30, 16) {real, imag} */,
  {32'h3c3ae68e, 32'h3d0609ba} /* (29, 30, 15) {real, imag} */,
  {32'h3cfc7e2c, 32'hbbeaa073} /* (29, 30, 14) {real, imag} */,
  {32'hbd160790, 32'hbda3006c} /* (29, 30, 13) {real, imag} */,
  {32'h3bf1cc70, 32'hbdeca77b} /* (29, 30, 12) {real, imag} */,
  {32'h3d903195, 32'hbda01d23} /* (29, 30, 11) {real, imag} */,
  {32'h3d8d78e7, 32'h3daf453f} /* (29, 30, 10) {real, imag} */,
  {32'hbc3979e4, 32'hbce18d41} /* (29, 30, 9) {real, imag} */,
  {32'h3c06d10a, 32'hbdc25920} /* (29, 30, 8) {real, imag} */,
  {32'h3d758a93, 32'hbcb7dcb0} /* (29, 30, 7) {real, imag} */,
  {32'hbd80d100, 32'h3d14cc8c} /* (29, 30, 6) {real, imag} */,
  {32'hbe301171, 32'hbe2a965e} /* (29, 30, 5) {real, imag} */,
  {32'h3e2d71d0, 32'hbdebc1de} /* (29, 30, 4) {real, imag} */,
  {32'hbd8609cd, 32'h3c022a70} /* (29, 30, 3) {real, imag} */,
  {32'hbf4c31f6, 32'hbef868eb} /* (29, 30, 2) {real, imag} */,
  {32'h3fb3033e, 32'h3edb3d88} /* (29, 30, 1) {real, imag} */,
  {32'h3f369d61, 32'h00000000} /* (29, 30, 0) {real, imag} */,
  {32'h3fd4ee18, 32'hbe891154} /* (29, 29, 31) {real, imag} */,
  {32'hbf895838, 32'h3eae5637} /* (29, 29, 30) {real, imag} */,
  {32'h3b799620, 32'hbd82f6b3} /* (29, 29, 29) {real, imag} */,
  {32'h3e78fd13, 32'h3d40fd9c} /* (29, 29, 28) {real, imag} */,
  {32'hbe63610a, 32'hbdf15cbd} /* (29, 29, 27) {real, imag} */,
  {32'h3d1a293c, 32'hbda2bcc0} /* (29, 29, 26) {real, imag} */,
  {32'hbcc3e5a6, 32'hbd7de5d6} /* (29, 29, 25) {real, imag} */,
  {32'hbc2644de, 32'hbddf3221} /* (29, 29, 24) {real, imag} */,
  {32'hbdaeb6d8, 32'h3da323bf} /* (29, 29, 23) {real, imag} */,
  {32'hbbe503e0, 32'hbe04aeaf} /* (29, 29, 22) {real, imag} */,
  {32'hbd052712, 32'h3ddea344} /* (29, 29, 21) {real, imag} */,
  {32'h3d55115c, 32'hbd188eae} /* (29, 29, 20) {real, imag} */,
  {32'hbe045b94, 32'h3d64c46e} /* (29, 29, 19) {real, imag} */,
  {32'hbc74c3d6, 32'h3dc7260c} /* (29, 29, 18) {real, imag} */,
  {32'h3d1b30ac, 32'hbd905be5} /* (29, 29, 17) {real, imag} */,
  {32'hbdba6b90, 32'h00000000} /* (29, 29, 16) {real, imag} */,
  {32'h3d1b30ac, 32'h3d905be5} /* (29, 29, 15) {real, imag} */,
  {32'hbc74c3d6, 32'hbdc7260c} /* (29, 29, 14) {real, imag} */,
  {32'hbe045b94, 32'hbd64c46e} /* (29, 29, 13) {real, imag} */,
  {32'h3d55115c, 32'h3d188eae} /* (29, 29, 12) {real, imag} */,
  {32'hbd052712, 32'hbddea344} /* (29, 29, 11) {real, imag} */,
  {32'hbbe503e0, 32'h3e04aeaf} /* (29, 29, 10) {real, imag} */,
  {32'hbdaeb6d8, 32'hbda323bf} /* (29, 29, 9) {real, imag} */,
  {32'hbc2644de, 32'h3ddf3221} /* (29, 29, 8) {real, imag} */,
  {32'hbcc3e5a6, 32'h3d7de5d6} /* (29, 29, 7) {real, imag} */,
  {32'h3d1a293c, 32'h3da2bcc0} /* (29, 29, 6) {real, imag} */,
  {32'hbe63610a, 32'h3df15cbd} /* (29, 29, 5) {real, imag} */,
  {32'h3e78fd13, 32'hbd40fd9c} /* (29, 29, 4) {real, imag} */,
  {32'h3b799620, 32'h3d82f6b3} /* (29, 29, 3) {real, imag} */,
  {32'hbf895838, 32'hbeae5637} /* (29, 29, 2) {real, imag} */,
  {32'h3fd4ee18, 32'h3e891154} /* (29, 29, 1) {real, imag} */,
  {32'h3f1d77a4, 32'h00000000} /* (29, 29, 0) {real, imag} */,
  {32'h3fcae112, 32'hbdc14650} /* (29, 28, 31) {real, imag} */,
  {32'hbf8c409c, 32'h3e9a1c8c} /* (29, 28, 30) {real, imag} */,
  {32'hbbacd4a8, 32'hbe834130} /* (29, 28, 29) {real, imag} */,
  {32'h3e593aca, 32'hbd49ae6c} /* (29, 28, 28) {real, imag} */,
  {32'hbe4b8a56, 32'h3dd915de} /* (29, 28, 27) {real, imag} */,
  {32'h3d3b1904, 32'hbd8315fb} /* (29, 28, 26) {real, imag} */,
  {32'hbdce4658, 32'hbd8dde02} /* (29, 28, 25) {real, imag} */,
  {32'hbb9a5af0, 32'h3d3d77fc} /* (29, 28, 24) {real, imag} */,
  {32'h3d45e309, 32'h3d28c204} /* (29, 28, 23) {real, imag} */,
  {32'h3d51e9e6, 32'h3cfdc703} /* (29, 28, 22) {real, imag} */,
  {32'hbcdff779, 32'h3d3f9513} /* (29, 28, 21) {real, imag} */,
  {32'h3d29abab, 32'hbcab110c} /* (29, 28, 20) {real, imag} */,
  {32'h3c43d7f8, 32'hbd692e54} /* (29, 28, 19) {real, imag} */,
  {32'h3db59938, 32'h3d84232b} /* (29, 28, 18) {real, imag} */,
  {32'h3b1dbb22, 32'hbbfc2db6} /* (29, 28, 17) {real, imag} */,
  {32'h3d4ab333, 32'h00000000} /* (29, 28, 16) {real, imag} */,
  {32'h3b1dbb22, 32'h3bfc2db6} /* (29, 28, 15) {real, imag} */,
  {32'h3db59938, 32'hbd84232b} /* (29, 28, 14) {real, imag} */,
  {32'h3c43d7f8, 32'h3d692e54} /* (29, 28, 13) {real, imag} */,
  {32'h3d29abab, 32'h3cab110c} /* (29, 28, 12) {real, imag} */,
  {32'hbcdff779, 32'hbd3f9513} /* (29, 28, 11) {real, imag} */,
  {32'h3d51e9e6, 32'hbcfdc703} /* (29, 28, 10) {real, imag} */,
  {32'h3d45e309, 32'hbd28c204} /* (29, 28, 9) {real, imag} */,
  {32'hbb9a5af0, 32'hbd3d77fc} /* (29, 28, 8) {real, imag} */,
  {32'hbdce4658, 32'h3d8dde02} /* (29, 28, 7) {real, imag} */,
  {32'h3d3b1904, 32'h3d8315fb} /* (29, 28, 6) {real, imag} */,
  {32'hbe4b8a56, 32'hbdd915de} /* (29, 28, 5) {real, imag} */,
  {32'h3e593aca, 32'h3d49ae6c} /* (29, 28, 4) {real, imag} */,
  {32'hbbacd4a8, 32'h3e834130} /* (29, 28, 3) {real, imag} */,
  {32'hbf8c409c, 32'hbe9a1c8c} /* (29, 28, 2) {real, imag} */,
  {32'h3fcae112, 32'h3dc14650} /* (29, 28, 1) {real, imag} */,
  {32'h3f5479fb, 32'h00000000} /* (29, 28, 0) {real, imag} */,
  {32'h3fd16735, 32'h3d6d2620} /* (29, 27, 31) {real, imag} */,
  {32'hbfa09dae, 32'h3e7358dc} /* (29, 27, 30) {real, imag} */,
  {32'hbdbb4225, 32'hbe028a7a} /* (29, 27, 29) {real, imag} */,
  {32'h3e5d8032, 32'hbc3a681e} /* (29, 27, 28) {real, imag} */,
  {32'hbe3a61e6, 32'h3e02d3aa} /* (29, 27, 27) {real, imag} */,
  {32'h3d944ae4, 32'hbd80c477} /* (29, 27, 26) {real, imag} */,
  {32'hbdde821c, 32'hbe069df3} /* (29, 27, 25) {real, imag} */,
  {32'hbd12993e, 32'h3d2e6f80} /* (29, 27, 24) {real, imag} */,
  {32'h3d04f61e, 32'hbd649748} /* (29, 27, 23) {real, imag} */,
  {32'hbc9735e0, 32'hbd9e4387} /* (29, 27, 22) {real, imag} */,
  {32'h3d84f248, 32'h3d94a0fc} /* (29, 27, 21) {real, imag} */,
  {32'h3c2778f4, 32'h3da2c654} /* (29, 27, 20) {real, imag} */,
  {32'h3d84908b, 32'h3d11bc59} /* (29, 27, 19) {real, imag} */,
  {32'hbca36d02, 32'h3c89c72c} /* (29, 27, 18) {real, imag} */,
  {32'hbd63dfdc, 32'h3b03d220} /* (29, 27, 17) {real, imag} */,
  {32'hbd11d460, 32'h00000000} /* (29, 27, 16) {real, imag} */,
  {32'hbd63dfdc, 32'hbb03d220} /* (29, 27, 15) {real, imag} */,
  {32'hbca36d02, 32'hbc89c72c} /* (29, 27, 14) {real, imag} */,
  {32'h3d84908b, 32'hbd11bc59} /* (29, 27, 13) {real, imag} */,
  {32'h3c2778f4, 32'hbda2c654} /* (29, 27, 12) {real, imag} */,
  {32'h3d84f248, 32'hbd94a0fc} /* (29, 27, 11) {real, imag} */,
  {32'hbc9735e0, 32'h3d9e4387} /* (29, 27, 10) {real, imag} */,
  {32'h3d04f61e, 32'h3d649748} /* (29, 27, 9) {real, imag} */,
  {32'hbd12993e, 32'hbd2e6f80} /* (29, 27, 8) {real, imag} */,
  {32'hbdde821c, 32'h3e069df3} /* (29, 27, 7) {real, imag} */,
  {32'h3d944ae4, 32'h3d80c477} /* (29, 27, 6) {real, imag} */,
  {32'hbe3a61e6, 32'hbe02d3aa} /* (29, 27, 5) {real, imag} */,
  {32'h3e5d8032, 32'h3c3a681e} /* (29, 27, 4) {real, imag} */,
  {32'hbdbb4225, 32'h3e028a7a} /* (29, 27, 3) {real, imag} */,
  {32'hbfa09dae, 32'hbe7358dc} /* (29, 27, 2) {real, imag} */,
  {32'h3fd16735, 32'hbd6d2620} /* (29, 27, 1) {real, imag} */,
  {32'h3f85efa3, 32'h00000000} /* (29, 27, 0) {real, imag} */,
  {32'h3fd7a119, 32'hbca3f9c0} /* (29, 26, 31) {real, imag} */,
  {32'hbf94dd02, 32'h3e4da46c} /* (29, 26, 30) {real, imag} */,
  {32'hbd9e90a2, 32'hbd46d657} /* (29, 26, 29) {real, imag} */,
  {32'h3decbf1e, 32'hbb618080} /* (29, 26, 28) {real, imag} */,
  {32'hbe341fac, 32'h3cf79554} /* (29, 26, 27) {real, imag} */,
  {32'hbd11a991, 32'h3ca9cfb4} /* (29, 26, 26) {real, imag} */,
  {32'h3d1beb30, 32'hbd0cc3ce} /* (29, 26, 25) {real, imag} */,
  {32'h3c0173bc, 32'h3c1f7d88} /* (29, 26, 24) {real, imag} */,
  {32'h3d72556f, 32'hbcebb39a} /* (29, 26, 23) {real, imag} */,
  {32'hbc657c1b, 32'h3d038178} /* (29, 26, 22) {real, imag} */,
  {32'h3d919fa4, 32'h3ca86f6a} /* (29, 26, 21) {real, imag} */,
  {32'h3de3bc08, 32'hbc3c74ca} /* (29, 26, 20) {real, imag} */,
  {32'hbcabeb60, 32'hbd0fdb50} /* (29, 26, 19) {real, imag} */,
  {32'hbcf43e4c, 32'h3cc8e4dc} /* (29, 26, 18) {real, imag} */,
  {32'h3c077510, 32'h3cf946a8} /* (29, 26, 17) {real, imag} */,
  {32'hbd9d7199, 32'h00000000} /* (29, 26, 16) {real, imag} */,
  {32'h3c077510, 32'hbcf946a8} /* (29, 26, 15) {real, imag} */,
  {32'hbcf43e4c, 32'hbcc8e4dc} /* (29, 26, 14) {real, imag} */,
  {32'hbcabeb60, 32'h3d0fdb50} /* (29, 26, 13) {real, imag} */,
  {32'h3de3bc08, 32'h3c3c74ca} /* (29, 26, 12) {real, imag} */,
  {32'h3d919fa4, 32'hbca86f6a} /* (29, 26, 11) {real, imag} */,
  {32'hbc657c1b, 32'hbd038178} /* (29, 26, 10) {real, imag} */,
  {32'h3d72556f, 32'h3cebb39a} /* (29, 26, 9) {real, imag} */,
  {32'h3c0173bc, 32'hbc1f7d88} /* (29, 26, 8) {real, imag} */,
  {32'h3d1beb30, 32'h3d0cc3ce} /* (29, 26, 7) {real, imag} */,
  {32'hbd11a991, 32'hbca9cfb4} /* (29, 26, 6) {real, imag} */,
  {32'hbe341fac, 32'hbcf79554} /* (29, 26, 5) {real, imag} */,
  {32'h3decbf1e, 32'h3b618080} /* (29, 26, 4) {real, imag} */,
  {32'hbd9e90a2, 32'h3d46d657} /* (29, 26, 3) {real, imag} */,
  {32'hbf94dd02, 32'hbe4da46c} /* (29, 26, 2) {real, imag} */,
  {32'h3fd7a119, 32'h3ca3f9c0} /* (29, 26, 1) {real, imag} */,
  {32'h3f63d032, 32'h00000000} /* (29, 26, 0) {real, imag} */,
  {32'h3fd39b92, 32'hbdbebe30} /* (29, 25, 31) {real, imag} */,
  {32'hbf9907a6, 32'h3e8ee525} /* (29, 25, 30) {real, imag} */,
  {32'hbdb58dd4, 32'hbe38a05a} /* (29, 25, 29) {real, imag} */,
  {32'h3e217aa6, 32'h3ca941c9} /* (29, 25, 28) {real, imag} */,
  {32'hbe17a475, 32'hbcb42d72} /* (29, 25, 27) {real, imag} */,
  {32'h3cd6dc76, 32'hbbe98078} /* (29, 25, 26) {real, imag} */,
  {32'hbc318340, 32'hbe09a476} /* (29, 25, 25) {real, imag} */,
  {32'h3d82b3e2, 32'h3d895083} /* (29, 25, 24) {real, imag} */,
  {32'hbd864b86, 32'h3d81ca2d} /* (29, 25, 23) {real, imag} */,
  {32'h3d9b7503, 32'hbc291d16} /* (29, 25, 22) {real, imag} */,
  {32'hbc849de0, 32'h3cd92628} /* (29, 25, 21) {real, imag} */,
  {32'hbd335672, 32'h3cbca24e} /* (29, 25, 20) {real, imag} */,
  {32'hbd478944, 32'hbdd120b3} /* (29, 25, 19) {real, imag} */,
  {32'hbc51e9c0, 32'hbc0e3590} /* (29, 25, 18) {real, imag} */,
  {32'h3d05eae3, 32'hbd5efb8c} /* (29, 25, 17) {real, imag} */,
  {32'h3c281a2c, 32'h00000000} /* (29, 25, 16) {real, imag} */,
  {32'h3d05eae3, 32'h3d5efb8c} /* (29, 25, 15) {real, imag} */,
  {32'hbc51e9c0, 32'h3c0e3590} /* (29, 25, 14) {real, imag} */,
  {32'hbd478944, 32'h3dd120b3} /* (29, 25, 13) {real, imag} */,
  {32'hbd335672, 32'hbcbca24e} /* (29, 25, 12) {real, imag} */,
  {32'hbc849de0, 32'hbcd92628} /* (29, 25, 11) {real, imag} */,
  {32'h3d9b7503, 32'h3c291d16} /* (29, 25, 10) {real, imag} */,
  {32'hbd864b86, 32'hbd81ca2d} /* (29, 25, 9) {real, imag} */,
  {32'h3d82b3e2, 32'hbd895083} /* (29, 25, 8) {real, imag} */,
  {32'hbc318340, 32'h3e09a476} /* (29, 25, 7) {real, imag} */,
  {32'h3cd6dc76, 32'h3be98078} /* (29, 25, 6) {real, imag} */,
  {32'hbe17a475, 32'h3cb42d72} /* (29, 25, 5) {real, imag} */,
  {32'h3e217aa6, 32'hbca941c9} /* (29, 25, 4) {real, imag} */,
  {32'hbdb58dd4, 32'h3e38a05a} /* (29, 25, 3) {real, imag} */,
  {32'hbf9907a6, 32'hbe8ee525} /* (29, 25, 2) {real, imag} */,
  {32'h3fd39b92, 32'h3dbebe30} /* (29, 25, 1) {real, imag} */,
  {32'h3f671a75, 32'h00000000} /* (29, 25, 0) {real, imag} */,
  {32'h3fca382e, 32'h3ce47380} /* (29, 24, 31) {real, imag} */,
  {32'hbfa52f32, 32'h3e976100} /* (29, 24, 30) {real, imag} */,
  {32'hbd2cc8f3, 32'h3bd58a56} /* (29, 24, 29) {real, imag} */,
  {32'h3e8a3a4a, 32'hbc9d89b8} /* (29, 24, 28) {real, imag} */,
  {32'hbd460d54, 32'h3d809ee2} /* (29, 24, 27) {real, imag} */,
  {32'hbcda5384, 32'hba89eec0} /* (29, 24, 26) {real, imag} */,
  {32'hbe23501a, 32'hbddc37e4} /* (29, 24, 25) {real, imag} */,
  {32'hbd8a0fa1, 32'h3d4b3c9e} /* (29, 24, 24) {real, imag} */,
  {32'hbcbd8c2f, 32'hbd313d7a} /* (29, 24, 23) {real, imag} */,
  {32'hbaba2580, 32'hbe197aac} /* (29, 24, 22) {real, imag} */,
  {32'hbd034c74, 32'h3d7fcf15} /* (29, 24, 21) {real, imag} */,
  {32'hbcabdd9e, 32'h3ceae93e} /* (29, 24, 20) {real, imag} */,
  {32'h3ca92bd9, 32'h3d303ca8} /* (29, 24, 19) {real, imag} */,
  {32'h3ba76e20, 32'h3d073bd0} /* (29, 24, 18) {real, imag} */,
  {32'h3d83424f, 32'hbd81e2a0} /* (29, 24, 17) {real, imag} */,
  {32'hbc8ff57a, 32'h00000000} /* (29, 24, 16) {real, imag} */,
  {32'h3d83424f, 32'h3d81e2a0} /* (29, 24, 15) {real, imag} */,
  {32'h3ba76e20, 32'hbd073bd0} /* (29, 24, 14) {real, imag} */,
  {32'h3ca92bd9, 32'hbd303ca8} /* (29, 24, 13) {real, imag} */,
  {32'hbcabdd9e, 32'hbceae93e} /* (29, 24, 12) {real, imag} */,
  {32'hbd034c74, 32'hbd7fcf15} /* (29, 24, 11) {real, imag} */,
  {32'hbaba2580, 32'h3e197aac} /* (29, 24, 10) {real, imag} */,
  {32'hbcbd8c2f, 32'h3d313d7a} /* (29, 24, 9) {real, imag} */,
  {32'hbd8a0fa1, 32'hbd4b3c9e} /* (29, 24, 8) {real, imag} */,
  {32'hbe23501a, 32'h3ddc37e4} /* (29, 24, 7) {real, imag} */,
  {32'hbcda5384, 32'h3a89eec0} /* (29, 24, 6) {real, imag} */,
  {32'hbd460d54, 32'hbd809ee2} /* (29, 24, 5) {real, imag} */,
  {32'h3e8a3a4a, 32'h3c9d89b8} /* (29, 24, 4) {real, imag} */,
  {32'hbd2cc8f3, 32'hbbd58a56} /* (29, 24, 3) {real, imag} */,
  {32'hbfa52f32, 32'hbe976100} /* (29, 24, 2) {real, imag} */,
  {32'h3fca382e, 32'hbce47380} /* (29, 24, 1) {real, imag} */,
  {32'h3f8632e0, 32'h00000000} /* (29, 24, 0) {real, imag} */,
  {32'h3fa2ce2a, 32'h3dd7c63c} /* (29, 23, 31) {real, imag} */,
  {32'hbf76a35e, 32'h3e75ead2} /* (29, 23, 30) {real, imag} */,
  {32'hbc96e636, 32'h3d90ad77} /* (29, 23, 29) {real, imag} */,
  {32'h3dee87c6, 32'hbe22ea03} /* (29, 23, 28) {real, imag} */,
  {32'hbda16afa, 32'h3e0b71c6} /* (29, 23, 27) {real, imag} */,
  {32'h3d5b9f75, 32'hbd576fa5} /* (29, 23, 26) {real, imag} */,
  {32'hbe02c16e, 32'hbdf0c9f2} /* (29, 23, 25) {real, imag} */,
  {32'hbc63c4a6, 32'h3c3fe8a2} /* (29, 23, 24) {real, imag} */,
  {32'hbc9a270c, 32'h3d0fd621} /* (29, 23, 23) {real, imag} */,
  {32'h3d64aac4, 32'h3c82b148} /* (29, 23, 22) {real, imag} */,
  {32'h3a34f800, 32'hbdc0c5a9} /* (29, 23, 21) {real, imag} */,
  {32'hbc9aea8a, 32'h3ca1dacc} /* (29, 23, 20) {real, imag} */,
  {32'hbc516b0e, 32'hbb9dc88e} /* (29, 23, 19) {real, imag} */,
  {32'hbdecb644, 32'h3cd9e2c0} /* (29, 23, 18) {real, imag} */,
  {32'h3cacf5ca, 32'hbc7412dc} /* (29, 23, 17) {real, imag} */,
  {32'hbd882122, 32'h00000000} /* (29, 23, 16) {real, imag} */,
  {32'h3cacf5ca, 32'h3c7412dc} /* (29, 23, 15) {real, imag} */,
  {32'hbdecb644, 32'hbcd9e2c0} /* (29, 23, 14) {real, imag} */,
  {32'hbc516b0e, 32'h3b9dc88e} /* (29, 23, 13) {real, imag} */,
  {32'hbc9aea8a, 32'hbca1dacc} /* (29, 23, 12) {real, imag} */,
  {32'h3a34f800, 32'h3dc0c5a9} /* (29, 23, 11) {real, imag} */,
  {32'h3d64aac4, 32'hbc82b148} /* (29, 23, 10) {real, imag} */,
  {32'hbc9a270c, 32'hbd0fd621} /* (29, 23, 9) {real, imag} */,
  {32'hbc63c4a6, 32'hbc3fe8a2} /* (29, 23, 8) {real, imag} */,
  {32'hbe02c16e, 32'h3df0c9f2} /* (29, 23, 7) {real, imag} */,
  {32'h3d5b9f75, 32'h3d576fa5} /* (29, 23, 6) {real, imag} */,
  {32'hbda16afa, 32'hbe0b71c6} /* (29, 23, 5) {real, imag} */,
  {32'h3dee87c6, 32'h3e22ea03} /* (29, 23, 4) {real, imag} */,
  {32'hbc96e636, 32'hbd90ad77} /* (29, 23, 3) {real, imag} */,
  {32'hbf76a35e, 32'hbe75ead2} /* (29, 23, 2) {real, imag} */,
  {32'h3fa2ce2a, 32'hbdd7c63c} /* (29, 23, 1) {real, imag} */,
  {32'h3f5a93b0, 32'h00000000} /* (29, 23, 0) {real, imag} */,
  {32'h3f574720, 32'h3d328392} /* (29, 22, 31) {real, imag} */,
  {32'hbf08deb6, 32'h3ea8a094} /* (29, 22, 30) {real, imag} */,
  {32'h392b3e00, 32'h3dec719f} /* (29, 22, 29) {real, imag} */,
  {32'h3e00d624, 32'hbd2fad4c} /* (29, 22, 28) {real, imag} */,
  {32'hbdd807f5, 32'h3d60a7a9} /* (29, 22, 27) {real, imag} */,
  {32'hbb399d30, 32'h3dc300b4} /* (29, 22, 26) {real, imag} */,
  {32'h3b251a20, 32'hbb09e3a8} /* (29, 22, 25) {real, imag} */,
  {32'hbdcd5bc8, 32'h3c7662d8} /* (29, 22, 24) {real, imag} */,
  {32'h3b71a2d8, 32'h3d6b4bd1} /* (29, 22, 23) {real, imag} */,
  {32'hbc4ef357, 32'hbd4b40e8} /* (29, 22, 22) {real, imag} */,
  {32'hbd51fb5f, 32'hbce07448} /* (29, 22, 21) {real, imag} */,
  {32'h3aebbf80, 32'hbde11e6a} /* (29, 22, 20) {real, imag} */,
  {32'hbd86e720, 32'hbd8d90ce} /* (29, 22, 19) {real, imag} */,
  {32'hbca48168, 32'h3dc72fad} /* (29, 22, 18) {real, imag} */,
  {32'h3b17db72, 32'hbd367810} /* (29, 22, 17) {real, imag} */,
  {32'hbd4700c5, 32'h00000000} /* (29, 22, 16) {real, imag} */,
  {32'h3b17db72, 32'h3d367810} /* (29, 22, 15) {real, imag} */,
  {32'hbca48168, 32'hbdc72fad} /* (29, 22, 14) {real, imag} */,
  {32'hbd86e720, 32'h3d8d90ce} /* (29, 22, 13) {real, imag} */,
  {32'h3aebbf80, 32'h3de11e6a} /* (29, 22, 12) {real, imag} */,
  {32'hbd51fb5f, 32'h3ce07448} /* (29, 22, 11) {real, imag} */,
  {32'hbc4ef357, 32'h3d4b40e8} /* (29, 22, 10) {real, imag} */,
  {32'h3b71a2d8, 32'hbd6b4bd1} /* (29, 22, 9) {real, imag} */,
  {32'hbdcd5bc8, 32'hbc7662d8} /* (29, 22, 8) {real, imag} */,
  {32'h3b251a20, 32'h3b09e3a8} /* (29, 22, 7) {real, imag} */,
  {32'hbb399d30, 32'hbdc300b4} /* (29, 22, 6) {real, imag} */,
  {32'hbdd807f5, 32'hbd60a7a9} /* (29, 22, 5) {real, imag} */,
  {32'h3e00d624, 32'h3d2fad4c} /* (29, 22, 4) {real, imag} */,
  {32'h392b3e00, 32'hbdec719f} /* (29, 22, 3) {real, imag} */,
  {32'hbf08deb6, 32'hbea8a094} /* (29, 22, 2) {real, imag} */,
  {32'h3f574720, 32'hbd328392} /* (29, 22, 1) {real, imag} */,
  {32'h3f3eaf6a, 32'h00000000} /* (29, 22, 0) {real, imag} */,
  {32'h3cedcce0, 32'h3e1c67a9} /* (29, 21, 31) {real, imag} */,
  {32'hbe20d0e2, 32'hbb3c20c0} /* (29, 21, 30) {real, imag} */,
  {32'h3e6c8412, 32'hbcd746be} /* (29, 21, 29) {real, imag} */,
  {32'hbc8f1908, 32'h3d193122} /* (29, 21, 28) {real, imag} */,
  {32'hbd875b40, 32'hbd930abc} /* (29, 21, 27) {real, imag} */,
  {32'hbd7e70d6, 32'h3d904ef3} /* (29, 21, 26) {real, imag} */,
  {32'hbd939a10, 32'hbcfc14c2} /* (29, 21, 25) {real, imag} */,
  {32'h3c6517e8, 32'h3cf0fef2} /* (29, 21, 24) {real, imag} */,
  {32'h3ce11733, 32'hbd372d3e} /* (29, 21, 23) {real, imag} */,
  {32'hbc659659, 32'hba28bfa0} /* (29, 21, 22) {real, imag} */,
  {32'hbd3c7b58, 32'h3dcb9c54} /* (29, 21, 21) {real, imag} */,
  {32'h3ca3a28a, 32'hbc8dee18} /* (29, 21, 20) {real, imag} */,
  {32'h3d051ad1, 32'hbda3b696} /* (29, 21, 19) {real, imag} */,
  {32'h3cbae354, 32'h3c155e1e} /* (29, 21, 18) {real, imag} */,
  {32'hbd382f88, 32'h3d516944} /* (29, 21, 17) {real, imag} */,
  {32'h3cfd2d2c, 32'h00000000} /* (29, 21, 16) {real, imag} */,
  {32'hbd382f88, 32'hbd516944} /* (29, 21, 15) {real, imag} */,
  {32'h3cbae354, 32'hbc155e1e} /* (29, 21, 14) {real, imag} */,
  {32'h3d051ad1, 32'h3da3b696} /* (29, 21, 13) {real, imag} */,
  {32'h3ca3a28a, 32'h3c8dee18} /* (29, 21, 12) {real, imag} */,
  {32'hbd3c7b58, 32'hbdcb9c54} /* (29, 21, 11) {real, imag} */,
  {32'hbc659659, 32'h3a28bfa0} /* (29, 21, 10) {real, imag} */,
  {32'h3ce11733, 32'h3d372d3e} /* (29, 21, 9) {real, imag} */,
  {32'h3c6517e8, 32'hbcf0fef2} /* (29, 21, 8) {real, imag} */,
  {32'hbd939a10, 32'h3cfc14c2} /* (29, 21, 7) {real, imag} */,
  {32'hbd7e70d6, 32'hbd904ef3} /* (29, 21, 6) {real, imag} */,
  {32'hbd875b40, 32'h3d930abc} /* (29, 21, 5) {real, imag} */,
  {32'hbc8f1908, 32'hbd193122} /* (29, 21, 4) {real, imag} */,
  {32'h3e6c8412, 32'h3cd746be} /* (29, 21, 3) {real, imag} */,
  {32'hbe20d0e2, 32'h3b3c20c0} /* (29, 21, 2) {real, imag} */,
  {32'h3cedcce0, 32'hbe1c67a9} /* (29, 21, 1) {real, imag} */,
  {32'h3d02dc38, 32'h00000000} /* (29, 21, 0) {real, imag} */,
  {32'hbf921729, 32'h3e0c3b3a} /* (29, 20, 31) {real, imag} */,
  {32'h3eec5354, 32'hbe522cda} /* (29, 20, 30) {real, imag} */,
  {32'h3e2cda50, 32'hbdba58e0} /* (29, 20, 29) {real, imag} */,
  {32'hbd1d5f46, 32'hbcd47822} /* (29, 20, 28) {real, imag} */,
  {32'h3e266592, 32'hbd65d79c} /* (29, 20, 27) {real, imag} */,
  {32'h3b7e5000, 32'hbd1a5ade} /* (29, 20, 26) {real, imag} */,
  {32'h3d1618da, 32'hbd8f6420} /* (29, 20, 25) {real, imag} */,
  {32'h3d133064, 32'hba5c2700} /* (29, 20, 24) {real, imag} */,
  {32'h3d2b2bfb, 32'h3d9021bc} /* (29, 20, 23) {real, imag} */,
  {32'hbc9a39c0, 32'h3de046b3} /* (29, 20, 22) {real, imag} */,
  {32'hbd029965, 32'h3cae269e} /* (29, 20, 21) {real, imag} */,
  {32'hb909fe00, 32'hbcc88e24} /* (29, 20, 20) {real, imag} */,
  {32'h3c9bbf91, 32'h3c67b07c} /* (29, 20, 19) {real, imag} */,
  {32'h3d4dbbf5, 32'hbd765d52} /* (29, 20, 18) {real, imag} */,
  {32'h3cc686da, 32'hbcd1a30d} /* (29, 20, 17) {real, imag} */,
  {32'h3ccd30f2, 32'h00000000} /* (29, 20, 16) {real, imag} */,
  {32'h3cc686da, 32'h3cd1a30d} /* (29, 20, 15) {real, imag} */,
  {32'h3d4dbbf5, 32'h3d765d52} /* (29, 20, 14) {real, imag} */,
  {32'h3c9bbf91, 32'hbc67b07c} /* (29, 20, 13) {real, imag} */,
  {32'hb909fe00, 32'h3cc88e24} /* (29, 20, 12) {real, imag} */,
  {32'hbd029965, 32'hbcae269e} /* (29, 20, 11) {real, imag} */,
  {32'hbc9a39c0, 32'hbde046b3} /* (29, 20, 10) {real, imag} */,
  {32'h3d2b2bfb, 32'hbd9021bc} /* (29, 20, 9) {real, imag} */,
  {32'h3d133064, 32'h3a5c2700} /* (29, 20, 8) {real, imag} */,
  {32'h3d1618da, 32'h3d8f6420} /* (29, 20, 7) {real, imag} */,
  {32'h3b7e5000, 32'h3d1a5ade} /* (29, 20, 6) {real, imag} */,
  {32'h3e266592, 32'h3d65d79c} /* (29, 20, 5) {real, imag} */,
  {32'hbd1d5f46, 32'h3cd47822} /* (29, 20, 4) {real, imag} */,
  {32'h3e2cda50, 32'h3dba58e0} /* (29, 20, 3) {real, imag} */,
  {32'h3eec5354, 32'h3e522cda} /* (29, 20, 2) {real, imag} */,
  {32'hbf921729, 32'hbe0c3b3a} /* (29, 20, 1) {real, imag} */,
  {32'hbf49d366, 32'h00000000} /* (29, 20, 0) {real, imag} */,
  {32'hbfd9eb0c, 32'h3e1d5264} /* (29, 19, 31) {real, imag} */,
  {32'h3f2a07c0, 32'hbe814b15} /* (29, 19, 30) {real, imag} */,
  {32'h3d1e1a54, 32'h3df68766} /* (29, 19, 29) {real, imag} */,
  {32'hbe6320e5, 32'h3de54c10} /* (29, 19, 28) {real, imag} */,
  {32'h3e56da7e, 32'hbe0d4d4c} /* (29, 19, 27) {real, imag} */,
  {32'h3d1ca7ac, 32'hbd80b600} /* (29, 19, 26) {real, imag} */,
  {32'hbd63fb96, 32'h3cf9396e} /* (29, 19, 25) {real, imag} */,
  {32'h3d712cc2, 32'hbc6f708c} /* (29, 19, 24) {real, imag} */,
  {32'hbd329eb0, 32'hbe1749e8} /* (29, 19, 23) {real, imag} */,
  {32'h3b1a22b8, 32'h3d938346} /* (29, 19, 22) {real, imag} */,
  {32'h3e0f562c, 32'h3d1a3a8c} /* (29, 19, 21) {real, imag} */,
  {32'h3ce9e9e9, 32'h3d9037fa} /* (29, 19, 20) {real, imag} */,
  {32'hbd531efa, 32'h3d5d4500} /* (29, 19, 19) {real, imag} */,
  {32'h3c9cc444, 32'h3db598f3} /* (29, 19, 18) {real, imag} */,
  {32'h3d981289, 32'h3bb46cf6} /* (29, 19, 17) {real, imag} */,
  {32'h3cc193be, 32'h00000000} /* (29, 19, 16) {real, imag} */,
  {32'h3d981289, 32'hbbb46cf6} /* (29, 19, 15) {real, imag} */,
  {32'h3c9cc444, 32'hbdb598f3} /* (29, 19, 14) {real, imag} */,
  {32'hbd531efa, 32'hbd5d4500} /* (29, 19, 13) {real, imag} */,
  {32'h3ce9e9e9, 32'hbd9037fa} /* (29, 19, 12) {real, imag} */,
  {32'h3e0f562c, 32'hbd1a3a8c} /* (29, 19, 11) {real, imag} */,
  {32'h3b1a22b8, 32'hbd938346} /* (29, 19, 10) {real, imag} */,
  {32'hbd329eb0, 32'h3e1749e8} /* (29, 19, 9) {real, imag} */,
  {32'h3d712cc2, 32'h3c6f708c} /* (29, 19, 8) {real, imag} */,
  {32'hbd63fb96, 32'hbcf9396e} /* (29, 19, 7) {real, imag} */,
  {32'h3d1ca7ac, 32'h3d80b600} /* (29, 19, 6) {real, imag} */,
  {32'h3e56da7e, 32'h3e0d4d4c} /* (29, 19, 5) {real, imag} */,
  {32'hbe6320e5, 32'hbde54c10} /* (29, 19, 4) {real, imag} */,
  {32'h3d1e1a54, 32'hbdf68766} /* (29, 19, 3) {real, imag} */,
  {32'h3f2a07c0, 32'h3e814b15} /* (29, 19, 2) {real, imag} */,
  {32'hbfd9eb0c, 32'hbe1d5264} /* (29, 19, 1) {real, imag} */,
  {32'hbf8aba4b, 32'h00000000} /* (29, 19, 0) {real, imag} */,
  {32'hbfff1691, 32'h3e698cbc} /* (29, 18, 31) {real, imag} */,
  {32'h3f524b60, 32'hbe5c0e04} /* (29, 18, 30) {real, imag} */,
  {32'hbdcfa414, 32'hbcb21764} /* (29, 18, 29) {real, imag} */,
  {32'hbe276999, 32'h3d461ce6} /* (29, 18, 28) {real, imag} */,
  {32'h3e8148bd, 32'hbe33965d} /* (29, 18, 27) {real, imag} */,
  {32'hbdae142e, 32'h3cc94320} /* (29, 18, 26) {real, imag} */,
  {32'hbdfac06a, 32'h3dbaf9b0} /* (29, 18, 25) {real, imag} */,
  {32'h3b88b200, 32'hbd620d0a} /* (29, 18, 24) {real, imag} */,
  {32'h3d7fdc7c, 32'h3d3cb5b6} /* (29, 18, 23) {real, imag} */,
  {32'hbdba65b9, 32'hbd0e7a7e} /* (29, 18, 22) {real, imag} */,
  {32'hbd4762b6, 32'h3acf8240} /* (29, 18, 21) {real, imag} */,
  {32'h3d357502, 32'hbd84d870} /* (29, 18, 20) {real, imag} */,
  {32'hbbc1e8d0, 32'h3d3455e2} /* (29, 18, 19) {real, imag} */,
  {32'h3cb7deb6, 32'hbcd5837d} /* (29, 18, 18) {real, imag} */,
  {32'hbd5a8148, 32'h3cd9ca2c} /* (29, 18, 17) {real, imag} */,
  {32'h3d850449, 32'h00000000} /* (29, 18, 16) {real, imag} */,
  {32'hbd5a8148, 32'hbcd9ca2c} /* (29, 18, 15) {real, imag} */,
  {32'h3cb7deb6, 32'h3cd5837d} /* (29, 18, 14) {real, imag} */,
  {32'hbbc1e8d0, 32'hbd3455e2} /* (29, 18, 13) {real, imag} */,
  {32'h3d357502, 32'h3d84d870} /* (29, 18, 12) {real, imag} */,
  {32'hbd4762b6, 32'hbacf8240} /* (29, 18, 11) {real, imag} */,
  {32'hbdba65b9, 32'h3d0e7a7e} /* (29, 18, 10) {real, imag} */,
  {32'h3d7fdc7c, 32'hbd3cb5b6} /* (29, 18, 9) {real, imag} */,
  {32'h3b88b200, 32'h3d620d0a} /* (29, 18, 8) {real, imag} */,
  {32'hbdfac06a, 32'hbdbaf9b0} /* (29, 18, 7) {real, imag} */,
  {32'hbdae142e, 32'hbcc94320} /* (29, 18, 6) {real, imag} */,
  {32'h3e8148bd, 32'h3e33965d} /* (29, 18, 5) {real, imag} */,
  {32'hbe276999, 32'hbd461ce6} /* (29, 18, 4) {real, imag} */,
  {32'hbdcfa414, 32'h3cb21764} /* (29, 18, 3) {real, imag} */,
  {32'h3f524b60, 32'h3e5c0e04} /* (29, 18, 2) {real, imag} */,
  {32'hbfff1691, 32'hbe698cbc} /* (29, 18, 1) {real, imag} */,
  {32'hbfbf409e, 32'h00000000} /* (29, 18, 0) {real, imag} */,
  {32'hc003f884, 32'h3eb51874} /* (29, 17, 31) {real, imag} */,
  {32'h3f7d692d, 32'hbe44ec4e} /* (29, 17, 30) {real, imag} */,
  {32'hbdaedc81, 32'h3dbbf7a3} /* (29, 17, 29) {real, imag} */,
  {32'h3c91df28, 32'h3dd85064} /* (29, 17, 28) {real, imag} */,
  {32'h3e19f445, 32'hbe2464aa} /* (29, 17, 27) {real, imag} */,
  {32'h3ce3fe6c, 32'h3a81e670} /* (29, 17, 26) {real, imag} */,
  {32'h3d81a2ae, 32'h3d9ae334} /* (29, 17, 25) {real, imag} */,
  {32'h3ca97602, 32'h3d3595f7} /* (29, 17, 24) {real, imag} */,
  {32'h3d350ed4, 32'hbc35d736} /* (29, 17, 23) {real, imag} */,
  {32'h3c81ed95, 32'h3b0f8558} /* (29, 17, 22) {real, imag} */,
  {32'h3d21c177, 32'hbdb81252} /* (29, 17, 21) {real, imag} */,
  {32'hbd0b99e2, 32'h3d93ddb6} /* (29, 17, 20) {real, imag} */,
  {32'h3dd8dca8, 32'hbe09088f} /* (29, 17, 19) {real, imag} */,
  {32'hbccd4e51, 32'hbc48631c} /* (29, 17, 18) {real, imag} */,
  {32'hbd1b577e, 32'hbd2bbbfc} /* (29, 17, 17) {real, imag} */,
  {32'hbd9b1c01, 32'h00000000} /* (29, 17, 16) {real, imag} */,
  {32'hbd1b577e, 32'h3d2bbbfc} /* (29, 17, 15) {real, imag} */,
  {32'hbccd4e51, 32'h3c48631c} /* (29, 17, 14) {real, imag} */,
  {32'h3dd8dca8, 32'h3e09088f} /* (29, 17, 13) {real, imag} */,
  {32'hbd0b99e2, 32'hbd93ddb6} /* (29, 17, 12) {real, imag} */,
  {32'h3d21c177, 32'h3db81252} /* (29, 17, 11) {real, imag} */,
  {32'h3c81ed95, 32'hbb0f8558} /* (29, 17, 10) {real, imag} */,
  {32'h3d350ed4, 32'h3c35d736} /* (29, 17, 9) {real, imag} */,
  {32'h3ca97602, 32'hbd3595f7} /* (29, 17, 8) {real, imag} */,
  {32'h3d81a2ae, 32'hbd9ae334} /* (29, 17, 7) {real, imag} */,
  {32'h3ce3fe6c, 32'hba81e670} /* (29, 17, 6) {real, imag} */,
  {32'h3e19f445, 32'h3e2464aa} /* (29, 17, 5) {real, imag} */,
  {32'h3c91df28, 32'hbdd85064} /* (29, 17, 4) {real, imag} */,
  {32'hbdaedc81, 32'hbdbbf7a3} /* (29, 17, 3) {real, imag} */,
  {32'h3f7d692d, 32'h3e44ec4e} /* (29, 17, 2) {real, imag} */,
  {32'hc003f884, 32'hbeb51874} /* (29, 17, 1) {real, imag} */,
  {32'hbfd71924, 32'h00000000} /* (29, 17, 0) {real, imag} */,
  {32'hc0041544, 32'h3e4878c0} /* (29, 16, 31) {real, imag} */,
  {32'h3f80bc8d, 32'hbe548854} /* (29, 16, 30) {real, imag} */,
  {32'hbd5e1ca2, 32'h3d25569a} /* (29, 16, 29) {real, imag} */,
  {32'hbd854d6e, 32'h3d3369f0} /* (29, 16, 28) {real, imag} */,
  {32'h3e04350b, 32'hbd99d78c} /* (29, 16, 27) {real, imag} */,
  {32'h3d552700, 32'hbde97066} /* (29, 16, 26) {real, imag} */,
  {32'hbaceb830, 32'h3d669506} /* (29, 16, 25) {real, imag} */,
  {32'hbc209f8b, 32'hbd1de6b8} /* (29, 16, 24) {real, imag} */,
  {32'hba1413e0, 32'h3d026fe8} /* (29, 16, 23) {real, imag} */,
  {32'h3e0b3037, 32'hbcb84003} /* (29, 16, 22) {real, imag} */,
  {32'h3cd60336, 32'hbdff448b} /* (29, 16, 21) {real, imag} */,
  {32'hbdaf3dfc, 32'hbdb7203a} /* (29, 16, 20) {real, imag} */,
  {32'h3c7a2fa2, 32'hbd7c12fa} /* (29, 16, 19) {real, imag} */,
  {32'h3cb792a0, 32'hbcb4f8db} /* (29, 16, 18) {real, imag} */,
  {32'h3d38eff8, 32'h3d9c1f42} /* (29, 16, 17) {real, imag} */,
  {32'h3ba6d684, 32'h00000000} /* (29, 16, 16) {real, imag} */,
  {32'h3d38eff8, 32'hbd9c1f42} /* (29, 16, 15) {real, imag} */,
  {32'h3cb792a0, 32'h3cb4f8db} /* (29, 16, 14) {real, imag} */,
  {32'h3c7a2fa2, 32'h3d7c12fa} /* (29, 16, 13) {real, imag} */,
  {32'hbdaf3dfc, 32'h3db7203a} /* (29, 16, 12) {real, imag} */,
  {32'h3cd60336, 32'h3dff448b} /* (29, 16, 11) {real, imag} */,
  {32'h3e0b3037, 32'h3cb84003} /* (29, 16, 10) {real, imag} */,
  {32'hba1413e0, 32'hbd026fe8} /* (29, 16, 9) {real, imag} */,
  {32'hbc209f8b, 32'h3d1de6b8} /* (29, 16, 8) {real, imag} */,
  {32'hbaceb830, 32'hbd669506} /* (29, 16, 7) {real, imag} */,
  {32'h3d552700, 32'h3de97066} /* (29, 16, 6) {real, imag} */,
  {32'h3e04350b, 32'h3d99d78c} /* (29, 16, 5) {real, imag} */,
  {32'hbd854d6e, 32'hbd3369f0} /* (29, 16, 4) {real, imag} */,
  {32'hbd5e1ca2, 32'hbd25569a} /* (29, 16, 3) {real, imag} */,
  {32'h3f80bc8d, 32'h3e548854} /* (29, 16, 2) {real, imag} */,
  {32'hc0041544, 32'hbe4878c0} /* (29, 16, 1) {real, imag} */,
  {32'hbfd97e25, 32'h00000000} /* (29, 16, 0) {real, imag} */,
  {32'hbffd72dd, 32'h3cc4a3c8} /* (29, 15, 31) {real, imag} */,
  {32'h3f897c78, 32'hbe680632} /* (29, 15, 30) {real, imag} */,
  {32'h3c8973e8, 32'h3e49abaa} /* (29, 15, 29) {real, imag} */,
  {32'hbe5b1381, 32'h3bf3ace0} /* (29, 15, 28) {real, imag} */,
  {32'h3d8315f8, 32'h3cdb98a0} /* (29, 15, 27) {real, imag} */,
  {32'h3d82dfff, 32'hbd2ad1d0} /* (29, 15, 26) {real, imag} */,
  {32'h3d7488a8, 32'h3c93783e} /* (29, 15, 25) {real, imag} */,
  {32'h3dd5763a, 32'hbd2405ed} /* (29, 15, 24) {real, imag} */,
  {32'hbda2ac9c, 32'h3cff1985} /* (29, 15, 23) {real, imag} */,
  {32'hbc131ba2, 32'hbd7813ce} /* (29, 15, 22) {real, imag} */,
  {32'h3e0740d6, 32'hbc38b7a4} /* (29, 15, 21) {real, imag} */,
  {32'h3c630481, 32'h3c8ee6d0} /* (29, 15, 20) {real, imag} */,
  {32'hbd8780d0, 32'h3d47521c} /* (29, 15, 19) {real, imag} */,
  {32'hbc71944a, 32'hbd7439ef} /* (29, 15, 18) {real, imag} */,
  {32'hbd598598, 32'hbcfd4664} /* (29, 15, 17) {real, imag} */,
  {32'h3dd24b2b, 32'h00000000} /* (29, 15, 16) {real, imag} */,
  {32'hbd598598, 32'h3cfd4664} /* (29, 15, 15) {real, imag} */,
  {32'hbc71944a, 32'h3d7439ef} /* (29, 15, 14) {real, imag} */,
  {32'hbd8780d0, 32'hbd47521c} /* (29, 15, 13) {real, imag} */,
  {32'h3c630481, 32'hbc8ee6d0} /* (29, 15, 12) {real, imag} */,
  {32'h3e0740d6, 32'h3c38b7a4} /* (29, 15, 11) {real, imag} */,
  {32'hbc131ba2, 32'h3d7813ce} /* (29, 15, 10) {real, imag} */,
  {32'hbda2ac9c, 32'hbcff1985} /* (29, 15, 9) {real, imag} */,
  {32'h3dd5763a, 32'h3d2405ed} /* (29, 15, 8) {real, imag} */,
  {32'h3d7488a8, 32'hbc93783e} /* (29, 15, 7) {real, imag} */,
  {32'h3d82dfff, 32'h3d2ad1d0} /* (29, 15, 6) {real, imag} */,
  {32'h3d8315f8, 32'hbcdb98a0} /* (29, 15, 5) {real, imag} */,
  {32'hbe5b1381, 32'hbbf3ace0} /* (29, 15, 4) {real, imag} */,
  {32'h3c8973e8, 32'hbe49abaa} /* (29, 15, 3) {real, imag} */,
  {32'h3f897c78, 32'h3e680632} /* (29, 15, 2) {real, imag} */,
  {32'hbffd72dd, 32'hbcc4a3c8} /* (29, 15, 1) {real, imag} */,
  {32'hbfbe78c8, 32'h00000000} /* (29, 15, 0) {real, imag} */,
  {32'hbff2a10b, 32'h3e129de8} /* (29, 14, 31) {real, imag} */,
  {32'h3f821706, 32'hbe84f118} /* (29, 14, 30) {real, imag} */,
  {32'hbd8a6f42, 32'h3dbdafef} /* (29, 14, 29) {real, imag} */,
  {32'hbe54c12d, 32'h3dfa9a0d} /* (29, 14, 28) {real, imag} */,
  {32'h3e568b3f, 32'h3cf02478} /* (29, 14, 27) {real, imag} */,
  {32'h3e24dd13, 32'hbcb43188} /* (29, 14, 26) {real, imag} */,
  {32'hbd614b94, 32'h3d656fff} /* (29, 14, 25) {real, imag} */,
  {32'h3da4dd22, 32'hbd9649bd} /* (29, 14, 24) {real, imag} */,
  {32'h3d869aea, 32'h3c2624ec} /* (29, 14, 23) {real, imag} */,
  {32'hbd4f489e, 32'h3df094b3} /* (29, 14, 22) {real, imag} */,
  {32'hbd154c8e, 32'hbdba3261} /* (29, 14, 21) {real, imag} */,
  {32'hbdb4cead, 32'h3d227b34} /* (29, 14, 20) {real, imag} */,
  {32'hbdc0f595, 32'h3c7238b6} /* (29, 14, 19) {real, imag} */,
  {32'hbb7bdf34, 32'h3bcb3fac} /* (29, 14, 18) {real, imag} */,
  {32'hbc97ea10, 32'hbdbaaafb} /* (29, 14, 17) {real, imag} */,
  {32'h3d8bd94b, 32'h00000000} /* (29, 14, 16) {real, imag} */,
  {32'hbc97ea10, 32'h3dbaaafb} /* (29, 14, 15) {real, imag} */,
  {32'hbb7bdf34, 32'hbbcb3fac} /* (29, 14, 14) {real, imag} */,
  {32'hbdc0f595, 32'hbc7238b6} /* (29, 14, 13) {real, imag} */,
  {32'hbdb4cead, 32'hbd227b34} /* (29, 14, 12) {real, imag} */,
  {32'hbd154c8e, 32'h3dba3261} /* (29, 14, 11) {real, imag} */,
  {32'hbd4f489e, 32'hbdf094b3} /* (29, 14, 10) {real, imag} */,
  {32'h3d869aea, 32'hbc2624ec} /* (29, 14, 9) {real, imag} */,
  {32'h3da4dd22, 32'h3d9649bd} /* (29, 14, 8) {real, imag} */,
  {32'hbd614b94, 32'hbd656fff} /* (29, 14, 7) {real, imag} */,
  {32'h3e24dd13, 32'h3cb43188} /* (29, 14, 6) {real, imag} */,
  {32'h3e568b3f, 32'hbcf02478} /* (29, 14, 5) {real, imag} */,
  {32'hbe54c12d, 32'hbdfa9a0d} /* (29, 14, 4) {real, imag} */,
  {32'hbd8a6f42, 32'hbdbdafef} /* (29, 14, 3) {real, imag} */,
  {32'h3f821706, 32'h3e84f118} /* (29, 14, 2) {real, imag} */,
  {32'hbff2a10b, 32'hbe129de8} /* (29, 14, 1) {real, imag} */,
  {32'hbfc4df0e, 32'h00000000} /* (29, 14, 0) {real, imag} */,
  {32'hbfe1bee2, 32'h3e2a7014} /* (29, 13, 31) {real, imag} */,
  {32'h3f74df0c, 32'hbe1d230a} /* (29, 13, 30) {real, imag} */,
  {32'hbd42621c, 32'hbd0eb58f} /* (29, 13, 29) {real, imag} */,
  {32'hbe531b27, 32'h3dee22ec} /* (29, 13, 28) {real, imag} */,
  {32'h3e8cd8e1, 32'hbe1775b4} /* (29, 13, 27) {real, imag} */,
  {32'h3de60748, 32'h3de94ffe} /* (29, 13, 26) {real, imag} */,
  {32'hbbb910cc, 32'h3cb1e822} /* (29, 13, 25) {real, imag} */,
  {32'hbc27f05a, 32'hbdd097a4} /* (29, 13, 24) {real, imag} */,
  {32'hbdd76482, 32'h3dc24a86} /* (29, 13, 23) {real, imag} */,
  {32'h3d768b20, 32'h3d2573d9} /* (29, 13, 22) {real, imag} */,
  {32'h3d3a95e7, 32'h3d7d31bc} /* (29, 13, 21) {real, imag} */,
  {32'hbc946cc1, 32'hbc4dfb98} /* (29, 13, 20) {real, imag} */,
  {32'hbd6c3b6e, 32'hbd44a7a4} /* (29, 13, 19) {real, imag} */,
  {32'h3dedca6f, 32'hbd2e1b4a} /* (29, 13, 18) {real, imag} */,
  {32'h3c98163c, 32'hbc54f7c5} /* (29, 13, 17) {real, imag} */,
  {32'hbd684b15, 32'h00000000} /* (29, 13, 16) {real, imag} */,
  {32'h3c98163c, 32'h3c54f7c5} /* (29, 13, 15) {real, imag} */,
  {32'h3dedca6f, 32'h3d2e1b4a} /* (29, 13, 14) {real, imag} */,
  {32'hbd6c3b6e, 32'h3d44a7a4} /* (29, 13, 13) {real, imag} */,
  {32'hbc946cc1, 32'h3c4dfb98} /* (29, 13, 12) {real, imag} */,
  {32'h3d3a95e7, 32'hbd7d31bc} /* (29, 13, 11) {real, imag} */,
  {32'h3d768b20, 32'hbd2573d9} /* (29, 13, 10) {real, imag} */,
  {32'hbdd76482, 32'hbdc24a86} /* (29, 13, 9) {real, imag} */,
  {32'hbc27f05a, 32'h3dd097a4} /* (29, 13, 8) {real, imag} */,
  {32'hbbb910cc, 32'hbcb1e822} /* (29, 13, 7) {real, imag} */,
  {32'h3de60748, 32'hbde94ffe} /* (29, 13, 6) {real, imag} */,
  {32'h3e8cd8e1, 32'h3e1775b4} /* (29, 13, 5) {real, imag} */,
  {32'hbe531b27, 32'hbdee22ec} /* (29, 13, 4) {real, imag} */,
  {32'hbd42621c, 32'h3d0eb58f} /* (29, 13, 3) {real, imag} */,
  {32'h3f74df0c, 32'h3e1d230a} /* (29, 13, 2) {real, imag} */,
  {32'hbfe1bee2, 32'hbe2a7014} /* (29, 13, 1) {real, imag} */,
  {32'hbfc48d93, 32'h00000000} /* (29, 13, 0) {real, imag} */,
  {32'hbfc5a03d, 32'h3dcac73c} /* (29, 12, 31) {real, imag} */,
  {32'h3f38d5ee, 32'hbd685028} /* (29, 12, 30) {real, imag} */,
  {32'h3acb95c0, 32'hbe038b7a} /* (29, 12, 29) {real, imag} */,
  {32'hbe692c0a, 32'h3c2f757c} /* (29, 12, 28) {real, imag} */,
  {32'h3de33637, 32'hbeb4fca4} /* (29, 12, 27) {real, imag} */,
  {32'hbda9d120, 32'hbdc7a309} /* (29, 12, 26) {real, imag} */,
  {32'hbcf2bdc9, 32'hbb7ceff0} /* (29, 12, 25) {real, imag} */,
  {32'hbc8b6f11, 32'hbe2d66a4} /* (29, 12, 24) {real, imag} */,
  {32'h3d64f50d, 32'h3d8342e4} /* (29, 12, 23) {real, imag} */,
  {32'h3e6b550e, 32'h3c994f44} /* (29, 12, 22) {real, imag} */,
  {32'h3d338fbd, 32'hbdaa11c4} /* (29, 12, 21) {real, imag} */,
  {32'h3d1501be, 32'h3c3f134b} /* (29, 12, 20) {real, imag} */,
  {32'hbd835dde, 32'hbd6279a5} /* (29, 12, 19) {real, imag} */,
  {32'h3d2ce591, 32'h3cf763c3} /* (29, 12, 18) {real, imag} */,
  {32'h3ccc9168, 32'h3c9f1cef} /* (29, 12, 17) {real, imag} */,
  {32'h3c34d0e4, 32'h00000000} /* (29, 12, 16) {real, imag} */,
  {32'h3ccc9168, 32'hbc9f1cef} /* (29, 12, 15) {real, imag} */,
  {32'h3d2ce591, 32'hbcf763c3} /* (29, 12, 14) {real, imag} */,
  {32'hbd835dde, 32'h3d6279a5} /* (29, 12, 13) {real, imag} */,
  {32'h3d1501be, 32'hbc3f134b} /* (29, 12, 12) {real, imag} */,
  {32'h3d338fbd, 32'h3daa11c4} /* (29, 12, 11) {real, imag} */,
  {32'h3e6b550e, 32'hbc994f44} /* (29, 12, 10) {real, imag} */,
  {32'h3d64f50d, 32'hbd8342e4} /* (29, 12, 9) {real, imag} */,
  {32'hbc8b6f11, 32'h3e2d66a4} /* (29, 12, 8) {real, imag} */,
  {32'hbcf2bdc9, 32'h3b7ceff0} /* (29, 12, 7) {real, imag} */,
  {32'hbda9d120, 32'h3dc7a309} /* (29, 12, 6) {real, imag} */,
  {32'h3de33637, 32'h3eb4fca4} /* (29, 12, 5) {real, imag} */,
  {32'hbe692c0a, 32'hbc2f757c} /* (29, 12, 4) {real, imag} */,
  {32'h3acb95c0, 32'h3e038b7a} /* (29, 12, 3) {real, imag} */,
  {32'h3f38d5ee, 32'h3d685028} /* (29, 12, 2) {real, imag} */,
  {32'hbfc5a03d, 32'hbdcac73c} /* (29, 12, 1) {real, imag} */,
  {32'hbf959e46, 32'h00000000} /* (29, 12, 0) {real, imag} */,
  {32'hbf5c9a5b, 32'h3d5e8914} /* (29, 11, 31) {real, imag} */,
  {32'h3ed67563, 32'hbc275f50} /* (29, 11, 30) {real, imag} */,
  {32'hbdce521c, 32'hbdbe18e8} /* (29, 11, 29) {real, imag} */,
  {32'hbad27380, 32'hbd9afcc7} /* (29, 11, 28) {real, imag} */,
  {32'h3d2f8fe0, 32'hbeae5b63} /* (29, 11, 27) {real, imag} */,
  {32'hbdc5159d, 32'hbc915984} /* (29, 11, 26) {real, imag} */,
  {32'h3dd2e654, 32'hbd368087} /* (29, 11, 25) {real, imag} */,
  {32'h3d088f16, 32'h3d7f87df} /* (29, 11, 24) {real, imag} */,
  {32'h3d1c0556, 32'h3daf06b1} /* (29, 11, 23) {real, imag} */,
  {32'h3bbc310e, 32'h3a5a7ee0} /* (29, 11, 22) {real, imag} */,
  {32'hbda6e4b6, 32'hbdc42a34} /* (29, 11, 21) {real, imag} */,
  {32'h3bd46518, 32'hbd6cd6ec} /* (29, 11, 20) {real, imag} */,
  {32'hba44dbc0, 32'h3d468b98} /* (29, 11, 19) {real, imag} */,
  {32'hbdbc4313, 32'hbd3345d4} /* (29, 11, 18) {real, imag} */,
  {32'h3bf48468, 32'h3a9ee9f0} /* (29, 11, 17) {real, imag} */,
  {32'h3d725a7c, 32'h00000000} /* (29, 11, 16) {real, imag} */,
  {32'h3bf48468, 32'hba9ee9f0} /* (29, 11, 15) {real, imag} */,
  {32'hbdbc4313, 32'h3d3345d4} /* (29, 11, 14) {real, imag} */,
  {32'hba44dbc0, 32'hbd468b98} /* (29, 11, 13) {real, imag} */,
  {32'h3bd46518, 32'h3d6cd6ec} /* (29, 11, 12) {real, imag} */,
  {32'hbda6e4b6, 32'h3dc42a34} /* (29, 11, 11) {real, imag} */,
  {32'h3bbc310e, 32'hba5a7ee0} /* (29, 11, 10) {real, imag} */,
  {32'h3d1c0556, 32'hbdaf06b1} /* (29, 11, 9) {real, imag} */,
  {32'h3d088f16, 32'hbd7f87df} /* (29, 11, 8) {real, imag} */,
  {32'h3dd2e654, 32'h3d368087} /* (29, 11, 7) {real, imag} */,
  {32'hbdc5159d, 32'h3c915984} /* (29, 11, 6) {real, imag} */,
  {32'h3d2f8fe0, 32'h3eae5b63} /* (29, 11, 5) {real, imag} */,
  {32'hbad27380, 32'h3d9afcc7} /* (29, 11, 4) {real, imag} */,
  {32'hbdce521c, 32'h3dbe18e8} /* (29, 11, 3) {real, imag} */,
  {32'h3ed67563, 32'h3c275f50} /* (29, 11, 2) {real, imag} */,
  {32'hbf5c9a5b, 32'hbd5e8914} /* (29, 11, 1) {real, imag} */,
  {32'hbf5e227c, 32'h00000000} /* (29, 11, 0) {real, imag} */,
  {32'h3f17f932, 32'hbdbe4df5} /* (29, 10, 31) {real, imag} */,
  {32'hbd465698, 32'h3c137100} /* (29, 10, 30) {real, imag} */,
  {32'hbe13365e, 32'h3dbff9c5} /* (29, 10, 29) {real, imag} */,
  {32'h3d12fb08, 32'hbd356436} /* (29, 10, 28) {real, imag} */,
  {32'hbd7351b6, 32'hbc7a8e4c} /* (29, 10, 27) {real, imag} */,
  {32'h3d44b53f, 32'h3b4e57c0} /* (29, 10, 26) {real, imag} */,
  {32'h3dff0a73, 32'h3d6faaca} /* (29, 10, 25) {real, imag} */,
  {32'hbcb5af16, 32'hbd0417e2} /* (29, 10, 24) {real, imag} */,
  {32'h3cdb93dd, 32'h3c8b30e2} /* (29, 10, 23) {real, imag} */,
  {32'hbd054f3f, 32'hbc91e27d} /* (29, 10, 22) {real, imag} */,
  {32'hbe0241d7, 32'h3dc1a84c} /* (29, 10, 21) {real, imag} */,
  {32'h3dff75ac, 32'h3cd13828} /* (29, 10, 20) {real, imag} */,
  {32'h3b8ada70, 32'hbbefa2e4} /* (29, 10, 19) {real, imag} */,
  {32'h3da0a9d1, 32'hbdf7e9f7} /* (29, 10, 18) {real, imag} */,
  {32'h3c164b7a, 32'hbd2d8e20} /* (29, 10, 17) {real, imag} */,
  {32'hbd133327, 32'h00000000} /* (29, 10, 16) {real, imag} */,
  {32'h3c164b7a, 32'h3d2d8e20} /* (29, 10, 15) {real, imag} */,
  {32'h3da0a9d1, 32'h3df7e9f7} /* (29, 10, 14) {real, imag} */,
  {32'h3b8ada70, 32'h3befa2e4} /* (29, 10, 13) {real, imag} */,
  {32'h3dff75ac, 32'hbcd13828} /* (29, 10, 12) {real, imag} */,
  {32'hbe0241d7, 32'hbdc1a84c} /* (29, 10, 11) {real, imag} */,
  {32'hbd054f3f, 32'h3c91e27d} /* (29, 10, 10) {real, imag} */,
  {32'h3cdb93dd, 32'hbc8b30e2} /* (29, 10, 9) {real, imag} */,
  {32'hbcb5af16, 32'h3d0417e2} /* (29, 10, 8) {real, imag} */,
  {32'h3dff0a73, 32'hbd6faaca} /* (29, 10, 7) {real, imag} */,
  {32'h3d44b53f, 32'hbb4e57c0} /* (29, 10, 6) {real, imag} */,
  {32'hbd7351b6, 32'h3c7a8e4c} /* (29, 10, 5) {real, imag} */,
  {32'h3d12fb08, 32'h3d356436} /* (29, 10, 4) {real, imag} */,
  {32'hbe13365e, 32'hbdbff9c5} /* (29, 10, 3) {real, imag} */,
  {32'hbd465698, 32'hbc137100} /* (29, 10, 2) {real, imag} */,
  {32'h3f17f932, 32'h3dbe4df5} /* (29, 10, 1) {real, imag} */,
  {32'h3d98e2d0, 32'h00000000} /* (29, 10, 0) {real, imag} */,
  {32'h3fb6cba4, 32'hbe780ca4} /* (29, 9, 31) {real, imag} */,
  {32'hbedac215, 32'h3e55f0ac} /* (29, 9, 30) {real, imag} */,
  {32'hbde6199e, 32'hbce07478} /* (29, 9, 29) {real, imag} */,
  {32'h3d1daca7, 32'hbdf772ae} /* (29, 9, 28) {real, imag} */,
  {32'hbe6da061, 32'hbcb6d00c} /* (29, 9, 27) {real, imag} */,
  {32'hbe057635, 32'h3ce9fb4e} /* (29, 9, 26) {real, imag} */,
  {32'h3de5a67c, 32'h3b63b7b0} /* (29, 9, 25) {real, imag} */,
  {32'hbd938e4c, 32'h3c85a42d} /* (29, 9, 24) {real, imag} */,
  {32'h3de78151, 32'hbd365637} /* (29, 9, 23) {real, imag} */,
  {32'h3e185995, 32'h3dd3c6e8} /* (29, 9, 22) {real, imag} */,
  {32'hbd7393b0, 32'hbc363bb8} /* (29, 9, 21) {real, imag} */,
  {32'h3d8003e8, 32'h3c8751b0} /* (29, 9, 20) {real, imag} */,
  {32'hbc4ced1e, 32'hbc9d4ca8} /* (29, 9, 19) {real, imag} */,
  {32'h3c85246e, 32'h3c56de11} /* (29, 9, 18) {real, imag} */,
  {32'hbc884052, 32'h3d67b48d} /* (29, 9, 17) {real, imag} */,
  {32'hbc6cbd7c, 32'h00000000} /* (29, 9, 16) {real, imag} */,
  {32'hbc884052, 32'hbd67b48d} /* (29, 9, 15) {real, imag} */,
  {32'h3c85246e, 32'hbc56de11} /* (29, 9, 14) {real, imag} */,
  {32'hbc4ced1e, 32'h3c9d4ca8} /* (29, 9, 13) {real, imag} */,
  {32'h3d8003e8, 32'hbc8751b0} /* (29, 9, 12) {real, imag} */,
  {32'hbd7393b0, 32'h3c363bb8} /* (29, 9, 11) {real, imag} */,
  {32'h3e185995, 32'hbdd3c6e8} /* (29, 9, 10) {real, imag} */,
  {32'h3de78151, 32'h3d365637} /* (29, 9, 9) {real, imag} */,
  {32'hbd938e4c, 32'hbc85a42d} /* (29, 9, 8) {real, imag} */,
  {32'h3de5a67c, 32'hbb63b7b0} /* (29, 9, 7) {real, imag} */,
  {32'hbe057635, 32'hbce9fb4e} /* (29, 9, 6) {real, imag} */,
  {32'hbe6da061, 32'h3cb6d00c} /* (29, 9, 5) {real, imag} */,
  {32'h3d1daca7, 32'h3df772ae} /* (29, 9, 4) {real, imag} */,
  {32'hbde6199e, 32'h3ce07478} /* (29, 9, 3) {real, imag} */,
  {32'hbedac215, 32'hbe55f0ac} /* (29, 9, 2) {real, imag} */,
  {32'h3fb6cba4, 32'h3e780ca4} /* (29, 9, 1) {real, imag} */,
  {32'h3f0cf812, 32'h00000000} /* (29, 9, 0) {real, imag} */,
  {32'h3fcf5a30, 32'hbe859354} /* (29, 8, 31) {real, imag} */,
  {32'hbee9e048, 32'h3eec9c90} /* (29, 8, 30) {real, imag} */,
  {32'h3c3233ec, 32'h3cb93c6e} /* (29, 8, 29) {real, imag} */,
  {32'h3dee2f76, 32'hbdd1f58f} /* (29, 8, 28) {real, imag} */,
  {32'hbe939ab0, 32'h3ba97b78} /* (29, 8, 27) {real, imag} */,
  {32'h3c37edbc, 32'hba8a2b80} /* (29, 8, 26) {real, imag} */,
  {32'hbd3fa0a4, 32'hbde747c4} /* (29, 8, 25) {real, imag} */,
  {32'hbd609657, 32'h3d889d01} /* (29, 8, 24) {real, imag} */,
  {32'hbda6d594, 32'h3dde58d1} /* (29, 8, 23) {real, imag} */,
  {32'h3d2690a5, 32'h3cc7b4f8} /* (29, 8, 22) {real, imag} */,
  {32'h3c82c7f6, 32'h3de2c866} /* (29, 8, 21) {real, imag} */,
  {32'hbd0b5751, 32'hbc3444dc} /* (29, 8, 20) {real, imag} */,
  {32'hbccc2bab, 32'h3d52802c} /* (29, 8, 19) {real, imag} */,
  {32'hbd81180a, 32'hbd0e4df2} /* (29, 8, 18) {real, imag} */,
  {32'hba6b5b80, 32'hbd96ee2e} /* (29, 8, 17) {real, imag} */,
  {32'hbb19040e, 32'h00000000} /* (29, 8, 16) {real, imag} */,
  {32'hba6b5b80, 32'h3d96ee2e} /* (29, 8, 15) {real, imag} */,
  {32'hbd81180a, 32'h3d0e4df2} /* (29, 8, 14) {real, imag} */,
  {32'hbccc2bab, 32'hbd52802c} /* (29, 8, 13) {real, imag} */,
  {32'hbd0b5751, 32'h3c3444dc} /* (29, 8, 12) {real, imag} */,
  {32'h3c82c7f6, 32'hbde2c866} /* (29, 8, 11) {real, imag} */,
  {32'h3d2690a5, 32'hbcc7b4f8} /* (29, 8, 10) {real, imag} */,
  {32'hbda6d594, 32'hbdde58d1} /* (29, 8, 9) {real, imag} */,
  {32'hbd609657, 32'hbd889d01} /* (29, 8, 8) {real, imag} */,
  {32'hbd3fa0a4, 32'h3de747c4} /* (29, 8, 7) {real, imag} */,
  {32'h3c37edbc, 32'h3a8a2b80} /* (29, 8, 6) {real, imag} */,
  {32'hbe939ab0, 32'hbba97b78} /* (29, 8, 5) {real, imag} */,
  {32'h3dee2f76, 32'h3dd1f58f} /* (29, 8, 4) {real, imag} */,
  {32'h3c3233ec, 32'hbcb93c6e} /* (29, 8, 3) {real, imag} */,
  {32'hbee9e048, 32'hbeec9c90} /* (29, 8, 2) {real, imag} */,
  {32'h3fcf5a30, 32'h3e859354} /* (29, 8, 1) {real, imag} */,
  {32'h3f38ab54, 32'h00000000} /* (29, 8, 0) {real, imag} */,
  {32'h3fce65e8, 32'hbe86c533} /* (29, 7, 31) {real, imag} */,
  {32'hbf1c637c, 32'h3edd5147} /* (29, 7, 30) {real, imag} */,
  {32'h3cddcffe, 32'h3e09917a} /* (29, 7, 29) {real, imag} */,
  {32'h3d7ea625, 32'hbd06e6fc} /* (29, 7, 28) {real, imag} */,
  {32'hbe887c0a, 32'h3d943a5a} /* (29, 7, 27) {real, imag} */,
  {32'h3c9a1292, 32'hbddf410a} /* (29, 7, 26) {real, imag} */,
  {32'hbe07c5cc, 32'hbd40baaf} /* (29, 7, 25) {real, imag} */,
  {32'hbcaa381a, 32'h3d8283f9} /* (29, 7, 24) {real, imag} */,
  {32'hbda89a92, 32'h3d50be5e} /* (29, 7, 23) {real, imag} */,
  {32'hbdc77785, 32'hbb9b7a6c} /* (29, 7, 22) {real, imag} */,
  {32'h3dc4c874, 32'h39d5b200} /* (29, 7, 21) {real, imag} */,
  {32'hbcc0fdc4, 32'hbd34e207} /* (29, 7, 20) {real, imag} */,
  {32'h3d7c984e, 32'h3db8f729} /* (29, 7, 19) {real, imag} */,
  {32'hbccdf5d4, 32'hbbc263a3} /* (29, 7, 18) {real, imag} */,
  {32'h3d041ded, 32'hbccf45d4} /* (29, 7, 17) {real, imag} */,
  {32'h3d36b301, 32'h00000000} /* (29, 7, 16) {real, imag} */,
  {32'h3d041ded, 32'h3ccf45d4} /* (29, 7, 15) {real, imag} */,
  {32'hbccdf5d4, 32'h3bc263a3} /* (29, 7, 14) {real, imag} */,
  {32'h3d7c984e, 32'hbdb8f729} /* (29, 7, 13) {real, imag} */,
  {32'hbcc0fdc4, 32'h3d34e207} /* (29, 7, 12) {real, imag} */,
  {32'h3dc4c874, 32'hb9d5b200} /* (29, 7, 11) {real, imag} */,
  {32'hbdc77785, 32'h3b9b7a6c} /* (29, 7, 10) {real, imag} */,
  {32'hbda89a92, 32'hbd50be5e} /* (29, 7, 9) {real, imag} */,
  {32'hbcaa381a, 32'hbd8283f9} /* (29, 7, 8) {real, imag} */,
  {32'hbe07c5cc, 32'h3d40baaf} /* (29, 7, 7) {real, imag} */,
  {32'h3c9a1292, 32'h3ddf410a} /* (29, 7, 6) {real, imag} */,
  {32'hbe887c0a, 32'hbd943a5a} /* (29, 7, 5) {real, imag} */,
  {32'h3d7ea625, 32'h3d06e6fc} /* (29, 7, 4) {real, imag} */,
  {32'h3cddcffe, 32'hbe09917a} /* (29, 7, 3) {real, imag} */,
  {32'hbf1c637c, 32'hbedd5147} /* (29, 7, 2) {real, imag} */,
  {32'h3fce65e8, 32'h3e86c533} /* (29, 7, 1) {real, imag} */,
  {32'h3f495449, 32'h00000000} /* (29, 7, 0) {real, imag} */,
  {32'h3fc74bf7, 32'hbf0713ce} /* (29, 6, 31) {real, imag} */,
  {32'hbefdbe0a, 32'h3f0dd4af} /* (29, 6, 30) {real, imag} */,
  {32'h3c4e2724, 32'h3c5e6594} /* (29, 6, 29) {real, imag} */,
  {32'hba8ed960, 32'hbd164e16} /* (29, 6, 28) {real, imag} */,
  {32'hbdddcdd0, 32'hbcc1af04} /* (29, 6, 27) {real, imag} */,
  {32'hbd8616ae, 32'hbd90a6df} /* (29, 6, 26) {real, imag} */,
  {32'h3d94d9a2, 32'hba034ee0} /* (29, 6, 25) {real, imag} */,
  {32'hbdaca3e2, 32'h3e132e3a} /* (29, 6, 24) {real, imag} */,
  {32'hbd62cd45, 32'hbafc5be0} /* (29, 6, 23) {real, imag} */,
  {32'hbcbf53cc, 32'h3d93779d} /* (29, 6, 22) {real, imag} */,
  {32'hbc3ef64c, 32'h3c3e7620} /* (29, 6, 21) {real, imag} */,
  {32'hbd2f9c34, 32'hbd0640e6} /* (29, 6, 20) {real, imag} */,
  {32'h3badf2c2, 32'hbd975a3e} /* (29, 6, 19) {real, imag} */,
  {32'h3c53edbf, 32'h3d453856} /* (29, 6, 18) {real, imag} */,
  {32'hbc036896, 32'hbc94413e} /* (29, 6, 17) {real, imag} */,
  {32'hbd974b17, 32'h00000000} /* (29, 6, 16) {real, imag} */,
  {32'hbc036896, 32'h3c94413e} /* (29, 6, 15) {real, imag} */,
  {32'h3c53edbf, 32'hbd453856} /* (29, 6, 14) {real, imag} */,
  {32'h3badf2c2, 32'h3d975a3e} /* (29, 6, 13) {real, imag} */,
  {32'hbd2f9c34, 32'h3d0640e6} /* (29, 6, 12) {real, imag} */,
  {32'hbc3ef64c, 32'hbc3e7620} /* (29, 6, 11) {real, imag} */,
  {32'hbcbf53cc, 32'hbd93779d} /* (29, 6, 10) {real, imag} */,
  {32'hbd62cd45, 32'h3afc5be0} /* (29, 6, 9) {real, imag} */,
  {32'hbdaca3e2, 32'hbe132e3a} /* (29, 6, 8) {real, imag} */,
  {32'h3d94d9a2, 32'h3a034ee0} /* (29, 6, 7) {real, imag} */,
  {32'hbd8616ae, 32'h3d90a6df} /* (29, 6, 6) {real, imag} */,
  {32'hbdddcdd0, 32'h3cc1af04} /* (29, 6, 5) {real, imag} */,
  {32'hba8ed960, 32'h3d164e16} /* (29, 6, 4) {real, imag} */,
  {32'h3c4e2724, 32'hbc5e6594} /* (29, 6, 3) {real, imag} */,
  {32'hbefdbe0a, 32'hbf0dd4af} /* (29, 6, 2) {real, imag} */,
  {32'h3fc74bf7, 32'h3f0713ce} /* (29, 6, 1) {real, imag} */,
  {32'h3f3d85ba, 32'h00000000} /* (29, 6, 0) {real, imag} */,
  {32'h3f9f0de9, 32'hbf87b207} /* (29, 5, 31) {real, imag} */,
  {32'hbe0f2fd4, 32'h3f5a93b9} /* (29, 5, 30) {real, imag} */,
  {32'hbd2eefb6, 32'hbd205258} /* (29, 5, 29) {real, imag} */,
  {32'hbd68a38e, 32'hbd2865a4} /* (29, 5, 28) {real, imag} */,
  {32'hbe21dda4, 32'h3da91dd4} /* (29, 5, 27) {real, imag} */,
  {32'hbc9e6b56, 32'hbd974843} /* (29, 5, 26) {real, imag} */,
  {32'hbceacfb0, 32'hbd9f258e} /* (29, 5, 25) {real, imag} */,
  {32'h3d10e8da, 32'h3e33572a} /* (29, 5, 24) {real, imag} */,
  {32'h3d0819ce, 32'h3cb7ea91} /* (29, 5, 23) {real, imag} */,
  {32'h3d2e9d76, 32'h3dea0515} /* (29, 5, 22) {real, imag} */,
  {32'hbd986632, 32'h3d8776d0} /* (29, 5, 21) {real, imag} */,
  {32'hbbc30cc1, 32'hbbd67da0} /* (29, 5, 20) {real, imag} */,
  {32'h3cbfac90, 32'hbd926e98} /* (29, 5, 19) {real, imag} */,
  {32'hbc8aaf10, 32'h3da6bbe9} /* (29, 5, 18) {real, imag} */,
  {32'hbc1d2ac2, 32'hbdb54b1f} /* (29, 5, 17) {real, imag} */,
  {32'h3d6a9a6a, 32'h00000000} /* (29, 5, 16) {real, imag} */,
  {32'hbc1d2ac2, 32'h3db54b1f} /* (29, 5, 15) {real, imag} */,
  {32'hbc8aaf10, 32'hbda6bbe9} /* (29, 5, 14) {real, imag} */,
  {32'h3cbfac90, 32'h3d926e98} /* (29, 5, 13) {real, imag} */,
  {32'hbbc30cc1, 32'h3bd67da0} /* (29, 5, 12) {real, imag} */,
  {32'hbd986632, 32'hbd8776d0} /* (29, 5, 11) {real, imag} */,
  {32'h3d2e9d76, 32'hbdea0515} /* (29, 5, 10) {real, imag} */,
  {32'h3d0819ce, 32'hbcb7ea91} /* (29, 5, 9) {real, imag} */,
  {32'h3d10e8da, 32'hbe33572a} /* (29, 5, 8) {real, imag} */,
  {32'hbceacfb0, 32'h3d9f258e} /* (29, 5, 7) {real, imag} */,
  {32'hbc9e6b56, 32'h3d974843} /* (29, 5, 6) {real, imag} */,
  {32'hbe21dda4, 32'hbda91dd4} /* (29, 5, 5) {real, imag} */,
  {32'hbd68a38e, 32'h3d2865a4} /* (29, 5, 4) {real, imag} */,
  {32'hbd2eefb6, 32'h3d205258} /* (29, 5, 3) {real, imag} */,
  {32'hbe0f2fd4, 32'hbf5a93b9} /* (29, 5, 2) {real, imag} */,
  {32'h3f9f0de9, 32'h3f87b207} /* (29, 5, 1) {real, imag} */,
  {32'h3f6f288e, 32'h00000000} /* (29, 5, 0) {real, imag} */,
  {32'h3f573440, 32'hbfa54443} /* (29, 4, 31) {real, imag} */,
  {32'h3e13c2fa, 32'h3f6ec296} /* (29, 4, 30) {real, imag} */,
  {32'hbdcfc438, 32'hbdbe323e} /* (29, 4, 29) {real, imag} */,
  {32'hbe6d5216, 32'h3e3d0ef1} /* (29, 4, 28) {real, imag} */,
  {32'hbd8dedd0, 32'h3ce86c32} /* (29, 4, 27) {real, imag} */,
  {32'hbd39ec44, 32'hbc5cad26} /* (29, 4, 26) {real, imag} */,
  {32'hbc20f054, 32'hbdbeb622} /* (29, 4, 25) {real, imag} */,
  {32'h3e12e682, 32'h3de559c4} /* (29, 4, 24) {real, imag} */,
  {32'hbd7d7809, 32'hbce70467} /* (29, 4, 23) {real, imag} */,
  {32'hbd4311d4, 32'h3ce2ff79} /* (29, 4, 22) {real, imag} */,
  {32'h3d336cfe, 32'hbd429a93} /* (29, 4, 21) {real, imag} */,
  {32'hbd8ac309, 32'hbd536118} /* (29, 4, 20) {real, imag} */,
  {32'hbd1277e9, 32'h3ac07480} /* (29, 4, 19) {real, imag} */,
  {32'h3d619b3c, 32'hbd9ab4b3} /* (29, 4, 18) {real, imag} */,
  {32'hbb9b2309, 32'hbc86b576} /* (29, 4, 17) {real, imag} */,
  {32'h3d7a0373, 32'h00000000} /* (29, 4, 16) {real, imag} */,
  {32'hbb9b2309, 32'h3c86b576} /* (29, 4, 15) {real, imag} */,
  {32'h3d619b3c, 32'h3d9ab4b3} /* (29, 4, 14) {real, imag} */,
  {32'hbd1277e9, 32'hbac07480} /* (29, 4, 13) {real, imag} */,
  {32'hbd8ac309, 32'h3d536118} /* (29, 4, 12) {real, imag} */,
  {32'h3d336cfe, 32'h3d429a93} /* (29, 4, 11) {real, imag} */,
  {32'hbd4311d4, 32'hbce2ff79} /* (29, 4, 10) {real, imag} */,
  {32'hbd7d7809, 32'h3ce70467} /* (29, 4, 9) {real, imag} */,
  {32'h3e12e682, 32'hbde559c4} /* (29, 4, 8) {real, imag} */,
  {32'hbc20f054, 32'h3dbeb622} /* (29, 4, 7) {real, imag} */,
  {32'hbd39ec44, 32'h3c5cad26} /* (29, 4, 6) {real, imag} */,
  {32'hbd8dedd0, 32'hbce86c32} /* (29, 4, 5) {real, imag} */,
  {32'hbe6d5216, 32'hbe3d0ef1} /* (29, 4, 4) {real, imag} */,
  {32'hbdcfc438, 32'h3dbe323e} /* (29, 4, 3) {real, imag} */,
  {32'h3e13c2fa, 32'hbf6ec296} /* (29, 4, 2) {real, imag} */,
  {32'h3f573440, 32'h3fa54443} /* (29, 4, 1) {real, imag} */,
  {32'h3f563e5f, 32'h00000000} /* (29, 4, 0) {real, imag} */,
  {32'h3f124b7d, 32'hbfab91be} /* (29, 3, 31) {real, imag} */,
  {32'h3e9c16e7, 32'h3f3b3ce8} /* (29, 3, 30) {real, imag} */,
  {32'hbe1372d2, 32'hbdea62d9} /* (29, 3, 29) {real, imag} */,
  {32'hbe0c5b6b, 32'h3e54ffdd} /* (29, 3, 28) {real, imag} */,
  {32'hbdd4f13c, 32'hbd3cdb86} /* (29, 3, 27) {real, imag} */,
  {32'hbd89fd74, 32'h3cd2ec1a} /* (29, 3, 26) {real, imag} */,
  {32'hbd0a3708, 32'hbdddebff} /* (29, 3, 25) {real, imag} */,
  {32'h3d782408, 32'h3d0a26c2} /* (29, 3, 24) {real, imag} */,
  {32'hbc87a258, 32'h3bb3f850} /* (29, 3, 23) {real, imag} */,
  {32'hbb08f890, 32'h3c2357ec} /* (29, 3, 22) {real, imag} */,
  {32'h3d9cd9ea, 32'h3d8cdd34} /* (29, 3, 21) {real, imag} */,
  {32'hbc4bc350, 32'hbd51f9e8} /* (29, 3, 20) {real, imag} */,
  {32'h3d9aae67, 32'hbcb4a864} /* (29, 3, 19) {real, imag} */,
  {32'h3c3e7696, 32'hbd1aab48} /* (29, 3, 18) {real, imag} */,
  {32'h3be5377e, 32'h3c710080} /* (29, 3, 17) {real, imag} */,
  {32'h3c96013e, 32'h00000000} /* (29, 3, 16) {real, imag} */,
  {32'h3be5377e, 32'hbc710080} /* (29, 3, 15) {real, imag} */,
  {32'h3c3e7696, 32'h3d1aab48} /* (29, 3, 14) {real, imag} */,
  {32'h3d9aae67, 32'h3cb4a864} /* (29, 3, 13) {real, imag} */,
  {32'hbc4bc350, 32'h3d51f9e8} /* (29, 3, 12) {real, imag} */,
  {32'h3d9cd9ea, 32'hbd8cdd34} /* (29, 3, 11) {real, imag} */,
  {32'hbb08f890, 32'hbc2357ec} /* (29, 3, 10) {real, imag} */,
  {32'hbc87a258, 32'hbbb3f850} /* (29, 3, 9) {real, imag} */,
  {32'h3d782408, 32'hbd0a26c2} /* (29, 3, 8) {real, imag} */,
  {32'hbd0a3708, 32'h3dddebff} /* (29, 3, 7) {real, imag} */,
  {32'hbd89fd74, 32'hbcd2ec1a} /* (29, 3, 6) {real, imag} */,
  {32'hbdd4f13c, 32'h3d3cdb86} /* (29, 3, 5) {real, imag} */,
  {32'hbe0c5b6b, 32'hbe54ffdd} /* (29, 3, 4) {real, imag} */,
  {32'hbe1372d2, 32'h3dea62d9} /* (29, 3, 3) {real, imag} */,
  {32'h3e9c16e7, 32'hbf3b3ce8} /* (29, 3, 2) {real, imag} */,
  {32'h3f124b7d, 32'h3fab91be} /* (29, 3, 1) {real, imag} */,
  {32'h3f05d4d0, 32'h00000000} /* (29, 3, 0) {real, imag} */,
  {32'h3f0419d1, 32'hbfc10672} /* (29, 2, 31) {real, imag} */,
  {32'h3eb392d4, 32'h3f1a253a} /* (29, 2, 30) {real, imag} */,
  {32'hbd57c5c2, 32'hbdacea4a} /* (29, 2, 29) {real, imag} */,
  {32'hbd9b7680, 32'h3cc925e8} /* (29, 2, 28) {real, imag} */,
  {32'hbe29306f, 32'hbdb2b84b} /* (29, 2, 27) {real, imag} */,
  {32'hbd2404f3, 32'hb92e0800} /* (29, 2, 26) {real, imag} */,
  {32'hbd6c7aa5, 32'hbe43c39a} /* (29, 2, 25) {real, imag} */,
  {32'h3d22c19a, 32'h3d832c82} /* (29, 2, 24) {real, imag} */,
  {32'h3dcf7874, 32'h3d717388} /* (29, 2, 23) {real, imag} */,
  {32'hbd380816, 32'h3d23454e} /* (29, 2, 22) {real, imag} */,
  {32'hbcd779dc, 32'h3cd10745} /* (29, 2, 21) {real, imag} */,
  {32'hbdb23b8f, 32'h3d56749e} /* (29, 2, 20) {real, imag} */,
  {32'h3d1e5708, 32'h3c0a7d74} /* (29, 2, 19) {real, imag} */,
  {32'hbd159988, 32'h3c068504} /* (29, 2, 18) {real, imag} */,
  {32'h3d346dae, 32'h3c84298b} /* (29, 2, 17) {real, imag} */,
  {32'hbcd45f0e, 32'h00000000} /* (29, 2, 16) {real, imag} */,
  {32'h3d346dae, 32'hbc84298b} /* (29, 2, 15) {real, imag} */,
  {32'hbd159988, 32'hbc068504} /* (29, 2, 14) {real, imag} */,
  {32'h3d1e5708, 32'hbc0a7d74} /* (29, 2, 13) {real, imag} */,
  {32'hbdb23b8f, 32'hbd56749e} /* (29, 2, 12) {real, imag} */,
  {32'hbcd779dc, 32'hbcd10745} /* (29, 2, 11) {real, imag} */,
  {32'hbd380816, 32'hbd23454e} /* (29, 2, 10) {real, imag} */,
  {32'h3dcf7874, 32'hbd717388} /* (29, 2, 9) {real, imag} */,
  {32'h3d22c19a, 32'hbd832c82} /* (29, 2, 8) {real, imag} */,
  {32'hbd6c7aa5, 32'h3e43c39a} /* (29, 2, 7) {real, imag} */,
  {32'hbd2404f3, 32'h392e0800} /* (29, 2, 6) {real, imag} */,
  {32'hbe29306f, 32'h3db2b84b} /* (29, 2, 5) {real, imag} */,
  {32'hbd9b7680, 32'hbcc925e8} /* (29, 2, 4) {real, imag} */,
  {32'hbd57c5c2, 32'h3dacea4a} /* (29, 2, 3) {real, imag} */,
  {32'h3eb392d4, 32'hbf1a253a} /* (29, 2, 2) {real, imag} */,
  {32'h3f0419d1, 32'h3fc10672} /* (29, 2, 1) {real, imag} */,
  {32'h3f138b47, 32'h00000000} /* (29, 2, 0) {real, imag} */,
  {32'h3f1234e4, 32'hbfba2d6a} /* (29, 1, 31) {real, imag} */,
  {32'h3e2b0236, 32'h3f4f74c8} /* (29, 1, 30) {real, imag} */,
  {32'hbdeeaf3c, 32'hbcc4da00} /* (29, 1, 29) {real, imag} */,
  {32'hbc4639c8, 32'h3e515804} /* (29, 1, 28) {real, imag} */,
  {32'hbe5d3e6d, 32'hbbca86a4} /* (29, 1, 27) {real, imag} */,
  {32'hbd7586a8, 32'hbc28f706} /* (29, 1, 26) {real, imag} */,
  {32'h3bbc3ee4, 32'hbdc504a2} /* (29, 1, 25) {real, imag} */,
  {32'h3cbb55d0, 32'h3d0a18b6} /* (29, 1, 24) {real, imag} */,
  {32'h3c1b40fb, 32'hbdfd6545} /* (29, 1, 23) {real, imag} */,
  {32'h3c615976, 32'h3d09bb94} /* (29, 1, 22) {real, imag} */,
  {32'hbd35f841, 32'h3c41f784} /* (29, 1, 21) {real, imag} */,
  {32'hbd02de0c, 32'hbd66132a} /* (29, 1, 20) {real, imag} */,
  {32'h3c8d4537, 32'h3d1c9cbe} /* (29, 1, 19) {real, imag} */,
  {32'hbd2eba58, 32'h3d06b5dd} /* (29, 1, 18) {real, imag} */,
  {32'h3c46fb1e, 32'h3cac45d2} /* (29, 1, 17) {real, imag} */,
  {32'h3cebf630, 32'h00000000} /* (29, 1, 16) {real, imag} */,
  {32'h3c46fb1e, 32'hbcac45d2} /* (29, 1, 15) {real, imag} */,
  {32'hbd2eba58, 32'hbd06b5dd} /* (29, 1, 14) {real, imag} */,
  {32'h3c8d4537, 32'hbd1c9cbe} /* (29, 1, 13) {real, imag} */,
  {32'hbd02de0c, 32'h3d66132a} /* (29, 1, 12) {real, imag} */,
  {32'hbd35f841, 32'hbc41f784} /* (29, 1, 11) {real, imag} */,
  {32'h3c615976, 32'hbd09bb94} /* (29, 1, 10) {real, imag} */,
  {32'h3c1b40fb, 32'h3dfd6545} /* (29, 1, 9) {real, imag} */,
  {32'h3cbb55d0, 32'hbd0a18b6} /* (29, 1, 8) {real, imag} */,
  {32'h3bbc3ee4, 32'h3dc504a2} /* (29, 1, 7) {real, imag} */,
  {32'hbd7586a8, 32'h3c28f706} /* (29, 1, 6) {real, imag} */,
  {32'hbe5d3e6d, 32'h3bca86a4} /* (29, 1, 5) {real, imag} */,
  {32'hbc4639c8, 32'hbe515804} /* (29, 1, 4) {real, imag} */,
  {32'hbdeeaf3c, 32'h3cc4da00} /* (29, 1, 3) {real, imag} */,
  {32'h3e2b0236, 32'hbf4f74c8} /* (29, 1, 2) {real, imag} */,
  {32'h3f1234e4, 32'h3fba2d6a} /* (29, 1, 1) {real, imag} */,
  {32'h3f178606, 32'h00000000} /* (29, 1, 0) {real, imag} */,
  {32'h3f19a5fe, 32'hbf7400e8} /* (29, 0, 31) {real, imag} */,
  {32'hbc277780, 32'h3f356381} /* (29, 0, 30) {real, imag} */,
  {32'hbdaa0c03, 32'hbd17d734} /* (29, 0, 29) {real, imag} */,
  {32'h3cc618c6, 32'h3e268a50} /* (29, 0, 28) {real, imag} */,
  {32'hbe603c91, 32'hbd3122e1} /* (29, 0, 27) {real, imag} */,
  {32'hbd08921e, 32'hbc75c1b0} /* (29, 0, 26) {real, imag} */,
  {32'hbced9c25, 32'h3c87d9a1} /* (29, 0, 25) {real, imag} */,
  {32'hbc695899, 32'h3ce4369b} /* (29, 0, 24) {real, imag} */,
  {32'h3c263f42, 32'h3cdc6545} /* (29, 0, 23) {real, imag} */,
  {32'hbdbbab87, 32'h3d43c606} /* (29, 0, 22) {real, imag} */,
  {32'h3d133345, 32'hbd78b0e2} /* (29, 0, 21) {real, imag} */,
  {32'h3cc04872, 32'hbd5b5933} /* (29, 0, 20) {real, imag} */,
  {32'h3d98dd8c, 32'h3c950579} /* (29, 0, 19) {real, imag} */,
  {32'h3d401740, 32'h3cbc0b2d} /* (29, 0, 18) {real, imag} */,
  {32'hbcff4dc0, 32'hbc332040} /* (29, 0, 17) {real, imag} */,
  {32'h3b64ccd8, 32'h00000000} /* (29, 0, 16) {real, imag} */,
  {32'hbcff4dc0, 32'h3c332040} /* (29, 0, 15) {real, imag} */,
  {32'h3d401740, 32'hbcbc0b2d} /* (29, 0, 14) {real, imag} */,
  {32'h3d98dd8c, 32'hbc950579} /* (29, 0, 13) {real, imag} */,
  {32'h3cc04872, 32'h3d5b5933} /* (29, 0, 12) {real, imag} */,
  {32'h3d133345, 32'h3d78b0e2} /* (29, 0, 11) {real, imag} */,
  {32'hbdbbab87, 32'hbd43c606} /* (29, 0, 10) {real, imag} */,
  {32'h3c263f42, 32'hbcdc6545} /* (29, 0, 9) {real, imag} */,
  {32'hbc695899, 32'hbce4369b} /* (29, 0, 8) {real, imag} */,
  {32'hbced9c25, 32'hbc87d9a1} /* (29, 0, 7) {real, imag} */,
  {32'hbd08921e, 32'h3c75c1b0} /* (29, 0, 6) {real, imag} */,
  {32'hbe603c91, 32'h3d3122e1} /* (29, 0, 5) {real, imag} */,
  {32'h3cc618c6, 32'hbe268a50} /* (29, 0, 4) {real, imag} */,
  {32'hbdaa0c03, 32'h3d17d734} /* (29, 0, 3) {real, imag} */,
  {32'hbc277780, 32'hbf356381} /* (29, 0, 2) {real, imag} */,
  {32'h3f19a5fe, 32'h3f7400e8} /* (29, 0, 1) {real, imag} */,
  {32'h3ecdc3cc, 32'h00000000} /* (29, 0, 0) {real, imag} */,
  {32'h3f365d3a, 32'hbed04c52} /* (28, 31, 31) {real, imag} */,
  {32'hbeed51db, 32'h3eff2a52} /* (28, 31, 30) {real, imag} */,
  {32'hbde344e0, 32'h3ba517b4} /* (28, 31, 29) {real, imag} */,
  {32'h3d6dc76f, 32'h3e48ef09} /* (28, 31, 28) {real, imag} */,
  {32'hbe006a4f, 32'h3dd86c26} /* (28, 31, 27) {real, imag} */,
  {32'h3cd01ff7, 32'hbc6f4618} /* (28, 31, 26) {real, imag} */,
  {32'h3cbd2b9a, 32'hbd165512} /* (28, 31, 25) {real, imag} */,
  {32'hbd30b255, 32'hbc5702a4} /* (28, 31, 24) {real, imag} */,
  {32'h3c47ec46, 32'h3d7284db} /* (28, 31, 23) {real, imag} */,
  {32'hbc424d2c, 32'h3bd62734} /* (28, 31, 22) {real, imag} */,
  {32'hbd310634, 32'hbc00ae6a} /* (28, 31, 21) {real, imag} */,
  {32'hbcb7a544, 32'hbd396a37} /* (28, 31, 20) {real, imag} */,
  {32'hbd85b1f6, 32'hbd0801f3} /* (28, 31, 19) {real, imag} */,
  {32'h3c388db2, 32'hbc86a1d0} /* (28, 31, 18) {real, imag} */,
  {32'hbb4128ec, 32'h3c202cb8} /* (28, 31, 17) {real, imag} */,
  {32'h3c0c0fca, 32'h00000000} /* (28, 31, 16) {real, imag} */,
  {32'hbb4128ec, 32'hbc202cb8} /* (28, 31, 15) {real, imag} */,
  {32'h3c388db2, 32'h3c86a1d0} /* (28, 31, 14) {real, imag} */,
  {32'hbd85b1f6, 32'h3d0801f3} /* (28, 31, 13) {real, imag} */,
  {32'hbcb7a544, 32'h3d396a37} /* (28, 31, 12) {real, imag} */,
  {32'hbd310634, 32'h3c00ae6a} /* (28, 31, 11) {real, imag} */,
  {32'hbc424d2c, 32'hbbd62734} /* (28, 31, 10) {real, imag} */,
  {32'h3c47ec46, 32'hbd7284db} /* (28, 31, 9) {real, imag} */,
  {32'hbd30b255, 32'h3c5702a4} /* (28, 31, 8) {real, imag} */,
  {32'h3cbd2b9a, 32'h3d165512} /* (28, 31, 7) {real, imag} */,
  {32'h3cd01ff7, 32'h3c6f4618} /* (28, 31, 6) {real, imag} */,
  {32'hbe006a4f, 32'hbdd86c26} /* (28, 31, 5) {real, imag} */,
  {32'h3d6dc76f, 32'hbe48ef09} /* (28, 31, 4) {real, imag} */,
  {32'hbde344e0, 32'hbba517b4} /* (28, 31, 3) {real, imag} */,
  {32'hbeed51db, 32'hbeff2a52} /* (28, 31, 2) {real, imag} */,
  {32'h3f365d3a, 32'h3ed04c52} /* (28, 31, 1) {real, imag} */,
  {32'h3de55e54, 32'h00000000} /* (28, 31, 0) {real, imag} */,
  {32'h3f970e2d, 32'hbe751170} /* (28, 30, 31) {real, imag} */,
  {32'hbf71707f, 32'h3eeb0c90} /* (28, 30, 30) {real, imag} */,
  {32'hbe0154de, 32'h3c6e37d0} /* (28, 30, 29) {real, imag} */,
  {32'h3de7afda, 32'h3de3e924} /* (28, 30, 28) {real, imag} */,
  {32'hbe29f685, 32'h3e159042} /* (28, 30, 27) {real, imag} */,
  {32'hbd12c3a4, 32'hbdf489c0} /* (28, 30, 26) {real, imag} */,
  {32'h3da747a1, 32'hbd8b2e10} /* (28, 30, 25) {real, imag} */,
  {32'h3caa7eb4, 32'hbd8c4eec} /* (28, 30, 24) {real, imag} */,
  {32'hbd158316, 32'hbcca23c8} /* (28, 30, 23) {real, imag} */,
  {32'h3d4c84a2, 32'hbcde2418} /* (28, 30, 22) {real, imag} */,
  {32'hbd7214d0, 32'h3da7e5f9} /* (28, 30, 21) {real, imag} */,
  {32'hbd11d6d7, 32'hbd1021c0} /* (28, 30, 20) {real, imag} */,
  {32'hbd787619, 32'hbd35b981} /* (28, 30, 19) {real, imag} */,
  {32'h3cf1d281, 32'hbcc06b03} /* (28, 30, 18) {real, imag} */,
  {32'h3b62c900, 32'h3d0bf806} /* (28, 30, 17) {real, imag} */,
  {32'hbdae478b, 32'h00000000} /* (28, 30, 16) {real, imag} */,
  {32'h3b62c900, 32'hbd0bf806} /* (28, 30, 15) {real, imag} */,
  {32'h3cf1d281, 32'h3cc06b03} /* (28, 30, 14) {real, imag} */,
  {32'hbd787619, 32'h3d35b981} /* (28, 30, 13) {real, imag} */,
  {32'hbd11d6d7, 32'h3d1021c0} /* (28, 30, 12) {real, imag} */,
  {32'hbd7214d0, 32'hbda7e5f9} /* (28, 30, 11) {real, imag} */,
  {32'h3d4c84a2, 32'h3cde2418} /* (28, 30, 10) {real, imag} */,
  {32'hbd158316, 32'h3cca23c8} /* (28, 30, 9) {real, imag} */,
  {32'h3caa7eb4, 32'h3d8c4eec} /* (28, 30, 8) {real, imag} */,
  {32'h3da747a1, 32'h3d8b2e10} /* (28, 30, 7) {real, imag} */,
  {32'hbd12c3a4, 32'h3df489c0} /* (28, 30, 6) {real, imag} */,
  {32'hbe29f685, 32'hbe159042} /* (28, 30, 5) {real, imag} */,
  {32'h3de7afda, 32'hbde3e924} /* (28, 30, 4) {real, imag} */,
  {32'hbe0154de, 32'hbc6e37d0} /* (28, 30, 3) {real, imag} */,
  {32'hbf71707f, 32'hbeeb0c90} /* (28, 30, 2) {real, imag} */,
  {32'h3f970e2d, 32'h3e751170} /* (28, 30, 1) {real, imag} */,
  {32'h3e8abf02, 32'h00000000} /* (28, 30, 0) {real, imag} */,
  {32'h3fbace3e, 32'hbd95bae8} /* (28, 29, 31) {real, imag} */,
  {32'hbf82b72c, 32'h3e8116ed} /* (28, 29, 30) {real, imag} */,
  {32'hbe159429, 32'h3cceff40} /* (28, 29, 29) {real, imag} */,
  {32'h3e05689a, 32'h3c16ec80} /* (28, 29, 28) {real, imag} */,
  {32'hbe699dde, 32'h3c4dc170} /* (28, 29, 27) {real, imag} */,
  {32'h3b9da244, 32'hbbd54790} /* (28, 29, 26) {real, imag} */,
  {32'hbcf50dc4, 32'hbd5bcbb0} /* (28, 29, 25) {real, imag} */,
  {32'hbd50ce82, 32'h3d1e8fc9} /* (28, 29, 24) {real, imag} */,
  {32'h3dd546cb, 32'hbd4c2ed6} /* (28, 29, 23) {real, imag} */,
  {32'h3cb80fda, 32'hbda7d6c7} /* (28, 29, 22) {real, imag} */,
  {32'hbd929944, 32'h3b37b300} /* (28, 29, 21) {real, imag} */,
  {32'hbdc4aaa2, 32'hbd2029ea} /* (28, 29, 20) {real, imag} */,
  {32'h3d23aa9c, 32'h3d740d03} /* (28, 29, 19) {real, imag} */,
  {32'hba4ee1c0, 32'hbc79ef3e} /* (28, 29, 18) {real, imag} */,
  {32'h3d2d971b, 32'h3c0845de} /* (28, 29, 17) {real, imag} */,
  {32'hbc2b3414, 32'h00000000} /* (28, 29, 16) {real, imag} */,
  {32'h3d2d971b, 32'hbc0845de} /* (28, 29, 15) {real, imag} */,
  {32'hba4ee1c0, 32'h3c79ef3e} /* (28, 29, 14) {real, imag} */,
  {32'h3d23aa9c, 32'hbd740d03} /* (28, 29, 13) {real, imag} */,
  {32'hbdc4aaa2, 32'h3d2029ea} /* (28, 29, 12) {real, imag} */,
  {32'hbd929944, 32'hbb37b300} /* (28, 29, 11) {real, imag} */,
  {32'h3cb80fda, 32'h3da7d6c7} /* (28, 29, 10) {real, imag} */,
  {32'h3dd546cb, 32'h3d4c2ed6} /* (28, 29, 9) {real, imag} */,
  {32'hbd50ce82, 32'hbd1e8fc9} /* (28, 29, 8) {real, imag} */,
  {32'hbcf50dc4, 32'h3d5bcbb0} /* (28, 29, 7) {real, imag} */,
  {32'h3b9da244, 32'h3bd54790} /* (28, 29, 6) {real, imag} */,
  {32'hbe699dde, 32'hbc4dc170} /* (28, 29, 5) {real, imag} */,
  {32'h3e05689a, 32'hbc16ec80} /* (28, 29, 4) {real, imag} */,
  {32'hbe159429, 32'hbcceff40} /* (28, 29, 3) {real, imag} */,
  {32'hbf82b72c, 32'hbe8116ed} /* (28, 29, 2) {real, imag} */,
  {32'h3fbace3e, 32'h3d95bae8} /* (28, 29, 1) {real, imag} */,
  {32'h3e649846, 32'h00000000} /* (28, 29, 0) {real, imag} */,
  {32'h3fbd3a62, 32'h3dad5c70} /* (28, 28, 31) {real, imag} */,
  {32'hbf9992ce, 32'h3e875e6e} /* (28, 28, 30) {real, imag} */,
  {32'hbd0ad1cf, 32'hbcb38dab} /* (28, 28, 29) {real, imag} */,
  {32'h3e113822, 32'hbd12c5dd} /* (28, 28, 28) {real, imag} */,
  {32'hbebcc3a6, 32'h3e1b1a43} /* (28, 28, 27) {real, imag} */,
  {32'h3cc67a8f, 32'hbd2c89c6} /* (28, 28, 26) {real, imag} */,
  {32'h3c89c07c, 32'hbdfcb1ab} /* (28, 28, 25) {real, imag} */,
  {32'hbd74a0a9, 32'h3db9f786} /* (28, 28, 24) {real, imag} */,
  {32'h3d785214, 32'hbd4578c6} /* (28, 28, 23) {real, imag} */,
  {32'h3cee89ba, 32'hbda6b48c} /* (28, 28, 22) {real, imag} */,
  {32'hbc696f60, 32'h3d89276f} /* (28, 28, 21) {real, imag} */,
  {32'hbcff94a5, 32'hbddd5d4c} /* (28, 28, 20) {real, imag} */,
  {32'hbd45e0be, 32'h3d77b96a} /* (28, 28, 19) {real, imag} */,
  {32'hbc21c348, 32'hbd204c2c} /* (28, 28, 18) {real, imag} */,
  {32'h3c900398, 32'h3cf615e0} /* (28, 28, 17) {real, imag} */,
  {32'h3ddb37de, 32'h00000000} /* (28, 28, 16) {real, imag} */,
  {32'h3c900398, 32'hbcf615e0} /* (28, 28, 15) {real, imag} */,
  {32'hbc21c348, 32'h3d204c2c} /* (28, 28, 14) {real, imag} */,
  {32'hbd45e0be, 32'hbd77b96a} /* (28, 28, 13) {real, imag} */,
  {32'hbcff94a5, 32'h3ddd5d4c} /* (28, 28, 12) {real, imag} */,
  {32'hbc696f60, 32'hbd89276f} /* (28, 28, 11) {real, imag} */,
  {32'h3cee89ba, 32'h3da6b48c} /* (28, 28, 10) {real, imag} */,
  {32'h3d785214, 32'h3d4578c6} /* (28, 28, 9) {real, imag} */,
  {32'hbd74a0a9, 32'hbdb9f786} /* (28, 28, 8) {real, imag} */,
  {32'h3c89c07c, 32'h3dfcb1ab} /* (28, 28, 7) {real, imag} */,
  {32'h3cc67a8f, 32'h3d2c89c6} /* (28, 28, 6) {real, imag} */,
  {32'hbebcc3a6, 32'hbe1b1a43} /* (28, 28, 5) {real, imag} */,
  {32'h3e113822, 32'h3d12c5dd} /* (28, 28, 4) {real, imag} */,
  {32'hbd0ad1cf, 32'h3cb38dab} /* (28, 28, 3) {real, imag} */,
  {32'hbf9992ce, 32'hbe875e6e} /* (28, 28, 2) {real, imag} */,
  {32'h3fbd3a62, 32'hbdad5c70} /* (28, 28, 1) {real, imag} */,
  {32'h3ee008e2, 32'h00000000} /* (28, 28, 0) {real, imag} */,
  {32'h3fb65eea, 32'h3e37d9b4} /* (28, 27, 31) {real, imag} */,
  {32'hbf91c7cc, 32'h3e96959a} /* (28, 27, 30) {real, imag} */,
  {32'hbc664230, 32'hbe3e2028} /* (28, 27, 29) {real, imag} */,
  {32'h3d858894, 32'hbe051ef8} /* (28, 27, 28) {real, imag} */,
  {32'hbe810036, 32'h3e3e6510} /* (28, 27, 27) {real, imag} */,
  {32'hbd0f5cfd, 32'hbc760ba8} /* (28, 27, 26) {real, imag} */,
  {32'h3c8ffcd2, 32'hba3db280} /* (28, 27, 25) {real, imag} */,
  {32'hbd64692e, 32'h3e230d8c} /* (28, 27, 24) {real, imag} */,
  {32'h3d841df4, 32'hbcbf6d7e} /* (28, 27, 23) {real, imag} */,
  {32'hbd2d19f8, 32'hbcc545a8} /* (28, 27, 22) {real, imag} */,
  {32'hbd81d7c4, 32'h3d200be0} /* (28, 27, 21) {real, imag} */,
  {32'hbc3ced18, 32'hbd917de4} /* (28, 27, 20) {real, imag} */,
  {32'h3d94d56c, 32'hbe11a7f0} /* (28, 27, 19) {real, imag} */,
  {32'h3c2b18f0, 32'h3d3ffa5c} /* (28, 27, 18) {real, imag} */,
  {32'h3d78c4ae, 32'h3da0fad3} /* (28, 27, 17) {real, imag} */,
  {32'hbdb99a08, 32'h00000000} /* (28, 27, 16) {real, imag} */,
  {32'h3d78c4ae, 32'hbda0fad3} /* (28, 27, 15) {real, imag} */,
  {32'h3c2b18f0, 32'hbd3ffa5c} /* (28, 27, 14) {real, imag} */,
  {32'h3d94d56c, 32'h3e11a7f0} /* (28, 27, 13) {real, imag} */,
  {32'hbc3ced18, 32'h3d917de4} /* (28, 27, 12) {real, imag} */,
  {32'hbd81d7c4, 32'hbd200be0} /* (28, 27, 11) {real, imag} */,
  {32'hbd2d19f8, 32'h3cc545a8} /* (28, 27, 10) {real, imag} */,
  {32'h3d841df4, 32'h3cbf6d7e} /* (28, 27, 9) {real, imag} */,
  {32'hbd64692e, 32'hbe230d8c} /* (28, 27, 8) {real, imag} */,
  {32'h3c8ffcd2, 32'h3a3db280} /* (28, 27, 7) {real, imag} */,
  {32'hbd0f5cfd, 32'h3c760ba8} /* (28, 27, 6) {real, imag} */,
  {32'hbe810036, 32'hbe3e6510} /* (28, 27, 5) {real, imag} */,
  {32'h3d858894, 32'h3e051ef8} /* (28, 27, 4) {real, imag} */,
  {32'hbc664230, 32'h3e3e2028} /* (28, 27, 3) {real, imag} */,
  {32'hbf91c7cc, 32'hbe96959a} /* (28, 27, 2) {real, imag} */,
  {32'h3fb65eea, 32'hbe37d9b4} /* (28, 27, 1) {real, imag} */,
  {32'h3f1befb2, 32'h00000000} /* (28, 27, 0) {real, imag} */,
  {32'h3fb1e26b, 32'h3dc7159c} /* (28, 26, 31) {real, imag} */,
  {32'hbf95b62c, 32'h3e7096b4} /* (28, 26, 30) {real, imag} */,
  {32'h3d96bfd2, 32'hbd3aad6a} /* (28, 26, 29) {real, imag} */,
  {32'h3e3a51be, 32'hbdca576c} /* (28, 26, 28) {real, imag} */,
  {32'hbdb4361e, 32'h3e45a722} /* (28, 26, 27) {real, imag} */,
  {32'hbc33e4a4, 32'hbd307a98} /* (28, 26, 26) {real, imag} */,
  {32'h3dad4a9e, 32'hbdf2b5d8} /* (28, 26, 25) {real, imag} */,
  {32'h3c3b33f9, 32'h3d9416db} /* (28, 26, 24) {real, imag} */,
  {32'hbcbdc854, 32'h3da1b72f} /* (28, 26, 23) {real, imag} */,
  {32'hbdbc9289, 32'hbcad6290} /* (28, 26, 22) {real, imag} */,
  {32'h3d4d30bc, 32'h3a5e5b5c} /* (28, 26, 21) {real, imag} */,
  {32'h3d52512e, 32'h3d441af4} /* (28, 26, 20) {real, imag} */,
  {32'hba5b42c0, 32'hbd18dcd1} /* (28, 26, 19) {real, imag} */,
  {32'hbdcd8b90, 32'h3ddb74d8} /* (28, 26, 18) {real, imag} */,
  {32'h3d4028a6, 32'hbd11363a} /* (28, 26, 17) {real, imag} */,
  {32'h3b219908, 32'h00000000} /* (28, 26, 16) {real, imag} */,
  {32'h3d4028a6, 32'h3d11363a} /* (28, 26, 15) {real, imag} */,
  {32'hbdcd8b90, 32'hbddb74d8} /* (28, 26, 14) {real, imag} */,
  {32'hba5b42c0, 32'h3d18dcd1} /* (28, 26, 13) {real, imag} */,
  {32'h3d52512e, 32'hbd441af4} /* (28, 26, 12) {real, imag} */,
  {32'h3d4d30bc, 32'hba5e5b5c} /* (28, 26, 11) {real, imag} */,
  {32'hbdbc9289, 32'h3cad6290} /* (28, 26, 10) {real, imag} */,
  {32'hbcbdc854, 32'hbda1b72f} /* (28, 26, 9) {real, imag} */,
  {32'h3c3b33f9, 32'hbd9416db} /* (28, 26, 8) {real, imag} */,
  {32'h3dad4a9e, 32'h3df2b5d8} /* (28, 26, 7) {real, imag} */,
  {32'hbc33e4a4, 32'h3d307a98} /* (28, 26, 6) {real, imag} */,
  {32'hbdb4361e, 32'hbe45a722} /* (28, 26, 5) {real, imag} */,
  {32'h3e3a51be, 32'h3dca576c} /* (28, 26, 4) {real, imag} */,
  {32'h3d96bfd2, 32'h3d3aad6a} /* (28, 26, 3) {real, imag} */,
  {32'hbf95b62c, 32'hbe7096b4} /* (28, 26, 2) {real, imag} */,
  {32'h3fb1e26b, 32'hbdc7159c} /* (28, 26, 1) {real, imag} */,
  {32'h3ecdc814, 32'h00000000} /* (28, 26, 0) {real, imag} */,
  {32'h3fa11918, 32'hbc155c90} /* (28, 25, 31) {real, imag} */,
  {32'hbf8a0f34, 32'h3e77453c} /* (28, 25, 30) {real, imag} */,
  {32'h3c9ec148, 32'hbd6cf162} /* (28, 25, 29) {real, imag} */,
  {32'h3e57f94d, 32'hbe1c07f3} /* (28, 25, 28) {real, imag} */,
  {32'hbe058dcf, 32'h3c8cacf8} /* (28, 25, 27) {real, imag} */,
  {32'h3d58d20d, 32'hbcef2507} /* (28, 25, 26) {real, imag} */,
  {32'h3dfd9b3a, 32'hbdd9d300} /* (28, 25, 25) {real, imag} */,
  {32'hbd0cd180, 32'h3d0bff98} /* (28, 25, 24) {real, imag} */,
  {32'hbbc33eb8, 32'h3dab2cc0} /* (28, 25, 23) {real, imag} */,
  {32'hbc884dbc, 32'hbd0ea075} /* (28, 25, 22) {real, imag} */,
  {32'hbdb55acd, 32'hbdd01700} /* (28, 25, 21) {real, imag} */,
  {32'h3d86cbba, 32'h3be3700c} /* (28, 25, 20) {real, imag} */,
  {32'h3d0172ec, 32'h3c4d3bc8} /* (28, 25, 19) {real, imag} */,
  {32'hba0a0e80, 32'h3cd4e0fd} /* (28, 25, 18) {real, imag} */,
  {32'hbaf319f0, 32'hbc822a96} /* (28, 25, 17) {real, imag} */,
  {32'hbcd31e6b, 32'h00000000} /* (28, 25, 16) {real, imag} */,
  {32'hbaf319f0, 32'h3c822a96} /* (28, 25, 15) {real, imag} */,
  {32'hba0a0e80, 32'hbcd4e0fd} /* (28, 25, 14) {real, imag} */,
  {32'h3d0172ec, 32'hbc4d3bc8} /* (28, 25, 13) {real, imag} */,
  {32'h3d86cbba, 32'hbbe3700c} /* (28, 25, 12) {real, imag} */,
  {32'hbdb55acd, 32'h3dd01700} /* (28, 25, 11) {real, imag} */,
  {32'hbc884dbc, 32'h3d0ea075} /* (28, 25, 10) {real, imag} */,
  {32'hbbc33eb8, 32'hbdab2cc0} /* (28, 25, 9) {real, imag} */,
  {32'hbd0cd180, 32'hbd0bff98} /* (28, 25, 8) {real, imag} */,
  {32'h3dfd9b3a, 32'h3dd9d300} /* (28, 25, 7) {real, imag} */,
  {32'h3d58d20d, 32'h3cef2507} /* (28, 25, 6) {real, imag} */,
  {32'hbe058dcf, 32'hbc8cacf8} /* (28, 25, 5) {real, imag} */,
  {32'h3e57f94d, 32'h3e1c07f3} /* (28, 25, 4) {real, imag} */,
  {32'h3c9ec148, 32'h3d6cf162} /* (28, 25, 3) {real, imag} */,
  {32'hbf8a0f34, 32'hbe77453c} /* (28, 25, 2) {real, imag} */,
  {32'h3fa11918, 32'h3c155c90} /* (28, 25, 1) {real, imag} */,
  {32'h3f1bcfa3, 32'h00000000} /* (28, 25, 0) {real, imag} */,
  {32'h3fa1267c, 32'hbd1e6ece} /* (28, 24, 31) {real, imag} */,
  {32'hbf99d6ca, 32'h3ea73b18} /* (28, 24, 30) {real, imag} */,
  {32'hbcc98e88, 32'hbe403452} /* (28, 24, 29) {real, imag} */,
  {32'h3e4d3346, 32'h3d526b68} /* (28, 24, 28) {real, imag} */,
  {32'hbd940552, 32'h3c5dcdf0} /* (28, 24, 27) {real, imag} */,
  {32'hbce62f41, 32'h3db6a532} /* (28, 24, 26) {real, imag} */,
  {32'hbd6bbdda, 32'hbe16963b} /* (28, 24, 25) {real, imag} */,
  {32'h3d7c8ca0, 32'h3d7ad9ce} /* (28, 24, 24) {real, imag} */,
  {32'hbdb10b73, 32'h3d1a82aa} /* (28, 24, 23) {real, imag} */,
  {32'hbc992642, 32'h3cb5fe28} /* (28, 24, 22) {real, imag} */,
  {32'hbd42792e, 32'h3d87cbbb} /* (28, 24, 21) {real, imag} */,
  {32'h3c12cd5c, 32'h3ccbd66a} /* (28, 24, 20) {real, imag} */,
  {32'h3dc2244d, 32'h3d925f98} /* (28, 24, 19) {real, imag} */,
  {32'h3bea06d8, 32'hbcc46e59} /* (28, 24, 18) {real, imag} */,
  {32'hbcb17048, 32'hbd863064} /* (28, 24, 17) {real, imag} */,
  {32'hbc92978b, 32'h00000000} /* (28, 24, 16) {real, imag} */,
  {32'hbcb17048, 32'h3d863064} /* (28, 24, 15) {real, imag} */,
  {32'h3bea06d8, 32'h3cc46e59} /* (28, 24, 14) {real, imag} */,
  {32'h3dc2244d, 32'hbd925f98} /* (28, 24, 13) {real, imag} */,
  {32'h3c12cd5c, 32'hbccbd66a} /* (28, 24, 12) {real, imag} */,
  {32'hbd42792e, 32'hbd87cbbb} /* (28, 24, 11) {real, imag} */,
  {32'hbc992642, 32'hbcb5fe28} /* (28, 24, 10) {real, imag} */,
  {32'hbdb10b73, 32'hbd1a82aa} /* (28, 24, 9) {real, imag} */,
  {32'h3d7c8ca0, 32'hbd7ad9ce} /* (28, 24, 8) {real, imag} */,
  {32'hbd6bbdda, 32'h3e16963b} /* (28, 24, 7) {real, imag} */,
  {32'hbce62f41, 32'hbdb6a532} /* (28, 24, 6) {real, imag} */,
  {32'hbd940552, 32'hbc5dcdf0} /* (28, 24, 5) {real, imag} */,
  {32'h3e4d3346, 32'hbd526b68} /* (28, 24, 4) {real, imag} */,
  {32'hbcc98e88, 32'h3e403452} /* (28, 24, 3) {real, imag} */,
  {32'hbf99d6ca, 32'hbea73b18} /* (28, 24, 2) {real, imag} */,
  {32'h3fa1267c, 32'h3d1e6ece} /* (28, 24, 1) {real, imag} */,
  {32'h3f32906c, 32'h00000000} /* (28, 24, 0) {real, imag} */,
  {32'h3f85969e, 32'hbdd5239a} /* (28, 23, 31) {real, imag} */,
  {32'hbf77d9f6, 32'h3e147a4f} /* (28, 23, 30) {real, imag} */,
  {32'hbc910422, 32'hbdc3737f} /* (28, 23, 29) {real, imag} */,
  {32'h3db34655, 32'hbd586a78} /* (28, 23, 28) {real, imag} */,
  {32'hbd3bf354, 32'h3e43817a} /* (28, 23, 27) {real, imag} */,
  {32'h3b237770, 32'h3d347ef6} /* (28, 23, 26) {real, imag} */,
  {32'hbd6bdece, 32'hbe3f38e4} /* (28, 23, 25) {real, imag} */,
  {32'hbcf6f299, 32'h3ddefbf8} /* (28, 23, 24) {real, imag} */,
  {32'hbdc4c674, 32'hbd8370ab} /* (28, 23, 23) {real, imag} */,
  {32'hbc9ebadc, 32'h3d21708c} /* (28, 23, 22) {real, imag} */,
  {32'h3da061b3, 32'h3d4c22cb} /* (28, 23, 21) {real, imag} */,
  {32'h3cfced74, 32'hbd5ee2dc} /* (28, 23, 20) {real, imag} */,
  {32'hbd23a1e2, 32'hbcc0c748} /* (28, 23, 19) {real, imag} */,
  {32'h3c82f90e, 32'h3d8008cb} /* (28, 23, 18) {real, imag} */,
  {32'h3d341ba9, 32'h3d6c9759} /* (28, 23, 17) {real, imag} */,
  {32'hbdd30014, 32'h00000000} /* (28, 23, 16) {real, imag} */,
  {32'h3d341ba9, 32'hbd6c9759} /* (28, 23, 15) {real, imag} */,
  {32'h3c82f90e, 32'hbd8008cb} /* (28, 23, 14) {real, imag} */,
  {32'hbd23a1e2, 32'h3cc0c748} /* (28, 23, 13) {real, imag} */,
  {32'h3cfced74, 32'h3d5ee2dc} /* (28, 23, 12) {real, imag} */,
  {32'h3da061b3, 32'hbd4c22cb} /* (28, 23, 11) {real, imag} */,
  {32'hbc9ebadc, 32'hbd21708c} /* (28, 23, 10) {real, imag} */,
  {32'hbdc4c674, 32'h3d8370ab} /* (28, 23, 9) {real, imag} */,
  {32'hbcf6f299, 32'hbddefbf8} /* (28, 23, 8) {real, imag} */,
  {32'hbd6bdece, 32'h3e3f38e4} /* (28, 23, 7) {real, imag} */,
  {32'h3b237770, 32'hbd347ef6} /* (28, 23, 6) {real, imag} */,
  {32'hbd3bf354, 32'hbe43817a} /* (28, 23, 5) {real, imag} */,
  {32'h3db34655, 32'h3d586a78} /* (28, 23, 4) {real, imag} */,
  {32'hbc910422, 32'h3dc3737f} /* (28, 23, 3) {real, imag} */,
  {32'hbf77d9f6, 32'hbe147a4f} /* (28, 23, 2) {real, imag} */,
  {32'h3f85969e, 32'h3dd5239a} /* (28, 23, 1) {real, imag} */,
  {32'h3f3b063a, 32'h00000000} /* (28, 23, 0) {real, imag} */,
  {32'h3f295648, 32'hbb639fa0} /* (28, 22, 31) {real, imag} */,
  {32'hbeeb1098, 32'h3d0393c5} /* (28, 22, 30) {real, imag} */,
  {32'h3d212e5a, 32'hbdcd7a91} /* (28, 22, 29) {real, imag} */,
  {32'hbbeecf90, 32'hbdcf0af8} /* (28, 22, 28) {real, imag} */,
  {32'hbe145658, 32'h3cffb712} /* (28, 22, 27) {real, imag} */,
  {32'hbd91d2cc, 32'h3d292486} /* (28, 22, 26) {real, imag} */,
  {32'hbcf5261a, 32'hbe166c28} /* (28, 22, 25) {real, imag} */,
  {32'hbd6c96e6, 32'h3c977f02} /* (28, 22, 24) {real, imag} */,
  {32'hbcab6fb7, 32'h3d9148ce} /* (28, 22, 23) {real, imag} */,
  {32'hbc69504e, 32'h3daedba7} /* (28, 22, 22) {real, imag} */,
  {32'h3d05a3b0, 32'h3d720685} /* (28, 22, 21) {real, imag} */,
  {32'hbc9f8c8c, 32'h3d9fc474} /* (28, 22, 20) {real, imag} */,
  {32'h3cfa46b5, 32'hbb1c2640} /* (28, 22, 19) {real, imag} */,
  {32'hbceffe33, 32'h3c91b284} /* (28, 22, 18) {real, imag} */,
  {32'h3caf401c, 32'h3b907248} /* (28, 22, 17) {real, imag} */,
  {32'h3ce21ee4, 32'h00000000} /* (28, 22, 16) {real, imag} */,
  {32'h3caf401c, 32'hbb907248} /* (28, 22, 15) {real, imag} */,
  {32'hbceffe33, 32'hbc91b284} /* (28, 22, 14) {real, imag} */,
  {32'h3cfa46b5, 32'h3b1c2640} /* (28, 22, 13) {real, imag} */,
  {32'hbc9f8c8c, 32'hbd9fc474} /* (28, 22, 12) {real, imag} */,
  {32'h3d05a3b0, 32'hbd720685} /* (28, 22, 11) {real, imag} */,
  {32'hbc69504e, 32'hbdaedba7} /* (28, 22, 10) {real, imag} */,
  {32'hbcab6fb7, 32'hbd9148ce} /* (28, 22, 9) {real, imag} */,
  {32'hbd6c96e6, 32'hbc977f02} /* (28, 22, 8) {real, imag} */,
  {32'hbcf5261a, 32'h3e166c28} /* (28, 22, 7) {real, imag} */,
  {32'hbd91d2cc, 32'hbd292486} /* (28, 22, 6) {real, imag} */,
  {32'hbe145658, 32'hbcffb712} /* (28, 22, 5) {real, imag} */,
  {32'hbbeecf90, 32'h3dcf0af8} /* (28, 22, 4) {real, imag} */,
  {32'h3d212e5a, 32'h3dcd7a91} /* (28, 22, 3) {real, imag} */,
  {32'hbeeb1098, 32'hbd0393c5} /* (28, 22, 2) {real, imag} */,
  {32'h3f295648, 32'h3b639fa0} /* (28, 22, 1) {real, imag} */,
  {32'h3f246f99, 32'h00000000} /* (28, 22, 0) {real, imag} */,
  {32'hbdc6581c, 32'h3d001a94} /* (28, 21, 31) {real, imag} */,
  {32'hbce6fbe8, 32'h3c33f540} /* (28, 21, 30) {real, imag} */,
  {32'h3d5ad882, 32'hbcc4b74c} /* (28, 21, 29) {real, imag} */,
  {32'hbd388ff4, 32'hbb849ae8} /* (28, 21, 28) {real, imag} */,
  {32'hbd56c3ff, 32'hbd0ee0e7} /* (28, 21, 27) {real, imag} */,
  {32'hbd62593d, 32'h3d18fc2a} /* (28, 21, 26) {real, imag} */,
  {32'h3d583076, 32'h3d2bb030} /* (28, 21, 25) {real, imag} */,
  {32'h3da5a0ca, 32'h3db4c6f9} /* (28, 21, 24) {real, imag} */,
  {32'h3d13526c, 32'hbd235060} /* (28, 21, 23) {real, imag} */,
  {32'h3d5fa561, 32'h3d5481ab} /* (28, 21, 22) {real, imag} */,
  {32'hbccba790, 32'h3dd9e1f0} /* (28, 21, 21) {real, imag} */,
  {32'hbcbd4b2c, 32'hbd60c016} /* (28, 21, 20) {real, imag} */,
  {32'hbca8772c, 32'hbbc8dba0} /* (28, 21, 19) {real, imag} */,
  {32'hbdca9278, 32'hbd141690} /* (28, 21, 18) {real, imag} */,
  {32'hba3ee9c0, 32'hbd408030} /* (28, 21, 17) {real, imag} */,
  {32'hbbaea170, 32'h00000000} /* (28, 21, 16) {real, imag} */,
  {32'hba3ee9c0, 32'h3d408030} /* (28, 21, 15) {real, imag} */,
  {32'hbdca9278, 32'h3d141690} /* (28, 21, 14) {real, imag} */,
  {32'hbca8772c, 32'h3bc8dba0} /* (28, 21, 13) {real, imag} */,
  {32'hbcbd4b2c, 32'h3d60c016} /* (28, 21, 12) {real, imag} */,
  {32'hbccba790, 32'hbdd9e1f0} /* (28, 21, 11) {real, imag} */,
  {32'h3d5fa561, 32'hbd5481ab} /* (28, 21, 10) {real, imag} */,
  {32'h3d13526c, 32'h3d235060} /* (28, 21, 9) {real, imag} */,
  {32'h3da5a0ca, 32'hbdb4c6f9} /* (28, 21, 8) {real, imag} */,
  {32'h3d583076, 32'hbd2bb030} /* (28, 21, 7) {real, imag} */,
  {32'hbd62593d, 32'hbd18fc2a} /* (28, 21, 6) {real, imag} */,
  {32'hbd56c3ff, 32'h3d0ee0e7} /* (28, 21, 5) {real, imag} */,
  {32'hbd388ff4, 32'h3b849ae8} /* (28, 21, 4) {real, imag} */,
  {32'h3d5ad882, 32'h3cc4b74c} /* (28, 21, 3) {real, imag} */,
  {32'hbce6fbe8, 32'hbc33f540} /* (28, 21, 2) {real, imag} */,
  {32'hbdc6581c, 32'hbd001a94} /* (28, 21, 1) {real, imag} */,
  {32'hb9f32c00, 32'h00000000} /* (28, 21, 0) {real, imag} */,
  {32'hbf92d9e6, 32'h3e663e28} /* (28, 20, 31) {real, imag} */,
  {32'h3f04c0a6, 32'hbe4948c5} /* (28, 20, 30) {real, imag} */,
  {32'h3e22e8d9, 32'hbdb0fa18} /* (28, 20, 29) {real, imag} */,
  {32'hbe39610a, 32'h3cf7beac} /* (28, 20, 28) {real, imag} */,
  {32'h3dc2c111, 32'hbcdbfda8} /* (28, 20, 27) {real, imag} */,
  {32'h3d0c139c, 32'hbd460f26} /* (28, 20, 26) {real, imag} */,
  {32'h3d099e0d, 32'h3d2a5907} /* (28, 20, 25) {real, imag} */,
  {32'h3c437336, 32'hbde34c18} /* (28, 20, 24) {real, imag} */,
  {32'h3d7c6ef8, 32'hbd7f7b30} /* (28, 20, 23) {real, imag} */,
  {32'h3e34135b, 32'h3d37d0de} /* (28, 20, 22) {real, imag} */,
  {32'h3e1980e9, 32'h3d761046} /* (28, 20, 21) {real, imag} */,
  {32'h3cabacea, 32'h3af6d280} /* (28, 20, 20) {real, imag} */,
  {32'hbd3d1232, 32'h3c926321} /* (28, 20, 19) {real, imag} */,
  {32'h3d035434, 32'hbae3ab00} /* (28, 20, 18) {real, imag} */,
  {32'h3c2ec2c0, 32'h3d7bb2c8} /* (28, 20, 17) {real, imag} */,
  {32'hbd8056c5, 32'h00000000} /* (28, 20, 16) {real, imag} */,
  {32'h3c2ec2c0, 32'hbd7bb2c8} /* (28, 20, 15) {real, imag} */,
  {32'h3d035434, 32'h3ae3ab00} /* (28, 20, 14) {real, imag} */,
  {32'hbd3d1232, 32'hbc926321} /* (28, 20, 13) {real, imag} */,
  {32'h3cabacea, 32'hbaf6d280} /* (28, 20, 12) {real, imag} */,
  {32'h3e1980e9, 32'hbd761046} /* (28, 20, 11) {real, imag} */,
  {32'h3e34135b, 32'hbd37d0de} /* (28, 20, 10) {real, imag} */,
  {32'h3d7c6ef8, 32'h3d7f7b30} /* (28, 20, 9) {real, imag} */,
  {32'h3c437336, 32'h3de34c18} /* (28, 20, 8) {real, imag} */,
  {32'h3d099e0d, 32'hbd2a5907} /* (28, 20, 7) {real, imag} */,
  {32'h3d0c139c, 32'h3d460f26} /* (28, 20, 6) {real, imag} */,
  {32'h3dc2c111, 32'h3cdbfda8} /* (28, 20, 5) {real, imag} */,
  {32'hbe39610a, 32'hbcf7beac} /* (28, 20, 4) {real, imag} */,
  {32'h3e22e8d9, 32'h3db0fa18} /* (28, 20, 3) {real, imag} */,
  {32'h3f04c0a6, 32'h3e4948c5} /* (28, 20, 2) {real, imag} */,
  {32'hbf92d9e6, 32'hbe663e28} /* (28, 20, 1) {real, imag} */,
  {32'hbf22adfe, 32'h00000000} /* (28, 20, 0) {real, imag} */,
  {32'hbfcd16d2, 32'h3e86ce36} /* (28, 19, 31) {real, imag} */,
  {32'h3f29588d, 32'hbe698e90} /* (28, 19, 30) {real, imag} */,
  {32'h3c969f38, 32'hbdea2df8} /* (28, 19, 29) {real, imag} */,
  {32'hbdfb0b68, 32'h3cf42046} /* (28, 19, 28) {real, imag} */,
  {32'h3d8d395a, 32'h3cc24978} /* (28, 19, 27) {real, imag} */,
  {32'hbd8a9825, 32'hbd3ccd73} /* (28, 19, 26) {real, imag} */,
  {32'hbd5f188e, 32'h3d2fece0} /* (28, 19, 25) {real, imag} */,
  {32'hbc32fc00, 32'hbddd023c} /* (28, 19, 24) {real, imag} */,
  {32'h3d56b3ec, 32'hbbf7c826} /* (28, 19, 23) {real, imag} */,
  {32'h3dc5b552, 32'hbc0c007c} /* (28, 19, 22) {real, imag} */,
  {32'hbd03bc13, 32'hbb2e8058} /* (28, 19, 21) {real, imag} */,
  {32'hbc610fe8, 32'h3aab3c64} /* (28, 19, 20) {real, imag} */,
  {32'hbd6c7eeb, 32'hbbaf3568} /* (28, 19, 19) {real, imag} */,
  {32'hbd8eb912, 32'hbd2e01dc} /* (28, 19, 18) {real, imag} */,
  {32'hbd2b69f5, 32'hbd0b2866} /* (28, 19, 17) {real, imag} */,
  {32'hbd61f6dc, 32'h00000000} /* (28, 19, 16) {real, imag} */,
  {32'hbd2b69f5, 32'h3d0b2866} /* (28, 19, 15) {real, imag} */,
  {32'hbd8eb912, 32'h3d2e01dc} /* (28, 19, 14) {real, imag} */,
  {32'hbd6c7eeb, 32'h3baf3568} /* (28, 19, 13) {real, imag} */,
  {32'hbc610fe8, 32'hbaab3c64} /* (28, 19, 12) {real, imag} */,
  {32'hbd03bc13, 32'h3b2e8058} /* (28, 19, 11) {real, imag} */,
  {32'h3dc5b552, 32'h3c0c007c} /* (28, 19, 10) {real, imag} */,
  {32'h3d56b3ec, 32'h3bf7c826} /* (28, 19, 9) {real, imag} */,
  {32'hbc32fc00, 32'h3ddd023c} /* (28, 19, 8) {real, imag} */,
  {32'hbd5f188e, 32'hbd2fece0} /* (28, 19, 7) {real, imag} */,
  {32'hbd8a9825, 32'h3d3ccd73} /* (28, 19, 6) {real, imag} */,
  {32'h3d8d395a, 32'hbcc24978} /* (28, 19, 5) {real, imag} */,
  {32'hbdfb0b68, 32'hbcf42046} /* (28, 19, 4) {real, imag} */,
  {32'h3c969f38, 32'h3dea2df8} /* (28, 19, 3) {real, imag} */,
  {32'h3f29588d, 32'h3e698e90} /* (28, 19, 2) {real, imag} */,
  {32'hbfcd16d2, 32'hbe86ce36} /* (28, 19, 1) {real, imag} */,
  {32'hbf8e4cc6, 32'h00000000} /* (28, 19, 0) {real, imag} */,
  {32'hbfe9aaab, 32'h3ec240e8} /* (28, 18, 31) {real, imag} */,
  {32'h3f63df0b, 32'hbeac505a} /* (28, 18, 30) {real, imag} */,
  {32'hbd81bb72, 32'hbba08d60} /* (28, 18, 29) {real, imag} */,
  {32'hbd8edc86, 32'h3e0c81a8} /* (28, 18, 28) {real, imag} */,
  {32'h3e474709, 32'hbdeda588} /* (28, 18, 27) {real, imag} */,
  {32'hbdfd11f6, 32'hbd0183b7} /* (28, 18, 26) {real, imag} */,
  {32'h3cc00045, 32'h3db41c7e} /* (28, 18, 25) {real, imag} */,
  {32'h3d52fa6b, 32'hbdc36303} /* (28, 18, 24) {real, imag} */,
  {32'h3bb23128, 32'hbddf202e} /* (28, 18, 23) {real, imag} */,
  {32'h3d8d588a, 32'h3bf85298} /* (28, 18, 22) {real, imag} */,
  {32'hbcc6fb08, 32'h3c221130} /* (28, 18, 21) {real, imag} */,
  {32'hbbebab40, 32'hbd14924e} /* (28, 18, 20) {real, imag} */,
  {32'hbd94fbeb, 32'h3d78ef70} /* (28, 18, 19) {real, imag} */,
  {32'hbcc6d14b, 32'hbd5822ae} /* (28, 18, 18) {real, imag} */,
  {32'hbd988a7b, 32'h3d3091fa} /* (28, 18, 17) {real, imag} */,
  {32'hbbfeba91, 32'h00000000} /* (28, 18, 16) {real, imag} */,
  {32'hbd988a7b, 32'hbd3091fa} /* (28, 18, 15) {real, imag} */,
  {32'hbcc6d14b, 32'h3d5822ae} /* (28, 18, 14) {real, imag} */,
  {32'hbd94fbeb, 32'hbd78ef70} /* (28, 18, 13) {real, imag} */,
  {32'hbbebab40, 32'h3d14924e} /* (28, 18, 12) {real, imag} */,
  {32'hbcc6fb08, 32'hbc221130} /* (28, 18, 11) {real, imag} */,
  {32'h3d8d588a, 32'hbbf85298} /* (28, 18, 10) {real, imag} */,
  {32'h3bb23128, 32'h3ddf202e} /* (28, 18, 9) {real, imag} */,
  {32'h3d52fa6b, 32'h3dc36303} /* (28, 18, 8) {real, imag} */,
  {32'h3cc00045, 32'hbdb41c7e} /* (28, 18, 7) {real, imag} */,
  {32'hbdfd11f6, 32'h3d0183b7} /* (28, 18, 6) {real, imag} */,
  {32'h3e474709, 32'h3deda588} /* (28, 18, 5) {real, imag} */,
  {32'hbd8edc86, 32'hbe0c81a8} /* (28, 18, 4) {real, imag} */,
  {32'hbd81bb72, 32'h3ba08d60} /* (28, 18, 3) {real, imag} */,
  {32'h3f63df0b, 32'h3eac505a} /* (28, 18, 2) {real, imag} */,
  {32'hbfe9aaab, 32'hbec240e8} /* (28, 18, 1) {real, imag} */,
  {32'hbfb7e1c5, 32'h00000000} /* (28, 18, 0) {real, imag} */,
  {32'hbff27d43, 32'h3ef8d990} /* (28, 17, 31) {real, imag} */,
  {32'h3f73e612, 32'hbe45f708} /* (28, 17, 30) {real, imag} */,
  {32'h3dcc1a0c, 32'hbd50e180} /* (28, 17, 29) {real, imag} */,
  {32'hbda071c5, 32'h3dc92f48} /* (28, 17, 28) {real, imag} */,
  {32'h3e412984, 32'hbd3004a2} /* (28, 17, 27) {real, imag} */,
  {32'h3c8bb190, 32'hbd16c8a1} /* (28, 17, 26) {real, imag} */,
  {32'h3ddd42c4, 32'h3d846666} /* (28, 17, 25) {real, imag} */,
  {32'h3d3fff44, 32'hbace0a90} /* (28, 17, 24) {real, imag} */,
  {32'h3cbde91e, 32'hbcb7f5ca} /* (28, 17, 23) {real, imag} */,
  {32'hbdf8020f, 32'hbda5e3d0} /* (28, 17, 22) {real, imag} */,
  {32'hbcecf772, 32'hbd1c1408} /* (28, 17, 21) {real, imag} */,
  {32'h3c1f148a, 32'h3c1bf754} /* (28, 17, 20) {real, imag} */,
  {32'h3cd363de, 32'hbd80f300} /* (28, 17, 19) {real, imag} */,
  {32'h3cce3728, 32'h3a80af00} /* (28, 17, 18) {real, imag} */,
  {32'hbd20e2a5, 32'h3d67a770} /* (28, 17, 17) {real, imag} */,
  {32'h3e1fff0e, 32'h00000000} /* (28, 17, 16) {real, imag} */,
  {32'hbd20e2a5, 32'hbd67a770} /* (28, 17, 15) {real, imag} */,
  {32'h3cce3728, 32'hba80af00} /* (28, 17, 14) {real, imag} */,
  {32'h3cd363de, 32'h3d80f300} /* (28, 17, 13) {real, imag} */,
  {32'h3c1f148a, 32'hbc1bf754} /* (28, 17, 12) {real, imag} */,
  {32'hbcecf772, 32'h3d1c1408} /* (28, 17, 11) {real, imag} */,
  {32'hbdf8020f, 32'h3da5e3d0} /* (28, 17, 10) {real, imag} */,
  {32'h3cbde91e, 32'h3cb7f5ca} /* (28, 17, 9) {real, imag} */,
  {32'h3d3fff44, 32'h3ace0a90} /* (28, 17, 8) {real, imag} */,
  {32'h3ddd42c4, 32'hbd846666} /* (28, 17, 7) {real, imag} */,
  {32'h3c8bb190, 32'h3d16c8a1} /* (28, 17, 6) {real, imag} */,
  {32'h3e412984, 32'h3d3004a2} /* (28, 17, 5) {real, imag} */,
  {32'hbda071c5, 32'hbdc92f48} /* (28, 17, 4) {real, imag} */,
  {32'h3dcc1a0c, 32'h3d50e180} /* (28, 17, 3) {real, imag} */,
  {32'h3f73e612, 32'h3e45f708} /* (28, 17, 2) {real, imag} */,
  {32'hbff27d43, 32'hbef8d990} /* (28, 17, 1) {real, imag} */,
  {32'hbfd094f4, 32'h00000000} /* (28, 17, 0) {real, imag} */,
  {32'hbff21890, 32'h3eafb89e} /* (28, 16, 31) {real, imag} */,
  {32'h3f7ecd50, 32'hbe45907a} /* (28, 16, 30) {real, imag} */,
  {32'h3d8e49e5, 32'h3c98ffd6} /* (28, 16, 29) {real, imag} */,
  {32'hbda7a401, 32'h3e20d283} /* (28, 16, 28) {real, imag} */,
  {32'h3cccc588, 32'hbd95669b} /* (28, 16, 27) {real, imag} */,
  {32'h3dee3bee, 32'h3c2859de} /* (28, 16, 26) {real, imag} */,
  {32'hbd0c563d, 32'hbb3fe1d8} /* (28, 16, 25) {real, imag} */,
  {32'hbbd65edc, 32'hbd488308} /* (28, 16, 24) {real, imag} */,
  {32'hbca5d242, 32'hbdca6807} /* (28, 16, 23) {real, imag} */,
  {32'h3d9f2a05, 32'h3c080124} /* (28, 16, 22) {real, imag} */,
  {32'h3d3f537d, 32'hbd88d8b7} /* (28, 16, 21) {real, imag} */,
  {32'h3d528722, 32'h3bdd7b5e} /* (28, 16, 20) {real, imag} */,
  {32'h3d77ce77, 32'hbd1c89b3} /* (28, 16, 19) {real, imag} */,
  {32'hbd50a208, 32'hbd870ea6} /* (28, 16, 18) {real, imag} */,
  {32'hbd7186d6, 32'h3d49323a} /* (28, 16, 17) {real, imag} */,
  {32'hbcc49701, 32'h00000000} /* (28, 16, 16) {real, imag} */,
  {32'hbd7186d6, 32'hbd49323a} /* (28, 16, 15) {real, imag} */,
  {32'hbd50a208, 32'h3d870ea6} /* (28, 16, 14) {real, imag} */,
  {32'h3d77ce77, 32'h3d1c89b3} /* (28, 16, 13) {real, imag} */,
  {32'h3d528722, 32'hbbdd7b5e} /* (28, 16, 12) {real, imag} */,
  {32'h3d3f537d, 32'h3d88d8b7} /* (28, 16, 11) {real, imag} */,
  {32'h3d9f2a05, 32'hbc080124} /* (28, 16, 10) {real, imag} */,
  {32'hbca5d242, 32'h3dca6807} /* (28, 16, 9) {real, imag} */,
  {32'hbbd65edc, 32'h3d488308} /* (28, 16, 8) {real, imag} */,
  {32'hbd0c563d, 32'h3b3fe1d8} /* (28, 16, 7) {real, imag} */,
  {32'h3dee3bee, 32'hbc2859de} /* (28, 16, 6) {real, imag} */,
  {32'h3cccc588, 32'h3d95669b} /* (28, 16, 5) {real, imag} */,
  {32'hbda7a401, 32'hbe20d283} /* (28, 16, 4) {real, imag} */,
  {32'h3d8e49e5, 32'hbc98ffd6} /* (28, 16, 3) {real, imag} */,
  {32'h3f7ecd50, 32'h3e45907a} /* (28, 16, 2) {real, imag} */,
  {32'hbff21890, 32'hbeafb89e} /* (28, 16, 1) {real, imag} */,
  {32'hbfc6dd09, 32'h00000000} /* (28, 16, 0) {real, imag} */,
  {32'hbfef3ebd, 32'h3e78e370} /* (28, 15, 31) {real, imag} */,
  {32'h3f837347, 32'hbe7478e8} /* (28, 15, 30) {real, imag} */,
  {32'h3d81cda4, 32'h3cc6104b} /* (28, 15, 29) {real, imag} */,
  {32'hbe810b81, 32'h3e218d38} /* (28, 15, 28) {real, imag} */,
  {32'h3dad7414, 32'hbd2840ea} /* (28, 15, 27) {real, imag} */,
  {32'h3de5cf20, 32'h3cc957b2} /* (28, 15, 26) {real, imag} */,
  {32'hbd5d6974, 32'h3cb99d05} /* (28, 15, 25) {real, imag} */,
  {32'h3e126c99, 32'hbd59f01e} /* (28, 15, 24) {real, imag} */,
  {32'hbce5475c, 32'hbcb90962} /* (28, 15, 23) {real, imag} */,
  {32'hbb803110, 32'hbd4d5688} /* (28, 15, 22) {real, imag} */,
  {32'h3d4f336f, 32'hbb294cb0} /* (28, 15, 21) {real, imag} */,
  {32'hbc7d3c1a, 32'hbd9f149c} /* (28, 15, 20) {real, imag} */,
  {32'hbbcfddd8, 32'hbd509315} /* (28, 15, 19) {real, imag} */,
  {32'hbc7df591, 32'hbdb0bba0} /* (28, 15, 18) {real, imag} */,
  {32'h3c99c662, 32'h3c918268} /* (28, 15, 17) {real, imag} */,
  {32'hbd3d4f56, 32'h00000000} /* (28, 15, 16) {real, imag} */,
  {32'h3c99c662, 32'hbc918268} /* (28, 15, 15) {real, imag} */,
  {32'hbc7df591, 32'h3db0bba0} /* (28, 15, 14) {real, imag} */,
  {32'hbbcfddd8, 32'h3d509315} /* (28, 15, 13) {real, imag} */,
  {32'hbc7d3c1a, 32'h3d9f149c} /* (28, 15, 12) {real, imag} */,
  {32'h3d4f336f, 32'h3b294cb0} /* (28, 15, 11) {real, imag} */,
  {32'hbb803110, 32'h3d4d5688} /* (28, 15, 10) {real, imag} */,
  {32'hbce5475c, 32'h3cb90962} /* (28, 15, 9) {real, imag} */,
  {32'h3e126c99, 32'h3d59f01e} /* (28, 15, 8) {real, imag} */,
  {32'hbd5d6974, 32'hbcb99d05} /* (28, 15, 7) {real, imag} */,
  {32'h3de5cf20, 32'hbcc957b2} /* (28, 15, 6) {real, imag} */,
  {32'h3dad7414, 32'h3d2840ea} /* (28, 15, 5) {real, imag} */,
  {32'hbe810b81, 32'hbe218d38} /* (28, 15, 4) {real, imag} */,
  {32'h3d81cda4, 32'hbcc6104b} /* (28, 15, 3) {real, imag} */,
  {32'h3f837347, 32'h3e7478e8} /* (28, 15, 2) {real, imag} */,
  {32'hbfef3ebd, 32'hbe78e370} /* (28, 15, 1) {real, imag} */,
  {32'hbfc03d80, 32'h00000000} /* (28, 15, 0) {real, imag} */,
  {32'hbfdf0181, 32'h3e8d7108} /* (28, 14, 31) {real, imag} */,
  {32'h3f78a265, 32'hbe534ee7} /* (28, 14, 30) {real, imag} */,
  {32'hbd5d6a8c, 32'hbd8f2214} /* (28, 14, 29) {real, imag} */,
  {32'hbe923126, 32'h3d27616f} /* (28, 14, 28) {real, imag} */,
  {32'h3e2cd11f, 32'hbdaedc40} /* (28, 14, 27) {real, imag} */,
  {32'h3e05a53f, 32'hbd30f939} /* (28, 14, 26) {real, imag} */,
  {32'h3c860b1d, 32'hbcc28d66} /* (28, 14, 25) {real, imag} */,
  {32'h3cf1236e, 32'hbb836c90} /* (28, 14, 24) {real, imag} */,
  {32'hbd173c07, 32'hbcfbfc06} /* (28, 14, 23) {real, imag} */,
  {32'h3d55b3f4, 32'hbcdc1836} /* (28, 14, 22) {real, imag} */,
  {32'hbd94f967, 32'h3cfc18e8} /* (28, 14, 21) {real, imag} */,
  {32'h3c63bfc0, 32'hbd17b84a} /* (28, 14, 20) {real, imag} */,
  {32'h3cf59c1c, 32'h3d055236} /* (28, 14, 19) {real, imag} */,
  {32'h3d54031e, 32'hbd17a7de} /* (28, 14, 18) {real, imag} */,
  {32'h3d22554a, 32'hbcd93da4} /* (28, 14, 17) {real, imag} */,
  {32'h3ca75a7c, 32'h00000000} /* (28, 14, 16) {real, imag} */,
  {32'h3d22554a, 32'h3cd93da4} /* (28, 14, 15) {real, imag} */,
  {32'h3d54031e, 32'h3d17a7de} /* (28, 14, 14) {real, imag} */,
  {32'h3cf59c1c, 32'hbd055236} /* (28, 14, 13) {real, imag} */,
  {32'h3c63bfc0, 32'h3d17b84a} /* (28, 14, 12) {real, imag} */,
  {32'hbd94f967, 32'hbcfc18e8} /* (28, 14, 11) {real, imag} */,
  {32'h3d55b3f4, 32'h3cdc1836} /* (28, 14, 10) {real, imag} */,
  {32'hbd173c07, 32'h3cfbfc06} /* (28, 14, 9) {real, imag} */,
  {32'h3cf1236e, 32'h3b836c90} /* (28, 14, 8) {real, imag} */,
  {32'h3c860b1d, 32'h3cc28d66} /* (28, 14, 7) {real, imag} */,
  {32'h3e05a53f, 32'h3d30f939} /* (28, 14, 6) {real, imag} */,
  {32'h3e2cd11f, 32'h3daedc40} /* (28, 14, 5) {real, imag} */,
  {32'hbe923126, 32'hbd27616f} /* (28, 14, 4) {real, imag} */,
  {32'hbd5d6a8c, 32'h3d8f2214} /* (28, 14, 3) {real, imag} */,
  {32'h3f78a265, 32'h3e534ee7} /* (28, 14, 2) {real, imag} */,
  {32'hbfdf0181, 32'hbe8d7108} /* (28, 14, 1) {real, imag} */,
  {32'hbfab78d7, 32'h00000000} /* (28, 14, 0) {real, imag} */,
  {32'hbfc7962a, 32'h3de8e5a2} /* (28, 13, 31) {real, imag} */,
  {32'h3f443763, 32'hbccc18e0} /* (28, 13, 30) {real, imag} */,
  {32'hbde36ba8, 32'h3c9a4cb0} /* (28, 13, 29) {real, imag} */,
  {32'hbe813238, 32'hbdc1970c} /* (28, 13, 28) {real, imag} */,
  {32'h3e35f20b, 32'hbdc84d8f} /* (28, 13, 27) {real, imag} */,
  {32'h3d9aed6b, 32'h3d4a7b39} /* (28, 13, 26) {real, imag} */,
  {32'h3cddb730, 32'hbcf09f90} /* (28, 13, 25) {real, imag} */,
  {32'h3c5c1efc, 32'hbdf55764} /* (28, 13, 24) {real, imag} */,
  {32'h3d46acc8, 32'h3c9bef12} /* (28, 13, 23) {real, imag} */,
  {32'hbd766c08, 32'h3d89ca7e} /* (28, 13, 22) {real, imag} */,
  {32'h3d6e5ef9, 32'h3bf9858c} /* (28, 13, 21) {real, imag} */,
  {32'hbd70530a, 32'hbc541578} /* (28, 13, 20) {real, imag} */,
  {32'h3d4e2ad7, 32'h3da85a06} /* (28, 13, 19) {real, imag} */,
  {32'hbcd90d4a, 32'h3c8ea850} /* (28, 13, 18) {real, imag} */,
  {32'h3c2c76ec, 32'hbb410090} /* (28, 13, 17) {real, imag} */,
  {32'h3bf07930, 32'h00000000} /* (28, 13, 16) {real, imag} */,
  {32'h3c2c76ec, 32'h3b410090} /* (28, 13, 15) {real, imag} */,
  {32'hbcd90d4a, 32'hbc8ea850} /* (28, 13, 14) {real, imag} */,
  {32'h3d4e2ad7, 32'hbda85a06} /* (28, 13, 13) {real, imag} */,
  {32'hbd70530a, 32'h3c541578} /* (28, 13, 12) {real, imag} */,
  {32'h3d6e5ef9, 32'hbbf9858c} /* (28, 13, 11) {real, imag} */,
  {32'hbd766c08, 32'hbd89ca7e} /* (28, 13, 10) {real, imag} */,
  {32'h3d46acc8, 32'hbc9bef12} /* (28, 13, 9) {real, imag} */,
  {32'h3c5c1efc, 32'h3df55764} /* (28, 13, 8) {real, imag} */,
  {32'h3cddb730, 32'h3cf09f90} /* (28, 13, 7) {real, imag} */,
  {32'h3d9aed6b, 32'hbd4a7b39} /* (28, 13, 6) {real, imag} */,
  {32'h3e35f20b, 32'h3dc84d8f} /* (28, 13, 5) {real, imag} */,
  {32'hbe813238, 32'h3dc1970c} /* (28, 13, 4) {real, imag} */,
  {32'hbde36ba8, 32'hbc9a4cb0} /* (28, 13, 3) {real, imag} */,
  {32'h3f443763, 32'h3ccc18e0} /* (28, 13, 2) {real, imag} */,
  {32'hbfc7962a, 32'hbde8e5a2} /* (28, 13, 1) {real, imag} */,
  {32'hbf976e22, 32'h00000000} /* (28, 13, 0) {real, imag} */,
  {32'hbfb4db04, 32'h3e07d650} /* (28, 12, 31) {real, imag} */,
  {32'h3f13bc86, 32'hbc15d170} /* (28, 12, 30) {real, imag} */,
  {32'hb98cf200, 32'hbe030e43} /* (28, 12, 29) {real, imag} */,
  {32'hbe0c745a, 32'hbd678978} /* (28, 12, 28) {real, imag} */,
  {32'h3e238b1c, 32'hbe35dbff} /* (28, 12, 27) {real, imag} */,
  {32'h3ca691c9, 32'h3c210eb6} /* (28, 12, 26) {real, imag} */,
  {32'h3d91d1d4, 32'h3d090661} /* (28, 12, 25) {real, imag} */,
  {32'h3d8cb1a6, 32'hbd982250} /* (28, 12, 24) {real, imag} */,
  {32'h3cdb282c, 32'hbdc2c39c} /* (28, 12, 23) {real, imag} */,
  {32'hbcc43e18, 32'hbd3ce560} /* (28, 12, 22) {real, imag} */,
  {32'hbb863060, 32'hbda69c13} /* (28, 12, 21) {real, imag} */,
  {32'hbc9a43ce, 32'hbd4d4afa} /* (28, 12, 20) {real, imag} */,
  {32'h3c6f1664, 32'hbd559726} /* (28, 12, 19) {real, imag} */,
  {32'h3d4657ec, 32'hbdf82a74} /* (28, 12, 18) {real, imag} */,
  {32'hbd1a1615, 32'hbcbe6ab4} /* (28, 12, 17) {real, imag} */,
  {32'h3c9f3d67, 32'h00000000} /* (28, 12, 16) {real, imag} */,
  {32'hbd1a1615, 32'h3cbe6ab4} /* (28, 12, 15) {real, imag} */,
  {32'h3d4657ec, 32'h3df82a74} /* (28, 12, 14) {real, imag} */,
  {32'h3c6f1664, 32'h3d559726} /* (28, 12, 13) {real, imag} */,
  {32'hbc9a43ce, 32'h3d4d4afa} /* (28, 12, 12) {real, imag} */,
  {32'hbb863060, 32'h3da69c13} /* (28, 12, 11) {real, imag} */,
  {32'hbcc43e18, 32'h3d3ce560} /* (28, 12, 10) {real, imag} */,
  {32'h3cdb282c, 32'h3dc2c39c} /* (28, 12, 9) {real, imag} */,
  {32'h3d8cb1a6, 32'h3d982250} /* (28, 12, 8) {real, imag} */,
  {32'h3d91d1d4, 32'hbd090661} /* (28, 12, 7) {real, imag} */,
  {32'h3ca691c9, 32'hbc210eb6} /* (28, 12, 6) {real, imag} */,
  {32'h3e238b1c, 32'h3e35dbff} /* (28, 12, 5) {real, imag} */,
  {32'hbe0c745a, 32'h3d678978} /* (28, 12, 4) {real, imag} */,
  {32'hb98cf200, 32'h3e030e43} /* (28, 12, 3) {real, imag} */,
  {32'h3f13bc86, 32'h3c15d170} /* (28, 12, 2) {real, imag} */,
  {32'hbfb4db04, 32'hbe07d650} /* (28, 12, 1) {real, imag} */,
  {32'hbf9b57a8, 32'h00000000} /* (28, 12, 0) {real, imag} */,
  {32'hbf3eb820, 32'h3da06d2a} /* (28, 11, 31) {real, imag} */,
  {32'h3ede82ce, 32'hbd8345b0} /* (28, 11, 30) {real, imag} */,
  {32'h3bdc3b9c, 32'hbd27308e} /* (28, 11, 29) {real, imag} */,
  {32'hbd859845, 32'hbd78c801} /* (28, 11, 28) {real, imag} */,
  {32'h3c953f4e, 32'hbd84e476} /* (28, 11, 27) {real, imag} */,
  {32'hbdbefd8a, 32'hbd50cd42} /* (28, 11, 26) {real, imag} */,
  {32'h3c94b5a8, 32'hbdbe9d58} /* (28, 11, 25) {real, imag} */,
  {32'h3dac4636, 32'h3d43bbc2} /* (28, 11, 24) {real, imag} */,
  {32'h3d7b2c22, 32'h3d323078} /* (28, 11, 23) {real, imag} */,
  {32'h3d74339b, 32'h3cc5f6f2} /* (28, 11, 22) {real, imag} */,
  {32'h3c38b741, 32'hbc1677b0} /* (28, 11, 21) {real, imag} */,
  {32'h3c14fbd4, 32'h3d967ecb} /* (28, 11, 20) {real, imag} */,
  {32'hbd74e0d8, 32'h3bbc5ee0} /* (28, 11, 19) {real, imag} */,
  {32'hbb75fd30, 32'hbb377bc0} /* (28, 11, 18) {real, imag} */,
  {32'h3d206d99, 32'hbb34d078} /* (28, 11, 17) {real, imag} */,
  {32'hbdc9a405, 32'h00000000} /* (28, 11, 16) {real, imag} */,
  {32'h3d206d99, 32'h3b34d078} /* (28, 11, 15) {real, imag} */,
  {32'hbb75fd30, 32'h3b377bc0} /* (28, 11, 14) {real, imag} */,
  {32'hbd74e0d8, 32'hbbbc5ee0} /* (28, 11, 13) {real, imag} */,
  {32'h3c14fbd4, 32'hbd967ecb} /* (28, 11, 12) {real, imag} */,
  {32'h3c38b741, 32'h3c1677b0} /* (28, 11, 11) {real, imag} */,
  {32'h3d74339b, 32'hbcc5f6f2} /* (28, 11, 10) {real, imag} */,
  {32'h3d7b2c22, 32'hbd323078} /* (28, 11, 9) {real, imag} */,
  {32'h3dac4636, 32'hbd43bbc2} /* (28, 11, 8) {real, imag} */,
  {32'h3c94b5a8, 32'h3dbe9d58} /* (28, 11, 7) {real, imag} */,
  {32'hbdbefd8a, 32'h3d50cd42} /* (28, 11, 6) {real, imag} */,
  {32'h3c953f4e, 32'h3d84e476} /* (28, 11, 5) {real, imag} */,
  {32'hbd859845, 32'h3d78c801} /* (28, 11, 4) {real, imag} */,
  {32'h3bdc3b9c, 32'h3d27308e} /* (28, 11, 3) {real, imag} */,
  {32'h3ede82ce, 32'h3d8345b0} /* (28, 11, 2) {real, imag} */,
  {32'hbf3eb820, 32'hbda06d2a} /* (28, 11, 1) {real, imag} */,
  {32'hbf60886c, 32'h00000000} /* (28, 11, 0) {real, imag} */,
  {32'h3ec9b7dc, 32'hbdc91ca1} /* (28, 10, 31) {real, imag} */,
  {32'hbe8e77e4, 32'h3dd50bd2} /* (28, 10, 30) {real, imag} */,
  {32'h3cb43350, 32'h3dc110b9} /* (28, 10, 29) {real, imag} */,
  {32'h3e53203c, 32'hbe3a4392} /* (28, 10, 28) {real, imag} */,
  {32'hbe0103f2, 32'hbd0778b1} /* (28, 10, 27) {real, imag} */,
  {32'hbce6e4e5, 32'hbbfecd7c} /* (28, 10, 26) {real, imag} */,
  {32'h3ddf19ec, 32'hbaabac00} /* (28, 10, 25) {real, imag} */,
  {32'hbc9af524, 32'h3cd5491e} /* (28, 10, 24) {real, imag} */,
  {32'hbcc57af5, 32'h3c6f731c} /* (28, 10, 23) {real, imag} */,
  {32'hbb9d405c, 32'hbdc4e615} /* (28, 10, 22) {real, imag} */,
  {32'hbe00e845, 32'h3d9ebc12} /* (28, 10, 21) {real, imag} */,
  {32'h3dcbc56b, 32'hbd4b2c8c} /* (28, 10, 20) {real, imag} */,
  {32'h3b962994, 32'h3c6168c0} /* (28, 10, 19) {real, imag} */,
  {32'hbcc59203, 32'hbc0b75a0} /* (28, 10, 18) {real, imag} */,
  {32'h3b836adc, 32'h3d2409a5} /* (28, 10, 17) {real, imag} */,
  {32'hbc01f1bc, 32'h00000000} /* (28, 10, 16) {real, imag} */,
  {32'h3b836adc, 32'hbd2409a5} /* (28, 10, 15) {real, imag} */,
  {32'hbcc59203, 32'h3c0b75a0} /* (28, 10, 14) {real, imag} */,
  {32'h3b962994, 32'hbc6168c0} /* (28, 10, 13) {real, imag} */,
  {32'h3dcbc56b, 32'h3d4b2c8c} /* (28, 10, 12) {real, imag} */,
  {32'hbe00e845, 32'hbd9ebc12} /* (28, 10, 11) {real, imag} */,
  {32'hbb9d405c, 32'h3dc4e615} /* (28, 10, 10) {real, imag} */,
  {32'hbcc57af5, 32'hbc6f731c} /* (28, 10, 9) {real, imag} */,
  {32'hbc9af524, 32'hbcd5491e} /* (28, 10, 8) {real, imag} */,
  {32'h3ddf19ec, 32'h3aabac00} /* (28, 10, 7) {real, imag} */,
  {32'hbce6e4e5, 32'h3bfecd7c} /* (28, 10, 6) {real, imag} */,
  {32'hbe0103f2, 32'h3d0778b1} /* (28, 10, 5) {real, imag} */,
  {32'h3e53203c, 32'h3e3a4392} /* (28, 10, 4) {real, imag} */,
  {32'h3cb43350, 32'hbdc110b9} /* (28, 10, 3) {real, imag} */,
  {32'hbe8e77e4, 32'hbdd50bd2} /* (28, 10, 2) {real, imag} */,
  {32'h3ec9b7dc, 32'h3dc91ca1} /* (28, 10, 1) {real, imag} */,
  {32'hbd9e9ec8, 32'h00000000} /* (28, 10, 0) {real, imag} */,
  {32'h3f8feaa6, 32'hbdfa4f92} /* (28, 9, 31) {real, imag} */,
  {32'hbf1fa5be, 32'h3e17a9df} /* (28, 9, 30) {real, imag} */,
  {32'h3dfa53d0, 32'h3dd17d4f} /* (28, 9, 29) {real, imag} */,
  {32'h3e17f8d5, 32'hbe327a1c} /* (28, 9, 28) {real, imag} */,
  {32'hbe569f8d, 32'h3d4a829c} /* (28, 9, 27) {real, imag} */,
  {32'hbdbdbd44, 32'hbe1e8720} /* (28, 9, 26) {real, imag} */,
  {32'h3db0eb49, 32'hbd652418} /* (28, 9, 25) {real, imag} */,
  {32'hbd90c9f6, 32'h3cee3b08} /* (28, 9, 24) {real, imag} */,
  {32'h3d35a4e1, 32'hbd27a0f8} /* (28, 9, 23) {real, imag} */,
  {32'hbad43cc0, 32'hbddb7d56} /* (28, 9, 22) {real, imag} */,
  {32'hbdb3ae2f, 32'h3e1cc365} /* (28, 9, 21) {real, imag} */,
  {32'h3bf28e20, 32'hbbce06fc} /* (28, 9, 20) {real, imag} */,
  {32'hbcdcb383, 32'hbc677d4c} /* (28, 9, 19) {real, imag} */,
  {32'h3cdba9fe, 32'hbd4fc501} /* (28, 9, 18) {real, imag} */,
  {32'hbced7876, 32'hbc12ac04} /* (28, 9, 17) {real, imag} */,
  {32'hbcc8e472, 32'h00000000} /* (28, 9, 16) {real, imag} */,
  {32'hbced7876, 32'h3c12ac04} /* (28, 9, 15) {real, imag} */,
  {32'h3cdba9fe, 32'h3d4fc501} /* (28, 9, 14) {real, imag} */,
  {32'hbcdcb383, 32'h3c677d4c} /* (28, 9, 13) {real, imag} */,
  {32'h3bf28e20, 32'h3bce06fc} /* (28, 9, 12) {real, imag} */,
  {32'hbdb3ae2f, 32'hbe1cc365} /* (28, 9, 11) {real, imag} */,
  {32'hbad43cc0, 32'h3ddb7d56} /* (28, 9, 10) {real, imag} */,
  {32'h3d35a4e1, 32'h3d27a0f8} /* (28, 9, 9) {real, imag} */,
  {32'hbd90c9f6, 32'hbcee3b08} /* (28, 9, 8) {real, imag} */,
  {32'h3db0eb49, 32'h3d652418} /* (28, 9, 7) {real, imag} */,
  {32'hbdbdbd44, 32'h3e1e8720} /* (28, 9, 6) {real, imag} */,
  {32'hbe569f8d, 32'hbd4a829c} /* (28, 9, 5) {real, imag} */,
  {32'h3e17f8d5, 32'h3e327a1c} /* (28, 9, 4) {real, imag} */,
  {32'h3dfa53d0, 32'hbdd17d4f} /* (28, 9, 3) {real, imag} */,
  {32'hbf1fa5be, 32'hbe17a9df} /* (28, 9, 2) {real, imag} */,
  {32'h3f8feaa6, 32'h3dfa4f92} /* (28, 9, 1) {real, imag} */,
  {32'h3effed35, 32'h00000000} /* (28, 9, 0) {real, imag} */,
  {32'h3fb1c2b4, 32'hbe38f064} /* (28, 8, 31) {real, imag} */,
  {32'hbf1b3104, 32'h3e93a8ea} /* (28, 8, 30) {real, imag} */,
  {32'h3e169538, 32'h3d5f7da0} /* (28, 8, 29) {real, imag} */,
  {32'h3e209392, 32'hbda8e2c8} /* (28, 8, 28) {real, imag} */,
  {32'hbe1a6813, 32'h3e39165b} /* (28, 8, 27) {real, imag} */,
  {32'h3d5051ac, 32'hbdcc033c} /* (28, 8, 26) {real, imag} */,
  {32'hbd446596, 32'h3cf97458} /* (28, 8, 25) {real, imag} */,
  {32'hbd65bf04, 32'h3c8d3fd4} /* (28, 8, 24) {real, imag} */,
  {32'hbdb480d1, 32'h3d4e49fa} /* (28, 8, 23) {real, imag} */,
  {32'h3de7094a, 32'hbbab2cae} /* (28, 8, 22) {real, imag} */,
  {32'hbaa21e80, 32'h3d103fa4} /* (28, 8, 21) {real, imag} */,
  {32'hbd37f355, 32'hbd5f984b} /* (28, 8, 20) {real, imag} */,
  {32'h3c8a59b0, 32'hbdbcfc58} /* (28, 8, 19) {real, imag} */,
  {32'hbdb792a2, 32'h3d712bd2} /* (28, 8, 18) {real, imag} */,
  {32'hbcf0c014, 32'h3b4bfc10} /* (28, 8, 17) {real, imag} */,
  {32'hbce35c03, 32'h00000000} /* (28, 8, 16) {real, imag} */,
  {32'hbcf0c014, 32'hbb4bfc10} /* (28, 8, 15) {real, imag} */,
  {32'hbdb792a2, 32'hbd712bd2} /* (28, 8, 14) {real, imag} */,
  {32'h3c8a59b0, 32'h3dbcfc58} /* (28, 8, 13) {real, imag} */,
  {32'hbd37f355, 32'h3d5f984b} /* (28, 8, 12) {real, imag} */,
  {32'hbaa21e80, 32'hbd103fa4} /* (28, 8, 11) {real, imag} */,
  {32'h3de7094a, 32'h3bab2cae} /* (28, 8, 10) {real, imag} */,
  {32'hbdb480d1, 32'hbd4e49fa} /* (28, 8, 9) {real, imag} */,
  {32'hbd65bf04, 32'hbc8d3fd4} /* (28, 8, 8) {real, imag} */,
  {32'hbd446596, 32'hbcf97458} /* (28, 8, 7) {real, imag} */,
  {32'h3d5051ac, 32'h3dcc033c} /* (28, 8, 6) {real, imag} */,
  {32'hbe1a6813, 32'hbe39165b} /* (28, 8, 5) {real, imag} */,
  {32'h3e209392, 32'h3da8e2c8} /* (28, 8, 4) {real, imag} */,
  {32'h3e169538, 32'hbd5f7da0} /* (28, 8, 3) {real, imag} */,
  {32'hbf1b3104, 32'hbe93a8ea} /* (28, 8, 2) {real, imag} */,
  {32'h3fb1c2b4, 32'h3e38f064} /* (28, 8, 1) {real, imag} */,
  {32'h3ef993e8, 32'h00000000} /* (28, 8, 0) {real, imag} */,
  {32'h3fba4d48, 32'hbe79e26d} /* (28, 7, 31) {real, imag} */,
  {32'hbf308cc3, 32'h3ed5dc22} /* (28, 7, 30) {real, imag} */,
  {32'h3bff50f0, 32'h3e3c75ce} /* (28, 7, 29) {real, imag} */,
  {32'h3e21db47, 32'hbd05613c} /* (28, 7, 28) {real, imag} */,
  {32'hbe144ffb, 32'h3bee7e80} /* (28, 7, 27) {real, imag} */,
  {32'hbd6fcee1, 32'hbd051b5e} /* (28, 7, 26) {real, imag} */,
  {32'hbd73d22d, 32'hbda9c3a0} /* (28, 7, 25) {real, imag} */,
  {32'hbc4b3cf2, 32'h3dd3890e} /* (28, 7, 24) {real, imag} */,
  {32'h3c8a9286, 32'hba3bd580} /* (28, 7, 23) {real, imag} */,
  {32'hbdf80265, 32'hbc31a52c} /* (28, 7, 22) {real, imag} */,
  {32'hbd49cd06, 32'h3d6e98df} /* (28, 7, 21) {real, imag} */,
  {32'h3dec69a6, 32'hbd429722} /* (28, 7, 20) {real, imag} */,
  {32'hbd996740, 32'hbc71788c} /* (28, 7, 19) {real, imag} */,
  {32'h3d83c608, 32'h3c1b606e} /* (28, 7, 18) {real, imag} */,
  {32'hbd5c313a, 32'h3ccbe8ee} /* (28, 7, 17) {real, imag} */,
  {32'h3dad69be, 32'h00000000} /* (28, 7, 16) {real, imag} */,
  {32'hbd5c313a, 32'hbccbe8ee} /* (28, 7, 15) {real, imag} */,
  {32'h3d83c608, 32'hbc1b606e} /* (28, 7, 14) {real, imag} */,
  {32'hbd996740, 32'h3c71788c} /* (28, 7, 13) {real, imag} */,
  {32'h3dec69a6, 32'h3d429722} /* (28, 7, 12) {real, imag} */,
  {32'hbd49cd06, 32'hbd6e98df} /* (28, 7, 11) {real, imag} */,
  {32'hbdf80265, 32'h3c31a52c} /* (28, 7, 10) {real, imag} */,
  {32'h3c8a9286, 32'h3a3bd580} /* (28, 7, 9) {real, imag} */,
  {32'hbc4b3cf2, 32'hbdd3890e} /* (28, 7, 8) {real, imag} */,
  {32'hbd73d22d, 32'h3da9c3a0} /* (28, 7, 7) {real, imag} */,
  {32'hbd6fcee1, 32'h3d051b5e} /* (28, 7, 6) {real, imag} */,
  {32'hbe144ffb, 32'hbbee7e80} /* (28, 7, 5) {real, imag} */,
  {32'h3e21db47, 32'h3d05613c} /* (28, 7, 4) {real, imag} */,
  {32'h3bff50f0, 32'hbe3c75ce} /* (28, 7, 3) {real, imag} */,
  {32'hbf308cc3, 32'hbed5dc22} /* (28, 7, 2) {real, imag} */,
  {32'h3fba4d48, 32'h3e79e26d} /* (28, 7, 1) {real, imag} */,
  {32'h3efc9073, 32'h00000000} /* (28, 7, 0) {real, imag} */,
  {32'h3fa9b921, 32'hbedc5ba1} /* (28, 6, 31) {real, imag} */,
  {32'hbf244ea2, 32'h3f09926d} /* (28, 6, 30) {real, imag} */,
  {32'hbdb670a6, 32'h3dcd7419} /* (28, 6, 29) {real, imag} */,
  {32'h3b787160, 32'hbb8e0410} /* (28, 6, 28) {real, imag} */,
  {32'hbe7ab7bf, 32'h3ce41880} /* (28, 6, 27) {real, imag} */,
  {32'h3dd85c96, 32'hbe0964ee} /* (28, 6, 26) {real, imag} */,
  {32'hbb8a5bb8, 32'hbe2e30f4} /* (28, 6, 25) {real, imag} */,
  {32'hbc03c025, 32'h3d2a498a} /* (28, 6, 24) {real, imag} */,
  {32'h3daea39f, 32'h3d649ddf} /* (28, 6, 23) {real, imag} */,
  {32'h3d44c35e, 32'h3d0ad18e} /* (28, 6, 22) {real, imag} */,
  {32'hbd0a4d7c, 32'hbb981d9c} /* (28, 6, 21) {real, imag} */,
  {32'hbd4aaffe, 32'hbb0d85f8} /* (28, 6, 20) {real, imag} */,
  {32'hbd034170, 32'hbcb78c2e} /* (28, 6, 19) {real, imag} */,
  {32'hbc990f98, 32'hbd59d0e7} /* (28, 6, 18) {real, imag} */,
  {32'h3c3bc7c0, 32'hbd163804} /* (28, 6, 17) {real, imag} */,
  {32'hbba48c44, 32'h00000000} /* (28, 6, 16) {real, imag} */,
  {32'h3c3bc7c0, 32'h3d163804} /* (28, 6, 15) {real, imag} */,
  {32'hbc990f98, 32'h3d59d0e7} /* (28, 6, 14) {real, imag} */,
  {32'hbd034170, 32'h3cb78c2e} /* (28, 6, 13) {real, imag} */,
  {32'hbd4aaffe, 32'h3b0d85f8} /* (28, 6, 12) {real, imag} */,
  {32'hbd0a4d7c, 32'h3b981d9c} /* (28, 6, 11) {real, imag} */,
  {32'h3d44c35e, 32'hbd0ad18e} /* (28, 6, 10) {real, imag} */,
  {32'h3daea39f, 32'hbd649ddf} /* (28, 6, 9) {real, imag} */,
  {32'hbc03c025, 32'hbd2a498a} /* (28, 6, 8) {real, imag} */,
  {32'hbb8a5bb8, 32'h3e2e30f4} /* (28, 6, 7) {real, imag} */,
  {32'h3dd85c96, 32'h3e0964ee} /* (28, 6, 6) {real, imag} */,
  {32'hbe7ab7bf, 32'hbce41880} /* (28, 6, 5) {real, imag} */,
  {32'h3b787160, 32'h3b8e0410} /* (28, 6, 4) {real, imag} */,
  {32'hbdb670a6, 32'hbdcd7419} /* (28, 6, 3) {real, imag} */,
  {32'hbf244ea2, 32'hbf09926d} /* (28, 6, 2) {real, imag} */,
  {32'h3fa9b921, 32'h3edc5ba1} /* (28, 6, 1) {real, imag} */,
  {32'h3f1b7c22, 32'h00000000} /* (28, 6, 0) {real, imag} */,
  {32'h3f72f530, 32'hbf6f78f7} /* (28, 5, 31) {real, imag} */,
  {32'hbe745edc, 32'h3f3a0623} /* (28, 5, 30) {real, imag} */,
  {32'hbe002d79, 32'h3d2ff21e} /* (28, 5, 29) {real, imag} */,
  {32'hbda00f74, 32'h3d07d995} /* (28, 5, 28) {real, imag} */,
  {32'hbdf7e18a, 32'h3d327eba} /* (28, 5, 27) {real, imag} */,
  {32'h3c676aac, 32'hbdcb9469} /* (28, 5, 26) {real, imag} */,
  {32'h3cabb09a, 32'hbd21de39} /* (28, 5, 25) {real, imag} */,
  {32'h3da823f3, 32'h3d52293e} /* (28, 5, 24) {real, imag} */,
  {32'hbd66b57e, 32'h3d1e7c71} /* (28, 5, 23) {real, imag} */,
  {32'hbda093b2, 32'hbd21ad58} /* (28, 5, 22) {real, imag} */,
  {32'h3db4aade, 32'h3d39f914} /* (28, 5, 21) {real, imag} */,
  {32'h3ae2b5dc, 32'hbcc0e5f8} /* (28, 5, 20) {real, imag} */,
  {32'h3d4278c6, 32'h3beb7940} /* (28, 5, 19) {real, imag} */,
  {32'h3c923a08, 32'h3d80bb48} /* (28, 5, 18) {real, imag} */,
  {32'hbd212d4a, 32'hbc2b2448} /* (28, 5, 17) {real, imag} */,
  {32'hbd108a04, 32'h00000000} /* (28, 5, 16) {real, imag} */,
  {32'hbd212d4a, 32'h3c2b2448} /* (28, 5, 15) {real, imag} */,
  {32'h3c923a08, 32'hbd80bb48} /* (28, 5, 14) {real, imag} */,
  {32'h3d4278c6, 32'hbbeb7940} /* (28, 5, 13) {real, imag} */,
  {32'h3ae2b5dc, 32'h3cc0e5f8} /* (28, 5, 12) {real, imag} */,
  {32'h3db4aade, 32'hbd39f914} /* (28, 5, 11) {real, imag} */,
  {32'hbda093b2, 32'h3d21ad58} /* (28, 5, 10) {real, imag} */,
  {32'hbd66b57e, 32'hbd1e7c71} /* (28, 5, 9) {real, imag} */,
  {32'h3da823f3, 32'hbd52293e} /* (28, 5, 8) {real, imag} */,
  {32'h3cabb09a, 32'h3d21de39} /* (28, 5, 7) {real, imag} */,
  {32'h3c676aac, 32'h3dcb9469} /* (28, 5, 6) {real, imag} */,
  {32'hbdf7e18a, 32'hbd327eba} /* (28, 5, 5) {real, imag} */,
  {32'hbda00f74, 32'hbd07d995} /* (28, 5, 4) {real, imag} */,
  {32'hbe002d79, 32'hbd2ff21e} /* (28, 5, 3) {real, imag} */,
  {32'hbe745edc, 32'hbf3a0623} /* (28, 5, 2) {real, imag} */,
  {32'h3f72f530, 32'h3f6f78f7} /* (28, 5, 1) {real, imag} */,
  {32'h3f371df0, 32'h00000000} /* (28, 5, 0) {real, imag} */,
  {32'h3f1481cf, 32'hbf7dd97e} /* (28, 4, 31) {real, imag} */,
  {32'h3e731362, 32'h3f417651} /* (28, 4, 30) {real, imag} */,
  {32'hbd92c620, 32'hbd850a8b} /* (28, 4, 29) {real, imag} */,
  {32'hbe0dce06, 32'h3dbfb086} /* (28, 4, 28) {real, imag} */,
  {32'hbe802238, 32'hbdc097e2} /* (28, 4, 27) {real, imag} */,
  {32'hbd9e7926, 32'h3dc6a92d} /* (28, 4, 26) {real, imag} */,
  {32'h3cb5559c, 32'hbd73288a} /* (28, 4, 25) {real, imag} */,
  {32'h3d41908f, 32'h3d442de5} /* (28, 4, 24) {real, imag} */,
  {32'hbd804763, 32'hbd0f2a1a} /* (28, 4, 23) {real, imag} */,
  {32'hbdd50bfa, 32'hbce8352c} /* (28, 4, 22) {real, imag} */,
  {32'h3cb4989c, 32'h3c7961b8} /* (28, 4, 21) {real, imag} */,
  {32'h3d13a655, 32'hbd0c23a7} /* (28, 4, 20) {real, imag} */,
  {32'hbcc2322d, 32'hbdd7d7e3} /* (28, 4, 19) {real, imag} */,
  {32'h3d855b2d, 32'h3d4924b0} /* (28, 4, 18) {real, imag} */,
  {32'h39b82580, 32'h3c077248} /* (28, 4, 17) {real, imag} */,
  {32'h3be1be68, 32'h00000000} /* (28, 4, 16) {real, imag} */,
  {32'h39b82580, 32'hbc077248} /* (28, 4, 15) {real, imag} */,
  {32'h3d855b2d, 32'hbd4924b0} /* (28, 4, 14) {real, imag} */,
  {32'hbcc2322d, 32'h3dd7d7e3} /* (28, 4, 13) {real, imag} */,
  {32'h3d13a655, 32'h3d0c23a7} /* (28, 4, 12) {real, imag} */,
  {32'h3cb4989c, 32'hbc7961b8} /* (28, 4, 11) {real, imag} */,
  {32'hbdd50bfa, 32'h3ce8352c} /* (28, 4, 10) {real, imag} */,
  {32'hbd804763, 32'h3d0f2a1a} /* (28, 4, 9) {real, imag} */,
  {32'h3d41908f, 32'hbd442de5} /* (28, 4, 8) {real, imag} */,
  {32'h3cb5559c, 32'h3d73288a} /* (28, 4, 7) {real, imag} */,
  {32'hbd9e7926, 32'hbdc6a92d} /* (28, 4, 6) {real, imag} */,
  {32'hbe802238, 32'h3dc097e2} /* (28, 4, 5) {real, imag} */,
  {32'hbe0dce06, 32'hbdbfb086} /* (28, 4, 4) {real, imag} */,
  {32'hbd92c620, 32'h3d850a8b} /* (28, 4, 3) {real, imag} */,
  {32'h3e731362, 32'hbf417651} /* (28, 4, 2) {real, imag} */,
  {32'h3f1481cf, 32'h3f7dd97e} /* (28, 4, 1) {real, imag} */,
  {32'h3eeab082, 32'h00000000} /* (28, 4, 0) {real, imag} */,
  {32'h3efc6528, 32'hbf9529fc} /* (28, 3, 31) {real, imag} */,
  {32'h3ed6ad28, 32'h3f23b55e} /* (28, 3, 30) {real, imag} */,
  {32'hbde4beb7, 32'hbe0a5510} /* (28, 3, 29) {real, imag} */,
  {32'hbdf7fd9b, 32'h3e8bfef8} /* (28, 3, 28) {real, imag} */,
  {32'hbe808ee1, 32'h3de1232d} /* (28, 3, 27) {real, imag} */,
  {32'hbc0f86fe, 32'h3e1a0b38} /* (28, 3, 26) {real, imag} */,
  {32'hbda9012e, 32'hbd40ec12} /* (28, 3, 25) {real, imag} */,
  {32'h3d0cbdda, 32'hbd462967} /* (28, 3, 24) {real, imag} */,
  {32'hbc81e1a4, 32'hbd2f88f6} /* (28, 3, 23) {real, imag} */,
  {32'hbc88d4dc, 32'h3d8f131f} /* (28, 3, 22) {real, imag} */,
  {32'hbda10e24, 32'hbd921858} /* (28, 3, 21) {real, imag} */,
  {32'hbccec0e2, 32'hbc87b56a} /* (28, 3, 20) {real, imag} */,
  {32'hbc8f1b73, 32'h3bd32c68} /* (28, 3, 19) {real, imag} */,
  {32'h3d9157d6, 32'hbc8a4fd9} /* (28, 3, 18) {real, imag} */,
  {32'hbc65541b, 32'h3d6548ce} /* (28, 3, 17) {real, imag} */,
  {32'h3c80b9ee, 32'h00000000} /* (28, 3, 16) {real, imag} */,
  {32'hbc65541b, 32'hbd6548ce} /* (28, 3, 15) {real, imag} */,
  {32'h3d9157d6, 32'h3c8a4fd9} /* (28, 3, 14) {real, imag} */,
  {32'hbc8f1b73, 32'hbbd32c68} /* (28, 3, 13) {real, imag} */,
  {32'hbccec0e2, 32'h3c87b56a} /* (28, 3, 12) {real, imag} */,
  {32'hbda10e24, 32'h3d921858} /* (28, 3, 11) {real, imag} */,
  {32'hbc88d4dc, 32'hbd8f131f} /* (28, 3, 10) {real, imag} */,
  {32'hbc81e1a4, 32'h3d2f88f6} /* (28, 3, 9) {real, imag} */,
  {32'h3d0cbdda, 32'h3d462967} /* (28, 3, 8) {real, imag} */,
  {32'hbda9012e, 32'h3d40ec12} /* (28, 3, 7) {real, imag} */,
  {32'hbc0f86fe, 32'hbe1a0b38} /* (28, 3, 6) {real, imag} */,
  {32'hbe808ee1, 32'hbde1232d} /* (28, 3, 5) {real, imag} */,
  {32'hbdf7fd9b, 32'hbe8bfef8} /* (28, 3, 4) {real, imag} */,
  {32'hbde4beb7, 32'h3e0a5510} /* (28, 3, 3) {real, imag} */,
  {32'h3ed6ad28, 32'hbf23b55e} /* (28, 3, 2) {real, imag} */,
  {32'h3efc6528, 32'h3f9529fc} /* (28, 3, 1) {real, imag} */,
  {32'h3eee52b9, 32'h00000000} /* (28, 3, 0) {real, imag} */,
  {32'h3ee045eb, 32'hbfb33540} /* (28, 2, 31) {real, imag} */,
  {32'h3ea24e4e, 32'h3f3a4f90} /* (28, 2, 30) {real, imag} */,
  {32'hbca1c890, 32'h3d690570} /* (28, 2, 29) {real, imag} */,
  {32'hbdf8d4fe, 32'h3e0aa7ce} /* (28, 2, 28) {real, imag} */,
  {32'hbd63d697, 32'hbd809f84} /* (28, 2, 27) {real, imag} */,
  {32'hbcf59fc8, 32'h3de7c2ec} /* (28, 2, 26) {real, imag} */,
  {32'hbe41f8a0, 32'hbcea8efa} /* (28, 2, 25) {real, imag} */,
  {32'h3e135e58, 32'hbdf49e50} /* (28, 2, 24) {real, imag} */,
  {32'hbd2fc5b4, 32'h3ba7d866} /* (28, 2, 23) {real, imag} */,
  {32'hbd0de586, 32'h3e0a3439} /* (28, 2, 22) {real, imag} */,
  {32'hbcdf5364, 32'hbd2e98fe} /* (28, 2, 21) {real, imag} */,
  {32'h3dd28704, 32'h3db5bed4} /* (28, 2, 20) {real, imag} */,
  {32'h3c84bd5e, 32'h3cabaf96} /* (28, 2, 19) {real, imag} */,
  {32'h3c33ac32, 32'h3aa131b0} /* (28, 2, 18) {real, imag} */,
  {32'hbd7c7400, 32'h3d01cba2} /* (28, 2, 17) {real, imag} */,
  {32'h3d9cf039, 32'h00000000} /* (28, 2, 16) {real, imag} */,
  {32'hbd7c7400, 32'hbd01cba2} /* (28, 2, 15) {real, imag} */,
  {32'h3c33ac32, 32'hbaa131b0} /* (28, 2, 14) {real, imag} */,
  {32'h3c84bd5e, 32'hbcabaf96} /* (28, 2, 13) {real, imag} */,
  {32'h3dd28704, 32'hbdb5bed4} /* (28, 2, 12) {real, imag} */,
  {32'hbcdf5364, 32'h3d2e98fe} /* (28, 2, 11) {real, imag} */,
  {32'hbd0de586, 32'hbe0a3439} /* (28, 2, 10) {real, imag} */,
  {32'hbd2fc5b4, 32'hbba7d866} /* (28, 2, 9) {real, imag} */,
  {32'h3e135e58, 32'h3df49e50} /* (28, 2, 8) {real, imag} */,
  {32'hbe41f8a0, 32'h3cea8efa} /* (28, 2, 7) {real, imag} */,
  {32'hbcf59fc8, 32'hbde7c2ec} /* (28, 2, 6) {real, imag} */,
  {32'hbd63d697, 32'h3d809f84} /* (28, 2, 5) {real, imag} */,
  {32'hbdf8d4fe, 32'hbe0aa7ce} /* (28, 2, 4) {real, imag} */,
  {32'hbca1c890, 32'hbd690570} /* (28, 2, 3) {real, imag} */,
  {32'h3ea24e4e, 32'hbf3a4f90} /* (28, 2, 2) {real, imag} */,
  {32'h3ee045eb, 32'h3fb33540} /* (28, 2, 1) {real, imag} */,
  {32'h3e7ff914, 32'h00000000} /* (28, 2, 0) {real, imag} */,
  {32'h3e7c1e36, 32'hbfa45798} /* (28, 1, 31) {real, imag} */,
  {32'h3e8e691d, 32'h3f5a6975} /* (28, 1, 30) {real, imag} */,
  {32'hbd9ca86c, 32'h3c666372} /* (28, 1, 29) {real, imag} */,
  {32'h3cfcee46, 32'h3d9caf3e} /* (28, 1, 28) {real, imag} */,
  {32'hbe539d83, 32'hbdf76442} /* (28, 1, 27) {real, imag} */,
  {32'hbc0ba4d6, 32'h3e32fd9c} /* (28, 1, 26) {real, imag} */,
  {32'hbd676a1b, 32'hbdb09d02} /* (28, 1, 25) {real, imag} */,
  {32'h3cf20306, 32'hbd9e6c5a} /* (28, 1, 24) {real, imag} */,
  {32'h3d23836c, 32'h3d669cff} /* (28, 1, 23) {real, imag} */,
  {32'hbdb2b54e, 32'h3d6197d0} /* (28, 1, 22) {real, imag} */,
  {32'h3c974e47, 32'hbd849da7} /* (28, 1, 21) {real, imag} */,
  {32'h3de2ac7b, 32'h3c140054} /* (28, 1, 20) {real, imag} */,
  {32'hbdca8720, 32'hbc94a3bf} /* (28, 1, 19) {real, imag} */,
  {32'h3ad92060, 32'hbca27e02} /* (28, 1, 18) {real, imag} */,
  {32'hbd02228e, 32'hbd78762a} /* (28, 1, 17) {real, imag} */,
  {32'hbc041756, 32'h00000000} /* (28, 1, 16) {real, imag} */,
  {32'hbd02228e, 32'h3d78762a} /* (28, 1, 15) {real, imag} */,
  {32'h3ad92060, 32'h3ca27e02} /* (28, 1, 14) {real, imag} */,
  {32'hbdca8720, 32'h3c94a3bf} /* (28, 1, 13) {real, imag} */,
  {32'h3de2ac7b, 32'hbc140054} /* (28, 1, 12) {real, imag} */,
  {32'h3c974e47, 32'h3d849da7} /* (28, 1, 11) {real, imag} */,
  {32'hbdb2b54e, 32'hbd6197d0} /* (28, 1, 10) {real, imag} */,
  {32'h3d23836c, 32'hbd669cff} /* (28, 1, 9) {real, imag} */,
  {32'h3cf20306, 32'h3d9e6c5a} /* (28, 1, 8) {real, imag} */,
  {32'hbd676a1b, 32'h3db09d02} /* (28, 1, 7) {real, imag} */,
  {32'hbc0ba4d6, 32'hbe32fd9c} /* (28, 1, 6) {real, imag} */,
  {32'hbe539d83, 32'h3df76442} /* (28, 1, 5) {real, imag} */,
  {32'h3cfcee46, 32'hbd9caf3e} /* (28, 1, 4) {real, imag} */,
  {32'hbd9ca86c, 32'hbc666372} /* (28, 1, 3) {real, imag} */,
  {32'h3e8e691d, 32'hbf5a6975} /* (28, 1, 2) {real, imag} */,
  {32'h3e7c1e36, 32'h3fa45798} /* (28, 1, 1) {real, imag} */,
  {32'h3e57346e, 32'h00000000} /* (28, 1, 0) {real, imag} */,
  {32'h3e9e1560, 32'hbf50d1c3} /* (28, 0, 31) {real, imag} */,
  {32'hbca37d10, 32'h3f287722} /* (28, 0, 30) {real, imag} */,
  {32'hbcf20efc, 32'hbd9f58e8} /* (28, 0, 29) {real, imag} */,
  {32'h3d49f8e6, 32'h3e05261b} /* (28, 0, 28) {real, imag} */,
  {32'hbe1fa41f, 32'hbc1d6fb0} /* (28, 0, 27) {real, imag} */,
  {32'hbd6d8f90, 32'hbd46fe7e} /* (28, 0, 26) {real, imag} */,
  {32'h3d4d3fdb, 32'h3c636396} /* (28, 0, 25) {real, imag} */,
  {32'h3b413740, 32'h3d9ce1f0} /* (28, 0, 24) {real, imag} */,
  {32'hbbcb0448, 32'hbd6eb256} /* (28, 0, 23) {real, imag} */,
  {32'h3d077988, 32'h3d328fa9} /* (28, 0, 22) {real, imag} */,
  {32'hbdaaecf2, 32'hbccb98b8} /* (28, 0, 21) {real, imag} */,
  {32'h3d5dabb8, 32'h3ad1ee48} /* (28, 0, 20) {real, imag} */,
  {32'hbc64ac54, 32'hbb659cd0} /* (28, 0, 19) {real, imag} */,
  {32'h3cca6c55, 32'h3c0bc596} /* (28, 0, 18) {real, imag} */,
  {32'h3bba24d0, 32'hbd24ab08} /* (28, 0, 17) {real, imag} */,
  {32'h3bb4754c, 32'h00000000} /* (28, 0, 16) {real, imag} */,
  {32'h3bba24d0, 32'h3d24ab08} /* (28, 0, 15) {real, imag} */,
  {32'h3cca6c55, 32'hbc0bc596} /* (28, 0, 14) {real, imag} */,
  {32'hbc64ac54, 32'h3b659cd0} /* (28, 0, 13) {real, imag} */,
  {32'h3d5dabb8, 32'hbad1ee48} /* (28, 0, 12) {real, imag} */,
  {32'hbdaaecf2, 32'h3ccb98b8} /* (28, 0, 11) {real, imag} */,
  {32'h3d077988, 32'hbd328fa9} /* (28, 0, 10) {real, imag} */,
  {32'hbbcb0448, 32'h3d6eb256} /* (28, 0, 9) {real, imag} */,
  {32'h3b413740, 32'hbd9ce1f0} /* (28, 0, 8) {real, imag} */,
  {32'h3d4d3fdb, 32'hbc636396} /* (28, 0, 7) {real, imag} */,
  {32'hbd6d8f90, 32'h3d46fe7e} /* (28, 0, 6) {real, imag} */,
  {32'hbe1fa41f, 32'h3c1d6fb0} /* (28, 0, 5) {real, imag} */,
  {32'h3d49f8e6, 32'hbe05261b} /* (28, 0, 4) {real, imag} */,
  {32'hbcf20efc, 32'h3d9f58e8} /* (28, 0, 3) {real, imag} */,
  {32'hbca37d10, 32'hbf287722} /* (28, 0, 2) {real, imag} */,
  {32'h3e9e1560, 32'h3f50d1c3} /* (28, 0, 1) {real, imag} */,
  {32'h3cb11a40, 32'h00000000} /* (28, 0, 0) {real, imag} */,
  {32'h3e1b5c29, 32'hbd752780} /* (27, 31, 31) {real, imag} */,
  {32'hbe90b6d6, 32'h3ed6fd1b} /* (27, 31, 30) {real, imag} */,
  {32'hbe182dd0, 32'hbb847204} /* (27, 31, 29) {real, imag} */,
  {32'h3e0529ec, 32'h3e3cb236} /* (27, 31, 28) {real, imag} */,
  {32'hbde7a235, 32'h3d43f234} /* (27, 31, 27) {real, imag} */,
  {32'h3d386360, 32'hbcda9e7d} /* (27, 31, 26) {real, imag} */,
  {32'h3b90ea78, 32'h3d825b28} /* (27, 31, 25) {real, imag} */,
  {32'h3b615340, 32'h3d579078} /* (27, 31, 24) {real, imag} */,
  {32'hbd1ce11e, 32'h3d2e3d53} /* (27, 31, 23) {real, imag} */,
  {32'hbda7cd1c, 32'hbd8987e8} /* (27, 31, 22) {real, imag} */,
  {32'hbd439bb6, 32'hbcbf1dae} /* (27, 31, 21) {real, imag} */,
  {32'hbda44412, 32'h3c4dbff0} /* (27, 31, 20) {real, imag} */,
  {32'h38e4ec00, 32'h39856da0} /* (27, 31, 19) {real, imag} */,
  {32'h3c46da00, 32'hbc71012a} /* (27, 31, 18) {real, imag} */,
  {32'h3c197e08, 32'hbdad5b7b} /* (27, 31, 17) {real, imag} */,
  {32'h3d53aaa8, 32'h00000000} /* (27, 31, 16) {real, imag} */,
  {32'h3c197e08, 32'h3dad5b7b} /* (27, 31, 15) {real, imag} */,
  {32'h3c46da00, 32'h3c71012a} /* (27, 31, 14) {real, imag} */,
  {32'h38e4ec00, 32'hb9856da0} /* (27, 31, 13) {real, imag} */,
  {32'hbda44412, 32'hbc4dbff0} /* (27, 31, 12) {real, imag} */,
  {32'hbd439bb6, 32'h3cbf1dae} /* (27, 31, 11) {real, imag} */,
  {32'hbda7cd1c, 32'h3d8987e8} /* (27, 31, 10) {real, imag} */,
  {32'hbd1ce11e, 32'hbd2e3d53} /* (27, 31, 9) {real, imag} */,
  {32'h3b615340, 32'hbd579078} /* (27, 31, 8) {real, imag} */,
  {32'h3b90ea78, 32'hbd825b28} /* (27, 31, 7) {real, imag} */,
  {32'h3d386360, 32'h3cda9e7d} /* (27, 31, 6) {real, imag} */,
  {32'hbde7a235, 32'hbd43f234} /* (27, 31, 5) {real, imag} */,
  {32'h3e0529ec, 32'hbe3cb236} /* (27, 31, 4) {real, imag} */,
  {32'hbe182dd0, 32'h3b847204} /* (27, 31, 3) {real, imag} */,
  {32'hbe90b6d6, 32'hbed6fd1b} /* (27, 31, 2) {real, imag} */,
  {32'h3e1b5c29, 32'h3d752780} /* (27, 31, 1) {real, imag} */,
  {32'hbf2613e8, 32'h00000000} /* (27, 31, 0) {real, imag} */,
  {32'h3f101014, 32'hbcb2d720} /* (27, 30, 31) {real, imag} */,
  {32'hbf266210, 32'h3ec6820e} /* (27, 30, 30) {real, imag} */,
  {32'hbe1dba3b, 32'hbcab0602} /* (27, 30, 29) {real, imag} */,
  {32'h3e1e913f, 32'h3e3c6807} /* (27, 30, 28) {real, imag} */,
  {32'hbe8bb51f, 32'h3d3e86b2} /* (27, 30, 27) {real, imag} */,
  {32'h3d70c5e6, 32'h3bb3e3c0} /* (27, 30, 26) {real, imag} */,
  {32'h3d9d7e38, 32'hbd3f3094} /* (27, 30, 25) {real, imag} */,
  {32'hbc6eff44, 32'h3b5e45f0} /* (27, 30, 24) {real, imag} */,
  {32'h3c635950, 32'hbc89f4cf} /* (27, 30, 23) {real, imag} */,
  {32'hbc3dc20a, 32'hbd753e21} /* (27, 30, 22) {real, imag} */,
  {32'hbd3fdecf, 32'hbd4b4e86} /* (27, 30, 21) {real, imag} */,
  {32'hbe288604, 32'hbc62992a} /* (27, 30, 20) {real, imag} */,
  {32'h3d88b7d0, 32'h3d5f0373} /* (27, 30, 19) {real, imag} */,
  {32'h3d8ea969, 32'hbb1d9680} /* (27, 30, 18) {real, imag} */,
  {32'h3d00efa8, 32'hbc9210d5} /* (27, 30, 17) {real, imag} */,
  {32'hbdc3eff6, 32'h00000000} /* (27, 30, 16) {real, imag} */,
  {32'h3d00efa8, 32'h3c9210d5} /* (27, 30, 15) {real, imag} */,
  {32'h3d8ea969, 32'h3b1d9680} /* (27, 30, 14) {real, imag} */,
  {32'h3d88b7d0, 32'hbd5f0373} /* (27, 30, 13) {real, imag} */,
  {32'hbe288604, 32'h3c62992a} /* (27, 30, 12) {real, imag} */,
  {32'hbd3fdecf, 32'h3d4b4e86} /* (27, 30, 11) {real, imag} */,
  {32'hbc3dc20a, 32'h3d753e21} /* (27, 30, 10) {real, imag} */,
  {32'h3c635950, 32'h3c89f4cf} /* (27, 30, 9) {real, imag} */,
  {32'hbc6eff44, 32'hbb5e45f0} /* (27, 30, 8) {real, imag} */,
  {32'h3d9d7e38, 32'h3d3f3094} /* (27, 30, 7) {real, imag} */,
  {32'h3d70c5e6, 32'hbbb3e3c0} /* (27, 30, 6) {real, imag} */,
  {32'hbe8bb51f, 32'hbd3e86b2} /* (27, 30, 5) {real, imag} */,
  {32'h3e1e913f, 32'hbe3c6807} /* (27, 30, 4) {real, imag} */,
  {32'hbe1dba3b, 32'h3cab0602} /* (27, 30, 3) {real, imag} */,
  {32'hbf266210, 32'hbec6820e} /* (27, 30, 2) {real, imag} */,
  {32'h3f101014, 32'h3cb2d720} /* (27, 30, 1) {real, imag} */,
  {32'hbf0a8758, 32'h00000000} /* (27, 30, 0) {real, imag} */,
  {32'h3f38fca0, 32'h3e374734} /* (27, 29, 31) {real, imag} */,
  {32'hbf44bec0, 32'h3e813b20} /* (27, 29, 30) {real, imag} */,
  {32'hbdcd4312, 32'h3b6f73b0} /* (27, 29, 29) {real, imag} */,
  {32'h3cf52a9e, 32'hba0a4a80} /* (27, 29, 28) {real, imag} */,
  {32'hbe933f55, 32'h3d6b2aaf} /* (27, 29, 27) {real, imag} */,
  {32'hbd93d2be, 32'hbd4338c2} /* (27, 29, 26) {real, imag} */,
  {32'h3d114325, 32'hbdc61461} /* (27, 29, 25) {real, imag} */,
  {32'h3de00add, 32'h3cd2c9de} /* (27, 29, 24) {real, imag} */,
  {32'h3d06843a, 32'hbdb6f9e4} /* (27, 29, 23) {real, imag} */,
  {32'h3c28aa08, 32'hbbd10a3c} /* (27, 29, 22) {real, imag} */,
  {32'hbd00058f, 32'h3d73f807} /* (27, 29, 21) {real, imag} */,
  {32'h3c3b67e4, 32'h3d4071f0} /* (27, 29, 20) {real, imag} */,
  {32'h3d03e5b6, 32'h3cfcf735} /* (27, 29, 19) {real, imag} */,
  {32'hbccfd6f2, 32'hbb542ab0} /* (27, 29, 18) {real, imag} */,
  {32'h3cd0d8f6, 32'hbd0d5baf} /* (27, 29, 17) {real, imag} */,
  {32'hbde16cc0, 32'h00000000} /* (27, 29, 16) {real, imag} */,
  {32'h3cd0d8f6, 32'h3d0d5baf} /* (27, 29, 15) {real, imag} */,
  {32'hbccfd6f2, 32'h3b542ab0} /* (27, 29, 14) {real, imag} */,
  {32'h3d03e5b6, 32'hbcfcf735} /* (27, 29, 13) {real, imag} */,
  {32'h3c3b67e4, 32'hbd4071f0} /* (27, 29, 12) {real, imag} */,
  {32'hbd00058f, 32'hbd73f807} /* (27, 29, 11) {real, imag} */,
  {32'h3c28aa08, 32'h3bd10a3c} /* (27, 29, 10) {real, imag} */,
  {32'h3d06843a, 32'h3db6f9e4} /* (27, 29, 9) {real, imag} */,
  {32'h3de00add, 32'hbcd2c9de} /* (27, 29, 8) {real, imag} */,
  {32'h3d114325, 32'h3dc61461} /* (27, 29, 7) {real, imag} */,
  {32'hbd93d2be, 32'h3d4338c2} /* (27, 29, 6) {real, imag} */,
  {32'hbe933f55, 32'hbd6b2aaf} /* (27, 29, 5) {real, imag} */,
  {32'h3cf52a9e, 32'h3a0a4a80} /* (27, 29, 4) {real, imag} */,
  {32'hbdcd4312, 32'hbb6f73b0} /* (27, 29, 3) {real, imag} */,
  {32'hbf44bec0, 32'hbe813b20} /* (27, 29, 2) {real, imag} */,
  {32'h3f38fca0, 32'hbe374734} /* (27, 29, 1) {real, imag} */,
  {32'hbed96505, 32'h00000000} /* (27, 29, 0) {real, imag} */,
  {32'h3f458346, 32'h3ea2976d} /* (27, 28, 31) {real, imag} */,
  {32'hbf4b13d2, 32'h3e15d25c} /* (27, 28, 30) {real, imag} */,
  {32'hb9f6c880, 32'hbd6d230e} /* (27, 28, 29) {real, imag} */,
  {32'h3e189c69, 32'hbcfb3ebf} /* (27, 28, 28) {real, imag} */,
  {32'hbe6fb0c8, 32'h3d4531b5} /* (27, 28, 27) {real, imag} */,
  {32'h3d53e553, 32'hbda5085a} /* (27, 28, 26) {real, imag} */,
  {32'h3d664564, 32'hbc9a8608} /* (27, 28, 25) {real, imag} */,
  {32'hbda38535, 32'h3e1bd6fc} /* (27, 28, 24) {real, imag} */,
  {32'hbe0fa2a0, 32'hbd4fee27} /* (27, 28, 23) {real, imag} */,
  {32'hbe33f676, 32'hbc07c9ca} /* (27, 28, 22) {real, imag} */,
  {32'h3dd10b16, 32'h3d8a9822} /* (27, 28, 21) {real, imag} */,
  {32'h3d83d59b, 32'hbdb8820d} /* (27, 28, 20) {real, imag} */,
  {32'h3b982d60, 32'hbd4f7bf2} /* (27, 28, 19) {real, imag} */,
  {32'h3da76e47, 32'h3d9378ae} /* (27, 28, 18) {real, imag} */,
  {32'h3d40ecf4, 32'h3ccf3d7a} /* (27, 28, 17) {real, imag} */,
  {32'hbcedd827, 32'h00000000} /* (27, 28, 16) {real, imag} */,
  {32'h3d40ecf4, 32'hbccf3d7a} /* (27, 28, 15) {real, imag} */,
  {32'h3da76e47, 32'hbd9378ae} /* (27, 28, 14) {real, imag} */,
  {32'h3b982d60, 32'h3d4f7bf2} /* (27, 28, 13) {real, imag} */,
  {32'h3d83d59b, 32'h3db8820d} /* (27, 28, 12) {real, imag} */,
  {32'h3dd10b16, 32'hbd8a9822} /* (27, 28, 11) {real, imag} */,
  {32'hbe33f676, 32'h3c07c9ca} /* (27, 28, 10) {real, imag} */,
  {32'hbe0fa2a0, 32'h3d4fee27} /* (27, 28, 9) {real, imag} */,
  {32'hbda38535, 32'hbe1bd6fc} /* (27, 28, 8) {real, imag} */,
  {32'h3d664564, 32'h3c9a8608} /* (27, 28, 7) {real, imag} */,
  {32'h3d53e553, 32'h3da5085a} /* (27, 28, 6) {real, imag} */,
  {32'hbe6fb0c8, 32'hbd4531b5} /* (27, 28, 5) {real, imag} */,
  {32'h3e189c69, 32'h3cfb3ebf} /* (27, 28, 4) {real, imag} */,
  {32'hb9f6c880, 32'h3d6d230e} /* (27, 28, 3) {real, imag} */,
  {32'hbf4b13d2, 32'hbe15d25c} /* (27, 28, 2) {real, imag} */,
  {32'h3f458346, 32'hbea2976d} /* (27, 28, 1) {real, imag} */,
  {32'hbeb696f0, 32'h00000000} /* (27, 28, 0) {real, imag} */,
  {32'h3f3ecbc7, 32'h3e6d7f8e} /* (27, 27, 31) {real, imag} */,
  {32'hbf51bf72, 32'h3e1e9910} /* (27, 27, 30) {real, imag} */,
  {32'h3b364000, 32'hbd624108} /* (27, 27, 29) {real, imag} */,
  {32'hbc07c915, 32'hbdfbafde} /* (27, 27, 28) {real, imag} */,
  {32'hbe07925c, 32'h3e71054c} /* (27, 27, 27) {real, imag} */,
  {32'h3cc56996, 32'hbd82c06d} /* (27, 27, 26) {real, imag} */,
  {32'h3dbe360e, 32'hbd0effe4} /* (27, 27, 25) {real, imag} */,
  {32'hbd69a326, 32'h3dce4618} /* (27, 27, 24) {real, imag} */,
  {32'hbd129415, 32'hbd07402c} /* (27, 27, 23) {real, imag} */,
  {32'h3c28d8ac, 32'hbc224d8c} /* (27, 27, 22) {real, imag} */,
  {32'h3bed2160, 32'h3d4ab3b1} /* (27, 27, 21) {real, imag} */,
  {32'h3cc5aeb9, 32'hbc89b90c} /* (27, 27, 20) {real, imag} */,
  {32'hbca99ec2, 32'h3c4d3620} /* (27, 27, 19) {real, imag} */,
  {32'h3cae3902, 32'h3d6f4c1c} /* (27, 27, 18) {real, imag} */,
  {32'h3cc3e826, 32'hbb45c5d0} /* (27, 27, 17) {real, imag} */,
  {32'hbc2cc226, 32'h00000000} /* (27, 27, 16) {real, imag} */,
  {32'h3cc3e826, 32'h3b45c5d0} /* (27, 27, 15) {real, imag} */,
  {32'h3cae3902, 32'hbd6f4c1c} /* (27, 27, 14) {real, imag} */,
  {32'hbca99ec2, 32'hbc4d3620} /* (27, 27, 13) {real, imag} */,
  {32'h3cc5aeb9, 32'h3c89b90c} /* (27, 27, 12) {real, imag} */,
  {32'h3bed2160, 32'hbd4ab3b1} /* (27, 27, 11) {real, imag} */,
  {32'h3c28d8ac, 32'h3c224d8c} /* (27, 27, 10) {real, imag} */,
  {32'hbd129415, 32'h3d07402c} /* (27, 27, 9) {real, imag} */,
  {32'hbd69a326, 32'hbdce4618} /* (27, 27, 8) {real, imag} */,
  {32'h3dbe360e, 32'h3d0effe4} /* (27, 27, 7) {real, imag} */,
  {32'h3cc56996, 32'h3d82c06d} /* (27, 27, 6) {real, imag} */,
  {32'hbe07925c, 32'hbe71054c} /* (27, 27, 5) {real, imag} */,
  {32'hbc07c915, 32'h3dfbafde} /* (27, 27, 4) {real, imag} */,
  {32'h3b364000, 32'h3d624108} /* (27, 27, 3) {real, imag} */,
  {32'hbf51bf72, 32'hbe1e9910} /* (27, 27, 2) {real, imag} */,
  {32'h3f3ecbc7, 32'hbe6d7f8e} /* (27, 27, 1) {real, imag} */,
  {32'hbeb3e658, 32'h00000000} /* (27, 27, 0) {real, imag} */,
  {32'h3f3c202d, 32'h3e02224c} /* (27, 26, 31) {real, imag} */,
  {32'hbf551e0a, 32'h3e618e23} /* (27, 26, 30) {real, imag} */,
  {32'h3d675408, 32'hbd1df60d} /* (27, 26, 29) {real, imag} */,
  {32'h3e0e4b0e, 32'hbda68b03} /* (27, 26, 28) {real, imag} */,
  {32'hbda5f138, 32'h3e25880e} /* (27, 26, 27) {real, imag} */,
  {32'hbc9d0f9c, 32'hbd4a083e} /* (27, 26, 26) {real, imag} */,
  {32'h3ca63ea8, 32'hbd62f67e} /* (27, 26, 25) {real, imag} */,
  {32'hbcfa0d2c, 32'h3dbbff0c} /* (27, 26, 24) {real, imag} */,
  {32'hbd9d20a8, 32'h3c344078} /* (27, 26, 23) {real, imag} */,
  {32'h3d33d6b1, 32'hbd0a9f38} /* (27, 26, 22) {real, imag} */,
  {32'hbd8c78b0, 32'hbcc1a44e} /* (27, 26, 21) {real, imag} */,
  {32'h3d1f4fbe, 32'h3d8ea5a2} /* (27, 26, 20) {real, imag} */,
  {32'hbd9f9570, 32'hbd933e89} /* (27, 26, 19) {real, imag} */,
  {32'h3cc4ffc6, 32'h3d66efdc} /* (27, 26, 18) {real, imag} */,
  {32'hbd6cff77, 32'hbc4601a8} /* (27, 26, 17) {real, imag} */,
  {32'hbba35520, 32'h00000000} /* (27, 26, 16) {real, imag} */,
  {32'hbd6cff77, 32'h3c4601a8} /* (27, 26, 15) {real, imag} */,
  {32'h3cc4ffc6, 32'hbd66efdc} /* (27, 26, 14) {real, imag} */,
  {32'hbd9f9570, 32'h3d933e89} /* (27, 26, 13) {real, imag} */,
  {32'h3d1f4fbe, 32'hbd8ea5a2} /* (27, 26, 12) {real, imag} */,
  {32'hbd8c78b0, 32'h3cc1a44e} /* (27, 26, 11) {real, imag} */,
  {32'h3d33d6b1, 32'h3d0a9f38} /* (27, 26, 10) {real, imag} */,
  {32'hbd9d20a8, 32'hbc344078} /* (27, 26, 9) {real, imag} */,
  {32'hbcfa0d2c, 32'hbdbbff0c} /* (27, 26, 8) {real, imag} */,
  {32'h3ca63ea8, 32'h3d62f67e} /* (27, 26, 7) {real, imag} */,
  {32'hbc9d0f9c, 32'h3d4a083e} /* (27, 26, 6) {real, imag} */,
  {32'hbda5f138, 32'hbe25880e} /* (27, 26, 5) {real, imag} */,
  {32'h3e0e4b0e, 32'h3da68b03} /* (27, 26, 4) {real, imag} */,
  {32'h3d675408, 32'h3d1df60d} /* (27, 26, 3) {real, imag} */,
  {32'hbf551e0a, 32'hbe618e23} /* (27, 26, 2) {real, imag} */,
  {32'h3f3c202d, 32'hbe02224c} /* (27, 26, 1) {real, imag} */,
  {32'hbf020968, 32'h00000000} /* (27, 26, 0) {real, imag} */,
  {32'h3f0c8318, 32'h3de5e564} /* (27, 25, 31) {real, imag} */,
  {32'hbf4bb554, 32'h3e655dc7} /* (27, 25, 30) {real, imag} */,
  {32'hbd4542ec, 32'hbe09c92e} /* (27, 25, 29) {real, imag} */,
  {32'h3e6ccc7d, 32'hbd624630} /* (27, 25, 28) {real, imag} */,
  {32'hbdb11f5e, 32'h3cb8bf1c} /* (27, 25, 27) {real, imag} */,
  {32'hbde77cad, 32'h3d418716} /* (27, 25, 26) {real, imag} */,
  {32'hbc9fbc3e, 32'hbe05ee10} /* (27, 25, 25) {real, imag} */,
  {32'h3b0a9438, 32'h39832740} /* (27, 25, 24) {real, imag} */,
  {32'hbded6a85, 32'h3cf10e38} /* (27, 25, 23) {real, imag} */,
  {32'hbcdff177, 32'h3b525e40} /* (27, 25, 22) {real, imag} */,
  {32'hbde4ed1f, 32'h3cf851c6} /* (27, 25, 21) {real, imag} */,
  {32'h3ded8bc9, 32'hbd892a5e} /* (27, 25, 20) {real, imag} */,
  {32'hbc864149, 32'hbc5a1cd5} /* (27, 25, 19) {real, imag} */,
  {32'hbd4b87cc, 32'hbd53b3a2} /* (27, 25, 18) {real, imag} */,
  {32'h3d1501ea, 32'h3c0c35b4} /* (27, 25, 17) {real, imag} */,
  {32'h3cb45679, 32'h00000000} /* (27, 25, 16) {real, imag} */,
  {32'h3d1501ea, 32'hbc0c35b4} /* (27, 25, 15) {real, imag} */,
  {32'hbd4b87cc, 32'h3d53b3a2} /* (27, 25, 14) {real, imag} */,
  {32'hbc864149, 32'h3c5a1cd5} /* (27, 25, 13) {real, imag} */,
  {32'h3ded8bc9, 32'h3d892a5e} /* (27, 25, 12) {real, imag} */,
  {32'hbde4ed1f, 32'hbcf851c6} /* (27, 25, 11) {real, imag} */,
  {32'hbcdff177, 32'hbb525e40} /* (27, 25, 10) {real, imag} */,
  {32'hbded6a85, 32'hbcf10e38} /* (27, 25, 9) {real, imag} */,
  {32'h3b0a9438, 32'hb9832740} /* (27, 25, 8) {real, imag} */,
  {32'hbc9fbc3e, 32'h3e05ee10} /* (27, 25, 7) {real, imag} */,
  {32'hbde77cad, 32'hbd418716} /* (27, 25, 6) {real, imag} */,
  {32'hbdb11f5e, 32'hbcb8bf1c} /* (27, 25, 5) {real, imag} */,
  {32'h3e6ccc7d, 32'h3d624630} /* (27, 25, 4) {real, imag} */,
  {32'hbd4542ec, 32'h3e09c92e} /* (27, 25, 3) {real, imag} */,
  {32'hbf4bb554, 32'hbe655dc7} /* (27, 25, 2) {real, imag} */,
  {32'h3f0c8318, 32'hbde5e564} /* (27, 25, 1) {real, imag} */,
  {32'hbeb2d5ac, 32'h00000000} /* (27, 25, 0) {real, imag} */,
  {32'h3f115f2b, 32'hbc041b34} /* (27, 24, 31) {real, imag} */,
  {32'hbf50b2b9, 32'h3e06328c} /* (27, 24, 30) {real, imag} */,
  {32'hbd1cb9ab, 32'hbe3b4fb5} /* (27, 24, 29) {real, imag} */,
  {32'h3e5732c0, 32'hbd87aff0} /* (27, 24, 28) {real, imag} */,
  {32'hbdd8ccff, 32'h3e398d5b} /* (27, 24, 27) {real, imag} */,
  {32'hbd57f6c7, 32'h3e055348} /* (27, 24, 26) {real, imag} */,
  {32'h3d544be0, 32'hbe3d54ba} /* (27, 24, 25) {real, imag} */,
  {32'hbc775a00, 32'h3e243988} /* (27, 24, 24) {real, imag} */,
  {32'hbdde0592, 32'hbd03cd77} /* (27, 24, 23) {real, imag} */,
  {32'h3d3c9ff9, 32'h3dcde882} /* (27, 24, 22) {real, imag} */,
  {32'h3d6faec5, 32'h3d12d88e} /* (27, 24, 21) {real, imag} */,
  {32'h3d723ae8, 32'hbaef8140} /* (27, 24, 20) {real, imag} */,
  {32'hbd9b0795, 32'h3da688c0} /* (27, 24, 19) {real, imag} */,
  {32'hbd552906, 32'h3c683274} /* (27, 24, 18) {real, imag} */,
  {32'h3d548ffe, 32'hbdaec486} /* (27, 24, 17) {real, imag} */,
  {32'hbca4d401, 32'h00000000} /* (27, 24, 16) {real, imag} */,
  {32'h3d548ffe, 32'h3daec486} /* (27, 24, 15) {real, imag} */,
  {32'hbd552906, 32'hbc683274} /* (27, 24, 14) {real, imag} */,
  {32'hbd9b0795, 32'hbda688c0} /* (27, 24, 13) {real, imag} */,
  {32'h3d723ae8, 32'h3aef8140} /* (27, 24, 12) {real, imag} */,
  {32'h3d6faec5, 32'hbd12d88e} /* (27, 24, 11) {real, imag} */,
  {32'h3d3c9ff9, 32'hbdcde882} /* (27, 24, 10) {real, imag} */,
  {32'hbdde0592, 32'h3d03cd77} /* (27, 24, 9) {real, imag} */,
  {32'hbc775a00, 32'hbe243988} /* (27, 24, 8) {real, imag} */,
  {32'h3d544be0, 32'h3e3d54ba} /* (27, 24, 7) {real, imag} */,
  {32'hbd57f6c7, 32'hbe055348} /* (27, 24, 6) {real, imag} */,
  {32'hbdd8ccff, 32'hbe398d5b} /* (27, 24, 5) {real, imag} */,
  {32'h3e5732c0, 32'h3d87aff0} /* (27, 24, 4) {real, imag} */,
  {32'hbd1cb9ab, 32'h3e3b4fb5} /* (27, 24, 3) {real, imag} */,
  {32'hbf50b2b9, 32'hbe06328c} /* (27, 24, 2) {real, imag} */,
  {32'h3f115f2b, 32'h3c041b34} /* (27, 24, 1) {real, imag} */,
  {32'hbd6dc6b2, 32'h00000000} /* (27, 24, 0) {real, imag} */,
  {32'h3f033fd0, 32'hbcbbecfa} /* (27, 23, 31) {real, imag} */,
  {32'hbf40b5d4, 32'h3d3d979e} /* (27, 23, 30) {real, imag} */,
  {32'h3d20c324, 32'hbe20fd98} /* (27, 23, 29) {real, imag} */,
  {32'h3e20d34d, 32'hbd7da526} /* (27, 23, 28) {real, imag} */,
  {32'hbe4daaaf, 32'h3e2b9236} /* (27, 23, 27) {real, imag} */,
  {32'h3c5f057c, 32'h3dd3ef1a} /* (27, 23, 26) {real, imag} */,
  {32'h3d5ffb8e, 32'hbddb164a} /* (27, 23, 25) {real, imag} */,
  {32'hbcc956f5, 32'hbc2862d4} /* (27, 23, 24) {real, imag} */,
  {32'hbde52675, 32'hbcf6536c} /* (27, 23, 23) {real, imag} */,
  {32'h3d3b855c, 32'h3d4e45fc} /* (27, 23, 22) {real, imag} */,
  {32'hbd3a9ee4, 32'h3da79cda} /* (27, 23, 21) {real, imag} */,
  {32'h3d3c8156, 32'hbd2baccc} /* (27, 23, 20) {real, imag} */,
  {32'h3da077f9, 32'h3d129754} /* (27, 23, 19) {real, imag} */,
  {32'hbb1bb740, 32'hbd4948f0} /* (27, 23, 18) {real, imag} */,
  {32'h3ce69cf6, 32'hbd976c14} /* (27, 23, 17) {real, imag} */,
  {32'h3d47cde3, 32'h00000000} /* (27, 23, 16) {real, imag} */,
  {32'h3ce69cf6, 32'h3d976c14} /* (27, 23, 15) {real, imag} */,
  {32'hbb1bb740, 32'h3d4948f0} /* (27, 23, 14) {real, imag} */,
  {32'h3da077f9, 32'hbd129754} /* (27, 23, 13) {real, imag} */,
  {32'h3d3c8156, 32'h3d2baccc} /* (27, 23, 12) {real, imag} */,
  {32'hbd3a9ee4, 32'hbda79cda} /* (27, 23, 11) {real, imag} */,
  {32'h3d3b855c, 32'hbd4e45fc} /* (27, 23, 10) {real, imag} */,
  {32'hbde52675, 32'h3cf6536c} /* (27, 23, 9) {real, imag} */,
  {32'hbcc956f5, 32'h3c2862d4} /* (27, 23, 8) {real, imag} */,
  {32'h3d5ffb8e, 32'h3ddb164a} /* (27, 23, 7) {real, imag} */,
  {32'h3c5f057c, 32'hbdd3ef1a} /* (27, 23, 6) {real, imag} */,
  {32'hbe4daaaf, 32'hbe2b9236} /* (27, 23, 5) {real, imag} */,
  {32'h3e20d34d, 32'h3d7da526} /* (27, 23, 4) {real, imag} */,
  {32'h3d20c324, 32'h3e20fd98} /* (27, 23, 3) {real, imag} */,
  {32'hbf40b5d4, 32'hbd3d979e} /* (27, 23, 2) {real, imag} */,
  {32'h3f033fd0, 32'h3cbbecfa} /* (27, 23, 1) {real, imag} */,
  {32'h3e67073b, 32'h00000000} /* (27, 23, 0) {real, imag} */,
  {32'h3ec97523, 32'h3e0f1908} /* (27, 22, 31) {real, imag} */,
  {32'hbea9a31c, 32'hbb040440} /* (27, 22, 30) {real, imag} */,
  {32'h3a966740, 32'hbd481836} /* (27, 22, 29) {real, imag} */,
  {32'h3d90917c, 32'hbd074fe4} /* (27, 22, 28) {real, imag} */,
  {32'hbdea90d2, 32'h3db7692a} /* (27, 22, 27) {real, imag} */,
  {32'h3d333042, 32'h3d097f44} /* (27, 22, 26) {real, imag} */,
  {32'hbc9fffec, 32'h3c8ad7ad} /* (27, 22, 25) {real, imag} */,
  {32'hbd93aff5, 32'hbd6ad622} /* (27, 22, 24) {real, imag} */,
  {32'h3d931156, 32'h3d50f48c} /* (27, 22, 23) {real, imag} */,
  {32'h3d4f8a02, 32'h3b49428c} /* (27, 22, 22) {real, imag} */,
  {32'h3c2863ae, 32'h3cf24cc3} /* (27, 22, 21) {real, imag} */,
  {32'h3d07138c, 32'h3c2f8db7} /* (27, 22, 20) {real, imag} */,
  {32'h3d126848, 32'hbd09dec1} /* (27, 22, 19) {real, imag} */,
  {32'h3cbd2696, 32'h3dccafa8} /* (27, 22, 18) {real, imag} */,
  {32'h38b3f7c0, 32'h3ce57986} /* (27, 22, 17) {real, imag} */,
  {32'h3d07f09f, 32'h00000000} /* (27, 22, 16) {real, imag} */,
  {32'h38b3f7c0, 32'hbce57986} /* (27, 22, 15) {real, imag} */,
  {32'h3cbd2696, 32'hbdccafa8} /* (27, 22, 14) {real, imag} */,
  {32'h3d126848, 32'h3d09dec1} /* (27, 22, 13) {real, imag} */,
  {32'h3d07138c, 32'hbc2f8db7} /* (27, 22, 12) {real, imag} */,
  {32'h3c2863ae, 32'hbcf24cc3} /* (27, 22, 11) {real, imag} */,
  {32'h3d4f8a02, 32'hbb49428c} /* (27, 22, 10) {real, imag} */,
  {32'h3d931156, 32'hbd50f48c} /* (27, 22, 9) {real, imag} */,
  {32'hbd93aff5, 32'h3d6ad622} /* (27, 22, 8) {real, imag} */,
  {32'hbc9fffec, 32'hbc8ad7ad} /* (27, 22, 7) {real, imag} */,
  {32'h3d333042, 32'hbd097f44} /* (27, 22, 6) {real, imag} */,
  {32'hbdea90d2, 32'hbdb7692a} /* (27, 22, 5) {real, imag} */,
  {32'h3d90917c, 32'h3d074fe4} /* (27, 22, 4) {real, imag} */,
  {32'h3a966740, 32'h3d481836} /* (27, 22, 3) {real, imag} */,
  {32'hbea9a31c, 32'h3b040440} /* (27, 22, 2) {real, imag} */,
  {32'h3ec97523, 32'hbe0f1908} /* (27, 22, 1) {real, imag} */,
  {32'h3e30c978, 32'h00000000} /* (27, 22, 0) {real, imag} */,
  {32'hbe2b0b03, 32'h3e5e448b} /* (27, 21, 31) {real, imag} */,
  {32'hbb21eb80, 32'h3b804a00} /* (27, 21, 30) {real, imag} */,
  {32'h3cc1206c, 32'hbe03d703} /* (27, 21, 29) {real, imag} */,
  {32'hbcf528e8, 32'h3deeaa96} /* (27, 21, 28) {real, imag} */,
  {32'hbc6c418c, 32'h3da71cdb} /* (27, 21, 27) {real, imag} */,
  {32'hbcb1cc8a, 32'hbd001030} /* (27, 21, 26) {real, imag} */,
  {32'h3dcdd7d2, 32'hbd68c4e1} /* (27, 21, 25) {real, imag} */,
  {32'hbe1c95c6, 32'h3c88d5ca} /* (27, 21, 24) {real, imag} */,
  {32'hbcc3c797, 32'hbdf10f8a} /* (27, 21, 23) {real, imag} */,
  {32'h3cfd20b4, 32'hbcc6cf20} /* (27, 21, 22) {real, imag} */,
  {32'h3ddf1ed0, 32'h3beb2aae} /* (27, 21, 21) {real, imag} */,
  {32'h3cc6d03e, 32'h3d8aab0f} /* (27, 21, 20) {real, imag} */,
  {32'hbc5d5f46, 32'hbc0b3bc2} /* (27, 21, 19) {real, imag} */,
  {32'hbcec2b30, 32'h3c9d20fd} /* (27, 21, 18) {real, imag} */,
  {32'h3cc7ccbc, 32'h3d1b7f25} /* (27, 21, 17) {real, imag} */,
  {32'hbdbbcec9, 32'h00000000} /* (27, 21, 16) {real, imag} */,
  {32'h3cc7ccbc, 32'hbd1b7f25} /* (27, 21, 15) {real, imag} */,
  {32'hbcec2b30, 32'hbc9d20fd} /* (27, 21, 14) {real, imag} */,
  {32'hbc5d5f46, 32'h3c0b3bc2} /* (27, 21, 13) {real, imag} */,
  {32'h3cc6d03e, 32'hbd8aab0f} /* (27, 21, 12) {real, imag} */,
  {32'h3ddf1ed0, 32'hbbeb2aae} /* (27, 21, 11) {real, imag} */,
  {32'h3cfd20b4, 32'h3cc6cf20} /* (27, 21, 10) {real, imag} */,
  {32'hbcc3c797, 32'h3df10f8a} /* (27, 21, 9) {real, imag} */,
  {32'hbe1c95c6, 32'hbc88d5ca} /* (27, 21, 8) {real, imag} */,
  {32'h3dcdd7d2, 32'h3d68c4e1} /* (27, 21, 7) {real, imag} */,
  {32'hbcb1cc8a, 32'h3d001030} /* (27, 21, 6) {real, imag} */,
  {32'hbc6c418c, 32'hbda71cdb} /* (27, 21, 5) {real, imag} */,
  {32'hbcf528e8, 32'hbdeeaa96} /* (27, 21, 4) {real, imag} */,
  {32'h3cc1206c, 32'h3e03d703} /* (27, 21, 3) {real, imag} */,
  {32'hbb21eb80, 32'hbb804a00} /* (27, 21, 2) {real, imag} */,
  {32'hbe2b0b03, 32'hbe5e448b} /* (27, 21, 1) {real, imag} */,
  {32'hbbdbbb00, 32'h00000000} /* (27, 21, 0) {real, imag} */,
  {32'hbf720e8f, 32'h3e32cfc3} /* (27, 20, 31) {real, imag} */,
  {32'h3ef65f8e, 32'hbdb5937c} /* (27, 20, 30) {real, imag} */,
  {32'hbcbc8ec7, 32'hbe0390ce} /* (27, 20, 29) {real, imag} */,
  {32'h3cc652e8, 32'h3d109720} /* (27, 20, 28) {real, imag} */,
  {32'h3d8744c4, 32'hbd9786cc} /* (27, 20, 27) {real, imag} */,
  {32'h3c9c2f36, 32'h3b7602e8} /* (27, 20, 26) {real, imag} */,
  {32'h3d760385, 32'hbde75346} /* (27, 20, 25) {real, imag} */,
  {32'hbd6f2113, 32'hbcd79b8c} /* (27, 20, 24) {real, imag} */,
  {32'hbdba39c2, 32'h3ce4e314} /* (27, 20, 23) {real, imag} */,
  {32'hbd2ab6cc, 32'h3dac13de} /* (27, 20, 22) {real, imag} */,
  {32'h3dab5ea1, 32'h3d54057d} /* (27, 20, 21) {real, imag} */,
  {32'h3d3a0da4, 32'hbd8d2d9c} /* (27, 20, 20) {real, imag} */,
  {32'hbd3f47b6, 32'hbc440bb4} /* (27, 20, 19) {real, imag} */,
  {32'h3d2dfec4, 32'hbd339d65} /* (27, 20, 18) {real, imag} */,
  {32'hbd47b529, 32'hbc64e1e0} /* (27, 20, 17) {real, imag} */,
  {32'h3d12f652, 32'h00000000} /* (27, 20, 16) {real, imag} */,
  {32'hbd47b529, 32'h3c64e1e0} /* (27, 20, 15) {real, imag} */,
  {32'h3d2dfec4, 32'h3d339d65} /* (27, 20, 14) {real, imag} */,
  {32'hbd3f47b6, 32'h3c440bb4} /* (27, 20, 13) {real, imag} */,
  {32'h3d3a0da4, 32'h3d8d2d9c} /* (27, 20, 12) {real, imag} */,
  {32'h3dab5ea1, 32'hbd54057d} /* (27, 20, 11) {real, imag} */,
  {32'hbd2ab6cc, 32'hbdac13de} /* (27, 20, 10) {real, imag} */,
  {32'hbdba39c2, 32'hbce4e314} /* (27, 20, 9) {real, imag} */,
  {32'hbd6f2113, 32'h3cd79b8c} /* (27, 20, 8) {real, imag} */,
  {32'h3d760385, 32'h3de75346} /* (27, 20, 7) {real, imag} */,
  {32'h3c9c2f36, 32'hbb7602e8} /* (27, 20, 6) {real, imag} */,
  {32'h3d8744c4, 32'h3d9786cc} /* (27, 20, 5) {real, imag} */,
  {32'h3cc652e8, 32'hbd109720} /* (27, 20, 4) {real, imag} */,
  {32'hbcbc8ec7, 32'h3e0390ce} /* (27, 20, 3) {real, imag} */,
  {32'h3ef65f8e, 32'h3db5937c} /* (27, 20, 2) {real, imag} */,
  {32'hbf720e8f, 32'hbe32cfc3} /* (27, 20, 1) {real, imag} */,
  {32'hbf0bb049, 32'h00000000} /* (27, 20, 0) {real, imag} */,
  {32'hbf95f8ca, 32'h3e73b1bd} /* (27, 19, 31) {real, imag} */,
  {32'h3f18a2dc, 32'hbe7631d0} /* (27, 19, 30) {real, imag} */,
  {32'h3bbb89c0, 32'hbe002b68} /* (27, 19, 29) {real, imag} */,
  {32'hbc734244, 32'hbd116ff8} /* (27, 19, 28) {real, imag} */,
  {32'h3e097302, 32'h3c38134c} /* (27, 19, 27) {real, imag} */,
  {32'h3d866972, 32'hbd877b67} /* (27, 19, 26) {real, imag} */,
  {32'hbc9be5c6, 32'h3d89df8e} /* (27, 19, 25) {real, imag} */,
  {32'h3cfd1f0a, 32'h3d075912} /* (27, 19, 24) {real, imag} */,
  {32'h3dc3cf6d, 32'h3c99d49e} /* (27, 19, 23) {real, imag} */,
  {32'h3db78f98, 32'h3d08db76} /* (27, 19, 22) {real, imag} */,
  {32'h3d8845fc, 32'h3d74772d} /* (27, 19, 21) {real, imag} */,
  {32'hbdaa9182, 32'h3db60b03} /* (27, 19, 20) {real, imag} */,
  {32'h3be69864, 32'h3dbf7a63} /* (27, 19, 19) {real, imag} */,
  {32'hbd62fe99, 32'hbccc083d} /* (27, 19, 18) {real, imag} */,
  {32'h3c1ae7bb, 32'h3cae7dda} /* (27, 19, 17) {real, imag} */,
  {32'hbc1c7744, 32'h00000000} /* (27, 19, 16) {real, imag} */,
  {32'h3c1ae7bb, 32'hbcae7dda} /* (27, 19, 15) {real, imag} */,
  {32'hbd62fe99, 32'h3ccc083d} /* (27, 19, 14) {real, imag} */,
  {32'h3be69864, 32'hbdbf7a63} /* (27, 19, 13) {real, imag} */,
  {32'hbdaa9182, 32'hbdb60b03} /* (27, 19, 12) {real, imag} */,
  {32'h3d8845fc, 32'hbd74772d} /* (27, 19, 11) {real, imag} */,
  {32'h3db78f98, 32'hbd08db76} /* (27, 19, 10) {real, imag} */,
  {32'h3dc3cf6d, 32'hbc99d49e} /* (27, 19, 9) {real, imag} */,
  {32'h3cfd1f0a, 32'hbd075912} /* (27, 19, 8) {real, imag} */,
  {32'hbc9be5c6, 32'hbd89df8e} /* (27, 19, 7) {real, imag} */,
  {32'h3d866972, 32'h3d877b67} /* (27, 19, 6) {real, imag} */,
  {32'h3e097302, 32'hbc38134c} /* (27, 19, 5) {real, imag} */,
  {32'hbc734244, 32'h3d116ff8} /* (27, 19, 4) {real, imag} */,
  {32'h3bbb89c0, 32'h3e002b68} /* (27, 19, 3) {real, imag} */,
  {32'h3f18a2dc, 32'h3e7631d0} /* (27, 19, 2) {real, imag} */,
  {32'hbf95f8ca, 32'hbe73b1bd} /* (27, 19, 1) {real, imag} */,
  {32'hbf267762, 32'h00000000} /* (27, 19, 0) {real, imag} */,
  {32'hbf9dd857, 32'h3eaf8800} /* (27, 18, 31) {real, imag} */,
  {32'h3f3ee154, 32'hbea1ab68} /* (27, 18, 30) {real, imag} */,
  {32'h3de20868, 32'hbc875a72} /* (27, 18, 29) {real, imag} */,
  {32'hbca74160, 32'h3e1493d7} /* (27, 18, 28) {real, imag} */,
  {32'h3d94f67b, 32'h3db451dc} /* (27, 18, 27) {real, imag} */,
  {32'hbba747d8, 32'h3d0979e2} /* (27, 18, 26) {real, imag} */,
  {32'hbc83f23d, 32'hbd93833c} /* (27, 18, 25) {real, imag} */,
  {32'h3d51680c, 32'h3ccd9968} /* (27, 18, 24) {real, imag} */,
  {32'h3d1f9b96, 32'h3ba44eaa} /* (27, 18, 23) {real, imag} */,
  {32'hbcb7f09d, 32'h3aea0680} /* (27, 18, 22) {real, imag} */,
  {32'hbd63ef74, 32'h3c962853} /* (27, 18, 21) {real, imag} */,
  {32'hbc45455c, 32'hbdbc932f} /* (27, 18, 20) {real, imag} */,
  {32'hbd14483e, 32'h3caa84f2} /* (27, 18, 19) {real, imag} */,
  {32'h3dd6fa0e, 32'hbd731224} /* (27, 18, 18) {real, imag} */,
  {32'h3da84736, 32'hbc0e85e2} /* (27, 18, 17) {real, imag} */,
  {32'hbd1304dc, 32'h00000000} /* (27, 18, 16) {real, imag} */,
  {32'h3da84736, 32'h3c0e85e2} /* (27, 18, 15) {real, imag} */,
  {32'h3dd6fa0e, 32'h3d731224} /* (27, 18, 14) {real, imag} */,
  {32'hbd14483e, 32'hbcaa84f2} /* (27, 18, 13) {real, imag} */,
  {32'hbc45455c, 32'h3dbc932f} /* (27, 18, 12) {real, imag} */,
  {32'hbd63ef74, 32'hbc962853} /* (27, 18, 11) {real, imag} */,
  {32'hbcb7f09d, 32'hbaea0680} /* (27, 18, 10) {real, imag} */,
  {32'h3d1f9b96, 32'hbba44eaa} /* (27, 18, 9) {real, imag} */,
  {32'h3d51680c, 32'hbccd9968} /* (27, 18, 8) {real, imag} */,
  {32'hbc83f23d, 32'h3d93833c} /* (27, 18, 7) {real, imag} */,
  {32'hbba747d8, 32'hbd0979e2} /* (27, 18, 6) {real, imag} */,
  {32'h3d94f67b, 32'hbdb451dc} /* (27, 18, 5) {real, imag} */,
  {32'hbca74160, 32'hbe1493d7} /* (27, 18, 4) {real, imag} */,
  {32'h3de20868, 32'h3c875a72} /* (27, 18, 3) {real, imag} */,
  {32'h3f3ee154, 32'h3ea1ab68} /* (27, 18, 2) {real, imag} */,
  {32'hbf9dd857, 32'hbeaf8800} /* (27, 18, 1) {real, imag} */,
  {32'hbf59088e, 32'h00000000} /* (27, 18, 0) {real, imag} */,
  {32'hbf9fade5, 32'h3ea721e4} /* (27, 17, 31) {real, imag} */,
  {32'h3f40c880, 32'hbe59a3e8} /* (27, 17, 30) {real, imag} */,
  {32'hba997050, 32'hbdb2c3b2} /* (27, 17, 29) {real, imag} */,
  {32'h3d2e3055, 32'h3e6074bb} /* (27, 17, 28) {real, imag} */,
  {32'h3e3a738e, 32'hbd8a56db} /* (27, 17, 27) {real, imag} */,
  {32'h3deea554, 32'h3c4a4812} /* (27, 17, 26) {real, imag} */,
  {32'h3d9052d7, 32'hbdec9c77} /* (27, 17, 25) {real, imag} */,
  {32'h3cc9e6b1, 32'hbc13f388} /* (27, 17, 24) {real, imag} */,
  {32'h3d9d21d1, 32'h3d10d7f5} /* (27, 17, 23) {real, imag} */,
  {32'h3d411766, 32'h3df542d9} /* (27, 17, 22) {real, imag} */,
  {32'hbc27d564, 32'hbdd1f185} /* (27, 17, 21) {real, imag} */,
  {32'h3b7f9190, 32'h3d654b49} /* (27, 17, 20) {real, imag} */,
  {32'h3c551f98, 32'h3c1a503c} /* (27, 17, 19) {real, imag} */,
  {32'hbd1e9dee, 32'h3d4cfd74} /* (27, 17, 18) {real, imag} */,
  {32'hbb549ee0, 32'h3dbb9f5a} /* (27, 17, 17) {real, imag} */,
  {32'hbd1f134c, 32'h00000000} /* (27, 17, 16) {real, imag} */,
  {32'hbb549ee0, 32'hbdbb9f5a} /* (27, 17, 15) {real, imag} */,
  {32'hbd1e9dee, 32'hbd4cfd74} /* (27, 17, 14) {real, imag} */,
  {32'h3c551f98, 32'hbc1a503c} /* (27, 17, 13) {real, imag} */,
  {32'h3b7f9190, 32'hbd654b49} /* (27, 17, 12) {real, imag} */,
  {32'hbc27d564, 32'h3dd1f185} /* (27, 17, 11) {real, imag} */,
  {32'h3d411766, 32'hbdf542d9} /* (27, 17, 10) {real, imag} */,
  {32'h3d9d21d1, 32'hbd10d7f5} /* (27, 17, 9) {real, imag} */,
  {32'h3cc9e6b1, 32'h3c13f388} /* (27, 17, 8) {real, imag} */,
  {32'h3d9052d7, 32'h3dec9c77} /* (27, 17, 7) {real, imag} */,
  {32'h3deea554, 32'hbc4a4812} /* (27, 17, 6) {real, imag} */,
  {32'h3e3a738e, 32'h3d8a56db} /* (27, 17, 5) {real, imag} */,
  {32'h3d2e3055, 32'hbe6074bb} /* (27, 17, 4) {real, imag} */,
  {32'hba997050, 32'h3db2c3b2} /* (27, 17, 3) {real, imag} */,
  {32'h3f40c880, 32'h3e59a3e8} /* (27, 17, 2) {real, imag} */,
  {32'hbf9fade5, 32'hbea721e4} /* (27, 17, 1) {real, imag} */,
  {32'hbf76fe8e, 32'h00000000} /* (27, 17, 0) {real, imag} */,
  {32'hbf9ebafa, 32'h3e8d8580} /* (27, 16, 31) {real, imag} */,
  {32'h3f2c113c, 32'hbdeefd58} /* (27, 16, 30) {real, imag} */,
  {32'h3d90fa18, 32'hbdb64edd} /* (27, 16, 29) {real, imag} */,
  {32'hbdec243f, 32'h3dc55686} /* (27, 16, 28) {real, imag} */,
  {32'h3e2ef188, 32'h3c495b8c} /* (27, 16, 27) {real, imag} */,
  {32'h3d67cd92, 32'h3a1ce550} /* (27, 16, 26) {real, imag} */,
  {32'h3b219370, 32'hbd36f3c3} /* (27, 16, 25) {real, imag} */,
  {32'h3d83ea7f, 32'hbd635194} /* (27, 16, 24) {real, imag} */,
  {32'hbd43c8dd, 32'hbc13c867} /* (27, 16, 23) {real, imag} */,
  {32'hbdbc56fc, 32'hbd80b1fa} /* (27, 16, 22) {real, imag} */,
  {32'h3c0db3aa, 32'hbd750cc8} /* (27, 16, 21) {real, imag} */,
  {32'h3bc1868c, 32'hbceeae29} /* (27, 16, 20) {real, imag} */,
  {32'hbc75ec42, 32'hbce47e2a} /* (27, 16, 19) {real, imag} */,
  {32'hbd7b0712, 32'h3ba4bb90} /* (27, 16, 18) {real, imag} */,
  {32'h3d0fd2be, 32'h3da8b736} /* (27, 16, 17) {real, imag} */,
  {32'hbcaba374, 32'h00000000} /* (27, 16, 16) {real, imag} */,
  {32'h3d0fd2be, 32'hbda8b736} /* (27, 16, 15) {real, imag} */,
  {32'hbd7b0712, 32'hbba4bb90} /* (27, 16, 14) {real, imag} */,
  {32'hbc75ec42, 32'h3ce47e2a} /* (27, 16, 13) {real, imag} */,
  {32'h3bc1868c, 32'h3ceeae29} /* (27, 16, 12) {real, imag} */,
  {32'h3c0db3aa, 32'h3d750cc8} /* (27, 16, 11) {real, imag} */,
  {32'hbdbc56fc, 32'h3d80b1fa} /* (27, 16, 10) {real, imag} */,
  {32'hbd43c8dd, 32'h3c13c867} /* (27, 16, 9) {real, imag} */,
  {32'h3d83ea7f, 32'h3d635194} /* (27, 16, 8) {real, imag} */,
  {32'h3b219370, 32'h3d36f3c3} /* (27, 16, 7) {real, imag} */,
  {32'h3d67cd92, 32'hba1ce550} /* (27, 16, 6) {real, imag} */,
  {32'h3e2ef188, 32'hbc495b8c} /* (27, 16, 5) {real, imag} */,
  {32'hbdec243f, 32'hbdc55686} /* (27, 16, 4) {real, imag} */,
  {32'h3d90fa18, 32'h3db64edd} /* (27, 16, 3) {real, imag} */,
  {32'h3f2c113c, 32'h3deefd58} /* (27, 16, 2) {real, imag} */,
  {32'hbf9ebafa, 32'hbe8d8580} /* (27, 16, 1) {real, imag} */,
  {32'hbf84ff20, 32'h00000000} /* (27, 16, 0) {real, imag} */,
  {32'hbf8c422f, 32'h3e923984} /* (27, 15, 31) {real, imag} */,
  {32'h3f38228a, 32'hbda87338} /* (27, 15, 30) {real, imag} */,
  {32'h3d29f956, 32'hbd4ed1dc} /* (27, 15, 29) {real, imag} */,
  {32'hbdc41b0c, 32'h3dec7ab2} /* (27, 15, 28) {real, imag} */,
  {32'h3da8ae8c, 32'hbda9b10d} /* (27, 15, 27) {real, imag} */,
  {32'hbd4c8681, 32'hbc88a6a3} /* (27, 15, 26) {real, imag} */,
  {32'hbd3c4f92, 32'h3db74e11} /* (27, 15, 25) {real, imag} */,
  {32'h3daa112a, 32'hbe0adbf2} /* (27, 15, 24) {real, imag} */,
  {32'hbcede169, 32'hbc82cf66} /* (27, 15, 23) {real, imag} */,
  {32'hbd7aa0da, 32'h3dd8770b} /* (27, 15, 22) {real, imag} */,
  {32'h3d185103, 32'hbd1efd8e} /* (27, 15, 21) {real, imag} */,
  {32'h3d271a25, 32'h39c55d80} /* (27, 15, 20) {real, imag} */,
  {32'hb9d17b40, 32'h3d53f90f} /* (27, 15, 19) {real, imag} */,
  {32'h3d692b96, 32'hbd94b422} /* (27, 15, 18) {real, imag} */,
  {32'h3dc3f64d, 32'hbd10b9f1} /* (27, 15, 17) {real, imag} */,
  {32'hbdabfdd2, 32'h00000000} /* (27, 15, 16) {real, imag} */,
  {32'h3dc3f64d, 32'h3d10b9f1} /* (27, 15, 15) {real, imag} */,
  {32'h3d692b96, 32'h3d94b422} /* (27, 15, 14) {real, imag} */,
  {32'hb9d17b40, 32'hbd53f90f} /* (27, 15, 13) {real, imag} */,
  {32'h3d271a25, 32'hb9c55d80} /* (27, 15, 12) {real, imag} */,
  {32'h3d185103, 32'h3d1efd8e} /* (27, 15, 11) {real, imag} */,
  {32'hbd7aa0da, 32'hbdd8770b} /* (27, 15, 10) {real, imag} */,
  {32'hbcede169, 32'h3c82cf66} /* (27, 15, 9) {real, imag} */,
  {32'h3daa112a, 32'h3e0adbf2} /* (27, 15, 8) {real, imag} */,
  {32'hbd3c4f92, 32'hbdb74e11} /* (27, 15, 7) {real, imag} */,
  {32'hbd4c8681, 32'h3c88a6a3} /* (27, 15, 6) {real, imag} */,
  {32'h3da8ae8c, 32'h3da9b10d} /* (27, 15, 5) {real, imag} */,
  {32'hbdc41b0c, 32'hbdec7ab2} /* (27, 15, 4) {real, imag} */,
  {32'h3d29f956, 32'h3d4ed1dc} /* (27, 15, 3) {real, imag} */,
  {32'h3f38228a, 32'h3da87338} /* (27, 15, 2) {real, imag} */,
  {32'hbf8c422f, 32'hbe923984} /* (27, 15, 1) {real, imag} */,
  {32'hbf988a5f, 32'h00000000} /* (27, 15, 0) {real, imag} */,
  {32'hbf84f901, 32'h3ea38156} /* (27, 14, 31) {real, imag} */,
  {32'h3f2d011c, 32'hbcff6808} /* (27, 14, 30) {real, imag} */,
  {32'hbbc00c38, 32'h3c245618} /* (27, 14, 29) {real, imag} */,
  {32'hbe3457f8, 32'h3dd626d3} /* (27, 14, 28) {real, imag} */,
  {32'h3e359a28, 32'hbde684a0} /* (27, 14, 27) {real, imag} */,
  {32'h3d9f129c, 32'hbce19c3a} /* (27, 14, 26) {real, imag} */,
  {32'hbb52f428, 32'h3d779a88} /* (27, 14, 25) {real, imag} */,
  {32'h3d613042, 32'hbcf41200} /* (27, 14, 24) {real, imag} */,
  {32'h3d401c9c, 32'h3c8c32e0} /* (27, 14, 23) {real, imag} */,
  {32'h3c98b283, 32'hbda7b803} /* (27, 14, 22) {real, imag} */,
  {32'h3e194f5d, 32'hbc81d9cf} /* (27, 14, 21) {real, imag} */,
  {32'h3d9f620e, 32'hbdae0141} /* (27, 14, 20) {real, imag} */,
  {32'hbbeccf74, 32'hbb88c6a6} /* (27, 14, 19) {real, imag} */,
  {32'h3c18c7b0, 32'hbce936ef} /* (27, 14, 18) {real, imag} */,
  {32'hbb997220, 32'hbd242398} /* (27, 14, 17) {real, imag} */,
  {32'h3cf944a0, 32'h00000000} /* (27, 14, 16) {real, imag} */,
  {32'hbb997220, 32'h3d242398} /* (27, 14, 15) {real, imag} */,
  {32'h3c18c7b0, 32'h3ce936ef} /* (27, 14, 14) {real, imag} */,
  {32'hbbeccf74, 32'h3b88c6a6} /* (27, 14, 13) {real, imag} */,
  {32'h3d9f620e, 32'h3dae0141} /* (27, 14, 12) {real, imag} */,
  {32'h3e194f5d, 32'h3c81d9cf} /* (27, 14, 11) {real, imag} */,
  {32'h3c98b283, 32'h3da7b803} /* (27, 14, 10) {real, imag} */,
  {32'h3d401c9c, 32'hbc8c32e0} /* (27, 14, 9) {real, imag} */,
  {32'h3d613042, 32'h3cf41200} /* (27, 14, 8) {real, imag} */,
  {32'hbb52f428, 32'hbd779a88} /* (27, 14, 7) {real, imag} */,
  {32'h3d9f129c, 32'h3ce19c3a} /* (27, 14, 6) {real, imag} */,
  {32'h3e359a28, 32'h3de684a0} /* (27, 14, 5) {real, imag} */,
  {32'hbe3457f8, 32'hbdd626d3} /* (27, 14, 4) {real, imag} */,
  {32'hbbc00c38, 32'hbc245618} /* (27, 14, 3) {real, imag} */,
  {32'h3f2d011c, 32'h3cff6808} /* (27, 14, 2) {real, imag} */,
  {32'hbf84f901, 32'hbea38156} /* (27, 14, 1) {real, imag} */,
  {32'hbf8f5b72, 32'h00000000} /* (27, 14, 0) {real, imag} */,
  {32'hbf6b0098, 32'h3e520d57} /* (27, 13, 31) {real, imag} */,
  {32'h3f0bd284, 32'hbd683660} /* (27, 13, 30) {real, imag} */,
  {32'hbd6407dc, 32'h3d8a91c4} /* (27, 13, 29) {real, imag} */,
  {32'hbe0258f6, 32'h3ddf06b6} /* (27, 13, 28) {real, imag} */,
  {32'h3dfaced8, 32'hbe0b201c} /* (27, 13, 27) {real, imag} */,
  {32'h3e1adc25, 32'h3d96c665} /* (27, 13, 26) {real, imag} */,
  {32'h3d6e4705, 32'hbbf2ab6c} /* (27, 13, 25) {real, imag} */,
  {32'h3cf290c0, 32'h3d5447ac} /* (27, 13, 24) {real, imag} */,
  {32'h39ee2d00, 32'h3dabc372} /* (27, 13, 23) {real, imag} */,
  {32'hbcdd1758, 32'hbb2bbe08} /* (27, 13, 22) {real, imag} */,
  {32'h3c3b2848, 32'hbdd96eb6} /* (27, 13, 21) {real, imag} */,
  {32'h3d4a55cc, 32'h3c83dfb0} /* (27, 13, 20) {real, imag} */,
  {32'hbca1ddd3, 32'h3c88027c} /* (27, 13, 19) {real, imag} */,
  {32'hbd317585, 32'hbc99e16b} /* (27, 13, 18) {real, imag} */,
  {32'hbbfa7a56, 32'h3c45fba3} /* (27, 13, 17) {real, imag} */,
  {32'h3df1454c, 32'h00000000} /* (27, 13, 16) {real, imag} */,
  {32'hbbfa7a56, 32'hbc45fba3} /* (27, 13, 15) {real, imag} */,
  {32'hbd317585, 32'h3c99e16b} /* (27, 13, 14) {real, imag} */,
  {32'hbca1ddd3, 32'hbc88027c} /* (27, 13, 13) {real, imag} */,
  {32'h3d4a55cc, 32'hbc83dfb0} /* (27, 13, 12) {real, imag} */,
  {32'h3c3b2848, 32'h3dd96eb6} /* (27, 13, 11) {real, imag} */,
  {32'hbcdd1758, 32'h3b2bbe08} /* (27, 13, 10) {real, imag} */,
  {32'h39ee2d00, 32'hbdabc372} /* (27, 13, 9) {real, imag} */,
  {32'h3cf290c0, 32'hbd5447ac} /* (27, 13, 8) {real, imag} */,
  {32'h3d6e4705, 32'h3bf2ab6c} /* (27, 13, 7) {real, imag} */,
  {32'h3e1adc25, 32'hbd96c665} /* (27, 13, 6) {real, imag} */,
  {32'h3dfaced8, 32'h3e0b201c} /* (27, 13, 5) {real, imag} */,
  {32'hbe0258f6, 32'hbddf06b6} /* (27, 13, 4) {real, imag} */,
  {32'hbd6407dc, 32'hbd8a91c4} /* (27, 13, 3) {real, imag} */,
  {32'h3f0bd284, 32'h3d683660} /* (27, 13, 2) {real, imag} */,
  {32'hbf6b0098, 32'hbe520d57} /* (27, 13, 1) {real, imag} */,
  {32'hbf845779, 32'h00000000} /* (27, 13, 0) {real, imag} */,
  {32'hbf4267a1, 32'h3e71be91} /* (27, 12, 31) {real, imag} */,
  {32'h3ed72910, 32'hbd0b3ff0} /* (27, 12, 30) {real, imag} */,
  {32'hbb4c9f28, 32'hbc3fd0e8} /* (27, 12, 29) {real, imag} */,
  {32'hbd0bca42, 32'h3d3d6d88} /* (27, 12, 28) {real, imag} */,
  {32'h3ca832d7, 32'hbd9f0b4c} /* (27, 12, 27) {real, imag} */,
  {32'hbcd7f8ca, 32'h3d032e48} /* (27, 12, 26) {real, imag} */,
  {32'h3d2a1e8b, 32'hbcd2b916} /* (27, 12, 25) {real, imag} */,
  {32'h3d4a6759, 32'h3c921604} /* (27, 12, 24) {real, imag} */,
  {32'h3dae0ffe, 32'hbccaed28} /* (27, 12, 23) {real, imag} */,
  {32'hbdc6f642, 32'h3e27c0ac} /* (27, 12, 22) {real, imag} */,
  {32'h3d32d6b2, 32'hbd078dbd} /* (27, 12, 21) {real, imag} */,
  {32'h3dda0344, 32'hbd6ce595} /* (27, 12, 20) {real, imag} */,
  {32'hbd890c85, 32'h3c622a66} /* (27, 12, 19) {real, imag} */,
  {32'hbc16692e, 32'hb87e3800} /* (27, 12, 18) {real, imag} */,
  {32'h3cd119f2, 32'hbca249d8} /* (27, 12, 17) {real, imag} */,
  {32'hbda7810b, 32'h00000000} /* (27, 12, 16) {real, imag} */,
  {32'h3cd119f2, 32'h3ca249d8} /* (27, 12, 15) {real, imag} */,
  {32'hbc16692e, 32'h387e3800} /* (27, 12, 14) {real, imag} */,
  {32'hbd890c85, 32'hbc622a66} /* (27, 12, 13) {real, imag} */,
  {32'h3dda0344, 32'h3d6ce595} /* (27, 12, 12) {real, imag} */,
  {32'h3d32d6b2, 32'h3d078dbd} /* (27, 12, 11) {real, imag} */,
  {32'hbdc6f642, 32'hbe27c0ac} /* (27, 12, 10) {real, imag} */,
  {32'h3dae0ffe, 32'h3ccaed28} /* (27, 12, 9) {real, imag} */,
  {32'h3d4a6759, 32'hbc921604} /* (27, 12, 8) {real, imag} */,
  {32'h3d2a1e8b, 32'h3cd2b916} /* (27, 12, 7) {real, imag} */,
  {32'hbcd7f8ca, 32'hbd032e48} /* (27, 12, 6) {real, imag} */,
  {32'h3ca832d7, 32'h3d9f0b4c} /* (27, 12, 5) {real, imag} */,
  {32'hbd0bca42, 32'hbd3d6d88} /* (27, 12, 4) {real, imag} */,
  {32'hbb4c9f28, 32'h3c3fd0e8} /* (27, 12, 3) {real, imag} */,
  {32'h3ed72910, 32'h3d0b3ff0} /* (27, 12, 2) {real, imag} */,
  {32'hbf4267a1, 32'hbe71be91} /* (27, 12, 1) {real, imag} */,
  {32'hbf664e41, 32'h00000000} /* (27, 12, 0) {real, imag} */,
  {32'hbf03ae97, 32'h3e2606b9} /* (27, 11, 31) {real, imag} */,
  {32'h3e9794eb, 32'h3d565470} /* (27, 11, 30) {real, imag} */,
  {32'hbcb50110, 32'hbcafbbd0} /* (27, 11, 29) {real, imag} */,
  {32'hbcaea29c, 32'hbdfd3e0e} /* (27, 11, 28) {real, imag} */,
  {32'h3d85f620, 32'hbd9e75f7} /* (27, 11, 27) {real, imag} */,
  {32'h3b266e50, 32'hbc24d038} /* (27, 11, 26) {real, imag} */,
  {32'h3d4d847d, 32'hbd7beef3} /* (27, 11, 25) {real, imag} */,
  {32'hbc95a17c, 32'h3c9b6dfa} /* (27, 11, 24) {real, imag} */,
  {32'h3c5480da, 32'hbd922242} /* (27, 11, 23) {real, imag} */,
  {32'hbe05a0b8, 32'h3e196c01} /* (27, 11, 22) {real, imag} */,
  {32'h3e0098fb, 32'hbc1da283} /* (27, 11, 21) {real, imag} */,
  {32'hbce54792, 32'hbd8142c7} /* (27, 11, 20) {real, imag} */,
  {32'h3d345c0e, 32'hbcfb8657} /* (27, 11, 19) {real, imag} */,
  {32'h3d26c280, 32'hbc284992} /* (27, 11, 18) {real, imag} */,
  {32'h3ca5c8be, 32'h3adb71e0} /* (27, 11, 17) {real, imag} */,
  {32'hbd313e66, 32'h00000000} /* (27, 11, 16) {real, imag} */,
  {32'h3ca5c8be, 32'hbadb71e0} /* (27, 11, 15) {real, imag} */,
  {32'h3d26c280, 32'h3c284992} /* (27, 11, 14) {real, imag} */,
  {32'h3d345c0e, 32'h3cfb8657} /* (27, 11, 13) {real, imag} */,
  {32'hbce54792, 32'h3d8142c7} /* (27, 11, 12) {real, imag} */,
  {32'h3e0098fb, 32'h3c1da283} /* (27, 11, 11) {real, imag} */,
  {32'hbe05a0b8, 32'hbe196c01} /* (27, 11, 10) {real, imag} */,
  {32'h3c5480da, 32'h3d922242} /* (27, 11, 9) {real, imag} */,
  {32'hbc95a17c, 32'hbc9b6dfa} /* (27, 11, 8) {real, imag} */,
  {32'h3d4d847d, 32'h3d7beef3} /* (27, 11, 7) {real, imag} */,
  {32'h3b266e50, 32'h3c24d038} /* (27, 11, 6) {real, imag} */,
  {32'h3d85f620, 32'h3d9e75f7} /* (27, 11, 5) {real, imag} */,
  {32'hbcaea29c, 32'h3dfd3e0e} /* (27, 11, 4) {real, imag} */,
  {32'hbcb50110, 32'h3cafbbd0} /* (27, 11, 3) {real, imag} */,
  {32'h3e9794eb, 32'hbd565470} /* (27, 11, 2) {real, imag} */,
  {32'hbf03ae97, 32'hbe2606b9} /* (27, 11, 1) {real, imag} */,
  {32'hbf0d43ae, 32'h00000000} /* (27, 11, 0) {real, imag} */,
  {32'h3e912615, 32'h3e1e40fc} /* (27, 10, 31) {real, imag} */,
  {32'hbe88d130, 32'h3e2f9c69} /* (27, 10, 30) {real, imag} */,
  {32'hbda55cc1, 32'h3b7a1b90} /* (27, 10, 29) {real, imag} */,
  {32'h3e361509, 32'hbea36414} /* (27, 10, 28) {real, imag} */,
  {32'h3cc15d78, 32'h3e02f1ab} /* (27, 10, 27) {real, imag} */,
  {32'h3ca9e87c, 32'h3cb42ea4} /* (27, 10, 26) {real, imag} */,
  {32'h3d76d426, 32'hbd95aa57} /* (27, 10, 25) {real, imag} */,
  {32'hbd90d42d, 32'h3d307aca} /* (27, 10, 24) {real, imag} */,
  {32'h3ccc29c6, 32'h3c9dfe6c} /* (27, 10, 23) {real, imag} */,
  {32'h3ce36bc8, 32'h3c99d27c} /* (27, 10, 22) {real, imag} */,
  {32'h3a9f5a94, 32'h3da22b10} /* (27, 10, 21) {real, imag} */,
  {32'hbdbba63f, 32'hbc882d8c} /* (27, 10, 20) {real, imag} */,
  {32'h3b966792, 32'hba266040} /* (27, 10, 19) {real, imag} */,
  {32'hbd4f295d, 32'h3b2fe640} /* (27, 10, 18) {real, imag} */,
  {32'hbc15a378, 32'hbc9b289c} /* (27, 10, 17) {real, imag} */,
  {32'h3daaf656, 32'h00000000} /* (27, 10, 16) {real, imag} */,
  {32'hbc15a378, 32'h3c9b289c} /* (27, 10, 15) {real, imag} */,
  {32'hbd4f295d, 32'hbb2fe640} /* (27, 10, 14) {real, imag} */,
  {32'h3b966792, 32'h3a266040} /* (27, 10, 13) {real, imag} */,
  {32'hbdbba63f, 32'h3c882d8c} /* (27, 10, 12) {real, imag} */,
  {32'h3a9f5a94, 32'hbda22b10} /* (27, 10, 11) {real, imag} */,
  {32'h3ce36bc8, 32'hbc99d27c} /* (27, 10, 10) {real, imag} */,
  {32'h3ccc29c6, 32'hbc9dfe6c} /* (27, 10, 9) {real, imag} */,
  {32'hbd90d42d, 32'hbd307aca} /* (27, 10, 8) {real, imag} */,
  {32'h3d76d426, 32'h3d95aa57} /* (27, 10, 7) {real, imag} */,
  {32'h3ca9e87c, 32'hbcb42ea4} /* (27, 10, 6) {real, imag} */,
  {32'h3cc15d78, 32'hbe02f1ab} /* (27, 10, 5) {real, imag} */,
  {32'h3e361509, 32'h3ea36414} /* (27, 10, 4) {real, imag} */,
  {32'hbda55cc1, 32'hbb7a1b90} /* (27, 10, 3) {real, imag} */,
  {32'hbe88d130, 32'hbe2f9c69} /* (27, 10, 2) {real, imag} */,
  {32'h3e912615, 32'hbe1e40fc} /* (27, 10, 1) {real, imag} */,
  {32'hbd71fb7e, 32'h00000000} /* (27, 10, 0) {real, imag} */,
  {32'h3f3b520a, 32'h3ded7cb2} /* (27, 9, 31) {real, imag} */,
  {32'hbf044530, 32'h3df68f23} /* (27, 9, 30) {real, imag} */,
  {32'h3e11542f, 32'hbd7a2952} /* (27, 9, 29) {real, imag} */,
  {32'h3e3c35d9, 32'hbe1e0422} /* (27, 9, 28) {real, imag} */,
  {32'hbe40bba9, 32'h3d77a3d6} /* (27, 9, 27) {real, imag} */,
  {32'h3d54afa5, 32'h3b6f67e0} /* (27, 9, 26) {real, imag} */,
  {32'h3d28839e, 32'hbcbe3e9e} /* (27, 9, 25) {real, imag} */,
  {32'hbd2be9ea, 32'h3dafb762} /* (27, 9, 24) {real, imag} */,
  {32'h3d8685ad, 32'hbc23f878} /* (27, 9, 23) {real, imag} */,
  {32'hbd444ea4, 32'hbd45e57a} /* (27, 9, 22) {real, imag} */,
  {32'h3d2d6cb8, 32'h3cd4a956} /* (27, 9, 21) {real, imag} */,
  {32'hbd052cba, 32'h3c8fe5ed} /* (27, 9, 20) {real, imag} */,
  {32'hbd2c95c6, 32'h3d0a29fa} /* (27, 9, 19) {real, imag} */,
  {32'h3d073c31, 32'h3d15bfa0} /* (27, 9, 18) {real, imag} */,
  {32'hbd61383b, 32'h3b310a10} /* (27, 9, 17) {real, imag} */,
  {32'h3d055efd, 32'h00000000} /* (27, 9, 16) {real, imag} */,
  {32'hbd61383b, 32'hbb310a10} /* (27, 9, 15) {real, imag} */,
  {32'h3d073c31, 32'hbd15bfa0} /* (27, 9, 14) {real, imag} */,
  {32'hbd2c95c6, 32'hbd0a29fa} /* (27, 9, 13) {real, imag} */,
  {32'hbd052cba, 32'hbc8fe5ed} /* (27, 9, 12) {real, imag} */,
  {32'h3d2d6cb8, 32'hbcd4a956} /* (27, 9, 11) {real, imag} */,
  {32'hbd444ea4, 32'h3d45e57a} /* (27, 9, 10) {real, imag} */,
  {32'h3d8685ad, 32'h3c23f878} /* (27, 9, 9) {real, imag} */,
  {32'hbd2be9ea, 32'hbdafb762} /* (27, 9, 8) {real, imag} */,
  {32'h3d28839e, 32'h3cbe3e9e} /* (27, 9, 7) {real, imag} */,
  {32'h3d54afa5, 32'hbb6f67e0} /* (27, 9, 6) {real, imag} */,
  {32'hbe40bba9, 32'hbd77a3d6} /* (27, 9, 5) {real, imag} */,
  {32'h3e3c35d9, 32'h3e1e0422} /* (27, 9, 4) {real, imag} */,
  {32'h3e11542f, 32'h3d7a2952} /* (27, 9, 3) {real, imag} */,
  {32'hbf044530, 32'hbdf68f23} /* (27, 9, 2) {real, imag} */,
  {32'h3f3b520a, 32'hbded7cb2} /* (27, 9, 1) {real, imag} */,
  {32'h3d5ed294, 32'h00000000} /* (27, 9, 0) {real, imag} */,
  {32'h3f63ca7f, 32'h3d03bafb} /* (27, 8, 31) {real, imag} */,
  {32'hbf2878df, 32'h3e8ee356} /* (27, 8, 30) {real, imag} */,
  {32'h3d75ac39, 32'hbd3c2c44} /* (27, 8, 29) {real, imag} */,
  {32'h3d95a7e1, 32'hbe47fff6} /* (27, 8, 28) {real, imag} */,
  {32'hbdfe36e3, 32'h3de697de} /* (27, 8, 27) {real, imag} */,
  {32'hbc3cd664, 32'h3b54e7c0} /* (27, 8, 26) {real, imag} */,
  {32'h3cdda460, 32'hbde34c94} /* (27, 8, 25) {real, imag} */,
  {32'hbd921118, 32'h3e2ef864} /* (27, 8, 24) {real, imag} */,
  {32'h3d701ffb, 32'hbb89ff88} /* (27, 8, 23) {real, imag} */,
  {32'h3e0b5356, 32'hbc797a64} /* (27, 8, 22) {real, imag} */,
  {32'h3ce11e8e, 32'hbbb1fe10} /* (27, 8, 21) {real, imag} */,
  {32'h3d233e60, 32'h3ddc0099} /* (27, 8, 20) {real, imag} */,
  {32'h3db509c9, 32'hbdeeec8e} /* (27, 8, 19) {real, imag} */,
  {32'hbdb99ff9, 32'hbce898d6} /* (27, 8, 18) {real, imag} */,
  {32'hbd6b8f72, 32'h3c2b80cc} /* (27, 8, 17) {real, imag} */,
  {32'h3c6a68e6, 32'h00000000} /* (27, 8, 16) {real, imag} */,
  {32'hbd6b8f72, 32'hbc2b80cc} /* (27, 8, 15) {real, imag} */,
  {32'hbdb99ff9, 32'h3ce898d6} /* (27, 8, 14) {real, imag} */,
  {32'h3db509c9, 32'h3deeec8e} /* (27, 8, 13) {real, imag} */,
  {32'h3d233e60, 32'hbddc0099} /* (27, 8, 12) {real, imag} */,
  {32'h3ce11e8e, 32'h3bb1fe10} /* (27, 8, 11) {real, imag} */,
  {32'h3e0b5356, 32'h3c797a64} /* (27, 8, 10) {real, imag} */,
  {32'h3d701ffb, 32'h3b89ff88} /* (27, 8, 9) {real, imag} */,
  {32'hbd921118, 32'hbe2ef864} /* (27, 8, 8) {real, imag} */,
  {32'h3cdda460, 32'h3de34c94} /* (27, 8, 7) {real, imag} */,
  {32'hbc3cd664, 32'hbb54e7c0} /* (27, 8, 6) {real, imag} */,
  {32'hbdfe36e3, 32'hbde697de} /* (27, 8, 5) {real, imag} */,
  {32'h3d95a7e1, 32'h3e47fff6} /* (27, 8, 4) {real, imag} */,
  {32'h3d75ac39, 32'h3d3c2c44} /* (27, 8, 3) {real, imag} */,
  {32'hbf2878df, 32'hbe8ee356} /* (27, 8, 2) {real, imag} */,
  {32'h3f63ca7f, 32'hbd03bafb} /* (27, 8, 1) {real, imag} */,
  {32'hbd4bb7ee, 32'h00000000} /* (27, 8, 0) {real, imag} */,
  {32'h3f5348ce, 32'h3d2e97c8} /* (27, 7, 31) {real, imag} */,
  {32'hbf1bb884, 32'h3eaec208} /* (27, 7, 30) {real, imag} */,
  {32'h3c5f7310, 32'h3dc41a6e} /* (27, 7, 29) {real, imag} */,
  {32'h3d53b3f4, 32'hbdc3aac2} /* (27, 7, 28) {real, imag} */,
  {32'hbd42ef45, 32'h3da551f1} /* (27, 7, 27) {real, imag} */,
  {32'h3cfe71ec, 32'hbc120fb0} /* (27, 7, 26) {real, imag} */,
  {32'h3c3c4bf8, 32'hbd3ce63d} /* (27, 7, 25) {real, imag} */,
  {32'h3d35cb14, 32'h3cc6cdc3} /* (27, 7, 24) {real, imag} */,
  {32'hbd2bac66, 32'h3da67210} /* (27, 7, 23) {real, imag} */,
  {32'hbda13d80, 32'hbdb7551b} /* (27, 7, 22) {real, imag} */,
  {32'hbd787d62, 32'h3c4973d4} /* (27, 7, 21) {real, imag} */,
  {32'hbd4a6d3e, 32'hbd3d6346} /* (27, 7, 20) {real, imag} */,
  {32'h3d384504, 32'h3cd4648e} /* (27, 7, 19) {real, imag} */,
  {32'h3dd87db4, 32'hbc3e9c78} /* (27, 7, 18) {real, imag} */,
  {32'hbca27700, 32'h3c1de454} /* (27, 7, 17) {real, imag} */,
  {32'hbd158052, 32'h00000000} /* (27, 7, 16) {real, imag} */,
  {32'hbca27700, 32'hbc1de454} /* (27, 7, 15) {real, imag} */,
  {32'h3dd87db4, 32'h3c3e9c78} /* (27, 7, 14) {real, imag} */,
  {32'h3d384504, 32'hbcd4648e} /* (27, 7, 13) {real, imag} */,
  {32'hbd4a6d3e, 32'h3d3d6346} /* (27, 7, 12) {real, imag} */,
  {32'hbd787d62, 32'hbc4973d4} /* (27, 7, 11) {real, imag} */,
  {32'hbda13d80, 32'h3db7551b} /* (27, 7, 10) {real, imag} */,
  {32'hbd2bac66, 32'hbda67210} /* (27, 7, 9) {real, imag} */,
  {32'h3d35cb14, 32'hbcc6cdc3} /* (27, 7, 8) {real, imag} */,
  {32'h3c3c4bf8, 32'h3d3ce63d} /* (27, 7, 7) {real, imag} */,
  {32'h3cfe71ec, 32'h3c120fb0} /* (27, 7, 6) {real, imag} */,
  {32'hbd42ef45, 32'hbda551f1} /* (27, 7, 5) {real, imag} */,
  {32'h3d53b3f4, 32'h3dc3aac2} /* (27, 7, 4) {real, imag} */,
  {32'h3c5f7310, 32'hbdc41a6e} /* (27, 7, 3) {real, imag} */,
  {32'hbf1bb884, 32'hbeaec208} /* (27, 7, 2) {real, imag} */,
  {32'h3f5348ce, 32'hbd2e97c8} /* (27, 7, 1) {real, imag} */,
  {32'hbd851d22, 32'h00000000} /* (27, 7, 0) {real, imag} */,
  {32'h3f2859eb, 32'h3c957d80} /* (27, 6, 31) {real, imag} */,
  {32'hbf0a8320, 32'h3ed162c2} /* (27, 6, 30) {real, imag} */,
  {32'hbab8b0f0, 32'h3ba96860} /* (27, 6, 29) {real, imag} */,
  {32'h3e041c7c, 32'h3d44de3e} /* (27, 6, 28) {real, imag} */,
  {32'hbe0ade04, 32'h3ddc0c10} /* (27, 6, 27) {real, imag} */,
  {32'h3e54c4ca, 32'hbd9df57d} /* (27, 6, 26) {real, imag} */,
  {32'hbd575d90, 32'h3c7c2056} /* (27, 6, 25) {real, imag} */,
  {32'hbc483939, 32'h3e153372} /* (27, 6, 24) {real, imag} */,
  {32'hbcc34f96, 32'h3d5a09b8} /* (27, 6, 23) {real, imag} */,
  {32'hbd087c17, 32'hbc00555e} /* (27, 6, 22) {real, imag} */,
  {32'hbceb949f, 32'h3dbd1762} /* (27, 6, 21) {real, imag} */,
  {32'hbd89fcf4, 32'h3d483ef4} /* (27, 6, 20) {real, imag} */,
  {32'h3b973810, 32'hbdb55e77} /* (27, 6, 19) {real, imag} */,
  {32'h3d19022b, 32'h3d913b88} /* (27, 6, 18) {real, imag} */,
  {32'hbd46043f, 32'hbc87e8f8} /* (27, 6, 17) {real, imag} */,
  {32'hbd87b651, 32'h00000000} /* (27, 6, 16) {real, imag} */,
  {32'hbd46043f, 32'h3c87e8f8} /* (27, 6, 15) {real, imag} */,
  {32'h3d19022b, 32'hbd913b88} /* (27, 6, 14) {real, imag} */,
  {32'h3b973810, 32'h3db55e77} /* (27, 6, 13) {real, imag} */,
  {32'hbd89fcf4, 32'hbd483ef4} /* (27, 6, 12) {real, imag} */,
  {32'hbceb949f, 32'hbdbd1762} /* (27, 6, 11) {real, imag} */,
  {32'hbd087c17, 32'h3c00555e} /* (27, 6, 10) {real, imag} */,
  {32'hbcc34f96, 32'hbd5a09b8} /* (27, 6, 9) {real, imag} */,
  {32'hbc483939, 32'hbe153372} /* (27, 6, 8) {real, imag} */,
  {32'hbd575d90, 32'hbc7c2056} /* (27, 6, 7) {real, imag} */,
  {32'h3e54c4ca, 32'h3d9df57d} /* (27, 6, 6) {real, imag} */,
  {32'hbe0ade04, 32'hbddc0c10} /* (27, 6, 5) {real, imag} */,
  {32'h3e041c7c, 32'hbd44de3e} /* (27, 6, 4) {real, imag} */,
  {32'hbab8b0f0, 32'hbba96860} /* (27, 6, 3) {real, imag} */,
  {32'hbf0a8320, 32'hbed162c2} /* (27, 6, 2) {real, imag} */,
  {32'h3f2859eb, 32'hbc957d80} /* (27, 6, 1) {real, imag} */,
  {32'h3d360520, 32'h00000000} /* (27, 6, 0) {real, imag} */,
  {32'h3ebd6982, 32'hbe99f415} /* (27, 5, 31) {real, imag} */,
  {32'hbe8596b9, 32'h3ee18222} /* (27, 5, 30) {real, imag} */,
  {32'h3c826b70, 32'hbc930627} /* (27, 5, 29) {real, imag} */,
  {32'hbc954aa2, 32'h3decbd56} /* (27, 5, 28) {real, imag} */,
  {32'hbdcf0fd0, 32'h3d1956ce} /* (27, 5, 27) {real, imag} */,
  {32'h3d88056e, 32'hbd91827f} /* (27, 5, 26) {real, imag} */,
  {32'hbdd5ec3e, 32'h3c89ff89} /* (27, 5, 25) {real, imag} */,
  {32'hbcc27db3, 32'h3e08cb82} /* (27, 5, 24) {real, imag} */,
  {32'hbbe6a9fe, 32'h3c3f79a8} /* (27, 5, 23) {real, imag} */,
  {32'h3d6d92a1, 32'hbd9e8cd0} /* (27, 5, 22) {real, imag} */,
  {32'hbcc62840, 32'h3cfd9656} /* (27, 5, 21) {real, imag} */,
  {32'hbd400858, 32'h3c77126c} /* (27, 5, 20) {real, imag} */,
  {32'h3db8f228, 32'h3ca73b30} /* (27, 5, 19) {real, imag} */,
  {32'hbc5fe3f7, 32'hbd282f48} /* (27, 5, 18) {real, imag} */,
  {32'h3d05df32, 32'h3d102ff9} /* (27, 5, 17) {real, imag} */,
  {32'h3c9aef7b, 32'h00000000} /* (27, 5, 16) {real, imag} */,
  {32'h3d05df32, 32'hbd102ff9} /* (27, 5, 15) {real, imag} */,
  {32'hbc5fe3f7, 32'h3d282f48} /* (27, 5, 14) {real, imag} */,
  {32'h3db8f228, 32'hbca73b30} /* (27, 5, 13) {real, imag} */,
  {32'hbd400858, 32'hbc77126c} /* (27, 5, 12) {real, imag} */,
  {32'hbcc62840, 32'hbcfd9656} /* (27, 5, 11) {real, imag} */,
  {32'h3d6d92a1, 32'h3d9e8cd0} /* (27, 5, 10) {real, imag} */,
  {32'hbbe6a9fe, 32'hbc3f79a8} /* (27, 5, 9) {real, imag} */,
  {32'hbcc27db3, 32'hbe08cb82} /* (27, 5, 8) {real, imag} */,
  {32'hbdd5ec3e, 32'hbc89ff89} /* (27, 5, 7) {real, imag} */,
  {32'h3d88056e, 32'h3d91827f} /* (27, 5, 6) {real, imag} */,
  {32'hbdcf0fd0, 32'hbd1956ce} /* (27, 5, 5) {real, imag} */,
  {32'hbc954aa2, 32'hbdecbd56} /* (27, 5, 4) {real, imag} */,
  {32'h3c826b70, 32'h3c930627} /* (27, 5, 3) {real, imag} */,
  {32'hbe8596b9, 32'hbee18222} /* (27, 5, 2) {real, imag} */,
  {32'h3ebd6982, 32'h3e99f415} /* (27, 5, 1) {real, imag} */,
  {32'hbca60960, 32'h00000000} /* (27, 5, 0) {real, imag} */,
  {32'h3d8e1dd0, 32'hbeb6797f} /* (27, 4, 31) {real, imag} */,
  {32'h3e171454, 32'h3f2dff03} /* (27, 4, 30) {real, imag} */,
  {32'hbdddbbe0, 32'hbbc1da70} /* (27, 4, 29) {real, imag} */,
  {32'hbdfec6a6, 32'h3d0485a8} /* (27, 4, 28) {real, imag} */,
  {32'hbe848578, 32'hbd540b79} /* (27, 4, 27) {real, imag} */,
  {32'h3d805696, 32'h3d262331} /* (27, 4, 26) {real, imag} */,
  {32'h3ccaafb8, 32'hbc3a4a38} /* (27, 4, 25) {real, imag} */,
  {32'h3de1bb0d, 32'h3cb32c5c} /* (27, 4, 24) {real, imag} */,
  {32'hbd938c6d, 32'hbd1dc577} /* (27, 4, 23) {real, imag} */,
  {32'hbd0257c6, 32'h3c3db4fa} /* (27, 4, 22) {real, imag} */,
  {32'hba1d5440, 32'hbd361dea} /* (27, 4, 21) {real, imag} */,
  {32'hbd4f183a, 32'h3b45c720} /* (27, 4, 20) {real, imag} */,
  {32'h3d82d7fe, 32'hbba61870} /* (27, 4, 19) {real, imag} */,
  {32'h3d747cda, 32'h3d00bb14} /* (27, 4, 18) {real, imag} */,
  {32'hbd5a6872, 32'h3dad6c10} /* (27, 4, 17) {real, imag} */,
  {32'h3bf59584, 32'h00000000} /* (27, 4, 16) {real, imag} */,
  {32'hbd5a6872, 32'hbdad6c10} /* (27, 4, 15) {real, imag} */,
  {32'h3d747cda, 32'hbd00bb14} /* (27, 4, 14) {real, imag} */,
  {32'h3d82d7fe, 32'h3ba61870} /* (27, 4, 13) {real, imag} */,
  {32'hbd4f183a, 32'hbb45c720} /* (27, 4, 12) {real, imag} */,
  {32'hba1d5440, 32'h3d361dea} /* (27, 4, 11) {real, imag} */,
  {32'hbd0257c6, 32'hbc3db4fa} /* (27, 4, 10) {real, imag} */,
  {32'hbd938c6d, 32'h3d1dc577} /* (27, 4, 9) {real, imag} */,
  {32'h3de1bb0d, 32'hbcb32c5c} /* (27, 4, 8) {real, imag} */,
  {32'h3ccaafb8, 32'h3c3a4a38} /* (27, 4, 7) {real, imag} */,
  {32'h3d805696, 32'hbd262331} /* (27, 4, 6) {real, imag} */,
  {32'hbe848578, 32'h3d540b79} /* (27, 4, 5) {real, imag} */,
  {32'hbdfec6a6, 32'hbd0485a8} /* (27, 4, 4) {real, imag} */,
  {32'hbdddbbe0, 32'h3bc1da70} /* (27, 4, 3) {real, imag} */,
  {32'h3e171454, 32'hbf2dff03} /* (27, 4, 2) {real, imag} */,
  {32'h3d8e1dd0, 32'h3eb6797f} /* (27, 4, 1) {real, imag} */,
  {32'hbe1be3c8, 32'h00000000} /* (27, 4, 0) {real, imag} */,
  {32'hbcecb570, 32'hbf111ea5} /* (27, 3, 31) {real, imag} */,
  {32'h3e943e09, 32'h3f1664c2} /* (27, 3, 30) {real, imag} */,
  {32'hbda30f74, 32'hbdc73a56} /* (27, 3, 29) {real, imag} */,
  {32'hbdd4971e, 32'h3db2ee87} /* (27, 3, 28) {real, imag} */,
  {32'hbe19b458, 32'h3d3bb877} /* (27, 3, 27) {real, imag} */,
  {32'hbd1e7b96, 32'h3ca0111c} /* (27, 3, 26) {real, imag} */,
  {32'h3b420f30, 32'h3d424dee} /* (27, 3, 25) {real, imag} */,
  {32'h3c6d41a8, 32'h3d42a7eb} /* (27, 3, 24) {real, imag} */,
  {32'hbca8ed6d, 32'h3caea8da} /* (27, 3, 23) {real, imag} */,
  {32'hbdb906fb, 32'h3d4d481a} /* (27, 3, 22) {real, imag} */,
  {32'h3c7c4b34, 32'hbcf06082} /* (27, 3, 21) {real, imag} */,
  {32'h3d05f899, 32'h3d8721bf} /* (27, 3, 20) {real, imag} */,
  {32'h3cc32bea, 32'hbd090726} /* (27, 3, 19) {real, imag} */,
  {32'h3d9a9f06, 32'h3d9b3a12} /* (27, 3, 18) {real, imag} */,
  {32'hbbc306e8, 32'hbd77bda7} /* (27, 3, 17) {real, imag} */,
  {32'h3d003a29, 32'h00000000} /* (27, 3, 16) {real, imag} */,
  {32'hbbc306e8, 32'h3d77bda7} /* (27, 3, 15) {real, imag} */,
  {32'h3d9a9f06, 32'hbd9b3a12} /* (27, 3, 14) {real, imag} */,
  {32'h3cc32bea, 32'h3d090726} /* (27, 3, 13) {real, imag} */,
  {32'h3d05f899, 32'hbd8721bf} /* (27, 3, 12) {real, imag} */,
  {32'h3c7c4b34, 32'h3cf06082} /* (27, 3, 11) {real, imag} */,
  {32'hbdb906fb, 32'hbd4d481a} /* (27, 3, 10) {real, imag} */,
  {32'hbca8ed6d, 32'hbcaea8da} /* (27, 3, 9) {real, imag} */,
  {32'h3c6d41a8, 32'hbd42a7eb} /* (27, 3, 8) {real, imag} */,
  {32'h3b420f30, 32'hbd424dee} /* (27, 3, 7) {real, imag} */,
  {32'hbd1e7b96, 32'hbca0111c} /* (27, 3, 6) {real, imag} */,
  {32'hbe19b458, 32'hbd3bb877} /* (27, 3, 5) {real, imag} */,
  {32'hbdd4971e, 32'hbdb2ee87} /* (27, 3, 4) {real, imag} */,
  {32'hbda30f74, 32'h3dc73a56} /* (27, 3, 3) {real, imag} */,
  {32'h3e943e09, 32'hbf1664c2} /* (27, 3, 2) {real, imag} */,
  {32'hbcecb570, 32'h3f111ea5} /* (27, 3, 1) {real, imag} */,
  {32'hbd9abbc4, 32'h00000000} /* (27, 3, 0) {real, imag} */,
  {32'hbdf9eaec, 32'hbf3e19e0} /* (27, 2, 31) {real, imag} */,
  {32'h3ebae610, 32'h3f2669c1} /* (27, 2, 30) {real, imag} */,
  {32'hbcc70c28, 32'hbc5da488} /* (27, 2, 29) {real, imag} */,
  {32'hbd8924ba, 32'h3e08cd05} /* (27, 2, 28) {real, imag} */,
  {32'hbd925bd9, 32'h3d8ce3be} /* (27, 2, 27) {real, imag} */,
  {32'hbd0c14de, 32'h3daac6be} /* (27, 2, 26) {real, imag} */,
  {32'hbddcf206, 32'hbcb590ff} /* (27, 2, 25) {real, imag} */,
  {32'h3d8d3ae2, 32'h3d838e00} /* (27, 2, 24) {real, imag} */,
  {32'hbd931d5f, 32'hbd3e0a0a} /* (27, 2, 23) {real, imag} */,
  {32'hbc759622, 32'h3de781f4} /* (27, 2, 22) {real, imag} */,
  {32'hbdc4c62e, 32'h3c1046ce} /* (27, 2, 21) {real, imag} */,
  {32'h3da2bb59, 32'h3d19a95a} /* (27, 2, 20) {real, imag} */,
  {32'hbd3d8530, 32'hbdb49d66} /* (27, 2, 19) {real, imag} */,
  {32'h3d1f8482, 32'h3ddaa3de} /* (27, 2, 18) {real, imag} */,
  {32'h3d4b1db8, 32'h3cd08bd3} /* (27, 2, 17) {real, imag} */,
  {32'hbcc00ec0, 32'h00000000} /* (27, 2, 16) {real, imag} */,
  {32'h3d4b1db8, 32'hbcd08bd3} /* (27, 2, 15) {real, imag} */,
  {32'h3d1f8482, 32'hbddaa3de} /* (27, 2, 14) {real, imag} */,
  {32'hbd3d8530, 32'h3db49d66} /* (27, 2, 13) {real, imag} */,
  {32'h3da2bb59, 32'hbd19a95a} /* (27, 2, 12) {real, imag} */,
  {32'hbdc4c62e, 32'hbc1046ce} /* (27, 2, 11) {real, imag} */,
  {32'hbc759622, 32'hbde781f4} /* (27, 2, 10) {real, imag} */,
  {32'hbd931d5f, 32'h3d3e0a0a} /* (27, 2, 9) {real, imag} */,
  {32'h3d8d3ae2, 32'hbd838e00} /* (27, 2, 8) {real, imag} */,
  {32'hbddcf206, 32'h3cb590ff} /* (27, 2, 7) {real, imag} */,
  {32'hbd0c14de, 32'hbdaac6be} /* (27, 2, 6) {real, imag} */,
  {32'hbd925bd9, 32'hbd8ce3be} /* (27, 2, 5) {real, imag} */,
  {32'hbd8924ba, 32'hbe08cd05} /* (27, 2, 4) {real, imag} */,
  {32'hbcc70c28, 32'h3c5da488} /* (27, 2, 3) {real, imag} */,
  {32'h3ebae610, 32'hbf2669c1} /* (27, 2, 2) {real, imag} */,
  {32'hbdf9eaec, 32'h3f3e19e0} /* (27, 2, 1) {real, imag} */,
  {32'hbe70427a, 32'h00000000} /* (27, 2, 0) {real, imag} */,
  {32'hbde45e12, 32'hbf56e2b8} /* (27, 1, 31) {real, imag} */,
  {32'h3ee5d5ea, 32'h3f2b7416} /* (27, 1, 30) {real, imag} */,
  {32'hbc0b85e8, 32'hbc40dcde} /* (27, 1, 29) {real, imag} */,
  {32'h3cea2a34, 32'h3ddcfacc} /* (27, 1, 28) {real, imag} */,
  {32'hbdd5b77d, 32'hbde1e79c} /* (27, 1, 27) {real, imag} */,
  {32'h3d1f323a, 32'h3d88ba94} /* (27, 1, 26) {real, imag} */,
  {32'hbd1a48d2, 32'hbc9d62ff} /* (27, 1, 25) {real, imag} */,
  {32'hbdb7bf3e, 32'h3d2b4dac} /* (27, 1, 24) {real, imag} */,
  {32'hbc6c2922, 32'h396ac700} /* (27, 1, 23) {real, imag} */,
  {32'h3d436009, 32'h3d0f9a78} /* (27, 1, 22) {real, imag} */,
  {32'hbe382c62, 32'h3dace78c} /* (27, 1, 21) {real, imag} */,
  {32'h3d3ba695, 32'h3d7a37b8} /* (27, 1, 20) {real, imag} */,
  {32'h3d6f1d80, 32'hbb0fec2c} /* (27, 1, 19) {real, imag} */,
  {32'h3daadf5e, 32'hbc4a831a} /* (27, 1, 18) {real, imag} */,
  {32'hbc6d72d8, 32'hbd3ea032} /* (27, 1, 17) {real, imag} */,
  {32'hbd6c3d1c, 32'h00000000} /* (27, 1, 16) {real, imag} */,
  {32'hbc6d72d8, 32'h3d3ea032} /* (27, 1, 15) {real, imag} */,
  {32'h3daadf5e, 32'h3c4a831a} /* (27, 1, 14) {real, imag} */,
  {32'h3d6f1d80, 32'h3b0fec2c} /* (27, 1, 13) {real, imag} */,
  {32'h3d3ba695, 32'hbd7a37b8} /* (27, 1, 12) {real, imag} */,
  {32'hbe382c62, 32'hbdace78c} /* (27, 1, 11) {real, imag} */,
  {32'h3d436009, 32'hbd0f9a78} /* (27, 1, 10) {real, imag} */,
  {32'hbc6c2922, 32'hb96ac700} /* (27, 1, 9) {real, imag} */,
  {32'hbdb7bf3e, 32'hbd2b4dac} /* (27, 1, 8) {real, imag} */,
  {32'hbd1a48d2, 32'h3c9d62ff} /* (27, 1, 7) {real, imag} */,
  {32'h3d1f323a, 32'hbd88ba94} /* (27, 1, 6) {real, imag} */,
  {32'hbdd5b77d, 32'h3de1e79c} /* (27, 1, 5) {real, imag} */,
  {32'h3cea2a34, 32'hbddcfacc} /* (27, 1, 4) {real, imag} */,
  {32'hbc0b85e8, 32'h3c40dcde} /* (27, 1, 3) {real, imag} */,
  {32'h3ee5d5ea, 32'hbf2b7416} /* (27, 1, 2) {real, imag} */,
  {32'hbde45e12, 32'h3f56e2b8} /* (27, 1, 1) {real, imag} */,
  {32'hbe988256, 32'h00000000} /* (27, 1, 0) {real, imag} */,
  {32'hbe5e3664, 32'hbec00c76} /* (27, 0, 31) {real, imag} */,
  {32'h3d9a2608, 32'h3eeee51a} /* (27, 0, 30) {real, imag} */,
  {32'h3bdfa408, 32'hbd14ea6e} /* (27, 0, 29) {real, imag} */,
  {32'hbba32db0, 32'h3e1bd077} /* (27, 0, 28) {real, imag} */,
  {32'hbe002aae, 32'hbda701bc} /* (27, 0, 27) {real, imag} */,
  {32'hbd8bd4e2, 32'h3c1c634b} /* (27, 0, 26) {real, imag} */,
  {32'h3d97f8e0, 32'hbd73b1cd} /* (27, 0, 25) {real, imag} */,
  {32'hbda3db55, 32'h3aebe300} /* (27, 0, 24) {real, imag} */,
  {32'h3d46ddd5, 32'h3d147a34} /* (27, 0, 23) {real, imag} */,
  {32'h3c202ea8, 32'hbd018563} /* (27, 0, 22) {real, imag} */,
  {32'h3ba86f44, 32'h3d229fc6} /* (27, 0, 21) {real, imag} */,
  {32'h3cb87dbb, 32'h3c8ac761} /* (27, 0, 20) {real, imag} */,
  {32'h3bf19d7d, 32'hbc0faf24} /* (27, 0, 19) {real, imag} */,
  {32'h3cb037c5, 32'hbc8f4794} /* (27, 0, 18) {real, imag} */,
  {32'hbcdd4e26, 32'h3d528134} /* (27, 0, 17) {real, imag} */,
  {32'hbc34c1eb, 32'h00000000} /* (27, 0, 16) {real, imag} */,
  {32'hbcdd4e26, 32'hbd528134} /* (27, 0, 15) {real, imag} */,
  {32'h3cb037c5, 32'h3c8f4794} /* (27, 0, 14) {real, imag} */,
  {32'h3bf19d7d, 32'h3c0faf24} /* (27, 0, 13) {real, imag} */,
  {32'h3cb87dbb, 32'hbc8ac761} /* (27, 0, 12) {real, imag} */,
  {32'h3ba86f44, 32'hbd229fc6} /* (27, 0, 11) {real, imag} */,
  {32'h3c202ea8, 32'h3d018563} /* (27, 0, 10) {real, imag} */,
  {32'h3d46ddd5, 32'hbd147a34} /* (27, 0, 9) {real, imag} */,
  {32'hbda3db55, 32'hbaebe300} /* (27, 0, 8) {real, imag} */,
  {32'h3d97f8e0, 32'h3d73b1cd} /* (27, 0, 7) {real, imag} */,
  {32'hbd8bd4e2, 32'hbc1c634b} /* (27, 0, 6) {real, imag} */,
  {32'hbe002aae, 32'h3da701bc} /* (27, 0, 5) {real, imag} */,
  {32'hbba32db0, 32'hbe1bd077} /* (27, 0, 4) {real, imag} */,
  {32'h3bdfa408, 32'h3d14ea6e} /* (27, 0, 3) {real, imag} */,
  {32'h3d9a2608, 32'hbeeee51a} /* (27, 0, 2) {real, imag} */,
  {32'hbe5e3664, 32'h3ec00c76} /* (27, 0, 1) {real, imag} */,
  {32'hbf1b3cfa, 32'h00000000} /* (27, 0, 0) {real, imag} */,
  {32'hbf52a408, 32'h3f0ba03f} /* (26, 31, 31) {real, imag} */,
  {32'h3d981b33, 32'h3dc49ad2} /* (26, 31, 30) {real, imag} */,
  {32'hbda1b7f2, 32'h3cf3116a} /* (26, 31, 29) {real, imag} */,
  {32'h3d53bfee, 32'h3e072451} /* (26, 31, 28) {real, imag} */,
  {32'h3d2832a8, 32'hbd1fb3ea} /* (26, 31, 27) {real, imag} */,
  {32'h3d978668, 32'h3dca170c} /* (26, 31, 26) {real, imag} */,
  {32'h3d4b0762, 32'h3c9f162e} /* (26, 31, 25) {real, imag} */,
  {32'hbc28c4c8, 32'hbb448d20} /* (26, 31, 24) {real, imag} */,
  {32'h3cbfafa2, 32'h3ca95af7} /* (26, 31, 23) {real, imag} */,
  {32'hbb8f5fc4, 32'hbdb28dc6} /* (26, 31, 22) {real, imag} */,
  {32'h3c87182c, 32'h3d6b9498} /* (26, 31, 21) {real, imag} */,
  {32'h3dba617b, 32'hbcf9f778} /* (26, 31, 20) {real, imag} */,
  {32'h3d8bcc14, 32'hbd8729de} /* (26, 31, 19) {real, imag} */,
  {32'hba9e61b0, 32'h3d83d30e} /* (26, 31, 18) {real, imag} */,
  {32'h3c469201, 32'h3b9d3844} /* (26, 31, 17) {real, imag} */,
  {32'hbd8a5019, 32'h00000000} /* (26, 31, 16) {real, imag} */,
  {32'h3c469201, 32'hbb9d3844} /* (26, 31, 15) {real, imag} */,
  {32'hba9e61b0, 32'hbd83d30e} /* (26, 31, 14) {real, imag} */,
  {32'h3d8bcc14, 32'h3d8729de} /* (26, 31, 13) {real, imag} */,
  {32'h3dba617b, 32'h3cf9f778} /* (26, 31, 12) {real, imag} */,
  {32'h3c87182c, 32'hbd6b9498} /* (26, 31, 11) {real, imag} */,
  {32'hbb8f5fc4, 32'h3db28dc6} /* (26, 31, 10) {real, imag} */,
  {32'h3cbfafa2, 32'hbca95af7} /* (26, 31, 9) {real, imag} */,
  {32'hbc28c4c8, 32'h3b448d20} /* (26, 31, 8) {real, imag} */,
  {32'h3d4b0762, 32'hbc9f162e} /* (26, 31, 7) {real, imag} */,
  {32'h3d978668, 32'hbdca170c} /* (26, 31, 6) {real, imag} */,
  {32'h3d2832a8, 32'h3d1fb3ea} /* (26, 31, 5) {real, imag} */,
  {32'h3d53bfee, 32'hbe072451} /* (26, 31, 4) {real, imag} */,
  {32'hbda1b7f2, 32'hbcf3116a} /* (26, 31, 3) {real, imag} */,
  {32'h3d981b33, 32'hbdc49ad2} /* (26, 31, 2) {real, imag} */,
  {32'hbf52a408, 32'hbf0ba03f} /* (26, 31, 1) {real, imag} */,
  {32'hbfe70ef1, 32'h00000000} /* (26, 31, 0) {real, imag} */,
  {32'hbf4a1c0b, 32'h3ef3b043} /* (26, 30, 31) {real, imag} */,
  {32'h3bc77e90, 32'h3e1ecf14} /* (26, 30, 30) {real, imag} */,
  {32'hbdf0fc6c, 32'hbc7b8ef6} /* (26, 30, 29) {real, imag} */,
  {32'hbdb4754c, 32'h3c1715c9} /* (26, 30, 28) {real, imag} */,
  {32'hbc010c60, 32'hbdbd318f} /* (26, 30, 27) {real, imag} */,
  {32'h3da0a660, 32'h3d11b2a6} /* (26, 30, 26) {real, imag} */,
  {32'h3d505db4, 32'h3d7285ce} /* (26, 30, 25) {real, imag} */,
  {32'hbd8fcb72, 32'hbda83490} /* (26, 30, 24) {real, imag} */,
  {32'hbce11a3e, 32'hbd23867a} /* (26, 30, 23) {real, imag} */,
  {32'h3a0b1b90, 32'hbc877898} /* (26, 30, 22) {real, imag} */,
  {32'h3c30ef74, 32'h3df9c3ee} /* (26, 30, 21) {real, imag} */,
  {32'h3c0ea896, 32'hbd9d5c26} /* (26, 30, 20) {real, imag} */,
  {32'h3c9f5c5d, 32'h3cf185e9} /* (26, 30, 19) {real, imag} */,
  {32'h3d0c60df, 32'hbd737058} /* (26, 30, 18) {real, imag} */,
  {32'hbcca1767, 32'hbd852262} /* (26, 30, 17) {real, imag} */,
  {32'h3d8d9922, 32'h00000000} /* (26, 30, 16) {real, imag} */,
  {32'hbcca1767, 32'h3d852262} /* (26, 30, 15) {real, imag} */,
  {32'h3d0c60df, 32'h3d737058} /* (26, 30, 14) {real, imag} */,
  {32'h3c9f5c5d, 32'hbcf185e9} /* (26, 30, 13) {real, imag} */,
  {32'h3c0ea896, 32'h3d9d5c26} /* (26, 30, 12) {real, imag} */,
  {32'h3c30ef74, 32'hbdf9c3ee} /* (26, 30, 11) {real, imag} */,
  {32'h3a0b1b90, 32'h3c877898} /* (26, 30, 10) {real, imag} */,
  {32'hbce11a3e, 32'h3d23867a} /* (26, 30, 9) {real, imag} */,
  {32'hbd8fcb72, 32'h3da83490} /* (26, 30, 8) {real, imag} */,
  {32'h3d505db4, 32'hbd7285ce} /* (26, 30, 7) {real, imag} */,
  {32'h3da0a660, 32'hbd11b2a6} /* (26, 30, 6) {real, imag} */,
  {32'hbc010c60, 32'h3dbd318f} /* (26, 30, 5) {real, imag} */,
  {32'hbdb4754c, 32'hbc1715c9} /* (26, 30, 4) {real, imag} */,
  {32'hbdf0fc6c, 32'h3c7b8ef6} /* (26, 30, 3) {real, imag} */,
  {32'h3bc77e90, 32'hbe1ecf14} /* (26, 30, 2) {real, imag} */,
  {32'hbf4a1c0b, 32'hbef3b043} /* (26, 30, 1) {real, imag} */,
  {32'hbfd7665c, 32'h00000000} /* (26, 30, 0) {real, imag} */,
  {32'hbf3132f3, 32'h3f0751f9} /* (26, 29, 31) {real, imag} */,
  {32'hbd4f7fc4, 32'h3e235a1a} /* (26, 29, 30) {real, imag} */,
  {32'hbd46a39e, 32'hbe1530b4} /* (26, 29, 29) {real, imag} */,
  {32'hbc8feea2, 32'hbd7bc4b3} /* (26, 29, 28) {real, imag} */,
  {32'hbd26e4af, 32'hbd19c4b3} /* (26, 29, 27) {real, imag} */,
  {32'h3bd30fe8, 32'hbe408204} /* (26, 29, 26) {real, imag} */,
  {32'h3e2e2964, 32'h3bb8a67c} /* (26, 29, 25) {real, imag} */,
  {32'hbd12c30d, 32'hbd4cffa8} /* (26, 29, 24) {real, imag} */,
  {32'hbe27881d, 32'hbdf78245} /* (26, 29, 23) {real, imag} */,
  {32'hbd677c6f, 32'hbd03a888} /* (26, 29, 22) {real, imag} */,
  {32'hbd33bfc4, 32'hbc154690} /* (26, 29, 21) {real, imag} */,
  {32'hbd3dc636, 32'hbcbfdefb} /* (26, 29, 20) {real, imag} */,
  {32'h3ccab38a, 32'hbc201268} /* (26, 29, 19) {real, imag} */,
  {32'h3c9540a0, 32'h3d247a21} /* (26, 29, 18) {real, imag} */,
  {32'h3cbf0c3a, 32'h3c067d88} /* (26, 29, 17) {real, imag} */,
  {32'h3c213c14, 32'h00000000} /* (26, 29, 16) {real, imag} */,
  {32'h3cbf0c3a, 32'hbc067d88} /* (26, 29, 15) {real, imag} */,
  {32'h3c9540a0, 32'hbd247a21} /* (26, 29, 14) {real, imag} */,
  {32'h3ccab38a, 32'h3c201268} /* (26, 29, 13) {real, imag} */,
  {32'hbd3dc636, 32'h3cbfdefb} /* (26, 29, 12) {real, imag} */,
  {32'hbd33bfc4, 32'h3c154690} /* (26, 29, 11) {real, imag} */,
  {32'hbd677c6f, 32'h3d03a888} /* (26, 29, 10) {real, imag} */,
  {32'hbe27881d, 32'h3df78245} /* (26, 29, 9) {real, imag} */,
  {32'hbd12c30d, 32'h3d4cffa8} /* (26, 29, 8) {real, imag} */,
  {32'h3e2e2964, 32'hbbb8a67c} /* (26, 29, 7) {real, imag} */,
  {32'h3bd30fe8, 32'h3e408204} /* (26, 29, 6) {real, imag} */,
  {32'hbd26e4af, 32'h3d19c4b3} /* (26, 29, 5) {real, imag} */,
  {32'hbc8feea2, 32'h3d7bc4b3} /* (26, 29, 4) {real, imag} */,
  {32'hbd46a39e, 32'h3e1530b4} /* (26, 29, 3) {real, imag} */,
  {32'hbd4f7fc4, 32'hbe235a1a} /* (26, 29, 2) {real, imag} */,
  {32'hbf3132f3, 32'hbf0751f9} /* (26, 29, 1) {real, imag} */,
  {32'hbfe32cdb, 32'h00000000} /* (26, 29, 0) {real, imag} */,
  {32'hbf25bc40, 32'h3f0c1cdf} /* (26, 28, 31) {real, imag} */,
  {32'hbdd9a4bf, 32'h3e07b51e} /* (26, 28, 30) {real, imag} */,
  {32'h3da140f4, 32'hbe352b96} /* (26, 28, 29) {real, imag} */,
  {32'h3d699df1, 32'hbca6ceb6} /* (26, 28, 28) {real, imag} */,
  {32'h3d3fdaf3, 32'hbd851dee} /* (26, 28, 27) {real, imag} */,
  {32'h3db8c25b, 32'h3e34c8e8} /* (26, 28, 26) {real, imag} */,
  {32'h3e1125f0, 32'hbd005a54} /* (26, 28, 25) {real, imag} */,
  {32'h3a94b580, 32'h3c80f63c} /* (26, 28, 24) {real, imag} */,
  {32'hbcd56f90, 32'hbe0cd4a8} /* (26, 28, 23) {real, imag} */,
  {32'hbe178ae4, 32'h3d3a531a} /* (26, 28, 22) {real, imag} */,
  {32'h3d09a594, 32'h3b8a5638} /* (26, 28, 21) {real, imag} */,
  {32'h3c3d904e, 32'h3e073983} /* (26, 28, 20) {real, imag} */,
  {32'hbca7d5b4, 32'hbd7b4d69} /* (26, 28, 19) {real, imag} */,
  {32'h3cebcfd5, 32'h3d870926} /* (26, 28, 18) {real, imag} */,
  {32'h3d3a906f, 32'hbd651f14} /* (26, 28, 17) {real, imag} */,
  {32'h3dba4bc4, 32'h00000000} /* (26, 28, 16) {real, imag} */,
  {32'h3d3a906f, 32'h3d651f14} /* (26, 28, 15) {real, imag} */,
  {32'h3cebcfd5, 32'hbd870926} /* (26, 28, 14) {real, imag} */,
  {32'hbca7d5b4, 32'h3d7b4d69} /* (26, 28, 13) {real, imag} */,
  {32'h3c3d904e, 32'hbe073983} /* (26, 28, 12) {real, imag} */,
  {32'h3d09a594, 32'hbb8a5638} /* (26, 28, 11) {real, imag} */,
  {32'hbe178ae4, 32'hbd3a531a} /* (26, 28, 10) {real, imag} */,
  {32'hbcd56f90, 32'h3e0cd4a8} /* (26, 28, 9) {real, imag} */,
  {32'h3a94b580, 32'hbc80f63c} /* (26, 28, 8) {real, imag} */,
  {32'h3e1125f0, 32'h3d005a54} /* (26, 28, 7) {real, imag} */,
  {32'h3db8c25b, 32'hbe34c8e8} /* (26, 28, 6) {real, imag} */,
  {32'h3d3fdaf3, 32'h3d851dee} /* (26, 28, 5) {real, imag} */,
  {32'h3d699df1, 32'h3ca6ceb6} /* (26, 28, 4) {real, imag} */,
  {32'h3da140f4, 32'h3e352b96} /* (26, 28, 3) {real, imag} */,
  {32'hbdd9a4bf, 32'hbe07b51e} /* (26, 28, 2) {real, imag} */,
  {32'hbf25bc40, 32'hbf0c1cdf} /* (26, 28, 1) {real, imag} */,
  {32'hbfeecf4c, 32'h00000000} /* (26, 28, 0) {real, imag} */,
  {32'hbf3c529a, 32'h3ee5c2f2} /* (26, 27, 31) {real, imag} */,
  {32'hbe13a65a, 32'h3dda5524} /* (26, 27, 30) {real, imag} */,
  {32'h3de2b984, 32'h3c2ad4a4} /* (26, 27, 29) {real, imag} */,
  {32'hbcc6f309, 32'hbc5f8a80} /* (26, 27, 28) {real, imag} */,
  {32'h3cf74c48, 32'h3db7b664} /* (26, 27, 27) {real, imag} */,
  {32'h3e1e479a, 32'h3e177a5a} /* (26, 27, 26) {real, imag} */,
  {32'h3d1b15cb, 32'h3aad8b40} /* (26, 27, 25) {real, imag} */,
  {32'h3d31cac1, 32'hbe323976} /* (26, 27, 24) {real, imag} */,
  {32'h3bae6fd4, 32'hbdd1a580} /* (26, 27, 23) {real, imag} */,
  {32'h3c4f34b0, 32'h3d3d8faf} /* (26, 27, 22) {real, imag} */,
  {32'hbdd86e72, 32'hbd1c69d7} /* (26, 27, 21) {real, imag} */,
  {32'h3ddafc12, 32'h3c8c0c58} /* (26, 27, 20) {real, imag} */,
  {32'hbd59a958, 32'h3dc2b90c} /* (26, 27, 19) {real, imag} */,
  {32'h3cc735ee, 32'h3d73bbaa} /* (26, 27, 18) {real, imag} */,
  {32'hbd7b86b1, 32'hbda40bb7} /* (26, 27, 17) {real, imag} */,
  {32'h3d623b68, 32'h00000000} /* (26, 27, 16) {real, imag} */,
  {32'hbd7b86b1, 32'h3da40bb7} /* (26, 27, 15) {real, imag} */,
  {32'h3cc735ee, 32'hbd73bbaa} /* (26, 27, 14) {real, imag} */,
  {32'hbd59a958, 32'hbdc2b90c} /* (26, 27, 13) {real, imag} */,
  {32'h3ddafc12, 32'hbc8c0c58} /* (26, 27, 12) {real, imag} */,
  {32'hbdd86e72, 32'h3d1c69d7} /* (26, 27, 11) {real, imag} */,
  {32'h3c4f34b0, 32'hbd3d8faf} /* (26, 27, 10) {real, imag} */,
  {32'h3bae6fd4, 32'h3dd1a580} /* (26, 27, 9) {real, imag} */,
  {32'h3d31cac1, 32'h3e323976} /* (26, 27, 8) {real, imag} */,
  {32'h3d1b15cb, 32'hbaad8b40} /* (26, 27, 7) {real, imag} */,
  {32'h3e1e479a, 32'hbe177a5a} /* (26, 27, 6) {real, imag} */,
  {32'h3cf74c48, 32'hbdb7b664} /* (26, 27, 5) {real, imag} */,
  {32'hbcc6f309, 32'h3c5f8a80} /* (26, 27, 4) {real, imag} */,
  {32'h3de2b984, 32'hbc2ad4a4} /* (26, 27, 3) {real, imag} */,
  {32'hbe13a65a, 32'hbdda5524} /* (26, 27, 2) {real, imag} */,
  {32'hbf3c529a, 32'hbee5c2f2} /* (26, 27, 1) {real, imag} */,
  {32'hbfe29bb5, 32'h00000000} /* (26, 27, 0) {real, imag} */,
  {32'hbf451256, 32'h3eb50864} /* (26, 26, 31) {real, imag} */,
  {32'hbe087b43, 32'h3e392f52} /* (26, 26, 30) {real, imag} */,
  {32'hbd24ee06, 32'h3d7185ec} /* (26, 26, 29) {real, imag} */,
  {32'h3d401906, 32'hbd36ec02} /* (26, 26, 28) {real, imag} */,
  {32'hbc64b126, 32'hbd9f9d33} /* (26, 26, 27) {real, imag} */,
  {32'hbba5323e, 32'hbcc05444} /* (26, 26, 26) {real, imag} */,
  {32'h3c9a4609, 32'hbd74bf63} /* (26, 26, 25) {real, imag} */,
  {32'h3bedbd92, 32'hbd577b8b} /* (26, 26, 24) {real, imag} */,
  {32'hbdd71b93, 32'h3c3838d8} /* (26, 26, 23) {real, imag} */,
  {32'h3a9ca450, 32'hbd732ffe} /* (26, 26, 22) {real, imag} */,
  {32'hbcd14bd2, 32'hbd1f0bf0} /* (26, 26, 21) {real, imag} */,
  {32'h3d14918e, 32'hbd8dc008} /* (26, 26, 20) {real, imag} */,
  {32'h3be90af3, 32'h3ca302cc} /* (26, 26, 19) {real, imag} */,
  {32'h3d97cde1, 32'hbd71ec02} /* (26, 26, 18) {real, imag} */,
  {32'h3d48e643, 32'h3d88c817} /* (26, 26, 17) {real, imag} */,
  {32'hbd02dc58, 32'h00000000} /* (26, 26, 16) {real, imag} */,
  {32'h3d48e643, 32'hbd88c817} /* (26, 26, 15) {real, imag} */,
  {32'h3d97cde1, 32'h3d71ec02} /* (26, 26, 14) {real, imag} */,
  {32'h3be90af3, 32'hbca302cc} /* (26, 26, 13) {real, imag} */,
  {32'h3d14918e, 32'h3d8dc008} /* (26, 26, 12) {real, imag} */,
  {32'hbcd14bd2, 32'h3d1f0bf0} /* (26, 26, 11) {real, imag} */,
  {32'h3a9ca450, 32'h3d732ffe} /* (26, 26, 10) {real, imag} */,
  {32'hbdd71b93, 32'hbc3838d8} /* (26, 26, 9) {real, imag} */,
  {32'h3bedbd92, 32'h3d577b8b} /* (26, 26, 8) {real, imag} */,
  {32'h3c9a4609, 32'h3d74bf63} /* (26, 26, 7) {real, imag} */,
  {32'hbba5323e, 32'h3cc05444} /* (26, 26, 6) {real, imag} */,
  {32'hbc64b126, 32'h3d9f9d33} /* (26, 26, 5) {real, imag} */,
  {32'h3d401906, 32'h3d36ec02} /* (26, 26, 4) {real, imag} */,
  {32'hbd24ee06, 32'hbd7185ec} /* (26, 26, 3) {real, imag} */,
  {32'hbe087b43, 32'hbe392f52} /* (26, 26, 2) {real, imag} */,
  {32'hbf451256, 32'hbeb50864} /* (26, 26, 1) {real, imag} */,
  {32'hbffbdf3c, 32'h00000000} /* (26, 26, 0) {real, imag} */,
  {32'hbf440b99, 32'h3ea0a578} /* (26, 25, 31) {real, imag} */,
  {32'hbe10635c, 32'h3e5cb938} /* (26, 25, 30) {real, imag} */,
  {32'hbbe770a0, 32'hbd632145} /* (26, 25, 29) {real, imag} */,
  {32'hbcd4619e, 32'hbd8d68c9} /* (26, 25, 28) {real, imag} */,
  {32'h3ce43796, 32'h3d3d682e} /* (26, 25, 27) {real, imag} */,
  {32'hbcfb93ad, 32'h3c81a77e} /* (26, 25, 26) {real, imag} */,
  {32'h3cf99534, 32'h3b2b26c0} /* (26, 25, 25) {real, imag} */,
  {32'h3e1c8590, 32'h3d1eb82a} /* (26, 25, 24) {real, imag} */,
  {32'hbd1f0791, 32'h3d047680} /* (26, 25, 23) {real, imag} */,
  {32'h3df1535f, 32'hbc9a2939} /* (26, 25, 22) {real, imag} */,
  {32'hbd4bd5a7, 32'hbce9e9f0} /* (26, 25, 21) {real, imag} */,
  {32'h3c94070d, 32'hbc90c1a5} /* (26, 25, 20) {real, imag} */,
  {32'h3cad2dcf, 32'hbd488322} /* (26, 25, 19) {real, imag} */,
  {32'h3c33e618, 32'h3c0d63d2} /* (26, 25, 18) {real, imag} */,
  {32'hbd7722ca, 32'hbd9f573c} /* (26, 25, 17) {real, imag} */,
  {32'h3b86b3f0, 32'h00000000} /* (26, 25, 16) {real, imag} */,
  {32'hbd7722ca, 32'h3d9f573c} /* (26, 25, 15) {real, imag} */,
  {32'h3c33e618, 32'hbc0d63d2} /* (26, 25, 14) {real, imag} */,
  {32'h3cad2dcf, 32'h3d488322} /* (26, 25, 13) {real, imag} */,
  {32'h3c94070d, 32'h3c90c1a5} /* (26, 25, 12) {real, imag} */,
  {32'hbd4bd5a7, 32'h3ce9e9f0} /* (26, 25, 11) {real, imag} */,
  {32'h3df1535f, 32'h3c9a2939} /* (26, 25, 10) {real, imag} */,
  {32'hbd1f0791, 32'hbd047680} /* (26, 25, 9) {real, imag} */,
  {32'h3e1c8590, 32'hbd1eb82a} /* (26, 25, 8) {real, imag} */,
  {32'h3cf99534, 32'hbb2b26c0} /* (26, 25, 7) {real, imag} */,
  {32'hbcfb93ad, 32'hbc81a77e} /* (26, 25, 6) {real, imag} */,
  {32'h3ce43796, 32'hbd3d682e} /* (26, 25, 5) {real, imag} */,
  {32'hbcd4619e, 32'h3d8d68c9} /* (26, 25, 4) {real, imag} */,
  {32'hbbe770a0, 32'h3d632145} /* (26, 25, 3) {real, imag} */,
  {32'hbe10635c, 32'hbe5cb938} /* (26, 25, 2) {real, imag} */,
  {32'hbf440b99, 32'hbea0a578} /* (26, 25, 1) {real, imag} */,
  {32'hbfc9bf53, 32'h00000000} /* (26, 25, 0) {real, imag} */,
  {32'hbf37897a, 32'h3e0a6e54} /* (26, 24, 31) {real, imag} */,
  {32'hbdd806de, 32'h3c8ffe18} /* (26, 24, 30) {real, imag} */,
  {32'hbc03ca00, 32'hbe115f28} /* (26, 24, 29) {real, imag} */,
  {32'h3dda7bd0, 32'hba982300} /* (26, 24, 28) {real, imag} */,
  {32'h3cc5bdc8, 32'h3e2cb779} /* (26, 24, 27) {real, imag} */,
  {32'hbe240640, 32'hbd6b47d3} /* (26, 24, 26) {real, imag} */,
  {32'h3d52f18c, 32'h3d58fe56} /* (26, 24, 25) {real, imag} */,
  {32'hbd802810, 32'h3c692986} /* (26, 24, 24) {real, imag} */,
  {32'hbcc5fadd, 32'hbdc50628} /* (26, 24, 23) {real, imag} */,
  {32'hbbe8f010, 32'h3cdb0251} /* (26, 24, 22) {real, imag} */,
  {32'h3b746390, 32'h3d46273c} /* (26, 24, 21) {real, imag} */,
  {32'h3de76f38, 32'h3b53b8b0} /* (26, 24, 20) {real, imag} */,
  {32'h3c9725eb, 32'hbd03a6d7} /* (26, 24, 19) {real, imag} */,
  {32'hbd4dd33c, 32'hbde4c397} /* (26, 24, 18) {real, imag} */,
  {32'hbd8d78de, 32'h3da9856b} /* (26, 24, 17) {real, imag} */,
  {32'hbd28f64c, 32'h00000000} /* (26, 24, 16) {real, imag} */,
  {32'hbd8d78de, 32'hbda9856b} /* (26, 24, 15) {real, imag} */,
  {32'hbd4dd33c, 32'h3de4c397} /* (26, 24, 14) {real, imag} */,
  {32'h3c9725eb, 32'h3d03a6d7} /* (26, 24, 13) {real, imag} */,
  {32'h3de76f38, 32'hbb53b8b0} /* (26, 24, 12) {real, imag} */,
  {32'h3b746390, 32'hbd46273c} /* (26, 24, 11) {real, imag} */,
  {32'hbbe8f010, 32'hbcdb0251} /* (26, 24, 10) {real, imag} */,
  {32'hbcc5fadd, 32'h3dc50628} /* (26, 24, 9) {real, imag} */,
  {32'hbd802810, 32'hbc692986} /* (26, 24, 8) {real, imag} */,
  {32'h3d52f18c, 32'hbd58fe56} /* (26, 24, 7) {real, imag} */,
  {32'hbe240640, 32'h3d6b47d3} /* (26, 24, 6) {real, imag} */,
  {32'h3cc5bdc8, 32'hbe2cb779} /* (26, 24, 5) {real, imag} */,
  {32'h3dda7bd0, 32'h3a982300} /* (26, 24, 4) {real, imag} */,
  {32'hbc03ca00, 32'h3e115f28} /* (26, 24, 3) {real, imag} */,
  {32'hbdd806de, 32'hbc8ffe18} /* (26, 24, 2) {real, imag} */,
  {32'hbf37897a, 32'hbe0a6e54} /* (26, 24, 1) {real, imag} */,
  {32'hbfa13e26, 32'h00000000} /* (26, 24, 0) {real, imag} */,
  {32'hbf380274, 32'h3e053868} /* (26, 23, 31) {real, imag} */,
  {32'h3ca14518, 32'hbcc15e34} /* (26, 23, 30) {real, imag} */,
  {32'h3c552e80, 32'hbd8e6558} /* (26, 23, 29) {real, imag} */,
  {32'h3ddba475, 32'hbbf1cfb4} /* (26, 23, 28) {real, imag} */,
  {32'hbd27cafd, 32'h3e85bd65} /* (26, 23, 27) {real, imag} */,
  {32'hbd22ca6e, 32'hbca8ec36} /* (26, 23, 26) {real, imag} */,
  {32'hbc914228, 32'h3cd5cc94} /* (26, 23, 25) {real, imag} */,
  {32'hbdcb48b4, 32'hbe071056} /* (26, 23, 24) {real, imag} */,
  {32'hbca3e03c, 32'hba5e49d8} /* (26, 23, 23) {real, imag} */,
  {32'hbd3d3b58, 32'h3d3c4000} /* (26, 23, 22) {real, imag} */,
  {32'hbd06478f, 32'h3d4813f2} /* (26, 23, 21) {real, imag} */,
  {32'h3b40056c, 32'hbcccdf9d} /* (26, 23, 20) {real, imag} */,
  {32'h3da72df1, 32'h385b1200} /* (26, 23, 19) {real, imag} */,
  {32'hbdbdffc7, 32'hbd2283d0} /* (26, 23, 18) {real, imag} */,
  {32'h3d7f52f8, 32'hbb9737f6} /* (26, 23, 17) {real, imag} */,
  {32'hbd2ea0f0, 32'h00000000} /* (26, 23, 16) {real, imag} */,
  {32'h3d7f52f8, 32'h3b9737f6} /* (26, 23, 15) {real, imag} */,
  {32'hbdbdffc7, 32'h3d2283d0} /* (26, 23, 14) {real, imag} */,
  {32'h3da72df1, 32'hb85b1200} /* (26, 23, 13) {real, imag} */,
  {32'h3b40056c, 32'h3cccdf9d} /* (26, 23, 12) {real, imag} */,
  {32'hbd06478f, 32'hbd4813f2} /* (26, 23, 11) {real, imag} */,
  {32'hbd3d3b58, 32'hbd3c4000} /* (26, 23, 10) {real, imag} */,
  {32'hbca3e03c, 32'h3a5e49d8} /* (26, 23, 9) {real, imag} */,
  {32'hbdcb48b4, 32'h3e071056} /* (26, 23, 8) {real, imag} */,
  {32'hbc914228, 32'hbcd5cc94} /* (26, 23, 7) {real, imag} */,
  {32'hbd22ca6e, 32'h3ca8ec36} /* (26, 23, 6) {real, imag} */,
  {32'hbd27cafd, 32'hbe85bd65} /* (26, 23, 5) {real, imag} */,
  {32'h3ddba475, 32'h3bf1cfb4} /* (26, 23, 4) {real, imag} */,
  {32'h3c552e80, 32'h3d8e6558} /* (26, 23, 3) {real, imag} */,
  {32'h3ca14518, 32'h3cc15e34} /* (26, 23, 2) {real, imag} */,
  {32'hbf380274, 32'hbe053868} /* (26, 23, 1) {real, imag} */,
  {32'hbf8ad002, 32'h00000000} /* (26, 23, 0) {real, imag} */,
  {32'hbf05fb36, 32'h3e8b8853} /* (26, 22, 31) {real, imag} */,
  {32'h3d95af9d, 32'hbd8832ca} /* (26, 22, 30) {real, imag} */,
  {32'h3d3655c2, 32'h3d22eac4} /* (26, 22, 29) {real, imag} */,
  {32'h3de8303d, 32'hbc9d1104} /* (26, 22, 28) {real, imag} */,
  {32'hbd7a4ff6, 32'h3d14eabe} /* (26, 22, 27) {real, imag} */,
  {32'h3c523a70, 32'h3dcf31b4} /* (26, 22, 26) {real, imag} */,
  {32'hbda11ab8, 32'hbd8c9bd4} /* (26, 22, 25) {real, imag} */,
  {32'hbd99fbbd, 32'hbd559152} /* (26, 22, 24) {real, imag} */,
  {32'h3dc5bdb5, 32'h3d529b6c} /* (26, 22, 23) {real, imag} */,
  {32'hbc35fc44, 32'hbd2a21ca} /* (26, 22, 22) {real, imag} */,
  {32'h3c19259c, 32'hbc75c5d8} /* (26, 22, 21) {real, imag} */,
  {32'hbd553c76, 32'hbd3e9c86} /* (26, 22, 20) {real, imag} */,
  {32'h3c9b3621, 32'h3d921e73} /* (26, 22, 19) {real, imag} */,
  {32'hbc4094ee, 32'h3d08b1b8} /* (26, 22, 18) {real, imag} */,
  {32'hbcfb19cc, 32'hbd2e139e} /* (26, 22, 17) {real, imag} */,
  {32'h3d2feff2, 32'h00000000} /* (26, 22, 16) {real, imag} */,
  {32'hbcfb19cc, 32'h3d2e139e} /* (26, 22, 15) {real, imag} */,
  {32'hbc4094ee, 32'hbd08b1b8} /* (26, 22, 14) {real, imag} */,
  {32'h3c9b3621, 32'hbd921e73} /* (26, 22, 13) {real, imag} */,
  {32'hbd553c76, 32'h3d3e9c86} /* (26, 22, 12) {real, imag} */,
  {32'h3c19259c, 32'h3c75c5d8} /* (26, 22, 11) {real, imag} */,
  {32'hbc35fc44, 32'h3d2a21ca} /* (26, 22, 10) {real, imag} */,
  {32'h3dc5bdb5, 32'hbd529b6c} /* (26, 22, 9) {real, imag} */,
  {32'hbd99fbbd, 32'h3d559152} /* (26, 22, 8) {real, imag} */,
  {32'hbda11ab8, 32'h3d8c9bd4} /* (26, 22, 7) {real, imag} */,
  {32'h3c523a70, 32'hbdcf31b4} /* (26, 22, 6) {real, imag} */,
  {32'hbd7a4ff6, 32'hbd14eabe} /* (26, 22, 5) {real, imag} */,
  {32'h3de8303d, 32'h3c9d1104} /* (26, 22, 4) {real, imag} */,
  {32'h3d3655c2, 32'hbd22eac4} /* (26, 22, 3) {real, imag} */,
  {32'h3d95af9d, 32'h3d8832ca} /* (26, 22, 2) {real, imag} */,
  {32'hbf05fb36, 32'hbe8b8853} /* (26, 22, 1) {real, imag} */,
  {32'hbef01824, 32'h00000000} /* (26, 22, 0) {real, imag} */,
  {32'hbecbdf6a, 32'h3e8fc76e} /* (26, 21, 31) {real, imag} */,
  {32'h3e67fd9f, 32'h3dffa153} /* (26, 21, 30) {real, imag} */,
  {32'h3c667e94, 32'h3cb06dba} /* (26, 21, 29) {real, imag} */,
  {32'hbccbe894, 32'hbd95a00a} /* (26, 21, 28) {real, imag} */,
  {32'h3d5a5c5f, 32'hbd4338be} /* (26, 21, 27) {real, imag} */,
  {32'h3d1ed5ef, 32'h3d98050f} /* (26, 21, 26) {real, imag} */,
  {32'hbcbdbeba, 32'h3b147b60} /* (26, 21, 25) {real, imag} */,
  {32'hbe1d92a0, 32'h3db0ba1a} /* (26, 21, 24) {real, imag} */,
  {32'h3b0958b8, 32'hbd843f1e} /* (26, 21, 23) {real, imag} */,
  {32'h3cf33632, 32'hbd957fce} /* (26, 21, 22) {real, imag} */,
  {32'h3c407074, 32'h3de20958} /* (26, 21, 21) {real, imag} */,
  {32'h3d1b16ad, 32'hbd2ce66a} /* (26, 21, 20) {real, imag} */,
  {32'hbc9493e8, 32'hbbb91e44} /* (26, 21, 19) {real, imag} */,
  {32'h3d2c065e, 32'hbd31e4cd} /* (26, 21, 18) {real, imag} */,
  {32'hbbbd3d0a, 32'h3cb1f41e} /* (26, 21, 17) {real, imag} */,
  {32'h3dd03896, 32'h00000000} /* (26, 21, 16) {real, imag} */,
  {32'hbbbd3d0a, 32'hbcb1f41e} /* (26, 21, 15) {real, imag} */,
  {32'h3d2c065e, 32'h3d31e4cd} /* (26, 21, 14) {real, imag} */,
  {32'hbc9493e8, 32'h3bb91e44} /* (26, 21, 13) {real, imag} */,
  {32'h3d1b16ad, 32'h3d2ce66a} /* (26, 21, 12) {real, imag} */,
  {32'h3c407074, 32'hbde20958} /* (26, 21, 11) {real, imag} */,
  {32'h3cf33632, 32'h3d957fce} /* (26, 21, 10) {real, imag} */,
  {32'h3b0958b8, 32'h3d843f1e} /* (26, 21, 9) {real, imag} */,
  {32'hbe1d92a0, 32'hbdb0ba1a} /* (26, 21, 8) {real, imag} */,
  {32'hbcbdbeba, 32'hbb147b60} /* (26, 21, 7) {real, imag} */,
  {32'h3d1ed5ef, 32'hbd98050f} /* (26, 21, 6) {real, imag} */,
  {32'h3d5a5c5f, 32'h3d4338be} /* (26, 21, 5) {real, imag} */,
  {32'hbccbe894, 32'h3d95a00a} /* (26, 21, 4) {real, imag} */,
  {32'h3c667e94, 32'hbcb06dba} /* (26, 21, 3) {real, imag} */,
  {32'h3e67fd9f, 32'hbdffa153} /* (26, 21, 2) {real, imag} */,
  {32'hbecbdf6a, 32'hbe8fc76e} /* (26, 21, 1) {real, imag} */,
  {32'hbea2f3fe, 32'h00000000} /* (26, 21, 0) {real, imag} */,
  {32'hbe9fbed2, 32'hbc05ede4} /* (26, 20, 31) {real, imag} */,
  {32'h3e40896c, 32'hbcd908e9} /* (26, 20, 30) {real, imag} */,
  {32'h3d2e3511, 32'hbd992766} /* (26, 20, 29) {real, imag} */,
  {32'h3d8a5fac, 32'hbdbf372d} /* (26, 20, 28) {real, imag} */,
  {32'hbd8042d3, 32'h3d9aa6ad} /* (26, 20, 27) {real, imag} */,
  {32'hbd8719f6, 32'h3da1ce6e} /* (26, 20, 26) {real, imag} */,
  {32'h3b63c1f0, 32'hbd8bd2a8} /* (26, 20, 25) {real, imag} */,
  {32'h3d6516f9, 32'hbd5c0780} /* (26, 20, 24) {real, imag} */,
  {32'h3c970562, 32'h3be8e280} /* (26, 20, 23) {real, imag} */,
  {32'hbc2c9ece, 32'hbbf4a1b8} /* (26, 20, 22) {real, imag} */,
  {32'h3c5d51ce, 32'hbc297863} /* (26, 20, 21) {real, imag} */,
  {32'hbcefcfbd, 32'hbc17dd8c} /* (26, 20, 20) {real, imag} */,
  {32'hbdccbf10, 32'h3d1f2119} /* (26, 20, 19) {real, imag} */,
  {32'h39973ec0, 32'hbc57d766} /* (26, 20, 18) {real, imag} */,
  {32'h3cbdc3bc, 32'h3c1df496} /* (26, 20, 17) {real, imag} */,
  {32'h3d68ca20, 32'h00000000} /* (26, 20, 16) {real, imag} */,
  {32'h3cbdc3bc, 32'hbc1df496} /* (26, 20, 15) {real, imag} */,
  {32'h39973ec0, 32'h3c57d766} /* (26, 20, 14) {real, imag} */,
  {32'hbdccbf10, 32'hbd1f2119} /* (26, 20, 13) {real, imag} */,
  {32'hbcefcfbd, 32'h3c17dd8c} /* (26, 20, 12) {real, imag} */,
  {32'h3c5d51ce, 32'h3c297863} /* (26, 20, 11) {real, imag} */,
  {32'hbc2c9ece, 32'h3bf4a1b8} /* (26, 20, 10) {real, imag} */,
  {32'h3c970562, 32'hbbe8e280} /* (26, 20, 9) {real, imag} */,
  {32'h3d6516f9, 32'h3d5c0780} /* (26, 20, 8) {real, imag} */,
  {32'h3b63c1f0, 32'h3d8bd2a8} /* (26, 20, 7) {real, imag} */,
  {32'hbd8719f6, 32'hbda1ce6e} /* (26, 20, 6) {real, imag} */,
  {32'hbd8042d3, 32'hbd9aa6ad} /* (26, 20, 5) {real, imag} */,
  {32'h3d8a5fac, 32'h3dbf372d} /* (26, 20, 4) {real, imag} */,
  {32'h3d2e3511, 32'h3d992766} /* (26, 20, 3) {real, imag} */,
  {32'h3e40896c, 32'h3cd908e9} /* (26, 20, 2) {real, imag} */,
  {32'hbe9fbed2, 32'h3c05ede4} /* (26, 20, 1) {real, imag} */,
  {32'hbe8c6a42, 32'h00000000} /* (26, 20, 0) {real, imag} */,
  {32'hbe7f8a12, 32'h3d1ebac2} /* (26, 19, 31) {real, imag} */,
  {32'h3e0a1430, 32'hbe42db7a} /* (26, 19, 30) {real, imag} */,
  {32'h3d69c5dc, 32'hbd28fde8} /* (26, 19, 29) {real, imag} */,
  {32'h3e292aed, 32'hbd88701a} /* (26, 19, 28) {real, imag} */,
  {32'h3c698a38, 32'h3d86ff4e} /* (26, 19, 27) {real, imag} */,
  {32'h3d448a58, 32'hbc3d4914} /* (26, 19, 26) {real, imag} */,
  {32'hbd959086, 32'h3d4d5e46} /* (26, 19, 25) {real, imag} */,
  {32'h3c9845d2, 32'hbdc03baa} /* (26, 19, 24) {real, imag} */,
  {32'hbdc78ca6, 32'h3d3397b4} /* (26, 19, 23) {real, imag} */,
  {32'h3cb7c73e, 32'hbd51a0d8} /* (26, 19, 22) {real, imag} */,
  {32'hbd500e62, 32'hbce3db68} /* (26, 19, 21) {real, imag} */,
  {32'h3d783dce, 32'h3be8e016} /* (26, 19, 20) {real, imag} */,
  {32'hbdc6d3a2, 32'h3dc24de8} /* (26, 19, 19) {real, imag} */,
  {32'h3d295d1a, 32'h3d3e51f0} /* (26, 19, 18) {real, imag} */,
  {32'h3babcac0, 32'h3c96274f} /* (26, 19, 17) {real, imag} */,
  {32'h3d0b7f9c, 32'h00000000} /* (26, 19, 16) {real, imag} */,
  {32'h3babcac0, 32'hbc96274f} /* (26, 19, 15) {real, imag} */,
  {32'h3d295d1a, 32'hbd3e51f0} /* (26, 19, 14) {real, imag} */,
  {32'hbdc6d3a2, 32'hbdc24de8} /* (26, 19, 13) {real, imag} */,
  {32'h3d783dce, 32'hbbe8e016} /* (26, 19, 12) {real, imag} */,
  {32'hbd500e62, 32'h3ce3db68} /* (26, 19, 11) {real, imag} */,
  {32'h3cb7c73e, 32'h3d51a0d8} /* (26, 19, 10) {real, imag} */,
  {32'hbdc78ca6, 32'hbd3397b4} /* (26, 19, 9) {real, imag} */,
  {32'h3c9845d2, 32'h3dc03baa} /* (26, 19, 8) {real, imag} */,
  {32'hbd959086, 32'hbd4d5e46} /* (26, 19, 7) {real, imag} */,
  {32'h3d448a58, 32'h3c3d4914} /* (26, 19, 6) {real, imag} */,
  {32'h3c698a38, 32'hbd86ff4e} /* (26, 19, 5) {real, imag} */,
  {32'h3e292aed, 32'h3d88701a} /* (26, 19, 4) {real, imag} */,
  {32'h3d69c5dc, 32'h3d28fde8} /* (26, 19, 3) {real, imag} */,
  {32'h3e0a1430, 32'h3e42db7a} /* (26, 19, 2) {real, imag} */,
  {32'hbe7f8a12, 32'hbd1ebac2} /* (26, 19, 1) {real, imag} */,
  {32'hbd4f2cce, 32'h00000000} /* (26, 19, 0) {real, imag} */,
  {32'hbc4b41b0, 32'h3e15b7b6} /* (26, 18, 31) {real, imag} */,
  {32'h3e2f5602, 32'hbe25420a} /* (26, 18, 30) {real, imag} */,
  {32'h3b61a0f8, 32'hbe02bf5c} /* (26, 18, 29) {real, imag} */,
  {32'h3dee0968, 32'h3cd1b17e} /* (26, 18, 28) {real, imag} */,
  {32'h3ca3406a, 32'h3c888484} /* (26, 18, 27) {real, imag} */,
  {32'h3de96b2d, 32'hbdafb8c4} /* (26, 18, 26) {real, imag} */,
  {32'hbdb15c77, 32'h3dd5b624} /* (26, 18, 25) {real, imag} */,
  {32'hbd7a6935, 32'hbc108ba8} /* (26, 18, 24) {real, imag} */,
  {32'h3ce6c070, 32'h3c6a5ea5} /* (26, 18, 23) {real, imag} */,
  {32'hbd8abc54, 32'hbbda53a0} /* (26, 18, 22) {real, imag} */,
  {32'hbd88c2c6, 32'hbdaea71e} /* (26, 18, 21) {real, imag} */,
  {32'hbc1016c2, 32'hbc6744ca} /* (26, 18, 20) {real, imag} */,
  {32'hbd0cf760, 32'hbd3a52a4} /* (26, 18, 19) {real, imag} */,
  {32'hbd72cfc0, 32'h3c928647} /* (26, 18, 18) {real, imag} */,
  {32'h3c792552, 32'h3b45c9d8} /* (26, 18, 17) {real, imag} */,
  {32'hbd3dba8c, 32'h00000000} /* (26, 18, 16) {real, imag} */,
  {32'h3c792552, 32'hbb45c9d8} /* (26, 18, 15) {real, imag} */,
  {32'hbd72cfc0, 32'hbc928647} /* (26, 18, 14) {real, imag} */,
  {32'hbd0cf760, 32'h3d3a52a4} /* (26, 18, 13) {real, imag} */,
  {32'hbc1016c2, 32'h3c6744ca} /* (26, 18, 12) {real, imag} */,
  {32'hbd88c2c6, 32'h3daea71e} /* (26, 18, 11) {real, imag} */,
  {32'hbd8abc54, 32'h3bda53a0} /* (26, 18, 10) {real, imag} */,
  {32'h3ce6c070, 32'hbc6a5ea5} /* (26, 18, 9) {real, imag} */,
  {32'hbd7a6935, 32'h3c108ba8} /* (26, 18, 8) {real, imag} */,
  {32'hbdb15c77, 32'hbdd5b624} /* (26, 18, 7) {real, imag} */,
  {32'h3de96b2d, 32'h3dafb8c4} /* (26, 18, 6) {real, imag} */,
  {32'h3ca3406a, 32'hbc888484} /* (26, 18, 5) {real, imag} */,
  {32'h3dee0968, 32'hbcd1b17e} /* (26, 18, 4) {real, imag} */,
  {32'h3b61a0f8, 32'h3e02bf5c} /* (26, 18, 3) {real, imag} */,
  {32'h3e2f5602, 32'h3e25420a} /* (26, 18, 2) {real, imag} */,
  {32'hbc4b41b0, 32'hbe15b7b6} /* (26, 18, 1) {real, imag} */,
  {32'h3d124940, 32'h00000000} /* (26, 18, 0) {real, imag} */,
  {32'h3d647b58, 32'h3e43adac} /* (26, 17, 31) {real, imag} */,
  {32'h3d48a97f, 32'hbdca7066} /* (26, 17, 30) {real, imag} */,
  {32'hbe1130d5, 32'hbe130cce} /* (26, 17, 29) {real, imag} */,
  {32'h3e152bb8, 32'h3b960ac4} /* (26, 17, 28) {real, imag} */,
  {32'h3ca0caf9, 32'hbbb6a2cc} /* (26, 17, 27) {real, imag} */,
  {32'h3d953445, 32'hbc70c04c} /* (26, 17, 26) {real, imag} */,
  {32'h3b8a16d0, 32'hbbe89448} /* (26, 17, 25) {real, imag} */,
  {32'hbdb4ecd0, 32'hbce9721c} /* (26, 17, 24) {real, imag} */,
  {32'h3d945ab2, 32'h3d03d34d} /* (26, 17, 23) {real, imag} */,
  {32'h3d7288b1, 32'h3d6591ea} /* (26, 17, 22) {real, imag} */,
  {32'h3d98cb4e, 32'h3c3a5f56} /* (26, 17, 21) {real, imag} */,
  {32'hbd555128, 32'h3c893337} /* (26, 17, 20) {real, imag} */,
  {32'hbd9d735a, 32'hbdcb502b} /* (26, 17, 19) {real, imag} */,
  {32'hbd869f82, 32'hbbcebf80} /* (26, 17, 18) {real, imag} */,
  {32'hbcdb0d09, 32'h3cd38be8} /* (26, 17, 17) {real, imag} */,
  {32'h3cab6994, 32'h00000000} /* (26, 17, 16) {real, imag} */,
  {32'hbcdb0d09, 32'hbcd38be8} /* (26, 17, 15) {real, imag} */,
  {32'hbd869f82, 32'h3bcebf80} /* (26, 17, 14) {real, imag} */,
  {32'hbd9d735a, 32'h3dcb502b} /* (26, 17, 13) {real, imag} */,
  {32'hbd555128, 32'hbc893337} /* (26, 17, 12) {real, imag} */,
  {32'h3d98cb4e, 32'hbc3a5f56} /* (26, 17, 11) {real, imag} */,
  {32'h3d7288b1, 32'hbd6591ea} /* (26, 17, 10) {real, imag} */,
  {32'h3d945ab2, 32'hbd03d34d} /* (26, 17, 9) {real, imag} */,
  {32'hbdb4ecd0, 32'h3ce9721c} /* (26, 17, 8) {real, imag} */,
  {32'h3b8a16d0, 32'h3be89448} /* (26, 17, 7) {real, imag} */,
  {32'h3d953445, 32'h3c70c04c} /* (26, 17, 6) {real, imag} */,
  {32'h3ca0caf9, 32'h3bb6a2cc} /* (26, 17, 5) {real, imag} */,
  {32'h3e152bb8, 32'hbb960ac4} /* (26, 17, 4) {real, imag} */,
  {32'hbe1130d5, 32'h3e130cce} /* (26, 17, 3) {real, imag} */,
  {32'h3d48a97f, 32'h3dca7066} /* (26, 17, 2) {real, imag} */,
  {32'h3d647b58, 32'hbe43adac} /* (26, 17, 1) {real, imag} */,
  {32'h3da99c52, 32'h00000000} /* (26, 17, 0) {real, imag} */,
  {32'h3e1d8860, 32'h3e4c6e82} /* (26, 16, 31) {real, imag} */,
  {32'hbbad04b0, 32'hbd756e20} /* (26, 16, 30) {real, imag} */,
  {32'hbd2cf7f8, 32'hbe00fcbc} /* (26, 16, 29) {real, imag} */,
  {32'h3cc5a3b4, 32'hbd0f5bba} /* (26, 16, 28) {real, imag} */,
  {32'h3d3570c9, 32'hbd8aee3a} /* (26, 16, 27) {real, imag} */,
  {32'h3c0db194, 32'h3d8047bb} /* (26, 16, 26) {real, imag} */,
  {32'h3c97ab59, 32'h3dc15680} /* (26, 16, 25) {real, imag} */,
  {32'h3cd0ae6e, 32'hbc12b786} /* (26, 16, 24) {real, imag} */,
  {32'h3c41b806, 32'h3b836bb0} /* (26, 16, 23) {real, imag} */,
  {32'h3d988820, 32'hbcb2472a} /* (26, 16, 22) {real, imag} */,
  {32'h3db289e6, 32'h3dd5ab21} /* (26, 16, 21) {real, imag} */,
  {32'hbd71a44a, 32'hbd22561c} /* (26, 16, 20) {real, imag} */,
  {32'h3b19faf8, 32'hbc107d02} /* (26, 16, 19) {real, imag} */,
  {32'h3d4e9afd, 32'h3db64ef2} /* (26, 16, 18) {real, imag} */,
  {32'hbc9b73da, 32'hbcc0b847} /* (26, 16, 17) {real, imag} */,
  {32'h3dbc5798, 32'h00000000} /* (26, 16, 16) {real, imag} */,
  {32'hbc9b73da, 32'h3cc0b847} /* (26, 16, 15) {real, imag} */,
  {32'h3d4e9afd, 32'hbdb64ef2} /* (26, 16, 14) {real, imag} */,
  {32'h3b19faf8, 32'h3c107d02} /* (26, 16, 13) {real, imag} */,
  {32'hbd71a44a, 32'h3d22561c} /* (26, 16, 12) {real, imag} */,
  {32'h3db289e6, 32'hbdd5ab21} /* (26, 16, 11) {real, imag} */,
  {32'h3d988820, 32'h3cb2472a} /* (26, 16, 10) {real, imag} */,
  {32'h3c41b806, 32'hbb836bb0} /* (26, 16, 9) {real, imag} */,
  {32'h3cd0ae6e, 32'h3c12b786} /* (26, 16, 8) {real, imag} */,
  {32'h3c97ab59, 32'hbdc15680} /* (26, 16, 7) {real, imag} */,
  {32'h3c0db194, 32'hbd8047bb} /* (26, 16, 6) {real, imag} */,
  {32'h3d3570c9, 32'h3d8aee3a} /* (26, 16, 5) {real, imag} */,
  {32'h3cc5a3b4, 32'h3d0f5bba} /* (26, 16, 4) {real, imag} */,
  {32'hbd2cf7f8, 32'h3e00fcbc} /* (26, 16, 3) {real, imag} */,
  {32'hbbad04b0, 32'h3d756e20} /* (26, 16, 2) {real, imag} */,
  {32'h3e1d8860, 32'hbe4c6e82} /* (26, 16, 1) {real, imag} */,
  {32'h3e2db864, 32'h00000000} /* (26, 16, 0) {real, imag} */,
  {32'h3e53c446, 32'h3e0cc49c} /* (26, 15, 31) {real, imag} */,
  {32'hbd4c3d65, 32'hbdc73f7e} /* (26, 15, 30) {real, imag} */,
  {32'h3c365950, 32'h3db9d4d7} /* (26, 15, 29) {real, imag} */,
  {32'h3c0fa278, 32'hbd44bf12} /* (26, 15, 28) {real, imag} */,
  {32'h3d8c0e8a, 32'hbbeac1a4} /* (26, 15, 27) {real, imag} */,
  {32'h3da92063, 32'h3d29ca95} /* (26, 15, 26) {real, imag} */,
  {32'h3d70e0d2, 32'h3e013370} /* (26, 15, 25) {real, imag} */,
  {32'h3e241da9, 32'hbda0871b} /* (26, 15, 24) {real, imag} */,
  {32'hbdbba6b4, 32'hbd8721fc} /* (26, 15, 23) {real, imag} */,
  {32'hbd05615f, 32'hbcec79f4} /* (26, 15, 22) {real, imag} */,
  {32'h3ca4772e, 32'h3d8644a9} /* (26, 15, 21) {real, imag} */,
  {32'hbc889228, 32'hbd4d0a1a} /* (26, 15, 20) {real, imag} */,
  {32'hbe301e23, 32'h3d589dc2} /* (26, 15, 19) {real, imag} */,
  {32'h3c581fc0, 32'h3d297097} /* (26, 15, 18) {real, imag} */,
  {32'h3cb296cb, 32'h3d20d368} /* (26, 15, 17) {real, imag} */,
  {32'h3db44be2, 32'h00000000} /* (26, 15, 16) {real, imag} */,
  {32'h3cb296cb, 32'hbd20d368} /* (26, 15, 15) {real, imag} */,
  {32'h3c581fc0, 32'hbd297097} /* (26, 15, 14) {real, imag} */,
  {32'hbe301e23, 32'hbd589dc2} /* (26, 15, 13) {real, imag} */,
  {32'hbc889228, 32'h3d4d0a1a} /* (26, 15, 12) {real, imag} */,
  {32'h3ca4772e, 32'hbd8644a9} /* (26, 15, 11) {real, imag} */,
  {32'hbd05615f, 32'h3cec79f4} /* (26, 15, 10) {real, imag} */,
  {32'hbdbba6b4, 32'h3d8721fc} /* (26, 15, 9) {real, imag} */,
  {32'h3e241da9, 32'h3da0871b} /* (26, 15, 8) {real, imag} */,
  {32'h3d70e0d2, 32'hbe013370} /* (26, 15, 7) {real, imag} */,
  {32'h3da92063, 32'hbd29ca95} /* (26, 15, 6) {real, imag} */,
  {32'h3d8c0e8a, 32'h3beac1a4} /* (26, 15, 5) {real, imag} */,
  {32'h3c0fa278, 32'h3d44bf12} /* (26, 15, 4) {real, imag} */,
  {32'h3c365950, 32'hbdb9d4d7} /* (26, 15, 3) {real, imag} */,
  {32'hbd4c3d65, 32'h3dc73f7e} /* (26, 15, 2) {real, imag} */,
  {32'h3e53c446, 32'hbe0cc49c} /* (26, 15, 1) {real, imag} */,
  {32'hbe937288, 32'h00000000} /* (26, 15, 0) {real, imag} */,
  {32'h3e3e7d7b, 32'h3e673954} /* (26, 14, 31) {real, imag} */,
  {32'h3d68618e, 32'h3d929219} /* (26, 14, 30) {real, imag} */,
  {32'hbcc60bad, 32'h3b7b0fa0} /* (26, 14, 29) {real, imag} */,
  {32'hbcca1f8a, 32'h3cc97e1a} /* (26, 14, 28) {real, imag} */,
  {32'h3d5b351b, 32'hbc01c81c} /* (26, 14, 27) {real, imag} */,
  {32'hbb8988d0, 32'hbcb77048} /* (26, 14, 26) {real, imag} */,
  {32'h3d0e8450, 32'h3aef9100} /* (26, 14, 25) {real, imag} */,
  {32'h3da669c6, 32'hbe0271f0} /* (26, 14, 24) {real, imag} */,
  {32'h3d12424c, 32'hbc0afd2d} /* (26, 14, 23) {real, imag} */,
  {32'h3cd0d074, 32'h3d7e9b82} /* (26, 14, 22) {real, imag} */,
  {32'h3d32c91d, 32'h3d28a945} /* (26, 14, 21) {real, imag} */,
  {32'h3b81a59c, 32'h3bf094d4} /* (26, 14, 20) {real, imag} */,
  {32'hbd9587fc, 32'hbc3ef39a} /* (26, 14, 19) {real, imag} */,
  {32'hbd93b698, 32'h3d450170} /* (26, 14, 18) {real, imag} */,
  {32'hbba05a71, 32'h3d204b1a} /* (26, 14, 17) {real, imag} */,
  {32'h3c7dc03f, 32'h00000000} /* (26, 14, 16) {real, imag} */,
  {32'hbba05a71, 32'hbd204b1a} /* (26, 14, 15) {real, imag} */,
  {32'hbd93b698, 32'hbd450170} /* (26, 14, 14) {real, imag} */,
  {32'hbd9587fc, 32'h3c3ef39a} /* (26, 14, 13) {real, imag} */,
  {32'h3b81a59c, 32'hbbf094d4} /* (26, 14, 12) {real, imag} */,
  {32'h3d32c91d, 32'hbd28a945} /* (26, 14, 11) {real, imag} */,
  {32'h3cd0d074, 32'hbd7e9b82} /* (26, 14, 10) {real, imag} */,
  {32'h3d12424c, 32'h3c0afd2d} /* (26, 14, 9) {real, imag} */,
  {32'h3da669c6, 32'h3e0271f0} /* (26, 14, 8) {real, imag} */,
  {32'h3d0e8450, 32'hbaef9100} /* (26, 14, 7) {real, imag} */,
  {32'hbb8988d0, 32'h3cb77048} /* (26, 14, 6) {real, imag} */,
  {32'h3d5b351b, 32'h3c01c81c} /* (26, 14, 5) {real, imag} */,
  {32'hbcca1f8a, 32'hbcc97e1a} /* (26, 14, 4) {real, imag} */,
  {32'hbcc60bad, 32'hbb7b0fa0} /* (26, 14, 3) {real, imag} */,
  {32'h3d68618e, 32'hbd929219} /* (26, 14, 2) {real, imag} */,
  {32'h3e3e7d7b, 32'hbe673954} /* (26, 14, 1) {real, imag} */,
  {32'hbea19fc0, 32'h00000000} /* (26, 14, 0) {real, imag} */,
  {32'h3e5df242, 32'h3e423cd0} /* (26, 13, 31) {real, imag} */,
  {32'hbd20cd76, 32'h3d00f428} /* (26, 13, 30) {real, imag} */,
  {32'hbc6bb8b2, 32'hbd850a23} /* (26, 13, 29) {real, imag} */,
  {32'hbde948de, 32'h3e0f5740} /* (26, 13, 28) {real, imag} */,
  {32'h3cc0d37e, 32'hbdcd44fa} /* (26, 13, 27) {real, imag} */,
  {32'h3d1c167c, 32'hbcff7172} /* (26, 13, 26) {real, imag} */,
  {32'h3e0d7a31, 32'hbd95c476} /* (26, 13, 25) {real, imag} */,
  {32'h3d3383b5, 32'hbd5c180c} /* (26, 13, 24) {real, imag} */,
  {32'hbd20b768, 32'hbbab0d7c} /* (26, 13, 23) {real, imag} */,
  {32'hbcd90aea, 32'h3c759550} /* (26, 13, 22) {real, imag} */,
  {32'h3d4e3c2a, 32'h3c23e2df} /* (26, 13, 21) {real, imag} */,
  {32'hbcbb6e3c, 32'hbb0aed24} /* (26, 13, 20) {real, imag} */,
  {32'h3ca1703e, 32'h3d819a84} /* (26, 13, 19) {real, imag} */,
  {32'h3d1ac416, 32'hbd6bea44} /* (26, 13, 18) {real, imag} */,
  {32'hbd185eb2, 32'hbcd1228b} /* (26, 13, 17) {real, imag} */,
  {32'hbc6fcb26, 32'h00000000} /* (26, 13, 16) {real, imag} */,
  {32'hbd185eb2, 32'h3cd1228b} /* (26, 13, 15) {real, imag} */,
  {32'h3d1ac416, 32'h3d6bea44} /* (26, 13, 14) {real, imag} */,
  {32'h3ca1703e, 32'hbd819a84} /* (26, 13, 13) {real, imag} */,
  {32'hbcbb6e3c, 32'h3b0aed24} /* (26, 13, 12) {real, imag} */,
  {32'h3d4e3c2a, 32'hbc23e2df} /* (26, 13, 11) {real, imag} */,
  {32'hbcd90aea, 32'hbc759550} /* (26, 13, 10) {real, imag} */,
  {32'hbd20b768, 32'h3bab0d7c} /* (26, 13, 9) {real, imag} */,
  {32'h3d3383b5, 32'h3d5c180c} /* (26, 13, 8) {real, imag} */,
  {32'h3e0d7a31, 32'h3d95c476} /* (26, 13, 7) {real, imag} */,
  {32'h3d1c167c, 32'h3cff7172} /* (26, 13, 6) {real, imag} */,
  {32'h3cc0d37e, 32'h3dcd44fa} /* (26, 13, 5) {real, imag} */,
  {32'hbde948de, 32'hbe0f5740} /* (26, 13, 4) {real, imag} */,
  {32'hbc6bb8b2, 32'h3d850a23} /* (26, 13, 3) {real, imag} */,
  {32'hbd20cd76, 32'hbd00f428} /* (26, 13, 2) {real, imag} */,
  {32'h3e5df242, 32'hbe423cd0} /* (26, 13, 1) {real, imag} */,
  {32'hbe841026, 32'h00000000} /* (26, 13, 0) {real, imag} */,
  {32'h3dbb3e40, 32'h3d8ac1dc} /* (26, 12, 31) {real, imag} */,
  {32'hbd76f2ee, 32'hbd88646e} /* (26, 12, 30) {real, imag} */,
  {32'h3cab3bc2, 32'hbd72378c} /* (26, 12, 29) {real, imag} */,
  {32'hbc907da0, 32'hbd362d4e} /* (26, 12, 28) {real, imag} */,
  {32'hbd3cb4e8, 32'hbd907989} /* (26, 12, 27) {real, imag} */,
  {32'h3d801018, 32'h3bba9e78} /* (26, 12, 26) {real, imag} */,
  {32'h3d9c174c, 32'hbc5bc4d0} /* (26, 12, 25) {real, imag} */,
  {32'hbc650664, 32'hbac397f0} /* (26, 12, 24) {real, imag} */,
  {32'h3cc7ba08, 32'hbd1a1114} /* (26, 12, 23) {real, imag} */,
  {32'h3cec9caf, 32'h3b72c930} /* (26, 12, 22) {real, imag} */,
  {32'h3d58b178, 32'h3bf6b3f2} /* (26, 12, 21) {real, imag} */,
  {32'h3c2b7a62, 32'hbd7c283b} /* (26, 12, 20) {real, imag} */,
  {32'hbc73fa38, 32'hbcab5eea} /* (26, 12, 19) {real, imag} */,
  {32'h3d49e820, 32'hbd191a68} /* (26, 12, 18) {real, imag} */,
  {32'h3dc9f08d, 32'h3d2aa97e} /* (26, 12, 17) {real, imag} */,
  {32'h3d4a5922, 32'h00000000} /* (26, 12, 16) {real, imag} */,
  {32'h3dc9f08d, 32'hbd2aa97e} /* (26, 12, 15) {real, imag} */,
  {32'h3d49e820, 32'h3d191a68} /* (26, 12, 14) {real, imag} */,
  {32'hbc73fa38, 32'h3cab5eea} /* (26, 12, 13) {real, imag} */,
  {32'h3c2b7a62, 32'h3d7c283b} /* (26, 12, 12) {real, imag} */,
  {32'h3d58b178, 32'hbbf6b3f2} /* (26, 12, 11) {real, imag} */,
  {32'h3cec9caf, 32'hbb72c930} /* (26, 12, 10) {real, imag} */,
  {32'h3cc7ba08, 32'h3d1a1114} /* (26, 12, 9) {real, imag} */,
  {32'hbc650664, 32'h3ac397f0} /* (26, 12, 8) {real, imag} */,
  {32'h3d9c174c, 32'h3c5bc4d0} /* (26, 12, 7) {real, imag} */,
  {32'h3d801018, 32'hbbba9e78} /* (26, 12, 6) {real, imag} */,
  {32'hbd3cb4e8, 32'h3d907989} /* (26, 12, 5) {real, imag} */,
  {32'hbc907da0, 32'h3d362d4e} /* (26, 12, 4) {real, imag} */,
  {32'h3cab3bc2, 32'h3d72378c} /* (26, 12, 3) {real, imag} */,
  {32'hbd76f2ee, 32'h3d88646e} /* (26, 12, 2) {real, imag} */,
  {32'h3dbb3e40, 32'hbd8ac1dc} /* (26, 12, 1) {real, imag} */,
  {32'hbe6eb1cc, 32'h00000000} /* (26, 12, 0) {real, imag} */,
  {32'hbcc46b68, 32'h3e1649e6} /* (26, 11, 31) {real, imag} */,
  {32'hbe2f3e3d, 32'h3d8871c9} /* (26, 11, 30) {real, imag} */,
  {32'h3d80b844, 32'hbe01211d} /* (26, 11, 29) {real, imag} */,
  {32'h3e12fbd2, 32'hbe0139eb} /* (26, 11, 28) {real, imag} */,
  {32'hbd989d60, 32'hbcce86a9} /* (26, 11, 27) {real, imag} */,
  {32'h3d4ede01, 32'hbd02740e} /* (26, 11, 26) {real, imag} */,
  {32'hbd28a45b, 32'hbd9c3249} /* (26, 11, 25) {real, imag} */,
  {32'h3d33cd4a, 32'hbce5e19e} /* (26, 11, 24) {real, imag} */,
  {32'h3c4623f6, 32'hbcc94223} /* (26, 11, 23) {real, imag} */,
  {32'hbddef404, 32'h3d80b214} /* (26, 11, 22) {real, imag} */,
  {32'hbcb34f22, 32'h3d95244c} /* (26, 11, 21) {real, imag} */,
  {32'hbda2495a, 32'hbc2ff948} /* (26, 11, 20) {real, imag} */,
  {32'h3d8435de, 32'hbd5d9cc4} /* (26, 11, 19) {real, imag} */,
  {32'hbcd06c5c, 32'hbd386107} /* (26, 11, 18) {real, imag} */,
  {32'h3c33e401, 32'hbca95bd6} /* (26, 11, 17) {real, imag} */,
  {32'h3d054d00, 32'h00000000} /* (26, 11, 16) {real, imag} */,
  {32'h3c33e401, 32'h3ca95bd6} /* (26, 11, 15) {real, imag} */,
  {32'hbcd06c5c, 32'h3d386107} /* (26, 11, 14) {real, imag} */,
  {32'h3d8435de, 32'h3d5d9cc4} /* (26, 11, 13) {real, imag} */,
  {32'hbda2495a, 32'h3c2ff948} /* (26, 11, 12) {real, imag} */,
  {32'hbcb34f22, 32'hbd95244c} /* (26, 11, 11) {real, imag} */,
  {32'hbddef404, 32'hbd80b214} /* (26, 11, 10) {real, imag} */,
  {32'h3c4623f6, 32'h3cc94223} /* (26, 11, 9) {real, imag} */,
  {32'h3d33cd4a, 32'h3ce5e19e} /* (26, 11, 8) {real, imag} */,
  {32'hbd28a45b, 32'h3d9c3249} /* (26, 11, 7) {real, imag} */,
  {32'h3d4ede01, 32'h3d02740e} /* (26, 11, 6) {real, imag} */,
  {32'hbd989d60, 32'h3cce86a9} /* (26, 11, 5) {real, imag} */,
  {32'h3e12fbd2, 32'h3e0139eb} /* (26, 11, 4) {real, imag} */,
  {32'h3d80b844, 32'h3e01211d} /* (26, 11, 3) {real, imag} */,
  {32'hbe2f3e3d, 32'hbd8871c9} /* (26, 11, 2) {real, imag} */,
  {32'hbcc46b68, 32'hbe1649e6} /* (26, 11, 1) {real, imag} */,
  {32'hbd4ec1cc, 32'h00000000} /* (26, 11, 0) {real, imag} */,
  {32'h3dbdbf90, 32'h3e8c0e45} /* (26, 10, 31) {real, imag} */,
  {32'hbe1fbbda, 32'h3dc5ee18} /* (26, 10, 30) {real, imag} */,
  {32'h3cb66cfc, 32'hbd87ac5e} /* (26, 10, 29) {real, imag} */,
  {32'h3e1c7470, 32'hbdd3b99b} /* (26, 10, 28) {real, imag} */,
  {32'h3d524044, 32'h3c23647e} /* (26, 10, 27) {real, imag} */,
  {32'h3d976c56, 32'hbd151b94} /* (26, 10, 26) {real, imag} */,
  {32'h3b0f5480, 32'h3d3af489} /* (26, 10, 25) {real, imag} */,
  {32'h3dcdfc1b, 32'hbd04e488} /* (26, 10, 24) {real, imag} */,
  {32'hbe11752a, 32'h3d42a608} /* (26, 10, 23) {real, imag} */,
  {32'h3d9cf8c2, 32'h3dd826d3} /* (26, 10, 22) {real, imag} */,
  {32'hbc9d05e4, 32'h3dd7832b} /* (26, 10, 21) {real, imag} */,
  {32'hbd3275f2, 32'h3d033994} /* (26, 10, 20) {real, imag} */,
  {32'h3cb04d7b, 32'h3dcc358f} /* (26, 10, 19) {real, imag} */,
  {32'h3d51c4ac, 32'hbd791c1c} /* (26, 10, 18) {real, imag} */,
  {32'h3b5616c0, 32'h3cc49fd4} /* (26, 10, 17) {real, imag} */,
  {32'h3d9e4a2b, 32'h00000000} /* (26, 10, 16) {real, imag} */,
  {32'h3b5616c0, 32'hbcc49fd4} /* (26, 10, 15) {real, imag} */,
  {32'h3d51c4ac, 32'h3d791c1c} /* (26, 10, 14) {real, imag} */,
  {32'h3cb04d7b, 32'hbdcc358f} /* (26, 10, 13) {real, imag} */,
  {32'hbd3275f2, 32'hbd033994} /* (26, 10, 12) {real, imag} */,
  {32'hbc9d05e4, 32'hbdd7832b} /* (26, 10, 11) {real, imag} */,
  {32'h3d9cf8c2, 32'hbdd826d3} /* (26, 10, 10) {real, imag} */,
  {32'hbe11752a, 32'hbd42a608} /* (26, 10, 9) {real, imag} */,
  {32'h3dcdfc1b, 32'h3d04e488} /* (26, 10, 8) {real, imag} */,
  {32'h3b0f5480, 32'hbd3af489} /* (26, 10, 7) {real, imag} */,
  {32'h3d976c56, 32'h3d151b94} /* (26, 10, 6) {real, imag} */,
  {32'h3d524044, 32'hbc23647e} /* (26, 10, 5) {real, imag} */,
  {32'h3e1c7470, 32'h3dd3b99b} /* (26, 10, 4) {real, imag} */,
  {32'h3cb66cfc, 32'h3d87ac5e} /* (26, 10, 3) {real, imag} */,
  {32'hbe1fbbda, 32'hbdc5ee18} /* (26, 10, 2) {real, imag} */,
  {32'h3dbdbf90, 32'hbe8c0e45} /* (26, 10, 1) {real, imag} */,
  {32'hbe670cb1, 32'h00000000} /* (26, 10, 0) {real, imag} */,
  {32'h3d00fae0, 32'h3eaaa79f} /* (26, 9, 31) {real, imag} */,
  {32'hbe49e8c3, 32'h3de3576b} /* (26, 9, 30) {real, imag} */,
  {32'h3d3f8efe, 32'hbdbc90ac} /* (26, 9, 29) {real, imag} */,
  {32'h3dc252f7, 32'hbd8ba487} /* (26, 9, 28) {real, imag} */,
  {32'hbb11dd30, 32'hb72a8000} /* (26, 9, 27) {real, imag} */,
  {32'h3a9e7b30, 32'hbd562399} /* (26, 9, 26) {real, imag} */,
  {32'hbdaf6dce, 32'h3d3f39a8} /* (26, 9, 25) {real, imag} */,
  {32'h3b7c5d10, 32'h3c8fd734} /* (26, 9, 24) {real, imag} */,
  {32'hbbce7b4e, 32'hbc297a02} /* (26, 9, 23) {real, imag} */,
  {32'hbd71d9ec, 32'h3d9c8ee4} /* (26, 9, 22) {real, imag} */,
  {32'h3c7dda74, 32'h3c0bafee} /* (26, 9, 21) {real, imag} */,
  {32'h3ca3291c, 32'h3ce47381} /* (26, 9, 20) {real, imag} */,
  {32'hbdc5f8df, 32'hbd566494} /* (26, 9, 19) {real, imag} */,
  {32'hbd7c634a, 32'h3bb43064} /* (26, 9, 18) {real, imag} */,
  {32'h3b201c38, 32'h3c9480fc} /* (26, 9, 17) {real, imag} */,
  {32'h3dc00884, 32'h00000000} /* (26, 9, 16) {real, imag} */,
  {32'h3b201c38, 32'hbc9480fc} /* (26, 9, 15) {real, imag} */,
  {32'hbd7c634a, 32'hbbb43064} /* (26, 9, 14) {real, imag} */,
  {32'hbdc5f8df, 32'h3d566494} /* (26, 9, 13) {real, imag} */,
  {32'h3ca3291c, 32'hbce47381} /* (26, 9, 12) {real, imag} */,
  {32'h3c7dda74, 32'hbc0bafee} /* (26, 9, 11) {real, imag} */,
  {32'hbd71d9ec, 32'hbd9c8ee4} /* (26, 9, 10) {real, imag} */,
  {32'hbbce7b4e, 32'h3c297a02} /* (26, 9, 9) {real, imag} */,
  {32'h3b7c5d10, 32'hbc8fd734} /* (26, 9, 8) {real, imag} */,
  {32'hbdaf6dce, 32'hbd3f39a8} /* (26, 9, 7) {real, imag} */,
  {32'h3a9e7b30, 32'h3d562399} /* (26, 9, 6) {real, imag} */,
  {32'hbb11dd30, 32'h372a8000} /* (26, 9, 5) {real, imag} */,
  {32'h3dc252f7, 32'h3d8ba487} /* (26, 9, 4) {real, imag} */,
  {32'h3d3f8efe, 32'h3dbc90ac} /* (26, 9, 3) {real, imag} */,
  {32'hbe49e8c3, 32'hbde3576b} /* (26, 9, 2) {real, imag} */,
  {32'h3d00fae0, 32'hbeaaa79f} /* (26, 9, 1) {real, imag} */,
  {32'hbf01093c, 32'h00000000} /* (26, 9, 0) {real, imag} */,
  {32'hbdabcfac, 32'h3f01c748} /* (26, 8, 31) {real, imag} */,
  {32'hbe76ee8d, 32'h3e311949} /* (26, 8, 30) {real, imag} */,
  {32'h3d50c221, 32'hbdcf261e} /* (26, 8, 29) {real, imag} */,
  {32'h3d85aa46, 32'hbd5e7933} /* (26, 8, 28) {real, imag} */,
  {32'hbd4a18b4, 32'h3d124384} /* (26, 8, 27) {real, imag} */,
  {32'hbc83bebc, 32'hbceaa482} /* (26, 8, 26) {real, imag} */,
  {32'h3c15a348, 32'hbd0d4e0e} /* (26, 8, 25) {real, imag} */,
  {32'hbc77f294, 32'hbcc68e6d} /* (26, 8, 24) {real, imag} */,
  {32'hbda91809, 32'hbd26cc8f} /* (26, 8, 23) {real, imag} */,
  {32'hbc9d0264, 32'h3b9cf89c} /* (26, 8, 22) {real, imag} */,
  {32'hbd89ca2c, 32'h3d071e20} /* (26, 8, 21) {real, imag} */,
  {32'hbda7c8da, 32'h3d25c3d2} /* (26, 8, 20) {real, imag} */,
  {32'hbd606a28, 32'hbc30add0} /* (26, 8, 19) {real, imag} */,
  {32'hbccfcf28, 32'hbcade184} /* (26, 8, 18) {real, imag} */,
  {32'h3c2e0a4e, 32'hbc420798} /* (26, 8, 17) {real, imag} */,
  {32'hbc7df8df, 32'h00000000} /* (26, 8, 16) {real, imag} */,
  {32'h3c2e0a4e, 32'h3c420798} /* (26, 8, 15) {real, imag} */,
  {32'hbccfcf28, 32'h3cade184} /* (26, 8, 14) {real, imag} */,
  {32'hbd606a28, 32'h3c30add0} /* (26, 8, 13) {real, imag} */,
  {32'hbda7c8da, 32'hbd25c3d2} /* (26, 8, 12) {real, imag} */,
  {32'hbd89ca2c, 32'hbd071e20} /* (26, 8, 11) {real, imag} */,
  {32'hbc9d0264, 32'hbb9cf89c} /* (26, 8, 10) {real, imag} */,
  {32'hbda91809, 32'h3d26cc8f} /* (26, 8, 9) {real, imag} */,
  {32'hbc77f294, 32'h3cc68e6d} /* (26, 8, 8) {real, imag} */,
  {32'h3c15a348, 32'h3d0d4e0e} /* (26, 8, 7) {real, imag} */,
  {32'hbc83bebc, 32'h3ceaa482} /* (26, 8, 6) {real, imag} */,
  {32'hbd4a18b4, 32'hbd124384} /* (26, 8, 5) {real, imag} */,
  {32'h3d85aa46, 32'h3d5e7933} /* (26, 8, 4) {real, imag} */,
  {32'h3d50c221, 32'h3dcf261e} /* (26, 8, 3) {real, imag} */,
  {32'hbe76ee8d, 32'hbe311949} /* (26, 8, 2) {real, imag} */,
  {32'hbdabcfac, 32'hbf01c748} /* (26, 8, 1) {real, imag} */,
  {32'hbf6d2ab8, 32'h00000000} /* (26, 8, 0) {real, imag} */,
  {32'hbea98776, 32'h3f09d31e} /* (26, 7, 31) {real, imag} */,
  {32'hbe659f94, 32'h3e6dae10} /* (26, 7, 30) {real, imag} */,
  {32'h3dc7dbf1, 32'h3d9a1000} /* (26, 7, 29) {real, imag} */,
  {32'h3d96c414, 32'hbda13ae3} /* (26, 7, 28) {real, imag} */,
  {32'h3d125725, 32'h3c4647f8} /* (26, 7, 27) {real, imag} */,
  {32'hbc62c206, 32'hbddca0a4} /* (26, 7, 26) {real, imag} */,
  {32'h3dcd3855, 32'hbd58c8be} /* (26, 7, 25) {real, imag} */,
  {32'hbd8cefa4, 32'hbd54e7e2} /* (26, 7, 24) {real, imag} */,
  {32'hbda0b5e8, 32'h3d31f6dc} /* (26, 7, 23) {real, imag} */,
  {32'h3d9c3afb, 32'h3d9a982c} /* (26, 7, 22) {real, imag} */,
  {32'h3d37cc69, 32'h3ddb8bac} /* (26, 7, 21) {real, imag} */,
  {32'hbd5ebb7a, 32'h3d4fa38a} /* (26, 7, 20) {real, imag} */,
  {32'h3ce4621f, 32'hbc57fad6} /* (26, 7, 19) {real, imag} */,
  {32'h3c0a9bb0, 32'h3d185c72} /* (26, 7, 18) {real, imag} */,
  {32'h3ccb362c, 32'hbc44d8fc} /* (26, 7, 17) {real, imag} */,
  {32'h3d4b656e, 32'h00000000} /* (26, 7, 16) {real, imag} */,
  {32'h3ccb362c, 32'h3c44d8fc} /* (26, 7, 15) {real, imag} */,
  {32'h3c0a9bb0, 32'hbd185c72} /* (26, 7, 14) {real, imag} */,
  {32'h3ce4621f, 32'h3c57fad6} /* (26, 7, 13) {real, imag} */,
  {32'hbd5ebb7a, 32'hbd4fa38a} /* (26, 7, 12) {real, imag} */,
  {32'h3d37cc69, 32'hbddb8bac} /* (26, 7, 11) {real, imag} */,
  {32'h3d9c3afb, 32'hbd9a982c} /* (26, 7, 10) {real, imag} */,
  {32'hbda0b5e8, 32'hbd31f6dc} /* (26, 7, 9) {real, imag} */,
  {32'hbd8cefa4, 32'h3d54e7e2} /* (26, 7, 8) {real, imag} */,
  {32'h3dcd3855, 32'h3d58c8be} /* (26, 7, 7) {real, imag} */,
  {32'hbc62c206, 32'h3ddca0a4} /* (26, 7, 6) {real, imag} */,
  {32'h3d125725, 32'hbc4647f8} /* (26, 7, 5) {real, imag} */,
  {32'h3d96c414, 32'h3da13ae3} /* (26, 7, 4) {real, imag} */,
  {32'h3dc7dbf1, 32'hbd9a1000} /* (26, 7, 3) {real, imag} */,
  {32'hbe659f94, 32'hbe6dae10} /* (26, 7, 2) {real, imag} */,
  {32'hbea98776, 32'hbf09d31e} /* (26, 7, 1) {real, imag} */,
  {32'hbf8fb8a1, 32'h00000000} /* (26, 7, 0) {real, imag} */,
  {32'hbf06fcf4, 32'h3efe8648} /* (26, 6, 31) {real, imag} */,
  {32'hbe844aa0, 32'h3ddce53d} /* (26, 6, 30) {real, imag} */,
  {32'h3d714b32, 32'h3cc19379} /* (26, 6, 29) {real, imag} */,
  {32'h3d923531, 32'h3c5bd124} /* (26, 6, 28) {real, imag} */,
  {32'hbc7984c6, 32'h3d883e57} /* (26, 6, 27) {real, imag} */,
  {32'h3c7556cf, 32'hbde105b3} /* (26, 6, 26) {real, imag} */,
  {32'h3c873b1b, 32'hbda2b844} /* (26, 6, 25) {real, imag} */,
  {32'hbd1cd946, 32'h3c3c0b24} /* (26, 6, 24) {real, imag} */,
  {32'h3d5547aa, 32'h3dd271eb} /* (26, 6, 23) {real, imag} */,
  {32'h3c2ac11a, 32'hbd4eeece} /* (26, 6, 22) {real, imag} */,
  {32'hbbab72a0, 32'hbc91578f} /* (26, 6, 21) {real, imag} */,
  {32'hbcd51457, 32'hbda8ecec} /* (26, 6, 20) {real, imag} */,
  {32'h3ca9e4c3, 32'hbcf9ea04} /* (26, 6, 19) {real, imag} */,
  {32'h3d049486, 32'hbbbacf74} /* (26, 6, 18) {real, imag} */,
  {32'hbd1c7ca9, 32'hbdfe7215} /* (26, 6, 17) {real, imag} */,
  {32'h3cd24927, 32'h00000000} /* (26, 6, 16) {real, imag} */,
  {32'hbd1c7ca9, 32'h3dfe7215} /* (26, 6, 15) {real, imag} */,
  {32'h3d049486, 32'h3bbacf74} /* (26, 6, 14) {real, imag} */,
  {32'h3ca9e4c3, 32'h3cf9ea04} /* (26, 6, 13) {real, imag} */,
  {32'hbcd51457, 32'h3da8ecec} /* (26, 6, 12) {real, imag} */,
  {32'hbbab72a0, 32'h3c91578f} /* (26, 6, 11) {real, imag} */,
  {32'h3c2ac11a, 32'h3d4eeece} /* (26, 6, 10) {real, imag} */,
  {32'h3d5547aa, 32'hbdd271eb} /* (26, 6, 9) {real, imag} */,
  {32'hbd1cd946, 32'hbc3c0b24} /* (26, 6, 8) {real, imag} */,
  {32'h3c873b1b, 32'h3da2b844} /* (26, 6, 7) {real, imag} */,
  {32'h3c7556cf, 32'h3de105b3} /* (26, 6, 6) {real, imag} */,
  {32'hbc7984c6, 32'hbd883e57} /* (26, 6, 5) {real, imag} */,
  {32'h3d923531, 32'hbc5bd124} /* (26, 6, 4) {real, imag} */,
  {32'h3d714b32, 32'hbcc19379} /* (26, 6, 3) {real, imag} */,
  {32'hbe844aa0, 32'hbddce53d} /* (26, 6, 2) {real, imag} */,
  {32'hbf06fcf4, 32'hbefe8648} /* (26, 6, 1) {real, imag} */,
  {32'hbf948b00, 32'h00000000} /* (26, 6, 0) {real, imag} */,
  {32'hbf20634e, 32'h3f02ab2d} /* (26, 5, 31) {real, imag} */,
  {32'hbdf8fb91, 32'h3e136828} /* (26, 5, 30) {real, imag} */,
  {32'h3e0ff71e, 32'hbe088b26} /* (26, 5, 29) {real, imag} */,
  {32'h3d20c722, 32'h3da4ebf1} /* (26, 5, 28) {real, imag} */,
  {32'hbda5037e, 32'h3e2c4082} /* (26, 5, 27) {real, imag} */,
  {32'h3c0258c0, 32'h3c85bc6c} /* (26, 5, 26) {real, imag} */,
  {32'h3d09da75, 32'hbc6cae28} /* (26, 5, 25) {real, imag} */,
  {32'h3dc26dbe, 32'h3dd9d210} /* (26, 5, 24) {real, imag} */,
  {32'h3c52843a, 32'h3c61a4ec} /* (26, 5, 23) {real, imag} */,
  {32'hbca57394, 32'h3d9bae3a} /* (26, 5, 22) {real, imag} */,
  {32'h3d7653f5, 32'h3cc84eba} /* (26, 5, 21) {real, imag} */,
  {32'hbbdc7ed8, 32'h3ceab128} /* (26, 5, 20) {real, imag} */,
  {32'hb93c3000, 32'hbdaa9d3a} /* (26, 5, 19) {real, imag} */,
  {32'hbc833c36, 32'h3e25c61a} /* (26, 5, 18) {real, imag} */,
  {32'hbd0b0263, 32'hbc7b19a8} /* (26, 5, 17) {real, imag} */,
  {32'hbdcb8734, 32'h00000000} /* (26, 5, 16) {real, imag} */,
  {32'hbd0b0263, 32'h3c7b19a8} /* (26, 5, 15) {real, imag} */,
  {32'hbc833c36, 32'hbe25c61a} /* (26, 5, 14) {real, imag} */,
  {32'hb93c3000, 32'h3daa9d3a} /* (26, 5, 13) {real, imag} */,
  {32'hbbdc7ed8, 32'hbceab128} /* (26, 5, 12) {real, imag} */,
  {32'h3d7653f5, 32'hbcc84eba} /* (26, 5, 11) {real, imag} */,
  {32'hbca57394, 32'hbd9bae3a} /* (26, 5, 10) {real, imag} */,
  {32'h3c52843a, 32'hbc61a4ec} /* (26, 5, 9) {real, imag} */,
  {32'h3dc26dbe, 32'hbdd9d210} /* (26, 5, 8) {real, imag} */,
  {32'h3d09da75, 32'h3c6cae28} /* (26, 5, 7) {real, imag} */,
  {32'h3c0258c0, 32'hbc85bc6c} /* (26, 5, 6) {real, imag} */,
  {32'hbda5037e, 32'hbe2c4082} /* (26, 5, 5) {real, imag} */,
  {32'h3d20c722, 32'hbda4ebf1} /* (26, 5, 4) {real, imag} */,
  {32'h3e0ff71e, 32'h3e088b26} /* (26, 5, 3) {real, imag} */,
  {32'hbdf8fb91, 32'hbe136828} /* (26, 5, 2) {real, imag} */,
  {32'hbf20634e, 32'hbf02ab2d} /* (26, 5, 1) {real, imag} */,
  {32'hbfb7875f, 32'h00000000} /* (26, 5, 0) {real, imag} */,
  {32'hbf453b70, 32'h3f28806b} /* (26, 4, 31) {real, imag} */,
  {32'hbd0196be, 32'h3e8460fe} /* (26, 4, 30) {real, imag} */,
  {32'h3d87c1ec, 32'h3d3c265e} /* (26, 4, 29) {real, imag} */,
  {32'hbdabab9c, 32'hbd09e314} /* (26, 4, 28) {real, imag} */,
  {32'hbd1c5d3d, 32'h3d850e7c} /* (26, 4, 27) {real, imag} */,
  {32'h3e0eea84, 32'hbd42b306} /* (26, 4, 26) {real, imag} */,
  {32'hbd9ced9c, 32'hbdb3a374} /* (26, 4, 25) {real, imag} */,
  {32'h3d240274, 32'h3dc33eed} /* (26, 4, 24) {real, imag} */,
  {32'hbac5ace8, 32'h3dd34df6} /* (26, 4, 23) {real, imag} */,
  {32'hbd72724a, 32'h3c73fac0} /* (26, 4, 22) {real, imag} */,
  {32'hbd8df848, 32'h3b322fe5} /* (26, 4, 21) {real, imag} */,
  {32'h3d524acc, 32'hbe254b95} /* (26, 4, 20) {real, imag} */,
  {32'h3ca505f0, 32'h3cc12d52} /* (26, 4, 19) {real, imag} */,
  {32'h3bc3e42c, 32'hbc29f3d4} /* (26, 4, 18) {real, imag} */,
  {32'h3d2f7a91, 32'h3c37d8f6} /* (26, 4, 17) {real, imag} */,
  {32'hbc4b6144, 32'h00000000} /* (26, 4, 16) {real, imag} */,
  {32'h3d2f7a91, 32'hbc37d8f6} /* (26, 4, 15) {real, imag} */,
  {32'h3bc3e42c, 32'h3c29f3d4} /* (26, 4, 14) {real, imag} */,
  {32'h3ca505f0, 32'hbcc12d52} /* (26, 4, 13) {real, imag} */,
  {32'h3d524acc, 32'h3e254b95} /* (26, 4, 12) {real, imag} */,
  {32'hbd8df848, 32'hbb322fe5} /* (26, 4, 11) {real, imag} */,
  {32'hbd72724a, 32'hbc73fac0} /* (26, 4, 10) {real, imag} */,
  {32'hbac5ace8, 32'hbdd34df6} /* (26, 4, 9) {real, imag} */,
  {32'h3d240274, 32'hbdc33eed} /* (26, 4, 8) {real, imag} */,
  {32'hbd9ced9c, 32'h3db3a374} /* (26, 4, 7) {real, imag} */,
  {32'h3e0eea84, 32'h3d42b306} /* (26, 4, 6) {real, imag} */,
  {32'hbd1c5d3d, 32'hbd850e7c} /* (26, 4, 5) {real, imag} */,
  {32'hbdabab9c, 32'h3d09e314} /* (26, 4, 4) {real, imag} */,
  {32'h3d87c1ec, 32'hbd3c265e} /* (26, 4, 3) {real, imag} */,
  {32'hbd0196be, 32'hbe8460fe} /* (26, 4, 2) {real, imag} */,
  {32'hbf453b70, 32'hbf28806b} /* (26, 4, 1) {real, imag} */,
  {32'hbfac1a02, 32'h00000000} /* (26, 4, 0) {real, imag} */,
  {32'hbf51b1e5, 32'h3f33b479} /* (26, 3, 31) {real, imag} */,
  {32'h3dcca584, 32'h3e89e80b} /* (26, 3, 30) {real, imag} */,
  {32'hbc48e8c4, 32'hbc2b4b88} /* (26, 3, 29) {real, imag} */,
  {32'hbd40de5f, 32'h3c397ae4} /* (26, 3, 28) {real, imag} */,
  {32'h3c66db30, 32'hbc814e76} /* (26, 3, 27) {real, imag} */,
  {32'h3cd64fee, 32'h3ce23344} /* (26, 3, 26) {real, imag} */,
  {32'hbdf59ab1, 32'hbcdbb31d} /* (26, 3, 25) {real, imag} */,
  {32'hbd9e49ac, 32'hbdccbdf4} /* (26, 3, 24) {real, imag} */,
  {32'h3cd74170, 32'h3e1aa435} /* (26, 3, 23) {real, imag} */,
  {32'hbe039220, 32'hbd662e24} /* (26, 3, 22) {real, imag} */,
  {32'hbddfd85a, 32'hbcdc4d6c} /* (26, 3, 21) {real, imag} */,
  {32'h3c17a788, 32'hbc44a482} /* (26, 3, 20) {real, imag} */,
  {32'h3d45855f, 32'h3d223db2} /* (26, 3, 19) {real, imag} */,
  {32'h3defa126, 32'h3c86b054} /* (26, 3, 18) {real, imag} */,
  {32'h3b9c9650, 32'h3e0c8bea} /* (26, 3, 17) {real, imag} */,
  {32'h3dae06d8, 32'h00000000} /* (26, 3, 16) {real, imag} */,
  {32'h3b9c9650, 32'hbe0c8bea} /* (26, 3, 15) {real, imag} */,
  {32'h3defa126, 32'hbc86b054} /* (26, 3, 14) {real, imag} */,
  {32'h3d45855f, 32'hbd223db2} /* (26, 3, 13) {real, imag} */,
  {32'h3c17a788, 32'h3c44a482} /* (26, 3, 12) {real, imag} */,
  {32'hbddfd85a, 32'h3cdc4d6c} /* (26, 3, 11) {real, imag} */,
  {32'hbe039220, 32'h3d662e24} /* (26, 3, 10) {real, imag} */,
  {32'h3cd74170, 32'hbe1aa435} /* (26, 3, 9) {real, imag} */,
  {32'hbd9e49ac, 32'h3dccbdf4} /* (26, 3, 8) {real, imag} */,
  {32'hbdf59ab1, 32'h3cdbb31d} /* (26, 3, 7) {real, imag} */,
  {32'h3cd64fee, 32'hbce23344} /* (26, 3, 6) {real, imag} */,
  {32'h3c66db30, 32'h3c814e76} /* (26, 3, 5) {real, imag} */,
  {32'hbd40de5f, 32'hbc397ae4} /* (26, 3, 4) {real, imag} */,
  {32'hbc48e8c4, 32'h3c2b4b88} /* (26, 3, 3) {real, imag} */,
  {32'h3dcca584, 32'hbe89e80b} /* (26, 3, 2) {real, imag} */,
  {32'hbf51b1e5, 32'hbf33b479} /* (26, 3, 1) {real, imag} */,
  {32'hbfa6cb3b, 32'h00000000} /* (26, 3, 0) {real, imag} */,
  {32'hbf6b0f8b, 32'h3ef7262d} /* (26, 2, 31) {real, imag} */,
  {32'h3e48914e, 32'h3e44d468} /* (26, 2, 30) {real, imag} */,
  {32'h3ce359d0, 32'hbbd90814} /* (26, 2, 29) {real, imag} */,
  {32'h3e0ba30b, 32'hbac6c5b8} /* (26, 2, 28) {real, imag} */,
  {32'hbd9848bc, 32'hbc9e13f4} /* (26, 2, 27) {real, imag} */,
  {32'hbd80b7a6, 32'hbd4bd1fe} /* (26, 2, 26) {real, imag} */,
  {32'hbdd15d78, 32'hbd008d62} /* (26, 2, 25) {real, imag} */,
  {32'hbd801892, 32'h3c25889c} /* (26, 2, 24) {real, imag} */,
  {32'hbc599ffc, 32'hbdaa6742} /* (26, 2, 23) {real, imag} */,
  {32'hbc434317, 32'h3ced0608} /* (26, 2, 22) {real, imag} */,
  {32'hbba1d950, 32'h3db1237e} /* (26, 2, 21) {real, imag} */,
  {32'hbcd9ade5, 32'h3b2cb040} /* (26, 2, 20) {real, imag} */,
  {32'h3d08cc42, 32'hbd6dec86} /* (26, 2, 19) {real, imag} */,
  {32'h3cb428b6, 32'h3d7b3b94} /* (26, 2, 18) {real, imag} */,
  {32'h3d364a60, 32'h3c52296e} /* (26, 2, 17) {real, imag} */,
  {32'hbcb8ba92, 32'h00000000} /* (26, 2, 16) {real, imag} */,
  {32'h3d364a60, 32'hbc52296e} /* (26, 2, 15) {real, imag} */,
  {32'h3cb428b6, 32'hbd7b3b94} /* (26, 2, 14) {real, imag} */,
  {32'h3d08cc42, 32'h3d6dec86} /* (26, 2, 13) {real, imag} */,
  {32'hbcd9ade5, 32'hbb2cb040} /* (26, 2, 12) {real, imag} */,
  {32'hbba1d950, 32'hbdb1237e} /* (26, 2, 11) {real, imag} */,
  {32'hbc434317, 32'hbced0608} /* (26, 2, 10) {real, imag} */,
  {32'hbc599ffc, 32'h3daa6742} /* (26, 2, 9) {real, imag} */,
  {32'hbd801892, 32'hbc25889c} /* (26, 2, 8) {real, imag} */,
  {32'hbdd15d78, 32'h3d008d62} /* (26, 2, 7) {real, imag} */,
  {32'hbd80b7a6, 32'h3d4bd1fe} /* (26, 2, 6) {real, imag} */,
  {32'hbd9848bc, 32'h3c9e13f4} /* (26, 2, 5) {real, imag} */,
  {32'h3e0ba30b, 32'h3ac6c5b8} /* (26, 2, 4) {real, imag} */,
  {32'h3ce359d0, 32'h3bd90814} /* (26, 2, 3) {real, imag} */,
  {32'h3e48914e, 32'hbe44d468} /* (26, 2, 2) {real, imag} */,
  {32'hbf6b0f8b, 32'hbef7262d} /* (26, 2, 1) {real, imag} */,
  {32'hbfb5f61c, 32'h00000000} /* (26, 2, 0) {real, imag} */,
  {32'hbf6deb28, 32'h3ed6de96} /* (26, 1, 31) {real, imag} */,
  {32'h3de81329, 32'h3e4af277} /* (26, 1, 30) {real, imag} */,
  {32'hbc992480, 32'h3d81191a} /* (26, 1, 29) {real, imag} */,
  {32'h3c4d908a, 32'h3e23eef5} /* (26, 1, 28) {real, imag} */,
  {32'hbd599990, 32'hbdfa2f03} /* (26, 1, 27) {real, imag} */,
  {32'hbd997bfe, 32'hbce4808e} /* (26, 1, 26) {real, imag} */,
  {32'hbdaa9ebf, 32'hbe09fea2} /* (26, 1, 25) {real, imag} */,
  {32'h3e215784, 32'hbcf09c74} /* (26, 1, 24) {real, imag} */,
  {32'hbd31afc7, 32'hbc358602} /* (26, 1, 23) {real, imag} */,
  {32'hbd19a3d0, 32'h3e0c8458} /* (26, 1, 22) {real, imag} */,
  {32'hbd227382, 32'hbd230f88} /* (26, 1, 21) {real, imag} */,
  {32'h3cc5ae84, 32'h3d16be76} /* (26, 1, 20) {real, imag} */,
  {32'h3d47c1d8, 32'hbd5adef9} /* (26, 1, 19) {real, imag} */,
  {32'hbc5dde2a, 32'hbd6d5665} /* (26, 1, 18) {real, imag} */,
  {32'h3cb34e8e, 32'h3d1e6c20} /* (26, 1, 17) {real, imag} */,
  {32'h3c6faf30, 32'h00000000} /* (26, 1, 16) {real, imag} */,
  {32'h3cb34e8e, 32'hbd1e6c20} /* (26, 1, 15) {real, imag} */,
  {32'hbc5dde2a, 32'h3d6d5665} /* (26, 1, 14) {real, imag} */,
  {32'h3d47c1d8, 32'h3d5adef9} /* (26, 1, 13) {real, imag} */,
  {32'h3cc5ae84, 32'hbd16be76} /* (26, 1, 12) {real, imag} */,
  {32'hbd227382, 32'h3d230f88} /* (26, 1, 11) {real, imag} */,
  {32'hbd19a3d0, 32'hbe0c8458} /* (26, 1, 10) {real, imag} */,
  {32'hbd31afc7, 32'h3c358602} /* (26, 1, 9) {real, imag} */,
  {32'h3e215784, 32'h3cf09c74} /* (26, 1, 8) {real, imag} */,
  {32'hbdaa9ebf, 32'h3e09fea2} /* (26, 1, 7) {real, imag} */,
  {32'hbd997bfe, 32'h3ce4808e} /* (26, 1, 6) {real, imag} */,
  {32'hbd599990, 32'h3dfa2f03} /* (26, 1, 5) {real, imag} */,
  {32'h3c4d908a, 32'hbe23eef5} /* (26, 1, 4) {real, imag} */,
  {32'hbc992480, 32'hbd81191a} /* (26, 1, 3) {real, imag} */,
  {32'h3de81329, 32'hbe4af277} /* (26, 1, 2) {real, imag} */,
  {32'hbf6deb28, 32'hbed6de96} /* (26, 1, 1) {real, imag} */,
  {32'hbfcb48ff, 32'h00000000} /* (26, 1, 0) {real, imag} */,
  {32'hbf818b32, 32'h3ec2ade1} /* (26, 0, 31) {real, imag} */,
  {32'h3e1332fc, 32'h3e626c02} /* (26, 0, 30) {real, imag} */,
  {32'h3d4fde4c, 32'hbd857d43} /* (26, 0, 29) {real, imag} */,
  {32'hbd89d1f7, 32'h3db986e7} /* (26, 0, 28) {real, imag} */,
  {32'hba8fc5a0, 32'hbd9e6e62} /* (26, 0, 27) {real, imag} */,
  {32'hbd876c0e, 32'hbd97980d} /* (26, 0, 26) {real, imag} */,
  {32'h3d4d1946, 32'hbd0d00d8} /* (26, 0, 25) {real, imag} */,
  {32'h3d51f71b, 32'h3c58d362} /* (26, 0, 24) {real, imag} */,
  {32'hbcc3f209, 32'h3d59215b} /* (26, 0, 23) {real, imag} */,
  {32'hbd5dd3f8, 32'h3d9a9ae4} /* (26, 0, 22) {real, imag} */,
  {32'h3d865a02, 32'hbdc12f73} /* (26, 0, 21) {real, imag} */,
  {32'hbc78b6da, 32'h3d4b0150} /* (26, 0, 20) {real, imag} */,
  {32'h3cb0a887, 32'h3d4bdd1e} /* (26, 0, 19) {real, imag} */,
  {32'hbc8afd8e, 32'hbcd80ab8} /* (26, 0, 18) {real, imag} */,
  {32'h3cfe97e0, 32'h3c031bea} /* (26, 0, 17) {real, imag} */,
  {32'h3d0b125b, 32'h00000000} /* (26, 0, 16) {real, imag} */,
  {32'h3cfe97e0, 32'hbc031bea} /* (26, 0, 15) {real, imag} */,
  {32'hbc8afd8e, 32'h3cd80ab8} /* (26, 0, 14) {real, imag} */,
  {32'h3cb0a887, 32'hbd4bdd1e} /* (26, 0, 13) {real, imag} */,
  {32'hbc78b6da, 32'hbd4b0150} /* (26, 0, 12) {real, imag} */,
  {32'h3d865a02, 32'h3dc12f73} /* (26, 0, 11) {real, imag} */,
  {32'hbd5dd3f8, 32'hbd9a9ae4} /* (26, 0, 10) {real, imag} */,
  {32'hbcc3f209, 32'hbd59215b} /* (26, 0, 9) {real, imag} */,
  {32'h3d51f71b, 32'hbc58d362} /* (26, 0, 8) {real, imag} */,
  {32'h3d4d1946, 32'h3d0d00d8} /* (26, 0, 7) {real, imag} */,
  {32'hbd876c0e, 32'h3d97980d} /* (26, 0, 6) {real, imag} */,
  {32'hba8fc5a0, 32'h3d9e6e62} /* (26, 0, 5) {real, imag} */,
  {32'hbd89d1f7, 32'hbdb986e7} /* (26, 0, 4) {real, imag} */,
  {32'h3d4fde4c, 32'h3d857d43} /* (26, 0, 3) {real, imag} */,
  {32'h3e1332fc, 32'hbe626c02} /* (26, 0, 2) {real, imag} */,
  {32'hbf818b32, 32'hbec2ade1} /* (26, 0, 1) {real, imag} */,
  {32'hbfdc00a2, 32'h00000000} /* (26, 0, 0) {real, imag} */,
  {32'hc00961c9, 32'h3f8b1db2} /* (25, 31, 31) {real, imag} */,
  {32'h3eb05348, 32'hbda757a0} /* (25, 31, 30) {real, imag} */,
  {32'h3cc54dc8, 32'hbd61b76c} /* (25, 31, 29) {real, imag} */,
  {32'hbdcc5927, 32'h3d20f477} /* (25, 31, 28) {real, imag} */,
  {32'h3df5693e, 32'hbd535b12} /* (25, 31, 27) {real, imag} */,
  {32'hbd3c1afd, 32'hbcee7101} /* (25, 31, 26) {real, imag} */,
  {32'h3cbc4d13, 32'hbd008fc7} /* (25, 31, 25) {real, imag} */,
  {32'hbcb42420, 32'hbd0a042c} /* (25, 31, 24) {real, imag} */,
  {32'hbc40000e, 32'hbd6faca2} /* (25, 31, 23) {real, imag} */,
  {32'h3c900c16, 32'hbd0f15b0} /* (25, 31, 22) {real, imag} */,
  {32'h3ccebb23, 32'hbca33f70} /* (25, 31, 21) {real, imag} */,
  {32'h3d106217, 32'hbd28ffd8} /* (25, 31, 20) {real, imag} */,
  {32'h3c899754, 32'hbc810e68} /* (25, 31, 19) {real, imag} */,
  {32'hbd198a7e, 32'hbd9eab15} /* (25, 31, 18) {real, imag} */,
  {32'h3d35d1ab, 32'hbbfebde1} /* (25, 31, 17) {real, imag} */,
  {32'h3d900102, 32'h00000000} /* (25, 31, 16) {real, imag} */,
  {32'h3d35d1ab, 32'h3bfebde1} /* (25, 31, 15) {real, imag} */,
  {32'hbd198a7e, 32'h3d9eab15} /* (25, 31, 14) {real, imag} */,
  {32'h3c899754, 32'h3c810e68} /* (25, 31, 13) {real, imag} */,
  {32'h3d106217, 32'h3d28ffd8} /* (25, 31, 12) {real, imag} */,
  {32'h3ccebb23, 32'h3ca33f70} /* (25, 31, 11) {real, imag} */,
  {32'h3c900c16, 32'h3d0f15b0} /* (25, 31, 10) {real, imag} */,
  {32'hbc40000e, 32'h3d6faca2} /* (25, 31, 9) {real, imag} */,
  {32'hbcb42420, 32'h3d0a042c} /* (25, 31, 8) {real, imag} */,
  {32'h3cbc4d13, 32'h3d008fc7} /* (25, 31, 7) {real, imag} */,
  {32'hbd3c1afd, 32'h3cee7101} /* (25, 31, 6) {real, imag} */,
  {32'h3df5693e, 32'h3d535b12} /* (25, 31, 5) {real, imag} */,
  {32'hbdcc5927, 32'hbd20f477} /* (25, 31, 4) {real, imag} */,
  {32'h3cc54dc8, 32'h3d61b76c} /* (25, 31, 3) {real, imag} */,
  {32'h3eb05348, 32'h3da757a0} /* (25, 31, 2) {real, imag} */,
  {32'hc00961c9, 32'hbf8b1db2} /* (25, 31, 1) {real, imag} */,
  {32'hc042c599, 32'h00000000} /* (25, 31, 0) {real, imag} */,
  {32'hc01d84de, 32'h3f73df27} /* (25, 30, 31) {real, imag} */,
  {32'h3f2a8dc4, 32'hbdbdb9de} /* (25, 30, 30) {real, imag} */,
  {32'h3c2ec19c, 32'hbd9e42a6} /* (25, 30, 29) {real, imag} */,
  {32'hbe1b58ea, 32'h3d132898} /* (25, 30, 28) {real, imag} */,
  {32'h3db9cd31, 32'h3c9dde35} /* (25, 30, 27) {real, imag} */,
  {32'h3d2ac3b1, 32'hbd6db6d0} /* (25, 30, 26) {real, imag} */,
  {32'hbc887d86, 32'hbd8575be} /* (25, 30, 25) {real, imag} */,
  {32'hbbaa9000, 32'hbd233490} /* (25, 30, 24) {real, imag} */,
  {32'hbd14a523, 32'hbcc27966} /* (25, 30, 23) {real, imag} */,
  {32'hbc35aab0, 32'hbd35ea96} /* (25, 30, 22) {real, imag} */,
  {32'hbd2d3a9b, 32'hbd02a03a} /* (25, 30, 21) {real, imag} */,
  {32'h3cbf991d, 32'hbd074dca} /* (25, 30, 20) {real, imag} */,
  {32'h3d6eac27, 32'h3d6fbabe} /* (25, 30, 19) {real, imag} */,
  {32'h3ccc18cc, 32'hbdf098ec} /* (25, 30, 18) {real, imag} */,
  {32'hbc04d3ca, 32'h3c937209} /* (25, 30, 17) {real, imag} */,
  {32'hbbdb080c, 32'h00000000} /* (25, 30, 16) {real, imag} */,
  {32'hbc04d3ca, 32'hbc937209} /* (25, 30, 15) {real, imag} */,
  {32'h3ccc18cc, 32'h3df098ec} /* (25, 30, 14) {real, imag} */,
  {32'h3d6eac27, 32'hbd6fbabe} /* (25, 30, 13) {real, imag} */,
  {32'h3cbf991d, 32'h3d074dca} /* (25, 30, 12) {real, imag} */,
  {32'hbd2d3a9b, 32'h3d02a03a} /* (25, 30, 11) {real, imag} */,
  {32'hbc35aab0, 32'h3d35ea96} /* (25, 30, 10) {real, imag} */,
  {32'hbd14a523, 32'h3cc27966} /* (25, 30, 9) {real, imag} */,
  {32'hbbaa9000, 32'h3d233490} /* (25, 30, 8) {real, imag} */,
  {32'hbc887d86, 32'h3d8575be} /* (25, 30, 7) {real, imag} */,
  {32'h3d2ac3b1, 32'h3d6db6d0} /* (25, 30, 6) {real, imag} */,
  {32'h3db9cd31, 32'hbc9dde35} /* (25, 30, 5) {real, imag} */,
  {32'hbe1b58ea, 32'hbd132898} /* (25, 30, 4) {real, imag} */,
  {32'h3c2ec19c, 32'h3d9e42a6} /* (25, 30, 3) {real, imag} */,
  {32'h3f2a8dc4, 32'h3dbdb9de} /* (25, 30, 2) {real, imag} */,
  {32'hc01d84de, 32'hbf73df27} /* (25, 30, 1) {real, imag} */,
  {32'hc046139e, 32'h00000000} /* (25, 30, 0) {real, imag} */,
  {32'hc0189312, 32'h3f78aeba} /* (25, 29, 31) {real, imag} */,
  {32'h3f37246a, 32'h3cddd080} /* (25, 29, 30) {real, imag} */,
  {32'h3d0db360, 32'hbd99bbf2} /* (25, 29, 29) {real, imag} */,
  {32'hbe1202fb, 32'hbd2b796e} /* (25, 29, 28) {real, imag} */,
  {32'h3d99ba3a, 32'hbe560870} /* (25, 29, 27) {real, imag} */,
  {32'h3d1907de, 32'hbc6bbe30} /* (25, 29, 26) {real, imag} */,
  {32'h3e23807c, 32'h3dec21fc} /* (25, 29, 25) {real, imag} */,
  {32'h3e0185f6, 32'hbd0f8b82} /* (25, 29, 24) {real, imag} */,
  {32'h3bc90a28, 32'h3cf05e3a} /* (25, 29, 23) {real, imag} */,
  {32'hbc632fc0, 32'h3c319ab6} /* (25, 29, 22) {real, imag} */,
  {32'h3dcf4648, 32'hbdbb9e20} /* (25, 29, 21) {real, imag} */,
  {32'hbdb4e1d3, 32'h3d9336f3} /* (25, 29, 20) {real, imag} */,
  {32'h3c5cde76, 32'h3d166031} /* (25, 29, 19) {real, imag} */,
  {32'h3c89b7ec, 32'hbd945c67} /* (25, 29, 18) {real, imag} */,
  {32'hbb49d898, 32'h3d49428c} /* (25, 29, 17) {real, imag} */,
  {32'h3caaf559, 32'h00000000} /* (25, 29, 16) {real, imag} */,
  {32'hbb49d898, 32'hbd49428c} /* (25, 29, 15) {real, imag} */,
  {32'h3c89b7ec, 32'h3d945c67} /* (25, 29, 14) {real, imag} */,
  {32'h3c5cde76, 32'hbd166031} /* (25, 29, 13) {real, imag} */,
  {32'hbdb4e1d3, 32'hbd9336f3} /* (25, 29, 12) {real, imag} */,
  {32'h3dcf4648, 32'h3dbb9e20} /* (25, 29, 11) {real, imag} */,
  {32'hbc632fc0, 32'hbc319ab6} /* (25, 29, 10) {real, imag} */,
  {32'h3bc90a28, 32'hbcf05e3a} /* (25, 29, 9) {real, imag} */,
  {32'h3e0185f6, 32'h3d0f8b82} /* (25, 29, 8) {real, imag} */,
  {32'h3e23807c, 32'hbdec21fc} /* (25, 29, 7) {real, imag} */,
  {32'h3d1907de, 32'h3c6bbe30} /* (25, 29, 6) {real, imag} */,
  {32'h3d99ba3a, 32'h3e560870} /* (25, 29, 5) {real, imag} */,
  {32'hbe1202fb, 32'h3d2b796e} /* (25, 29, 4) {real, imag} */,
  {32'h3d0db360, 32'h3d99bbf2} /* (25, 29, 3) {real, imag} */,
  {32'h3f37246a, 32'hbcddd080} /* (25, 29, 2) {real, imag} */,
  {32'hc0189312, 32'hbf78aeba} /* (25, 29, 1) {real, imag} */,
  {32'hc052ed26, 32'h00000000} /* (25, 29, 0) {real, imag} */,
  {32'hc0245522, 32'h3f645b0f} /* (25, 28, 31) {real, imag} */,
  {32'h3f3d98c8, 32'hbd4ea7f4} /* (25, 28, 30) {real, imag} */,
  {32'h3c73c2f8, 32'hbe0a01ee} /* (25, 28, 29) {real, imag} */,
  {32'hbdc21e86, 32'h3dd328d6} /* (25, 28, 28) {real, imag} */,
  {32'h3deda673, 32'hbe62e26b} /* (25, 28, 27) {real, imag} */,
  {32'hbd43ce17, 32'h3dd27aac} /* (25, 28, 26) {real, imag} */,
  {32'h3d7ec37d, 32'h382ef100} /* (25, 28, 25) {real, imag} */,
  {32'h3cbae4e5, 32'hbe05f23d} /* (25, 28, 24) {real, imag} */,
  {32'h3d852fa4, 32'hbd0d159e} /* (25, 28, 23) {real, imag} */,
  {32'hbbc50308, 32'hbd8e2308} /* (25, 28, 22) {real, imag} */,
  {32'h3dbe1c9d, 32'hbd6d9291} /* (25, 28, 21) {real, imag} */,
  {32'hbdb7dcce, 32'hbc3ab70e} /* (25, 28, 20) {real, imag} */,
  {32'hbd076798, 32'hbd3d0aff} /* (25, 28, 19) {real, imag} */,
  {32'hbc9faa06, 32'hbdb3c804} /* (25, 28, 18) {real, imag} */,
  {32'hbd8bf7de, 32'h3d420dae} /* (25, 28, 17) {real, imag} */,
  {32'h3e1078eb, 32'h00000000} /* (25, 28, 16) {real, imag} */,
  {32'hbd8bf7de, 32'hbd420dae} /* (25, 28, 15) {real, imag} */,
  {32'hbc9faa06, 32'h3db3c804} /* (25, 28, 14) {real, imag} */,
  {32'hbd076798, 32'h3d3d0aff} /* (25, 28, 13) {real, imag} */,
  {32'hbdb7dcce, 32'h3c3ab70e} /* (25, 28, 12) {real, imag} */,
  {32'h3dbe1c9d, 32'h3d6d9291} /* (25, 28, 11) {real, imag} */,
  {32'hbbc50308, 32'h3d8e2308} /* (25, 28, 10) {real, imag} */,
  {32'h3d852fa4, 32'h3d0d159e} /* (25, 28, 9) {real, imag} */,
  {32'h3cbae4e5, 32'h3e05f23d} /* (25, 28, 8) {real, imag} */,
  {32'h3d7ec37d, 32'hb82ef100} /* (25, 28, 7) {real, imag} */,
  {32'hbd43ce17, 32'hbdd27aac} /* (25, 28, 6) {real, imag} */,
  {32'h3deda673, 32'h3e62e26b} /* (25, 28, 5) {real, imag} */,
  {32'hbdc21e86, 32'hbdd328d6} /* (25, 28, 4) {real, imag} */,
  {32'h3c73c2f8, 32'h3e0a01ee} /* (25, 28, 3) {real, imag} */,
  {32'h3f3d98c8, 32'h3d4ea7f4} /* (25, 28, 2) {real, imag} */,
  {32'hc0245522, 32'hbf645b0f} /* (25, 28, 1) {real, imag} */,
  {32'hc05d778a, 32'h00000000} /* (25, 28, 0) {real, imag} */,
  {32'hc024652c, 32'h3f29e4be} /* (25, 27, 31) {real, imag} */,
  {32'h3f60413c, 32'hbd0be5a0} /* (25, 27, 30) {real, imag} */,
  {32'h3d88f712, 32'hbe5aade8} /* (25, 27, 29) {real, imag} */,
  {32'hbc99afac, 32'hbcf0de7a} /* (25, 27, 28) {real, imag} */,
  {32'h3e20e3ea, 32'hbe5ec030} /* (25, 27, 27) {real, imag} */,
  {32'h3c841904, 32'h3e1bfa24} /* (25, 27, 26) {real, imag} */,
  {32'hbd655a32, 32'h3dd606f3} /* (25, 27, 25) {real, imag} */,
  {32'hbc8f89aa, 32'hbe0c3170} /* (25, 27, 24) {real, imag} */,
  {32'hbb88f9b8, 32'h3d802dde} /* (25, 27, 23) {real, imag} */,
  {32'hbd05d6ba, 32'h3d29069b} /* (25, 27, 22) {real, imag} */,
  {32'hbd560db1, 32'hbdceabd9} /* (25, 27, 21) {real, imag} */,
  {32'hbc722bc2, 32'hbe05ea78} /* (25, 27, 20) {real, imag} */,
  {32'h3bae075a, 32'h3d829cc7} /* (25, 27, 19) {real, imag} */,
  {32'hbcb6d184, 32'hbd4de5c3} /* (25, 27, 18) {real, imag} */,
  {32'h3c25d6cc, 32'hbc784d28} /* (25, 27, 17) {real, imag} */,
  {32'h3c741fbc, 32'h00000000} /* (25, 27, 16) {real, imag} */,
  {32'h3c25d6cc, 32'h3c784d28} /* (25, 27, 15) {real, imag} */,
  {32'hbcb6d184, 32'h3d4de5c3} /* (25, 27, 14) {real, imag} */,
  {32'h3bae075a, 32'hbd829cc7} /* (25, 27, 13) {real, imag} */,
  {32'hbc722bc2, 32'h3e05ea78} /* (25, 27, 12) {real, imag} */,
  {32'hbd560db1, 32'h3dceabd9} /* (25, 27, 11) {real, imag} */,
  {32'hbd05d6ba, 32'hbd29069b} /* (25, 27, 10) {real, imag} */,
  {32'hbb88f9b8, 32'hbd802dde} /* (25, 27, 9) {real, imag} */,
  {32'hbc8f89aa, 32'h3e0c3170} /* (25, 27, 8) {real, imag} */,
  {32'hbd655a32, 32'hbdd606f3} /* (25, 27, 7) {real, imag} */,
  {32'h3c841904, 32'hbe1bfa24} /* (25, 27, 6) {real, imag} */,
  {32'h3e20e3ea, 32'h3e5ec030} /* (25, 27, 5) {real, imag} */,
  {32'hbc99afac, 32'h3cf0de7a} /* (25, 27, 4) {real, imag} */,
  {32'h3d88f712, 32'h3e5aade8} /* (25, 27, 3) {real, imag} */,
  {32'h3f60413c, 32'h3d0be5a0} /* (25, 27, 2) {real, imag} */,
  {32'hc024652c, 32'hbf29e4be} /* (25, 27, 1) {real, imag} */,
  {32'hc05cb2b2, 32'h00000000} /* (25, 27, 0) {real, imag} */,
  {32'hc01c5f65, 32'h3f1056ec} /* (25, 26, 31) {real, imag} */,
  {32'h3f4332d5, 32'h3dfb15a9} /* (25, 26, 30) {real, imag} */,
  {32'h3c9c2794, 32'h3c533356} /* (25, 26, 29) {real, imag} */,
  {32'hbcfa292d, 32'h3cd61d71} /* (25, 26, 28) {real, imag} */,
  {32'h3e05285e, 32'hbe18affd} /* (25, 26, 27) {real, imag} */,
  {32'h3d53504a, 32'h3d31e150} /* (25, 26, 26) {real, imag} */,
  {32'h3d4f9932, 32'hbb90b6f8} /* (25, 26, 25) {real, imag} */,
  {32'hbc4b745d, 32'hbe4f1450} /* (25, 26, 24) {real, imag} */,
  {32'h39d23fc0, 32'h3bb362d4} /* (25, 26, 23) {real, imag} */,
  {32'h3855e500, 32'h3d46b5d2} /* (25, 26, 22) {real, imag} */,
  {32'hbd023045, 32'h3c178c42} /* (25, 26, 21) {real, imag} */,
  {32'h3d0d7f0c, 32'h3cbb44e8} /* (25, 26, 20) {real, imag} */,
  {32'hbd272328, 32'h3d00daf8} /* (25, 26, 19) {real, imag} */,
  {32'hbd34a3ee, 32'hbcc52eb1} /* (25, 26, 18) {real, imag} */,
  {32'hbc9948ec, 32'h3bcc3e80} /* (25, 26, 17) {real, imag} */,
  {32'h3dcc921b, 32'h00000000} /* (25, 26, 16) {real, imag} */,
  {32'hbc9948ec, 32'hbbcc3e80} /* (25, 26, 15) {real, imag} */,
  {32'hbd34a3ee, 32'h3cc52eb1} /* (25, 26, 14) {real, imag} */,
  {32'hbd272328, 32'hbd00daf8} /* (25, 26, 13) {real, imag} */,
  {32'h3d0d7f0c, 32'hbcbb44e8} /* (25, 26, 12) {real, imag} */,
  {32'hbd023045, 32'hbc178c42} /* (25, 26, 11) {real, imag} */,
  {32'h3855e500, 32'hbd46b5d2} /* (25, 26, 10) {real, imag} */,
  {32'h39d23fc0, 32'hbbb362d4} /* (25, 26, 9) {real, imag} */,
  {32'hbc4b745d, 32'h3e4f1450} /* (25, 26, 8) {real, imag} */,
  {32'h3d4f9932, 32'h3b90b6f8} /* (25, 26, 7) {real, imag} */,
  {32'h3d53504a, 32'hbd31e150} /* (25, 26, 6) {real, imag} */,
  {32'h3e05285e, 32'h3e18affd} /* (25, 26, 5) {real, imag} */,
  {32'hbcfa292d, 32'hbcd61d71} /* (25, 26, 4) {real, imag} */,
  {32'h3c9c2794, 32'hbc533356} /* (25, 26, 3) {real, imag} */,
  {32'h3f4332d5, 32'hbdfb15a9} /* (25, 26, 2) {real, imag} */,
  {32'hc01c5f65, 32'hbf1056ec} /* (25, 26, 1) {real, imag} */,
  {32'hc04b4993, 32'h00000000} /* (25, 26, 0) {real, imag} */,
  {32'hc01a50b5, 32'h3ed3fe31} /* (25, 25, 31) {real, imag} */,
  {32'h3f3ca530, 32'h3e023fdc} /* (25, 25, 30) {real, imag} */,
  {32'hbc2db634, 32'h3dd03591} /* (25, 25, 29) {real, imag} */,
  {32'hbe3db77a, 32'hbd7ddc5b} /* (25, 25, 28) {real, imag} */,
  {32'h3e580b20, 32'h3cd3ee94} /* (25, 25, 27) {real, imag} */,
  {32'hbaf68220, 32'hbc3fe390} /* (25, 25, 26) {real, imag} */,
  {32'hbd6b6e22, 32'h3cc40c88} /* (25, 25, 25) {real, imag} */,
  {32'h3d4b405f, 32'h3d27a7d0} /* (25, 25, 24) {real, imag} */,
  {32'h3c2aede6, 32'hbd9eb650} /* (25, 25, 23) {real, imag} */,
  {32'h3c4ebed0, 32'h3bdd6736} /* (25, 25, 22) {real, imag} */,
  {32'hbc10d0a0, 32'hbd312db0} /* (25, 25, 21) {real, imag} */,
  {32'hbdbc66b2, 32'hbd964198} /* (25, 25, 20) {real, imag} */,
  {32'hbd1f2b3e, 32'h3d9fe008} /* (25, 25, 19) {real, imag} */,
  {32'h3deec893, 32'hbd42ac86} /* (25, 25, 18) {real, imag} */,
  {32'hbd5f3fb1, 32'h3d6ce338} /* (25, 25, 17) {real, imag} */,
  {32'h3d3227d3, 32'h00000000} /* (25, 25, 16) {real, imag} */,
  {32'hbd5f3fb1, 32'hbd6ce338} /* (25, 25, 15) {real, imag} */,
  {32'h3deec893, 32'h3d42ac86} /* (25, 25, 14) {real, imag} */,
  {32'hbd1f2b3e, 32'hbd9fe008} /* (25, 25, 13) {real, imag} */,
  {32'hbdbc66b2, 32'h3d964198} /* (25, 25, 12) {real, imag} */,
  {32'hbc10d0a0, 32'h3d312db0} /* (25, 25, 11) {real, imag} */,
  {32'h3c4ebed0, 32'hbbdd6736} /* (25, 25, 10) {real, imag} */,
  {32'h3c2aede6, 32'h3d9eb650} /* (25, 25, 9) {real, imag} */,
  {32'h3d4b405f, 32'hbd27a7d0} /* (25, 25, 8) {real, imag} */,
  {32'hbd6b6e22, 32'hbcc40c88} /* (25, 25, 7) {real, imag} */,
  {32'hbaf68220, 32'h3c3fe390} /* (25, 25, 6) {real, imag} */,
  {32'h3e580b20, 32'hbcd3ee94} /* (25, 25, 5) {real, imag} */,
  {32'hbe3db77a, 32'h3d7ddc5b} /* (25, 25, 4) {real, imag} */,
  {32'hbc2db634, 32'hbdd03591} /* (25, 25, 3) {real, imag} */,
  {32'h3f3ca530, 32'hbe023fdc} /* (25, 25, 2) {real, imag} */,
  {32'hc01a50b5, 32'hbed3fe31} /* (25, 25, 1) {real, imag} */,
  {32'hc0391734, 32'h00000000} /* (25, 25, 0) {real, imag} */,
  {32'hc00a7fde, 32'h3ea08ec8} /* (25, 24, 31) {real, imag} */,
  {32'h3f32013a, 32'hbc075d10} /* (25, 24, 30) {real, imag} */,
  {32'hbdd4405c, 32'hbb3ccdb0} /* (25, 24, 29) {real, imag} */,
  {32'hbe362e9b, 32'hbddd0065} /* (25, 24, 28) {real, imag} */,
  {32'h3e45d0cd, 32'h3d48c136} /* (25, 24, 27) {real, imag} */,
  {32'hbd730c21, 32'h3bc8f920} /* (25, 24, 26) {real, imag} */,
  {32'h3d7fced0, 32'h3a61cc80} /* (25, 24, 25) {real, imag} */,
  {32'h3ca34327, 32'hbd961af0} /* (25, 24, 24) {real, imag} */,
  {32'h3ba7fe38, 32'hbc249ed2} /* (25, 24, 23) {real, imag} */,
  {32'hbd78bbdb, 32'h3d035de8} /* (25, 24, 22) {real, imag} */,
  {32'h3d60fe0e, 32'hbd654026} /* (25, 24, 21) {real, imag} */,
  {32'h3c9bbe7b, 32'hbdd24d4e} /* (25, 24, 20) {real, imag} */,
  {32'h3b7f7320, 32'hbc54d06a} /* (25, 24, 19) {real, imag} */,
  {32'h3cef9abc, 32'h3c6f54ac} /* (25, 24, 18) {real, imag} */,
  {32'h3b878b20, 32'hbc29b822} /* (25, 24, 17) {real, imag} */,
  {32'h3d070e08, 32'h00000000} /* (25, 24, 16) {real, imag} */,
  {32'h3b878b20, 32'h3c29b822} /* (25, 24, 15) {real, imag} */,
  {32'h3cef9abc, 32'hbc6f54ac} /* (25, 24, 14) {real, imag} */,
  {32'h3b7f7320, 32'h3c54d06a} /* (25, 24, 13) {real, imag} */,
  {32'h3c9bbe7b, 32'h3dd24d4e} /* (25, 24, 12) {real, imag} */,
  {32'h3d60fe0e, 32'h3d654026} /* (25, 24, 11) {real, imag} */,
  {32'hbd78bbdb, 32'hbd035de8} /* (25, 24, 10) {real, imag} */,
  {32'h3ba7fe38, 32'h3c249ed2} /* (25, 24, 9) {real, imag} */,
  {32'h3ca34327, 32'h3d961af0} /* (25, 24, 8) {real, imag} */,
  {32'h3d7fced0, 32'hba61cc80} /* (25, 24, 7) {real, imag} */,
  {32'hbd730c21, 32'hbbc8f920} /* (25, 24, 6) {real, imag} */,
  {32'h3e45d0cd, 32'hbd48c136} /* (25, 24, 5) {real, imag} */,
  {32'hbe362e9b, 32'h3ddd0065} /* (25, 24, 4) {real, imag} */,
  {32'hbdd4405c, 32'h3b3ccdb0} /* (25, 24, 3) {real, imag} */,
  {32'h3f32013a, 32'h3c075d10} /* (25, 24, 2) {real, imag} */,
  {32'hc00a7fde, 32'hbea08ec8} /* (25, 24, 1) {real, imag} */,
  {32'hc025242a, 32'h00000000} /* (25, 24, 0) {real, imag} */,
  {32'hc000cca2, 32'h3e9dabba} /* (25, 23, 31) {real, imag} */,
  {32'h3f3d60f9, 32'hbd2dc232} /* (25, 23, 30) {real, imag} */,
  {32'hbd2b8b86, 32'hbdbdfe11} /* (25, 23, 29) {real, imag} */,
  {32'hbca1437a, 32'hbceb9969} /* (25, 23, 28) {real, imag} */,
  {32'h3e03177b, 32'h3dac4fea} /* (25, 23, 27) {real, imag} */,
  {32'hbdc416ff, 32'hbde9aa46} /* (25, 23, 26) {real, imag} */,
  {32'hbde84aae, 32'hbd145216} /* (25, 23, 25) {real, imag} */,
  {32'h3d82fc14, 32'hbe247295} /* (25, 23, 24) {real, imag} */,
  {32'h3ab51ad0, 32'hbe09b8b6} /* (25, 23, 23) {real, imag} */,
  {32'hbe1c78ac, 32'h3d45f62e} /* (25, 23, 22) {real, imag} */,
  {32'h3dd1222c, 32'hbb3b2ac0} /* (25, 23, 21) {real, imag} */,
  {32'hbc8938b2, 32'hbc1e89e5} /* (25, 23, 20) {real, imag} */,
  {32'h3cfe8f4b, 32'hbd526232} /* (25, 23, 19) {real, imag} */,
  {32'hbcd6adf7, 32'h3d969464} /* (25, 23, 18) {real, imag} */,
  {32'h3d123fa2, 32'h3d85d482} /* (25, 23, 17) {real, imag} */,
  {32'h3c9eb672, 32'h00000000} /* (25, 23, 16) {real, imag} */,
  {32'h3d123fa2, 32'hbd85d482} /* (25, 23, 15) {real, imag} */,
  {32'hbcd6adf7, 32'hbd969464} /* (25, 23, 14) {real, imag} */,
  {32'h3cfe8f4b, 32'h3d526232} /* (25, 23, 13) {real, imag} */,
  {32'hbc8938b2, 32'h3c1e89e5} /* (25, 23, 12) {real, imag} */,
  {32'h3dd1222c, 32'h3b3b2ac0} /* (25, 23, 11) {real, imag} */,
  {32'hbe1c78ac, 32'hbd45f62e} /* (25, 23, 10) {real, imag} */,
  {32'h3ab51ad0, 32'h3e09b8b6} /* (25, 23, 9) {real, imag} */,
  {32'h3d82fc14, 32'h3e247295} /* (25, 23, 8) {real, imag} */,
  {32'hbde84aae, 32'h3d145216} /* (25, 23, 7) {real, imag} */,
  {32'hbdc416ff, 32'h3de9aa46} /* (25, 23, 6) {real, imag} */,
  {32'h3e03177b, 32'hbdac4fea} /* (25, 23, 5) {real, imag} */,
  {32'hbca1437a, 32'h3ceb9969} /* (25, 23, 4) {real, imag} */,
  {32'hbd2b8b86, 32'h3dbdfe11} /* (25, 23, 3) {real, imag} */,
  {32'h3f3d60f9, 32'h3d2dc232} /* (25, 23, 2) {real, imag} */,
  {32'hc000cca2, 32'hbe9dabba} /* (25, 23, 1) {real, imag} */,
  {32'hc0073a84, 32'h00000000} /* (25, 23, 0) {real, imag} */,
  {32'hbfd3ca33, 32'h3e38b5ad} /* (25, 22, 31) {real, imag} */,
  {32'h3f290569, 32'hbdef4ad7} /* (25, 22, 30) {real, imag} */,
  {32'h3d894273, 32'h3d3b1076} /* (25, 22, 29) {real, imag} */,
  {32'hbdeff18f, 32'h3df7fa28} /* (25, 22, 28) {real, imag} */,
  {32'h3e3ad70a, 32'hbb05f370} /* (25, 22, 27) {real, imag} */,
  {32'hbd090a14, 32'h3d676af6} /* (25, 22, 26) {real, imag} */,
  {32'hbc5eb0a2, 32'hbc13b21c} /* (25, 22, 25) {real, imag} */,
  {32'h3ba1498a, 32'hbc29e730} /* (25, 22, 24) {real, imag} */,
  {32'h3caf8ab9, 32'h3d474d02} /* (25, 22, 23) {real, imag} */,
  {32'hbc058d50, 32'h3d07ecc4} /* (25, 22, 22) {real, imag} */,
  {32'h3bfc6458, 32'h3d831f5e} /* (25, 22, 21) {real, imag} */,
  {32'hbb1d97bc, 32'hbc21181f} /* (25, 22, 20) {real, imag} */,
  {32'hbcd76e2c, 32'h3da2ada4} /* (25, 22, 19) {real, imag} */,
  {32'hbbc57a9b, 32'hbe23da24} /* (25, 22, 18) {real, imag} */,
  {32'hba97ad80, 32'hbd11b12f} /* (25, 22, 17) {real, imag} */,
  {32'hbcbaf0e2, 32'h00000000} /* (25, 22, 16) {real, imag} */,
  {32'hba97ad80, 32'h3d11b12f} /* (25, 22, 15) {real, imag} */,
  {32'hbbc57a9b, 32'h3e23da24} /* (25, 22, 14) {real, imag} */,
  {32'hbcd76e2c, 32'hbda2ada4} /* (25, 22, 13) {real, imag} */,
  {32'hbb1d97bc, 32'h3c21181f} /* (25, 22, 12) {real, imag} */,
  {32'h3bfc6458, 32'hbd831f5e} /* (25, 22, 11) {real, imag} */,
  {32'hbc058d50, 32'hbd07ecc4} /* (25, 22, 10) {real, imag} */,
  {32'h3caf8ab9, 32'hbd474d02} /* (25, 22, 9) {real, imag} */,
  {32'h3ba1498a, 32'h3c29e730} /* (25, 22, 8) {real, imag} */,
  {32'hbc5eb0a2, 32'h3c13b21c} /* (25, 22, 7) {real, imag} */,
  {32'hbd090a14, 32'hbd676af6} /* (25, 22, 6) {real, imag} */,
  {32'h3e3ad70a, 32'h3b05f370} /* (25, 22, 5) {real, imag} */,
  {32'hbdeff18f, 32'hbdf7fa28} /* (25, 22, 4) {real, imag} */,
  {32'h3d894273, 32'hbd3b1076} /* (25, 22, 3) {real, imag} */,
  {32'h3f290569, 32'h3def4ad7} /* (25, 22, 2) {real, imag} */,
  {32'hbfd3ca33, 32'hbe38b5ad} /* (25, 22, 1) {real, imag} */,
  {32'hbfc08995, 32'h00000000} /* (25, 22, 0) {real, imag} */,
  {32'hbf557486, 32'h3d25b850} /* (25, 21, 31) {real, imag} */,
  {32'h3ee0308b, 32'h3cf0a5d8} /* (25, 21, 30) {real, imag} */,
  {32'h3c9d84d8, 32'h3e88aec2} /* (25, 21, 29) {real, imag} */,
  {32'hbe3a9a70, 32'hbdb1bfa8} /* (25, 21, 28) {real, imag} */,
  {32'h3dd72307, 32'hbd7d84cc} /* (25, 21, 27) {real, imag} */,
  {32'h3dab7502, 32'h3e1f42fd} /* (25, 21, 26) {real, imag} */,
  {32'hbdae99bc, 32'h3c96d5ae} /* (25, 21, 25) {real, imag} */,
  {32'h3cff9706, 32'h3cfeaae8} /* (25, 21, 24) {real, imag} */,
  {32'h3df4255e, 32'hbc251810} /* (25, 21, 23) {real, imag} */,
  {32'h3adbcf10, 32'hbb0774bc} /* (25, 21, 22) {real, imag} */,
  {32'h3dae404c, 32'hbddd4d40} /* (25, 21, 21) {real, imag} */,
  {32'h3c4506f4, 32'hbbec3b1c} /* (25, 21, 20) {real, imag} */,
  {32'h3d53047e, 32'hbc4ebf40} /* (25, 21, 19) {real, imag} */,
  {32'hbdc838d1, 32'hbaa2d210} /* (25, 21, 18) {real, imag} */,
  {32'h3d6fe918, 32'hbd4e005a} /* (25, 21, 17) {real, imag} */,
  {32'h3e0e407e, 32'h00000000} /* (25, 21, 16) {real, imag} */,
  {32'h3d6fe918, 32'h3d4e005a} /* (25, 21, 15) {real, imag} */,
  {32'hbdc838d1, 32'h3aa2d210} /* (25, 21, 14) {real, imag} */,
  {32'h3d53047e, 32'h3c4ebf40} /* (25, 21, 13) {real, imag} */,
  {32'h3c4506f4, 32'h3bec3b1c} /* (25, 21, 12) {real, imag} */,
  {32'h3dae404c, 32'h3ddd4d40} /* (25, 21, 11) {real, imag} */,
  {32'h3adbcf10, 32'h3b0774bc} /* (25, 21, 10) {real, imag} */,
  {32'h3df4255e, 32'h3c251810} /* (25, 21, 9) {real, imag} */,
  {32'h3cff9706, 32'hbcfeaae8} /* (25, 21, 8) {real, imag} */,
  {32'hbdae99bc, 32'hbc96d5ae} /* (25, 21, 7) {real, imag} */,
  {32'h3dab7502, 32'hbe1f42fd} /* (25, 21, 6) {real, imag} */,
  {32'h3dd72307, 32'h3d7d84cc} /* (25, 21, 5) {real, imag} */,
  {32'hbe3a9a70, 32'h3db1bfa8} /* (25, 21, 4) {real, imag} */,
  {32'h3c9d84d8, 32'hbe88aec2} /* (25, 21, 3) {real, imag} */,
  {32'h3ee0308b, 32'hbcf0a5d8} /* (25, 21, 2) {real, imag} */,
  {32'hbf557486, 32'hbd25b850} /* (25, 21, 1) {real, imag} */,
  {32'hbf4d75e1, 32'h00000000} /* (25, 21, 0) {real, imag} */,
  {32'h3ea540c3, 32'hbdf9a600} /* (25, 20, 31) {real, imag} */,
  {32'hbe572a02, 32'h3dde6b47} /* (25, 20, 30) {real, imag} */,
  {32'h3d937ad7, 32'h3d21f3f1} /* (25, 20, 29) {real, imag} */,
  {32'h3bf7b6d0, 32'hbe246f21} /* (25, 20, 28) {real, imag} */,
  {32'hb9df2880, 32'h3d97f18c} /* (25, 20, 27) {real, imag} */,
  {32'h3ddc5198, 32'h3e5421e4} /* (25, 20, 26) {real, imag} */,
  {32'h3d3ae675, 32'hbd8815ac} /* (25, 20, 25) {real, imag} */,
  {32'hbc5c7088, 32'h3d8cc6e6} /* (25, 20, 24) {real, imag} */,
  {32'h3bb1ca58, 32'hbd5eeb8a} /* (25, 20, 23) {real, imag} */,
  {32'h3d8b096c, 32'h3d70818c} /* (25, 20, 22) {real, imag} */,
  {32'h3d68395e, 32'h3d3eb97a} /* (25, 20, 21) {real, imag} */,
  {32'h3c0de50c, 32'h3cd1267c} /* (25, 20, 20) {real, imag} */,
  {32'hbcd547e7, 32'h3d081c3a} /* (25, 20, 19) {real, imag} */,
  {32'hbd64c3cf, 32'h3bf25608} /* (25, 20, 18) {real, imag} */,
  {32'hbcaa032c, 32'hbdd62c29} /* (25, 20, 17) {real, imag} */,
  {32'h3c9e476e, 32'h00000000} /* (25, 20, 16) {real, imag} */,
  {32'hbcaa032c, 32'h3dd62c29} /* (25, 20, 15) {real, imag} */,
  {32'hbd64c3cf, 32'hbbf25608} /* (25, 20, 14) {real, imag} */,
  {32'hbcd547e7, 32'hbd081c3a} /* (25, 20, 13) {real, imag} */,
  {32'h3c0de50c, 32'hbcd1267c} /* (25, 20, 12) {real, imag} */,
  {32'h3d68395e, 32'hbd3eb97a} /* (25, 20, 11) {real, imag} */,
  {32'h3d8b096c, 32'hbd70818c} /* (25, 20, 10) {real, imag} */,
  {32'h3bb1ca58, 32'h3d5eeb8a} /* (25, 20, 9) {real, imag} */,
  {32'hbc5c7088, 32'hbd8cc6e6} /* (25, 20, 8) {real, imag} */,
  {32'h3d3ae675, 32'h3d8815ac} /* (25, 20, 7) {real, imag} */,
  {32'h3ddc5198, 32'hbe5421e4} /* (25, 20, 6) {real, imag} */,
  {32'hb9df2880, 32'hbd97f18c} /* (25, 20, 5) {real, imag} */,
  {32'h3bf7b6d0, 32'h3e246f21} /* (25, 20, 4) {real, imag} */,
  {32'h3d937ad7, 32'hbd21f3f1} /* (25, 20, 3) {real, imag} */,
  {32'hbe572a02, 32'hbdde6b47} /* (25, 20, 2) {real, imag} */,
  {32'h3ea540c3, 32'h3df9a600} /* (25, 20, 1) {real, imag} */,
  {32'h3e6e773c, 32'h00000000} /* (25, 20, 0) {real, imag} */,
  {32'h3f501dd3, 32'hbe28dd9a} /* (25, 19, 31) {real, imag} */,
  {32'hbedbadfc, 32'hbd14cfd2} /* (25, 19, 30) {real, imag} */,
  {32'h3c808e78, 32'hbda149fa} /* (25, 19, 29) {real, imag} */,
  {32'h3e176daf, 32'hbddda6a6} /* (25, 19, 28) {real, imag} */,
  {32'hbde7492a, 32'h3e0e09be} /* (25, 19, 27) {real, imag} */,
  {32'h3d8a17b4, 32'hbc6b9adc} /* (25, 19, 26) {real, imag} */,
  {32'h3dcc416a, 32'hbd7984d7} /* (25, 19, 25) {real, imag} */,
  {32'hbdf68fe1, 32'hbcc23691} /* (25, 19, 24) {real, imag} */,
  {32'h3d033af6, 32'h3a85dbe0} /* (25, 19, 23) {real, imag} */,
  {32'h3da99394, 32'h3d15d99c} /* (25, 19, 22) {real, imag} */,
  {32'hbdb23ee4, 32'h3da34434} /* (25, 19, 21) {real, imag} */,
  {32'hbc2d9556, 32'hbcffeea3} /* (25, 19, 20) {real, imag} */,
  {32'h3cedb574, 32'hbcd1cf24} /* (25, 19, 19) {real, imag} */,
  {32'hbc52a79e, 32'hbb0ea40c} /* (25, 19, 18) {real, imag} */,
  {32'h3c3a6cb2, 32'hbc36e4a6} /* (25, 19, 17) {real, imag} */,
  {32'hbd9f6069, 32'h00000000} /* (25, 19, 16) {real, imag} */,
  {32'h3c3a6cb2, 32'h3c36e4a6} /* (25, 19, 15) {real, imag} */,
  {32'hbc52a79e, 32'h3b0ea40c} /* (25, 19, 14) {real, imag} */,
  {32'h3cedb574, 32'h3cd1cf24} /* (25, 19, 13) {real, imag} */,
  {32'hbc2d9556, 32'h3cffeea3} /* (25, 19, 12) {real, imag} */,
  {32'hbdb23ee4, 32'hbda34434} /* (25, 19, 11) {real, imag} */,
  {32'h3da99394, 32'hbd15d99c} /* (25, 19, 10) {real, imag} */,
  {32'h3d033af6, 32'hba85dbe0} /* (25, 19, 9) {real, imag} */,
  {32'hbdf68fe1, 32'h3cc23691} /* (25, 19, 8) {real, imag} */,
  {32'h3dcc416a, 32'h3d7984d7} /* (25, 19, 7) {real, imag} */,
  {32'h3d8a17b4, 32'h3c6b9adc} /* (25, 19, 6) {real, imag} */,
  {32'hbde7492a, 32'hbe0e09be} /* (25, 19, 5) {real, imag} */,
  {32'h3e176daf, 32'h3ddda6a6} /* (25, 19, 4) {real, imag} */,
  {32'h3c808e78, 32'h3da149fa} /* (25, 19, 3) {real, imag} */,
  {32'hbedbadfc, 32'h3d14cfd2} /* (25, 19, 2) {real, imag} */,
  {32'h3f501dd3, 32'h3e28dd9a} /* (25, 19, 1) {real, imag} */,
  {32'h3f40d512, 32'h00000000} /* (25, 19, 0) {real, imag} */,
  {32'h3fa10cca, 32'hbdca50c8} /* (25, 18, 31) {real, imag} */,
  {32'hbf07810a, 32'h3d0136aa} /* (25, 18, 30) {real, imag} */,
  {32'hbb192d50, 32'hbbe3e038} /* (25, 18, 29) {real, imag} */,
  {32'h3e5d357e, 32'hbd8fba7c} /* (25, 18, 28) {real, imag} */,
  {32'h3c03169c, 32'h3da4c8e5} /* (25, 18, 27) {real, imag} */,
  {32'h3c655bee, 32'h3b51da28} /* (25, 18, 26) {real, imag} */,
  {32'hbcb7773e, 32'hbb93f218} /* (25, 18, 25) {real, imag} */,
  {32'hbd980f82, 32'hbd8443d4} /* (25, 18, 24) {real, imag} */,
  {32'hbe118a32, 32'hbc659938} /* (25, 18, 23) {real, imag} */,
  {32'hbdadedf4, 32'hbd193cf0} /* (25, 18, 22) {real, imag} */,
  {32'hbd296d15, 32'hbc13498c} /* (25, 18, 21) {real, imag} */,
  {32'h3bd8171c, 32'h3d155d6a} /* (25, 18, 20) {real, imag} */,
  {32'hbd3bfe29, 32'hbda8b482} /* (25, 18, 19) {real, imag} */,
  {32'h3d26b13b, 32'hbd8394ec} /* (25, 18, 18) {real, imag} */,
  {32'h3c24207e, 32'h3c06daca} /* (25, 18, 17) {real, imag} */,
  {32'h3d44df2f, 32'h00000000} /* (25, 18, 16) {real, imag} */,
  {32'h3c24207e, 32'hbc06daca} /* (25, 18, 15) {real, imag} */,
  {32'h3d26b13b, 32'h3d8394ec} /* (25, 18, 14) {real, imag} */,
  {32'hbd3bfe29, 32'h3da8b482} /* (25, 18, 13) {real, imag} */,
  {32'h3bd8171c, 32'hbd155d6a} /* (25, 18, 12) {real, imag} */,
  {32'hbd296d15, 32'h3c13498c} /* (25, 18, 11) {real, imag} */,
  {32'hbdadedf4, 32'h3d193cf0} /* (25, 18, 10) {real, imag} */,
  {32'hbe118a32, 32'h3c659938} /* (25, 18, 9) {real, imag} */,
  {32'hbd980f82, 32'h3d8443d4} /* (25, 18, 8) {real, imag} */,
  {32'hbcb7773e, 32'h3b93f218} /* (25, 18, 7) {real, imag} */,
  {32'h3c655bee, 32'hbb51da28} /* (25, 18, 6) {real, imag} */,
  {32'h3c03169c, 32'hbda4c8e5} /* (25, 18, 5) {real, imag} */,
  {32'h3e5d357e, 32'h3d8fba7c} /* (25, 18, 4) {real, imag} */,
  {32'hbb192d50, 32'h3be3e038} /* (25, 18, 3) {real, imag} */,
  {32'hbf07810a, 32'hbd0136aa} /* (25, 18, 2) {real, imag} */,
  {32'h3fa10cca, 32'h3dca50c8} /* (25, 18, 1) {real, imag} */,
  {32'h3f7a8d04, 32'h00000000} /* (25, 18, 0) {real, imag} */,
  {32'h3fc39ba2, 32'hbe4336e5} /* (25, 17, 31) {real, imag} */,
  {32'hbf45f14a, 32'h3da120c6} /* (25, 17, 30) {real, imag} */,
  {32'hbd9b7d5e, 32'hbd6d0752} /* (25, 17, 29) {real, imag} */,
  {32'h3e5e4f30, 32'hbd8d58f6} /* (25, 17, 28) {real, imag} */,
  {32'hbd7b919d, 32'h3da43691} /* (25, 17, 27) {real, imag} */,
  {32'hbd011020, 32'h3d9dcb9a} /* (25, 17, 26) {real, imag} */,
  {32'hbd066fa4, 32'h3c2c1bfa} /* (25, 17, 25) {real, imag} */,
  {32'hbbe8be68, 32'hbd9646ad} /* (25, 17, 24) {real, imag} */,
  {32'h3b7fdaf8, 32'hbce5d194} /* (25, 17, 23) {real, imag} */,
  {32'hbc3ee21f, 32'hbd0afbfc} /* (25, 17, 22) {real, imag} */,
  {32'hbc07efb0, 32'h3d6af270} /* (25, 17, 21) {real, imag} */,
  {32'h3d306848, 32'hbd7499b7} /* (25, 17, 20) {real, imag} */,
  {32'h3d74a3dc, 32'hbd45f596} /* (25, 17, 19) {real, imag} */,
  {32'h3c8029c8, 32'h3cc915d7} /* (25, 17, 18) {real, imag} */,
  {32'hbc7ffa56, 32'hbc1a131c} /* (25, 17, 17) {real, imag} */,
  {32'hbcd47347, 32'h00000000} /* (25, 17, 16) {real, imag} */,
  {32'hbc7ffa56, 32'h3c1a131c} /* (25, 17, 15) {real, imag} */,
  {32'h3c8029c8, 32'hbcc915d7} /* (25, 17, 14) {real, imag} */,
  {32'h3d74a3dc, 32'h3d45f596} /* (25, 17, 13) {real, imag} */,
  {32'h3d306848, 32'h3d7499b7} /* (25, 17, 12) {real, imag} */,
  {32'hbc07efb0, 32'hbd6af270} /* (25, 17, 11) {real, imag} */,
  {32'hbc3ee21f, 32'h3d0afbfc} /* (25, 17, 10) {real, imag} */,
  {32'h3b7fdaf8, 32'h3ce5d194} /* (25, 17, 9) {real, imag} */,
  {32'hbbe8be68, 32'h3d9646ad} /* (25, 17, 8) {real, imag} */,
  {32'hbd066fa4, 32'hbc2c1bfa} /* (25, 17, 7) {real, imag} */,
  {32'hbd011020, 32'hbd9dcb9a} /* (25, 17, 6) {real, imag} */,
  {32'hbd7b919d, 32'hbda43691} /* (25, 17, 5) {real, imag} */,
  {32'h3e5e4f30, 32'h3d8d58f6} /* (25, 17, 4) {real, imag} */,
  {32'hbd9b7d5e, 32'h3d6d0752} /* (25, 17, 3) {real, imag} */,
  {32'hbf45f14a, 32'hbda120c6} /* (25, 17, 2) {real, imag} */,
  {32'h3fc39ba2, 32'h3e4336e5} /* (25, 17, 1) {real, imag} */,
  {32'h3fa2e52d, 32'h00000000} /* (25, 17, 0) {real, imag} */,
  {32'h3fed3f81, 32'hbd2ebb10} /* (25, 16, 31) {real, imag} */,
  {32'hbf2810da, 32'h3e9bb818} /* (25, 16, 30) {real, imag} */,
  {32'hbe369933, 32'hbd9bdc8c} /* (25, 16, 29) {real, imag} */,
  {32'h3e2dbb53, 32'hbe2d734a} /* (25, 16, 28) {real, imag} */,
  {32'hbd1fc86a, 32'h3ce48eff} /* (25, 16, 27) {real, imag} */,
  {32'hbc6c1af4, 32'h3d8fdf38} /* (25, 16, 26) {real, imag} */,
  {32'hbc94a3cc, 32'h3db2415e} /* (25, 16, 25) {real, imag} */,
  {32'hbdcace42, 32'hbcd5061e} /* (25, 16, 24) {real, imag} */,
  {32'h3dbf5dae, 32'hbdd6dcba} /* (25, 16, 23) {real, imag} */,
  {32'h3e0afe26, 32'hbd9377c8} /* (25, 16, 22) {real, imag} */,
  {32'h3ce3feb0, 32'h3c54bbf4} /* (25, 16, 21) {real, imag} */,
  {32'hbdba3fe3, 32'h3d5dea0a} /* (25, 16, 20) {real, imag} */,
  {32'hbc16d99c, 32'h3de401ab} /* (25, 16, 19) {real, imag} */,
  {32'hbd20b36c, 32'hbc556146} /* (25, 16, 18) {real, imag} */,
  {32'h3da988d6, 32'hbd94e10c} /* (25, 16, 17) {real, imag} */,
  {32'h3da3991d, 32'h00000000} /* (25, 16, 16) {real, imag} */,
  {32'h3da988d6, 32'h3d94e10c} /* (25, 16, 15) {real, imag} */,
  {32'hbd20b36c, 32'h3c556146} /* (25, 16, 14) {real, imag} */,
  {32'hbc16d99c, 32'hbde401ab} /* (25, 16, 13) {real, imag} */,
  {32'hbdba3fe3, 32'hbd5dea0a} /* (25, 16, 12) {real, imag} */,
  {32'h3ce3feb0, 32'hbc54bbf4} /* (25, 16, 11) {real, imag} */,
  {32'h3e0afe26, 32'h3d9377c8} /* (25, 16, 10) {real, imag} */,
  {32'h3dbf5dae, 32'h3dd6dcba} /* (25, 16, 9) {real, imag} */,
  {32'hbdcace42, 32'h3cd5061e} /* (25, 16, 8) {real, imag} */,
  {32'hbc94a3cc, 32'hbdb2415e} /* (25, 16, 7) {real, imag} */,
  {32'hbc6c1af4, 32'hbd8fdf38} /* (25, 16, 6) {real, imag} */,
  {32'hbd1fc86a, 32'hbce48eff} /* (25, 16, 5) {real, imag} */,
  {32'h3e2dbb53, 32'h3e2d734a} /* (25, 16, 4) {real, imag} */,
  {32'hbe369933, 32'h3d9bdc8c} /* (25, 16, 3) {real, imag} */,
  {32'hbf2810da, 32'hbe9bb818} /* (25, 16, 2) {real, imag} */,
  {32'h3fed3f81, 32'h3d2ebb10} /* (25, 16, 1) {real, imag} */,
  {32'h3faed6c8, 32'h00000000} /* (25, 16, 0) {real, imag} */,
  {32'h3fe669fa, 32'hbcb0c298} /* (25, 15, 31) {real, imag} */,
  {32'hbf242b78, 32'h3e281d5d} /* (25, 15, 30) {real, imag} */,
  {32'h3d094f28, 32'hbd1b8226} /* (25, 15, 29) {real, imag} */,
  {32'h3beb36f0, 32'hbe12aecd} /* (25, 15, 28) {real, imag} */,
  {32'hbe2e0995, 32'hba87d540} /* (25, 15, 27) {real, imag} */,
  {32'hbcddc088, 32'h3d07a248} /* (25, 15, 26) {real, imag} */,
  {32'h3dc1bb5c, 32'hbd19846c} /* (25, 15, 25) {real, imag} */,
  {32'h3c780ba4, 32'hbbfd1db0} /* (25, 15, 24) {real, imag} */,
  {32'hbaf2e650, 32'hbc2ab628} /* (25, 15, 23) {real, imag} */,
  {32'h3c75dbfd, 32'hbc00eff3} /* (25, 15, 22) {real, imag} */,
  {32'hbc07b02c, 32'h3d0c4cf8} /* (25, 15, 21) {real, imag} */,
  {32'hbd4fec3c, 32'hbd545899} /* (25, 15, 20) {real, imag} */,
  {32'hbd32588c, 32'h3d2afe4a} /* (25, 15, 19) {real, imag} */,
  {32'h3cff6388, 32'hbbba92fc} /* (25, 15, 18) {real, imag} */,
  {32'h3cba6047, 32'h3c4ad582} /* (25, 15, 17) {real, imag} */,
  {32'h3d055eea, 32'h00000000} /* (25, 15, 16) {real, imag} */,
  {32'h3cba6047, 32'hbc4ad582} /* (25, 15, 15) {real, imag} */,
  {32'h3cff6388, 32'h3bba92fc} /* (25, 15, 14) {real, imag} */,
  {32'hbd32588c, 32'hbd2afe4a} /* (25, 15, 13) {real, imag} */,
  {32'hbd4fec3c, 32'h3d545899} /* (25, 15, 12) {real, imag} */,
  {32'hbc07b02c, 32'hbd0c4cf8} /* (25, 15, 11) {real, imag} */,
  {32'h3c75dbfd, 32'h3c00eff3} /* (25, 15, 10) {real, imag} */,
  {32'hbaf2e650, 32'h3c2ab628} /* (25, 15, 9) {real, imag} */,
  {32'h3c780ba4, 32'h3bfd1db0} /* (25, 15, 8) {real, imag} */,
  {32'h3dc1bb5c, 32'h3d19846c} /* (25, 15, 7) {real, imag} */,
  {32'hbcddc088, 32'hbd07a248} /* (25, 15, 6) {real, imag} */,
  {32'hbe2e0995, 32'h3a87d540} /* (25, 15, 5) {real, imag} */,
  {32'h3beb36f0, 32'h3e12aecd} /* (25, 15, 4) {real, imag} */,
  {32'h3d094f28, 32'h3d1b8226} /* (25, 15, 3) {real, imag} */,
  {32'hbf242b78, 32'hbe281d5d} /* (25, 15, 2) {real, imag} */,
  {32'h3fe669fa, 32'h3cb0c298} /* (25, 15, 1) {real, imag} */,
  {32'h3f91929b, 32'h00000000} /* (25, 15, 0) {real, imag} */,
  {32'h3fdeda42, 32'hbc01b1c0} /* (25, 14, 31) {real, imag} */,
  {32'hbf36137e, 32'h3e164948} /* (25, 14, 30) {real, imag} */,
  {32'hbcbdb2f6, 32'hbd35a6d9} /* (25, 14, 29) {real, imag} */,
  {32'h3d0a3184, 32'hbdaaf5a8} /* (25, 14, 28) {real, imag} */,
  {32'hbdb2cfd2, 32'h3d8c36af} /* (25, 14, 27) {real, imag} */,
  {32'h3c5404f8, 32'hbc312806} /* (25, 14, 26) {real, imag} */,
  {32'h3d281637, 32'hbc4404a8} /* (25, 14, 25) {real, imag} */,
  {32'hbc4d74c0, 32'h3b2e3440} /* (25, 14, 24) {real, imag} */,
  {32'hbb154c20, 32'h3c9b0778} /* (25, 14, 23) {real, imag} */,
  {32'hbd7ce399, 32'h3d8f405c} /* (25, 14, 22) {real, imag} */,
  {32'h3d389ac3, 32'h3cd57782} /* (25, 14, 21) {real, imag} */,
  {32'hbd556476, 32'hbb9f163c} /* (25, 14, 20) {real, imag} */,
  {32'h3cd1c31a, 32'hbd05ca54} /* (25, 14, 19) {real, imag} */,
  {32'hbc9d3d74, 32'h3ca91957} /* (25, 14, 18) {real, imag} */,
  {32'hbd3ab926, 32'hbcbe9ee3} /* (25, 14, 17) {real, imag} */,
  {32'hbd9534a0, 32'h00000000} /* (25, 14, 16) {real, imag} */,
  {32'hbd3ab926, 32'h3cbe9ee3} /* (25, 14, 15) {real, imag} */,
  {32'hbc9d3d74, 32'hbca91957} /* (25, 14, 14) {real, imag} */,
  {32'h3cd1c31a, 32'h3d05ca54} /* (25, 14, 13) {real, imag} */,
  {32'hbd556476, 32'h3b9f163c} /* (25, 14, 12) {real, imag} */,
  {32'h3d389ac3, 32'hbcd57782} /* (25, 14, 11) {real, imag} */,
  {32'hbd7ce399, 32'hbd8f405c} /* (25, 14, 10) {real, imag} */,
  {32'hbb154c20, 32'hbc9b0778} /* (25, 14, 9) {real, imag} */,
  {32'hbc4d74c0, 32'hbb2e3440} /* (25, 14, 8) {real, imag} */,
  {32'h3d281637, 32'h3c4404a8} /* (25, 14, 7) {real, imag} */,
  {32'h3c5404f8, 32'h3c312806} /* (25, 14, 6) {real, imag} */,
  {32'hbdb2cfd2, 32'hbd8c36af} /* (25, 14, 5) {real, imag} */,
  {32'h3d0a3184, 32'h3daaf5a8} /* (25, 14, 4) {real, imag} */,
  {32'hbcbdb2f6, 32'h3d35a6d9} /* (25, 14, 3) {real, imag} */,
  {32'hbf36137e, 32'hbe164948} /* (25, 14, 2) {real, imag} */,
  {32'h3fdeda42, 32'h3c01b1c0} /* (25, 14, 1) {real, imag} */,
  {32'h3f6e84a4, 32'h00000000} /* (25, 14, 0) {real, imag} */,
  {32'h3fccf586, 32'h3d1e9b28} /* (25, 13, 31) {real, imag} */,
  {32'hbf4a8096, 32'h3e1f4b84} /* (25, 13, 30) {real, imag} */,
  {32'hbd50b650, 32'hbc871f1e} /* (25, 13, 29) {real, imag} */,
  {32'hbcc13210, 32'hbde45b80} /* (25, 13, 28) {real, imag} */,
  {32'hbdc5af9e, 32'hbcb40144} /* (25, 13, 27) {real, imag} */,
  {32'hbd4888f8, 32'h3c32cc18} /* (25, 13, 26) {real, imag} */,
  {32'h3e372d59, 32'hbc158864} /* (25, 13, 25) {real, imag} */,
  {32'hbdb37f07, 32'h3b22ae10} /* (25, 13, 24) {real, imag} */,
  {32'h3d835ec8, 32'hbc9e5c84} /* (25, 13, 23) {real, imag} */,
  {32'hbcec4022, 32'h3c175e3a} /* (25, 13, 22) {real, imag} */,
  {32'hbd8d2db4, 32'h3da7ebe0} /* (25, 13, 21) {real, imag} */,
  {32'hbd4002bc, 32'h3c3c255a} /* (25, 13, 20) {real, imag} */,
  {32'h3d828db8, 32'h3cb5c198} /* (25, 13, 19) {real, imag} */,
  {32'h3c770f60, 32'h3ac814f8} /* (25, 13, 18) {real, imag} */,
  {32'h3d3cb420, 32'hbc963679} /* (25, 13, 17) {real, imag} */,
  {32'h3c6d9748, 32'h00000000} /* (25, 13, 16) {real, imag} */,
  {32'h3d3cb420, 32'h3c963679} /* (25, 13, 15) {real, imag} */,
  {32'h3c770f60, 32'hbac814f8} /* (25, 13, 14) {real, imag} */,
  {32'h3d828db8, 32'hbcb5c198} /* (25, 13, 13) {real, imag} */,
  {32'hbd4002bc, 32'hbc3c255a} /* (25, 13, 12) {real, imag} */,
  {32'hbd8d2db4, 32'hbda7ebe0} /* (25, 13, 11) {real, imag} */,
  {32'hbcec4022, 32'hbc175e3a} /* (25, 13, 10) {real, imag} */,
  {32'h3d835ec8, 32'h3c9e5c84} /* (25, 13, 9) {real, imag} */,
  {32'hbdb37f07, 32'hbb22ae10} /* (25, 13, 8) {real, imag} */,
  {32'h3e372d59, 32'h3c158864} /* (25, 13, 7) {real, imag} */,
  {32'hbd4888f8, 32'hbc32cc18} /* (25, 13, 6) {real, imag} */,
  {32'hbdc5af9e, 32'h3cb40144} /* (25, 13, 5) {real, imag} */,
  {32'hbcc13210, 32'h3de45b80} /* (25, 13, 4) {real, imag} */,
  {32'hbd50b650, 32'h3c871f1e} /* (25, 13, 3) {real, imag} */,
  {32'hbf4a8096, 32'hbe1f4b84} /* (25, 13, 2) {real, imag} */,
  {32'h3fccf586, 32'hbd1e9b28} /* (25, 13, 1) {real, imag} */,
  {32'h3f89f4cb, 32'h00000000} /* (25, 13, 0) {real, imag} */,
  {32'h3fa7e78d, 32'h3e436ab0} /* (25, 12, 31) {real, imag} */,
  {32'hbf3b368e, 32'hbc1fb568} /* (25, 12, 30) {real, imag} */,
  {32'h3c2f3f78, 32'h3bef3b10} /* (25, 12, 29) {real, imag} */,
  {32'h3e1c49e6, 32'hbe28c93d} /* (25, 12, 28) {real, imag} */,
  {32'hbdfa694a, 32'h3c7c1c70} /* (25, 12, 27) {real, imag} */,
  {32'hb98c2980, 32'hbcab359c} /* (25, 12, 26) {real, imag} */,
  {32'h3d185d2b, 32'h3ceb191a} /* (25, 12, 25) {real, imag} */,
  {32'hbde204b3, 32'h3dff09d0} /* (25, 12, 24) {real, imag} */,
  {32'hbd8eb9ee, 32'hbe1f81a4} /* (25, 12, 23) {real, imag} */,
  {32'hbc479d90, 32'hbb995a40} /* (25, 12, 22) {real, imag} */,
  {32'hbe14f41c, 32'h3dc19ec7} /* (25, 12, 21) {real, imag} */,
  {32'hbd680109, 32'hbcbe5148} /* (25, 12, 20) {real, imag} */,
  {32'h3d005e00, 32'h3cbad49b} /* (25, 12, 19) {real, imag} */,
  {32'hbc27ae64, 32'h3d88c0be} /* (25, 12, 18) {real, imag} */,
  {32'h3cb973c8, 32'hbd79c54a} /* (25, 12, 17) {real, imag} */,
  {32'h3c5b8c04, 32'h00000000} /* (25, 12, 16) {real, imag} */,
  {32'h3cb973c8, 32'h3d79c54a} /* (25, 12, 15) {real, imag} */,
  {32'hbc27ae64, 32'hbd88c0be} /* (25, 12, 14) {real, imag} */,
  {32'h3d005e00, 32'hbcbad49b} /* (25, 12, 13) {real, imag} */,
  {32'hbd680109, 32'h3cbe5148} /* (25, 12, 12) {real, imag} */,
  {32'hbe14f41c, 32'hbdc19ec7} /* (25, 12, 11) {real, imag} */,
  {32'hbc479d90, 32'h3b995a40} /* (25, 12, 10) {real, imag} */,
  {32'hbd8eb9ee, 32'h3e1f81a4} /* (25, 12, 9) {real, imag} */,
  {32'hbde204b3, 32'hbdff09d0} /* (25, 12, 8) {real, imag} */,
  {32'h3d185d2b, 32'hbceb191a} /* (25, 12, 7) {real, imag} */,
  {32'hb98c2980, 32'h3cab359c} /* (25, 12, 6) {real, imag} */,
  {32'hbdfa694a, 32'hbc7c1c70} /* (25, 12, 5) {real, imag} */,
  {32'h3e1c49e6, 32'h3e28c93d} /* (25, 12, 4) {real, imag} */,
  {32'h3c2f3f78, 32'hbbef3b10} /* (25, 12, 3) {real, imag} */,
  {32'hbf3b368e, 32'h3c1fb568} /* (25, 12, 2) {real, imag} */,
  {32'h3fa7e78d, 32'hbe436ab0} /* (25, 12, 1) {real, imag} */,
  {32'h3f3eb545, 32'h00000000} /* (25, 12, 0) {real, imag} */,
  {32'h3f3c549e, 32'h3e9e96ea} /* (25, 11, 31) {real, imag} */,
  {32'hbf10c71c, 32'h3d223f60} /* (25, 11, 30) {real, imag} */,
  {32'hbc1180fd, 32'h3b983020} /* (25, 11, 29) {real, imag} */,
  {32'h3e8af096, 32'hbe89c1f2} /* (25, 11, 28) {real, imag} */,
  {32'hbcf6d574, 32'h3e339d82} /* (25, 11, 27) {real, imag} */,
  {32'hbd09918d, 32'h3c866608} /* (25, 11, 26) {real, imag} */,
  {32'hb91f8100, 32'h3d2ac431} /* (25, 11, 25) {real, imag} */,
  {32'h3d14c1b9, 32'hbbd379a0} /* (25, 11, 24) {real, imag} */,
  {32'hbcc421ae, 32'h3d2fd960} /* (25, 11, 23) {real, imag} */,
  {32'h3d7b6bfc, 32'hbc0b2655} /* (25, 11, 22) {real, imag} */,
  {32'hbde071c4, 32'h3d6be768} /* (25, 11, 21) {real, imag} */,
  {32'h3ca94470, 32'h3ce559df} /* (25, 11, 20) {real, imag} */,
  {32'hbb0f15f8, 32'hbbf5c470} /* (25, 11, 19) {real, imag} */,
  {32'h3c475a60, 32'h3d6036f2} /* (25, 11, 18) {real, imag} */,
  {32'hbc7306d0, 32'h3c93e3ab} /* (25, 11, 17) {real, imag} */,
  {32'h3cd79996, 32'h00000000} /* (25, 11, 16) {real, imag} */,
  {32'hbc7306d0, 32'hbc93e3ab} /* (25, 11, 15) {real, imag} */,
  {32'h3c475a60, 32'hbd6036f2} /* (25, 11, 14) {real, imag} */,
  {32'hbb0f15f8, 32'h3bf5c470} /* (25, 11, 13) {real, imag} */,
  {32'h3ca94470, 32'hbce559df} /* (25, 11, 12) {real, imag} */,
  {32'hbde071c4, 32'hbd6be768} /* (25, 11, 11) {real, imag} */,
  {32'h3d7b6bfc, 32'h3c0b2655} /* (25, 11, 10) {real, imag} */,
  {32'hbcc421ae, 32'hbd2fd960} /* (25, 11, 9) {real, imag} */,
  {32'h3d14c1b9, 32'h3bd379a0} /* (25, 11, 8) {real, imag} */,
  {32'hb91f8100, 32'hbd2ac431} /* (25, 11, 7) {real, imag} */,
  {32'hbd09918d, 32'hbc866608} /* (25, 11, 6) {real, imag} */,
  {32'hbcf6d574, 32'hbe339d82} /* (25, 11, 5) {real, imag} */,
  {32'h3e8af096, 32'h3e89c1f2} /* (25, 11, 4) {real, imag} */,
  {32'hbc1180fd, 32'hbb983020} /* (25, 11, 3) {real, imag} */,
  {32'hbf10c71c, 32'hbd223f60} /* (25, 11, 2) {real, imag} */,
  {32'h3f3c549e, 32'hbe9e96ea} /* (25, 11, 1) {real, imag} */,
  {32'h3ec542d2, 32'h00000000} /* (25, 11, 0) {real, imag} */,
  {32'hbf050f12, 32'h3f0d852c} /* (25, 10, 31) {real, imag} */,
  {32'hbd1ac590, 32'h3c8b4054} /* (25, 10, 30) {real, imag} */,
  {32'hbd158c3e, 32'hbe01748c} /* (25, 10, 29) {real, imag} */,
  {32'h3df7fc51, 32'hbd91609c} /* (25, 10, 28) {real, imag} */,
  {32'hbc7e5f60, 32'hbdd8d3f0} /* (25, 10, 27) {real, imag} */,
  {32'h3d12ec60, 32'h3cd21759} /* (25, 10, 26) {real, imag} */,
  {32'hbd8aef2e, 32'h3c610924} /* (25, 10, 25) {real, imag} */,
  {32'hbc94d028, 32'hbe3b3eae} /* (25, 10, 24) {real, imag} */,
  {32'h3c2d6b36, 32'hbdbffa63} /* (25, 10, 23) {real, imag} */,
  {32'hbd869e3f, 32'h3d6899d4} /* (25, 10, 22) {real, imag} */,
  {32'hbd972fca, 32'hbd46f238} /* (25, 10, 21) {real, imag} */,
  {32'hbcbd8b9e, 32'hbc5d378f} /* (25, 10, 20) {real, imag} */,
  {32'h3d3eb314, 32'hbdf1c8a8} /* (25, 10, 19) {real, imag} */,
  {32'h3ca14ed0, 32'h3cc23868} /* (25, 10, 18) {real, imag} */,
  {32'h3da0f19d, 32'h3dc03a50} /* (25, 10, 17) {real, imag} */,
  {32'hbd1bbc51, 32'h00000000} /* (25, 10, 16) {real, imag} */,
  {32'h3da0f19d, 32'hbdc03a50} /* (25, 10, 15) {real, imag} */,
  {32'h3ca14ed0, 32'hbcc23868} /* (25, 10, 14) {real, imag} */,
  {32'h3d3eb314, 32'h3df1c8a8} /* (25, 10, 13) {real, imag} */,
  {32'hbcbd8b9e, 32'h3c5d378f} /* (25, 10, 12) {real, imag} */,
  {32'hbd972fca, 32'h3d46f238} /* (25, 10, 11) {real, imag} */,
  {32'hbd869e3f, 32'hbd6899d4} /* (25, 10, 10) {real, imag} */,
  {32'h3c2d6b36, 32'h3dbffa63} /* (25, 10, 9) {real, imag} */,
  {32'hbc94d028, 32'h3e3b3eae} /* (25, 10, 8) {real, imag} */,
  {32'hbd8aef2e, 32'hbc610924} /* (25, 10, 7) {real, imag} */,
  {32'h3d12ec60, 32'hbcd21759} /* (25, 10, 6) {real, imag} */,
  {32'hbc7e5f60, 32'h3dd8d3f0} /* (25, 10, 5) {real, imag} */,
  {32'h3df7fc51, 32'h3d91609c} /* (25, 10, 4) {real, imag} */,
  {32'hbd158c3e, 32'h3e01748c} /* (25, 10, 3) {real, imag} */,
  {32'hbd1ac590, 32'hbc8b4054} /* (25, 10, 2) {real, imag} */,
  {32'hbf050f12, 32'hbf0d852c} /* (25, 10, 1) {real, imag} */,
  {32'hbf14fe9e, 32'h00000000} /* (25, 10, 0) {real, imag} */,
  {32'hbf98875b, 32'h3f2f5b2e} /* (25, 9, 31) {real, imag} */,
  {32'h3e82e2e8, 32'hbdcaa217} /* (25, 9, 30) {real, imag} */,
  {32'h3d4abd54, 32'hbd42ebee} /* (25, 9, 29) {real, imag} */,
  {32'hbcaf85f2, 32'hbd7978bc} /* (25, 9, 28) {real, imag} */,
  {32'h3d7c523f, 32'hbdf47982} /* (25, 9, 27) {real, imag} */,
  {32'hbd634a7e, 32'h39e90100} /* (25, 9, 26) {real, imag} */,
  {32'hbc5361a0, 32'h3d873554} /* (25, 9, 25) {real, imag} */,
  {32'hbca67ca8, 32'hbd82ac54} /* (25, 9, 24) {real, imag} */,
  {32'h3d015b90, 32'hbd57d678} /* (25, 9, 23) {real, imag} */,
  {32'h3d1b822a, 32'hbad82a90} /* (25, 9, 22) {real, imag} */,
  {32'h3d11a99f, 32'hbda9d15b} /* (25, 9, 21) {real, imag} */,
  {32'hbd919826, 32'h3c92eb2a} /* (25, 9, 20) {real, imag} */,
  {32'hbc774cea, 32'h3a2734e0} /* (25, 9, 19) {real, imag} */,
  {32'h3d5e0442, 32'hbcb8783f} /* (25, 9, 18) {real, imag} */,
  {32'hbc9f7720, 32'hbbe5c684} /* (25, 9, 17) {real, imag} */,
  {32'h3d0bfa71, 32'h00000000} /* (25, 9, 16) {real, imag} */,
  {32'hbc9f7720, 32'h3be5c684} /* (25, 9, 15) {real, imag} */,
  {32'h3d5e0442, 32'h3cb8783f} /* (25, 9, 14) {real, imag} */,
  {32'hbc774cea, 32'hba2734e0} /* (25, 9, 13) {real, imag} */,
  {32'hbd919826, 32'hbc92eb2a} /* (25, 9, 12) {real, imag} */,
  {32'h3d11a99f, 32'h3da9d15b} /* (25, 9, 11) {real, imag} */,
  {32'h3d1b822a, 32'h3ad82a90} /* (25, 9, 10) {real, imag} */,
  {32'h3d015b90, 32'h3d57d678} /* (25, 9, 9) {real, imag} */,
  {32'hbca67ca8, 32'h3d82ac54} /* (25, 9, 8) {real, imag} */,
  {32'hbc5361a0, 32'hbd873554} /* (25, 9, 7) {real, imag} */,
  {32'hbd634a7e, 32'hb9e90100} /* (25, 9, 6) {real, imag} */,
  {32'h3d7c523f, 32'h3df47982} /* (25, 9, 5) {real, imag} */,
  {32'hbcaf85f2, 32'h3d7978bc} /* (25, 9, 4) {real, imag} */,
  {32'h3d4abd54, 32'h3d42ebee} /* (25, 9, 3) {real, imag} */,
  {32'h3e82e2e8, 32'h3dcaa217} /* (25, 9, 2) {real, imag} */,
  {32'hbf98875b, 32'hbf2f5b2e} /* (25, 9, 1) {real, imag} */,
  {32'hbfae249c, 32'h00000000} /* (25, 9, 0) {real, imag} */,
  {32'hbfc5deb3, 32'h3f569bae} /* (25, 8, 31) {real, imag} */,
  {32'h3ecbae23, 32'hbe0589df} /* (25, 8, 30) {real, imag} */,
  {32'h3d0200f7, 32'hbcabc3e6} /* (25, 8, 29) {real, imag} */,
  {32'hbda8870e, 32'h3c94deac} /* (25, 8, 28) {real, imag} */,
  {32'h3d01ab4c, 32'hbd5e7e7e} /* (25, 8, 27) {real, imag} */,
  {32'hbd65d837, 32'hbdd7a465} /* (25, 8, 26) {real, imag} */,
  {32'hbc5ee60e, 32'hbd9d5b88} /* (25, 8, 25) {real, imag} */,
  {32'hbb2618e8, 32'hbe1cdbf0} /* (25, 8, 24) {real, imag} */,
  {32'hbd800664, 32'hbcbb48fb} /* (25, 8, 23) {real, imag} */,
  {32'hbd744fcf, 32'h3d00d810} /* (25, 8, 22) {real, imag} */,
  {32'hbc650520, 32'hbba6bff0} /* (25, 8, 21) {real, imag} */,
  {32'hbc514f4a, 32'h3c22fdf0} /* (25, 8, 20) {real, imag} */,
  {32'hbcf60ce2, 32'h3d00f814} /* (25, 8, 19) {real, imag} */,
  {32'h3c214670, 32'hbd0faa91} /* (25, 8, 18) {real, imag} */,
  {32'h3c877030, 32'h3c1cb686} /* (25, 8, 17) {real, imag} */,
  {32'h3c03526c, 32'h00000000} /* (25, 8, 16) {real, imag} */,
  {32'h3c877030, 32'hbc1cb686} /* (25, 8, 15) {real, imag} */,
  {32'h3c214670, 32'h3d0faa91} /* (25, 8, 14) {real, imag} */,
  {32'hbcf60ce2, 32'hbd00f814} /* (25, 8, 13) {real, imag} */,
  {32'hbc514f4a, 32'hbc22fdf0} /* (25, 8, 12) {real, imag} */,
  {32'hbc650520, 32'h3ba6bff0} /* (25, 8, 11) {real, imag} */,
  {32'hbd744fcf, 32'hbd00d810} /* (25, 8, 10) {real, imag} */,
  {32'hbd800664, 32'h3cbb48fb} /* (25, 8, 9) {real, imag} */,
  {32'hbb2618e8, 32'h3e1cdbf0} /* (25, 8, 8) {real, imag} */,
  {32'hbc5ee60e, 32'h3d9d5b88} /* (25, 8, 7) {real, imag} */,
  {32'hbd65d837, 32'h3dd7a465} /* (25, 8, 6) {real, imag} */,
  {32'h3d01ab4c, 32'h3d5e7e7e} /* (25, 8, 5) {real, imag} */,
  {32'hbda8870e, 32'hbc94deac} /* (25, 8, 4) {real, imag} */,
  {32'h3d0200f7, 32'h3cabc3e6} /* (25, 8, 3) {real, imag} */,
  {32'h3ecbae23, 32'h3e0589df} /* (25, 8, 2) {real, imag} */,
  {32'hbfc5deb3, 32'hbf569bae} /* (25, 8, 1) {real, imag} */,
  {32'hbfe9802d, 32'h00000000} /* (25, 8, 0) {real, imag} */,
  {32'hbfe3784e, 32'h3f7daebc} /* (25, 7, 31) {real, imag} */,
  {32'h3ec5b2f8, 32'hbdc26112} /* (25, 7, 30) {real, imag} */,
  {32'h3d973084, 32'hbc92a1dc} /* (25, 7, 29) {real, imag} */,
  {32'hbd4e8af0, 32'h3d11a301} /* (25, 7, 28) {real, imag} */,
  {32'h3e5fc39c, 32'hbdcb5593} /* (25, 7, 27) {real, imag} */,
  {32'h3d1c087c, 32'hbe451a51} /* (25, 7, 26) {real, imag} */,
  {32'hbd6635aa, 32'hbdb036bb} /* (25, 7, 25) {real, imag} */,
  {32'hbd16d29d, 32'hbe2330e9} /* (25, 7, 24) {real, imag} */,
  {32'hbced63e7, 32'hbe1bbf9c} /* (25, 7, 23) {real, imag} */,
  {32'h3d50e09c, 32'h3b3b18e4} /* (25, 7, 22) {real, imag} */,
  {32'h3de43303, 32'h3b0d6e60} /* (25, 7, 21) {real, imag} */,
  {32'h3d33448f, 32'h3d0b72fe} /* (25, 7, 20) {real, imag} */,
  {32'h3c2acb8a, 32'h3cbc40a2} /* (25, 7, 19) {real, imag} */,
  {32'hbd49bf32, 32'hbc816d5d} /* (25, 7, 18) {real, imag} */,
  {32'h3c0b87fc, 32'h3d498bc4} /* (25, 7, 17) {real, imag} */,
  {32'h3b7219b0, 32'h00000000} /* (25, 7, 16) {real, imag} */,
  {32'h3c0b87fc, 32'hbd498bc4} /* (25, 7, 15) {real, imag} */,
  {32'hbd49bf32, 32'h3c816d5d} /* (25, 7, 14) {real, imag} */,
  {32'h3c2acb8a, 32'hbcbc40a2} /* (25, 7, 13) {real, imag} */,
  {32'h3d33448f, 32'hbd0b72fe} /* (25, 7, 12) {real, imag} */,
  {32'h3de43303, 32'hbb0d6e60} /* (25, 7, 11) {real, imag} */,
  {32'h3d50e09c, 32'hbb3b18e4} /* (25, 7, 10) {real, imag} */,
  {32'hbced63e7, 32'h3e1bbf9c} /* (25, 7, 9) {real, imag} */,
  {32'hbd16d29d, 32'h3e2330e9} /* (25, 7, 8) {real, imag} */,
  {32'hbd6635aa, 32'h3db036bb} /* (25, 7, 7) {real, imag} */,
  {32'h3d1c087c, 32'h3e451a51} /* (25, 7, 6) {real, imag} */,
  {32'h3e5fc39c, 32'h3dcb5593} /* (25, 7, 5) {real, imag} */,
  {32'hbd4e8af0, 32'hbd11a301} /* (25, 7, 4) {real, imag} */,
  {32'h3d973084, 32'h3c92a1dc} /* (25, 7, 3) {real, imag} */,
  {32'h3ec5b2f8, 32'h3dc26112} /* (25, 7, 2) {real, imag} */,
  {32'hbfe3784e, 32'hbf7daebc} /* (25, 7, 1) {real, imag} */,
  {32'hc01c7402, 32'h00000000} /* (25, 7, 0) {real, imag} */,
  {32'hbfeeb672, 32'h3f9f19ac} /* (25, 6, 31) {real, imag} */,
  {32'h3e8eabb2, 32'hbe61fde2} /* (25, 6, 30) {real, imag} */,
  {32'h3da760df, 32'h3b1a1018} /* (25, 6, 29) {real, imag} */,
  {32'h3b69d918, 32'hbb46eb78} /* (25, 6, 28) {real, imag} */,
  {32'h3e283f92, 32'h3d36c635} /* (25, 6, 27) {real, imag} */,
  {32'h3b9b52ec, 32'h3d49d98e} /* (25, 6, 26) {real, imag} */,
  {32'hbd26ce22, 32'hbd9a86c2} /* (25, 6, 25) {real, imag} */,
  {32'h3b5c539c, 32'hbd467c5e} /* (25, 6, 24) {real, imag} */,
  {32'hbcad2a3f, 32'h3d44b5dc} /* (25, 6, 23) {real, imag} */,
  {32'hbc921a72, 32'h3d3d6f8a} /* (25, 6, 22) {real, imag} */,
  {32'h3dcd441a, 32'hbd8bdec0} /* (25, 6, 21) {real, imag} */,
  {32'h3cc76219, 32'hbcaba3ac} /* (25, 6, 20) {real, imag} */,
  {32'h3d909947, 32'hbcc8f45d} /* (25, 6, 19) {real, imag} */,
  {32'h3b4d09c8, 32'hbcad2f29} /* (25, 6, 18) {real, imag} */,
  {32'hbd3ed11c, 32'h3d3721cc} /* (25, 6, 17) {real, imag} */,
  {32'h3d35dc02, 32'h00000000} /* (25, 6, 16) {real, imag} */,
  {32'hbd3ed11c, 32'hbd3721cc} /* (25, 6, 15) {real, imag} */,
  {32'h3b4d09c8, 32'h3cad2f29} /* (25, 6, 14) {real, imag} */,
  {32'h3d909947, 32'h3cc8f45d} /* (25, 6, 13) {real, imag} */,
  {32'h3cc76219, 32'h3caba3ac} /* (25, 6, 12) {real, imag} */,
  {32'h3dcd441a, 32'h3d8bdec0} /* (25, 6, 11) {real, imag} */,
  {32'hbc921a72, 32'hbd3d6f8a} /* (25, 6, 10) {real, imag} */,
  {32'hbcad2a3f, 32'hbd44b5dc} /* (25, 6, 9) {real, imag} */,
  {32'h3b5c539c, 32'h3d467c5e} /* (25, 6, 8) {real, imag} */,
  {32'hbd26ce22, 32'h3d9a86c2} /* (25, 6, 7) {real, imag} */,
  {32'h3b9b52ec, 32'hbd49d98e} /* (25, 6, 6) {real, imag} */,
  {32'h3e283f92, 32'hbd36c635} /* (25, 6, 5) {real, imag} */,
  {32'h3b69d918, 32'h3b46eb78} /* (25, 6, 4) {real, imag} */,
  {32'h3da760df, 32'hbb1a1018} /* (25, 6, 3) {real, imag} */,
  {32'h3e8eabb2, 32'h3e61fde2} /* (25, 6, 2) {real, imag} */,
  {32'hbfeeb672, 32'hbf9f19ac} /* (25, 6, 1) {real, imag} */,
  {32'hc021ac05, 32'h00000000} /* (25, 6, 0) {real, imag} */,
  {32'hbff131eb, 32'h3fd0a541} /* (25, 5, 31) {real, imag} */,
  {32'hbce27130, 32'hbe976bb2} /* (25, 5, 30) {real, imag} */,
  {32'h3b77d800, 32'hbcf33cc0} /* (25, 5, 29) {real, imag} */,
  {32'h3daa963d, 32'hbdbdf506} /* (25, 5, 28) {real, imag} */,
  {32'h3debc65c, 32'h3d9bde87} /* (25, 5, 27) {real, imag} */,
  {32'h3c87a070, 32'h3c7f1cc0} /* (25, 5, 26) {real, imag} */,
  {32'hbd16a22c, 32'hbdb7a825} /* (25, 5, 25) {real, imag} */,
  {32'h3d0b701d, 32'hbe36188a} /* (25, 5, 24) {real, imag} */,
  {32'h3c000b34, 32'h3c3bac4c} /* (25, 5, 23) {real, imag} */,
  {32'h3dac66d9, 32'h3ce9f4c2} /* (25, 5, 22) {real, imag} */,
  {32'h3d7b0e97, 32'h3d1dd6fe} /* (25, 5, 21) {real, imag} */,
  {32'hbbacfa2c, 32'hbda78f2d} /* (25, 5, 20) {real, imag} */,
  {32'h3c0963d7, 32'hbd993b99} /* (25, 5, 19) {real, imag} */,
  {32'h3d16fce8, 32'hbde8b816} /* (25, 5, 18) {real, imag} */,
  {32'h3d672e2d, 32'hbd77b9da} /* (25, 5, 17) {real, imag} */,
  {32'h3d575d11, 32'h00000000} /* (25, 5, 16) {real, imag} */,
  {32'h3d672e2d, 32'h3d77b9da} /* (25, 5, 15) {real, imag} */,
  {32'h3d16fce8, 32'h3de8b816} /* (25, 5, 14) {real, imag} */,
  {32'h3c0963d7, 32'h3d993b99} /* (25, 5, 13) {real, imag} */,
  {32'hbbacfa2c, 32'h3da78f2d} /* (25, 5, 12) {real, imag} */,
  {32'h3d7b0e97, 32'hbd1dd6fe} /* (25, 5, 11) {real, imag} */,
  {32'h3dac66d9, 32'hbce9f4c2} /* (25, 5, 10) {real, imag} */,
  {32'h3c000b34, 32'hbc3bac4c} /* (25, 5, 9) {real, imag} */,
  {32'h3d0b701d, 32'h3e36188a} /* (25, 5, 8) {real, imag} */,
  {32'hbd16a22c, 32'h3db7a825} /* (25, 5, 7) {real, imag} */,
  {32'h3c87a070, 32'hbc7f1cc0} /* (25, 5, 6) {real, imag} */,
  {32'h3debc65c, 32'hbd9bde87} /* (25, 5, 5) {real, imag} */,
  {32'h3daa963d, 32'h3dbdf506} /* (25, 5, 4) {real, imag} */,
  {32'h3b77d800, 32'h3cf33cc0} /* (25, 5, 3) {real, imag} */,
  {32'hbce27130, 32'h3e976bb2} /* (25, 5, 2) {real, imag} */,
  {32'hbff131eb, 32'hbfd0a541} /* (25, 5, 1) {real, imag} */,
  {32'hc0367f94, 32'h00000000} /* (25, 5, 0) {real, imag} */,
  {32'hbfd67225, 32'h400015eb} /* (25, 4, 31) {real, imag} */,
  {32'hbe33cd4a, 32'hbe86a0c4} /* (25, 4, 30) {real, imag} */,
  {32'h3e033608, 32'hbbcf0a50} /* (25, 4, 29) {real, imag} */,
  {32'h3dfc3fbc, 32'hbe144d43} /* (25, 4, 28) {real, imag} */,
  {32'h3e1a9f0f, 32'h3e09386d} /* (25, 4, 27) {real, imag} */,
  {32'h3ca0118a, 32'hbc4871ec} /* (25, 4, 26) {real, imag} */,
  {32'hbda9a06e, 32'h3cbb1912} /* (25, 4, 25) {real, imag} */,
  {32'hbd947c3f, 32'hbd38f019} /* (25, 4, 24) {real, imag} */,
  {32'h3dbe22d4, 32'h3d3f2f7e} /* (25, 4, 23) {real, imag} */,
  {32'h3a5bc280, 32'hbd9b7cf2} /* (25, 4, 22) {real, imag} */,
  {32'h3db36841, 32'hbd5f618f} /* (25, 4, 21) {real, imag} */,
  {32'hbbe140b8, 32'h3d06e078} /* (25, 4, 20) {real, imag} */,
  {32'hbcff360c, 32'h3d9b41be} /* (25, 4, 19) {real, imag} */,
  {32'hbdeb0c5a, 32'h3d2d0a7c} /* (25, 4, 18) {real, imag} */,
  {32'h3c6866e8, 32'h3cefe3db} /* (25, 4, 17) {real, imag} */,
  {32'h3cade03e, 32'h00000000} /* (25, 4, 16) {real, imag} */,
  {32'h3c6866e8, 32'hbcefe3db} /* (25, 4, 15) {real, imag} */,
  {32'hbdeb0c5a, 32'hbd2d0a7c} /* (25, 4, 14) {real, imag} */,
  {32'hbcff360c, 32'hbd9b41be} /* (25, 4, 13) {real, imag} */,
  {32'hbbe140b8, 32'hbd06e078} /* (25, 4, 12) {real, imag} */,
  {32'h3db36841, 32'h3d5f618f} /* (25, 4, 11) {real, imag} */,
  {32'h3a5bc280, 32'h3d9b7cf2} /* (25, 4, 10) {real, imag} */,
  {32'h3dbe22d4, 32'hbd3f2f7e} /* (25, 4, 9) {real, imag} */,
  {32'hbd947c3f, 32'h3d38f019} /* (25, 4, 8) {real, imag} */,
  {32'hbda9a06e, 32'hbcbb1912} /* (25, 4, 7) {real, imag} */,
  {32'h3ca0118a, 32'h3c4871ec} /* (25, 4, 6) {real, imag} */,
  {32'h3e1a9f0f, 32'hbe09386d} /* (25, 4, 5) {real, imag} */,
  {32'h3dfc3fbc, 32'h3e144d43} /* (25, 4, 4) {real, imag} */,
  {32'h3e033608, 32'h3bcf0a50} /* (25, 4, 3) {real, imag} */,
  {32'hbe33cd4a, 32'h3e86a0c4} /* (25, 4, 2) {real, imag} */,
  {32'hbfd67225, 32'hc00015eb} /* (25, 4, 1) {real, imag} */,
  {32'hc038b4a2, 32'h00000000} /* (25, 4, 0) {real, imag} */,
  {32'hbfe5f6e4, 32'h400a7f74} /* (25, 3, 31) {real, imag} */,
  {32'hbe82f857, 32'hbeb25250} /* (25, 3, 30) {real, imag} */,
  {32'h3e3f5137, 32'hbd96e75c} /* (25, 3, 29) {real, imag} */,
  {32'h3e07d455, 32'hbe343270} /* (25, 3, 28) {real, imag} */,
  {32'h3e653f7f, 32'hbcae7124} /* (25, 3, 27) {real, imag} */,
  {32'hbdc376df, 32'h3dab3066} /* (25, 3, 26) {real, imag} */,
  {32'hbda8a110, 32'hbcfb6c40} /* (25, 3, 25) {real, imag} */,
  {32'hbe437486, 32'hbc9d43b8} /* (25, 3, 24) {real, imag} */,
  {32'h3df60d9a, 32'hbcd2a4d4} /* (25, 3, 23) {real, imag} */,
  {32'hbc0a3668, 32'hbc3e552e} /* (25, 3, 22) {real, imag} */,
  {32'hbc8f1cce, 32'hbd3a3daf} /* (25, 3, 21) {real, imag} */,
  {32'h3d21dcaa, 32'hbddd5fe5} /* (25, 3, 20) {real, imag} */,
  {32'hbae2736c, 32'h3da58d88} /* (25, 3, 19) {real, imag} */,
  {32'hbbc932fc, 32'hbcdb000c} /* (25, 3, 18) {real, imag} */,
  {32'h3d497c6c, 32'h3d35188e} /* (25, 3, 17) {real, imag} */,
  {32'hbda0c2dc, 32'h00000000} /* (25, 3, 16) {real, imag} */,
  {32'h3d497c6c, 32'hbd35188e} /* (25, 3, 15) {real, imag} */,
  {32'hbbc932fc, 32'h3cdb000c} /* (25, 3, 14) {real, imag} */,
  {32'hbae2736c, 32'hbda58d88} /* (25, 3, 13) {real, imag} */,
  {32'h3d21dcaa, 32'h3ddd5fe5} /* (25, 3, 12) {real, imag} */,
  {32'hbc8f1cce, 32'h3d3a3daf} /* (25, 3, 11) {real, imag} */,
  {32'hbc0a3668, 32'h3c3e552e} /* (25, 3, 10) {real, imag} */,
  {32'h3df60d9a, 32'h3cd2a4d4} /* (25, 3, 9) {real, imag} */,
  {32'hbe437486, 32'h3c9d43b8} /* (25, 3, 8) {real, imag} */,
  {32'hbda8a110, 32'h3cfb6c40} /* (25, 3, 7) {real, imag} */,
  {32'hbdc376df, 32'hbdab3066} /* (25, 3, 6) {real, imag} */,
  {32'h3e653f7f, 32'h3cae7124} /* (25, 3, 5) {real, imag} */,
  {32'h3e07d455, 32'h3e343270} /* (25, 3, 4) {real, imag} */,
  {32'h3e3f5137, 32'h3d96e75c} /* (25, 3, 3) {real, imag} */,
  {32'hbe82f857, 32'h3eb25250} /* (25, 3, 2) {real, imag} */,
  {32'hbfe5f6e4, 32'hc00a7f74} /* (25, 3, 1) {real, imag} */,
  {32'hc0410144, 32'h00000000} /* (25, 3, 0) {real, imag} */,
  {32'hbfef53e8, 32'h40055565} /* (25, 2, 31) {real, imag} */,
  {32'hbe462532, 32'hbec65ede} /* (25, 2, 30) {real, imag} */,
  {32'h3ded09d0, 32'h3cb81324} /* (25, 2, 29) {real, imag} */,
  {32'h3e79712a, 32'hbe437902} /* (25, 2, 28) {real, imag} */,
  {32'h3e58bf9c, 32'hbbd9e1b4} /* (25, 2, 27) {real, imag} */,
  {32'h3d196829, 32'h3d1bbbcc} /* (25, 2, 26) {real, imag} */,
  {32'hbdfa8466, 32'h3d109b08} /* (25, 2, 25) {real, imag} */,
  {32'hbde3c692, 32'hbc5f2380} /* (25, 2, 24) {real, imag} */,
  {32'hbd1e6b4b, 32'hbc5967a4} /* (25, 2, 23) {real, imag} */,
  {32'h3df9a972, 32'hbe1e97ae} /* (25, 2, 22) {real, imag} */,
  {32'h3d87fb57, 32'h3d40e662} /* (25, 2, 21) {real, imag} */,
  {32'hbc82c281, 32'h3d7c336c} /* (25, 2, 20) {real, imag} */,
  {32'hbd4e7b53, 32'hbdb067c7} /* (25, 2, 19) {real, imag} */,
  {32'hbc88f25e, 32'hbc01bfd0} /* (25, 2, 18) {real, imag} */,
  {32'h3cc70b97, 32'hbc832c2f} /* (25, 2, 17) {real, imag} */,
  {32'hbd743cd0, 32'h00000000} /* (25, 2, 16) {real, imag} */,
  {32'h3cc70b97, 32'h3c832c2f} /* (25, 2, 15) {real, imag} */,
  {32'hbc88f25e, 32'h3c01bfd0} /* (25, 2, 14) {real, imag} */,
  {32'hbd4e7b53, 32'h3db067c7} /* (25, 2, 13) {real, imag} */,
  {32'hbc82c281, 32'hbd7c336c} /* (25, 2, 12) {real, imag} */,
  {32'h3d87fb57, 32'hbd40e662} /* (25, 2, 11) {real, imag} */,
  {32'h3df9a972, 32'h3e1e97ae} /* (25, 2, 10) {real, imag} */,
  {32'hbd1e6b4b, 32'h3c5967a4} /* (25, 2, 9) {real, imag} */,
  {32'hbde3c692, 32'h3c5f2380} /* (25, 2, 8) {real, imag} */,
  {32'hbdfa8466, 32'hbd109b08} /* (25, 2, 7) {real, imag} */,
  {32'h3d196829, 32'hbd1bbbcc} /* (25, 2, 6) {real, imag} */,
  {32'h3e58bf9c, 32'h3bd9e1b4} /* (25, 2, 5) {real, imag} */,
  {32'h3e79712a, 32'h3e437902} /* (25, 2, 4) {real, imag} */,
  {32'h3ded09d0, 32'hbcb81324} /* (25, 2, 3) {real, imag} */,
  {32'hbe462532, 32'h3ec65ede} /* (25, 2, 2) {real, imag} */,
  {32'hbfef53e8, 32'hc0055565} /* (25, 2, 1) {real, imag} */,
  {32'hc03aac66, 32'h00000000} /* (25, 2, 0) {real, imag} */,
  {32'hbfe4754a, 32'h3feb03be} /* (25, 1, 31) {real, imag} */,
  {32'hbdec5592, 32'hbe8d8dc2} /* (25, 1, 30) {real, imag} */,
  {32'h3e3f3ac8, 32'h3c8cc148} /* (25, 1, 29) {real, imag} */,
  {32'h3e3c6478, 32'hbdaf5062} /* (25, 1, 28) {real, imag} */,
  {32'h3d981e3e, 32'h3c9d3295} /* (25, 1, 27) {real, imag} */,
  {32'hbd64dff7, 32'hbd7d0008} /* (25, 1, 26) {real, imag} */,
  {32'h3d5bf5d2, 32'h3dd18242} /* (25, 1, 25) {real, imag} */,
  {32'hbda9907f, 32'hbd966ddc} /* (25, 1, 24) {real, imag} */,
  {32'h3d93138e, 32'h3dc3de0b} /* (25, 1, 23) {real, imag} */,
  {32'hbd3da8d5, 32'hbc4fd245} /* (25, 1, 22) {real, imag} */,
  {32'h3d9f2295, 32'hbda34f16} /* (25, 1, 21) {real, imag} */,
  {32'hbc873248, 32'h3c8c8ea0} /* (25, 1, 20) {real, imag} */,
  {32'h3daad471, 32'hbd13b165} /* (25, 1, 19) {real, imag} */,
  {32'hbd9606cd, 32'hbda3de5d} /* (25, 1, 18) {real, imag} */,
  {32'hbdd61a1e, 32'hbb9c69fd} /* (25, 1, 17) {real, imag} */,
  {32'h3bab7418, 32'h00000000} /* (25, 1, 16) {real, imag} */,
  {32'hbdd61a1e, 32'h3b9c69fd} /* (25, 1, 15) {real, imag} */,
  {32'hbd9606cd, 32'h3da3de5d} /* (25, 1, 14) {real, imag} */,
  {32'h3daad471, 32'h3d13b165} /* (25, 1, 13) {real, imag} */,
  {32'hbc873248, 32'hbc8c8ea0} /* (25, 1, 12) {real, imag} */,
  {32'h3d9f2295, 32'h3da34f16} /* (25, 1, 11) {real, imag} */,
  {32'hbd3da8d5, 32'h3c4fd245} /* (25, 1, 10) {real, imag} */,
  {32'h3d93138e, 32'hbdc3de0b} /* (25, 1, 9) {real, imag} */,
  {32'hbda9907f, 32'h3d966ddc} /* (25, 1, 8) {real, imag} */,
  {32'h3d5bf5d2, 32'hbdd18242} /* (25, 1, 7) {real, imag} */,
  {32'hbd64dff7, 32'h3d7d0008} /* (25, 1, 6) {real, imag} */,
  {32'h3d981e3e, 32'hbc9d3295} /* (25, 1, 5) {real, imag} */,
  {32'h3e3c6478, 32'h3daf5062} /* (25, 1, 4) {real, imag} */,
  {32'h3e3f3ac8, 32'hbc8cc148} /* (25, 1, 3) {real, imag} */,
  {32'hbdec5592, 32'h3e8d8dc2} /* (25, 1, 2) {real, imag} */,
  {32'hbfe4754a, 32'hbfeb03be} /* (25, 1, 1) {real, imag} */,
  {32'hc043edb7, 32'h00000000} /* (25, 1, 0) {real, imag} */,
  {32'hbfee5faf, 32'h3fb34140} /* (25, 0, 31) {real, imag} */,
  {32'h3d849714, 32'hbe2c8d2d} /* (25, 0, 30) {real, imag} */,
  {32'h3dd944ce, 32'hbd8f699c} /* (25, 0, 29) {real, imag} */,
  {32'h3d4c616f, 32'hbdcbb264} /* (25, 0, 28) {real, imag} */,
  {32'h3dc7db05, 32'hbdae9e5c} /* (25, 0, 27) {real, imag} */,
  {32'hbcde39ce, 32'hbcf9812c} /* (25, 0, 26) {real, imag} */,
  {32'h3ba3b3a2, 32'h3ce20e5e} /* (25, 0, 25) {real, imag} */,
  {32'h3d6c90ec, 32'hbd32bdd1} /* (25, 0, 24) {real, imag} */,
  {32'h3d25d5dc, 32'h3b934a68} /* (25, 0, 23) {real, imag} */,
  {32'h3d430a5e, 32'h3ae9b800} /* (25, 0, 22) {real, imag} */,
  {32'h3bf91300, 32'h3ced8f0e} /* (25, 0, 21) {real, imag} */,
  {32'h3cfe72a5, 32'h3c50f398} /* (25, 0, 20) {real, imag} */,
  {32'h3d16a5e4, 32'h3d29477a} /* (25, 0, 19) {real, imag} */,
  {32'h3d373990, 32'h3c286952} /* (25, 0, 18) {real, imag} */,
  {32'hbc1fe97c, 32'hbcb564d8} /* (25, 0, 17) {real, imag} */,
  {32'h3c0a4638, 32'h00000000} /* (25, 0, 16) {real, imag} */,
  {32'hbc1fe97c, 32'h3cb564d8} /* (25, 0, 15) {real, imag} */,
  {32'h3d373990, 32'hbc286952} /* (25, 0, 14) {real, imag} */,
  {32'h3d16a5e4, 32'hbd29477a} /* (25, 0, 13) {real, imag} */,
  {32'h3cfe72a5, 32'hbc50f398} /* (25, 0, 12) {real, imag} */,
  {32'h3bf91300, 32'hbced8f0e} /* (25, 0, 11) {real, imag} */,
  {32'h3d430a5e, 32'hbae9b800} /* (25, 0, 10) {real, imag} */,
  {32'h3d25d5dc, 32'hbb934a68} /* (25, 0, 9) {real, imag} */,
  {32'h3d6c90ec, 32'h3d32bdd1} /* (25, 0, 8) {real, imag} */,
  {32'h3ba3b3a2, 32'hbce20e5e} /* (25, 0, 7) {real, imag} */,
  {32'hbcde39ce, 32'h3cf9812c} /* (25, 0, 6) {real, imag} */,
  {32'h3dc7db05, 32'h3dae9e5c} /* (25, 0, 5) {real, imag} */,
  {32'h3d4c616f, 32'h3dcbb264} /* (25, 0, 4) {real, imag} */,
  {32'h3dd944ce, 32'h3d8f699c} /* (25, 0, 3) {real, imag} */,
  {32'h3d849714, 32'h3e2c8d2d} /* (25, 0, 2) {real, imag} */,
  {32'hbfee5faf, 32'hbfb34140} /* (25, 0, 1) {real, imag} */,
  {32'hc03f26a0, 32'h00000000} /* (25, 0, 0) {real, imag} */,
  {32'hc03fc377, 32'h3fd32d0c} /* (24, 31, 31) {real, imag} */,
  {32'h3f14a04e, 32'hbe1e99e5} /* (24, 31, 30) {real, imag} */,
  {32'h3d9f7337, 32'hb9982ea0} /* (24, 31, 29) {real, imag} */,
  {32'hbd14feee, 32'h3baa92a0} /* (24, 31, 28) {real, imag} */,
  {32'h3e306db6, 32'hbd1f25e4} /* (24, 31, 27) {real, imag} */,
  {32'hbd85f85e, 32'hbc925e98} /* (24, 31, 26) {real, imag} */,
  {32'hbd442882, 32'h3c0d6210} /* (24, 31, 25) {real, imag} */,
  {32'h3d7eb2e6, 32'hbd994b8e} /* (24, 31, 24) {real, imag} */,
  {32'h3cc1bb11, 32'h3cc563f5} /* (24, 31, 23) {real, imag} */,
  {32'h3db8033a, 32'hbcc8be61} /* (24, 31, 22) {real, imag} */,
  {32'h3c6771cb, 32'hbd54c01e} /* (24, 31, 21) {real, imag} */,
  {32'hbd22fa68, 32'h3ad6c000} /* (24, 31, 20) {real, imag} */,
  {32'hbdb51c7a, 32'hbd12b79f} /* (24, 31, 19) {real, imag} */,
  {32'h3d81f771, 32'h3cceadaa} /* (24, 31, 18) {real, imag} */,
  {32'h3cf35b58, 32'h3d307912} /* (24, 31, 17) {real, imag} */,
  {32'hbd71e948, 32'h00000000} /* (24, 31, 16) {real, imag} */,
  {32'h3cf35b58, 32'hbd307912} /* (24, 31, 15) {real, imag} */,
  {32'h3d81f771, 32'hbcceadaa} /* (24, 31, 14) {real, imag} */,
  {32'hbdb51c7a, 32'h3d12b79f} /* (24, 31, 13) {real, imag} */,
  {32'hbd22fa68, 32'hbad6c000} /* (24, 31, 12) {real, imag} */,
  {32'h3c6771cb, 32'h3d54c01e} /* (24, 31, 11) {real, imag} */,
  {32'h3db8033a, 32'h3cc8be61} /* (24, 31, 10) {real, imag} */,
  {32'h3cc1bb11, 32'hbcc563f5} /* (24, 31, 9) {real, imag} */,
  {32'h3d7eb2e6, 32'h3d994b8e} /* (24, 31, 8) {real, imag} */,
  {32'hbd442882, 32'hbc0d6210} /* (24, 31, 7) {real, imag} */,
  {32'hbd85f85e, 32'h3c925e98} /* (24, 31, 6) {real, imag} */,
  {32'h3e306db6, 32'h3d1f25e4} /* (24, 31, 5) {real, imag} */,
  {32'hbd14feee, 32'hbbaa92a0} /* (24, 31, 4) {real, imag} */,
  {32'h3d9f7337, 32'h39982ea0} /* (24, 31, 3) {real, imag} */,
  {32'h3f14a04e, 32'h3e1e99e5} /* (24, 31, 2) {real, imag} */,
  {32'hc03fc377, 32'hbfd32d0c} /* (24, 31, 1) {real, imag} */,
  {32'hc08502ae, 32'h00000000} /* (24, 31, 0) {real, imag} */,
  {32'hc05bd0bd, 32'h3fae15cc} /* (24, 30, 31) {real, imag} */,
  {32'h3f70354b, 32'hbe54e104} /* (24, 30, 30) {real, imag} */,
  {32'h3dc57a62, 32'hbcde4250} /* (24, 30, 29) {real, imag} */,
  {32'hbdc3dd1c, 32'h3dec1666} /* (24, 30, 28) {real, imag} */,
  {32'h3e255736, 32'hbdfe7f18} /* (24, 30, 27) {real, imag} */,
  {32'h3c468c2c, 32'h3b6a0898} /* (24, 30, 26) {real, imag} */,
  {32'hbd16560d, 32'h3d89df1b} /* (24, 30, 25) {real, imag} */,
  {32'h3ddb5479, 32'hbd601416} /* (24, 30, 24) {real, imag} */,
  {32'h3ca2099d, 32'hbc8a4342} /* (24, 30, 23) {real, imag} */,
  {32'hbd2e486c, 32'h3debd3e8} /* (24, 30, 22) {real, imag} */,
  {32'h3dcc9068, 32'hbd858edc} /* (24, 30, 21) {real, imag} */,
  {32'hbd774e6c, 32'hbd1a9b30} /* (24, 30, 20) {real, imag} */,
  {32'hbdd578e5, 32'hbd068806} /* (24, 30, 19) {real, imag} */,
  {32'h3d63c3c7, 32'hbceadc94} /* (24, 30, 18) {real, imag} */,
  {32'hbbcb6ba8, 32'h3d68b330} /* (24, 30, 17) {real, imag} */,
  {32'h3c460f00, 32'h00000000} /* (24, 30, 16) {real, imag} */,
  {32'hbbcb6ba8, 32'hbd68b330} /* (24, 30, 15) {real, imag} */,
  {32'h3d63c3c7, 32'h3ceadc94} /* (24, 30, 14) {real, imag} */,
  {32'hbdd578e5, 32'h3d068806} /* (24, 30, 13) {real, imag} */,
  {32'hbd774e6c, 32'h3d1a9b30} /* (24, 30, 12) {real, imag} */,
  {32'h3dcc9068, 32'h3d858edc} /* (24, 30, 11) {real, imag} */,
  {32'hbd2e486c, 32'hbdebd3e8} /* (24, 30, 10) {real, imag} */,
  {32'h3ca2099d, 32'h3c8a4342} /* (24, 30, 9) {real, imag} */,
  {32'h3ddb5479, 32'h3d601416} /* (24, 30, 8) {real, imag} */,
  {32'hbd16560d, 32'hbd89df1b} /* (24, 30, 7) {real, imag} */,
  {32'h3c468c2c, 32'hbb6a0898} /* (24, 30, 6) {real, imag} */,
  {32'h3e255736, 32'h3dfe7f18} /* (24, 30, 5) {real, imag} */,
  {32'hbdc3dd1c, 32'hbdec1666} /* (24, 30, 4) {real, imag} */,
  {32'h3dc57a62, 32'h3cde4250} /* (24, 30, 3) {real, imag} */,
  {32'h3f70354b, 32'h3e54e104} /* (24, 30, 2) {real, imag} */,
  {32'hc05bd0bd, 32'hbfae15cc} /* (24, 30, 1) {real, imag} */,
  {32'hc085ed5b, 32'h00000000} /* (24, 30, 0) {real, imag} */,
  {32'hc06818bc, 32'h3f9ceaea} /* (24, 29, 31) {real, imag} */,
  {32'h3f80848d, 32'hbdfa18dc} /* (24, 29, 30) {real, imag} */,
  {32'h3d384fc8, 32'h3c2a08f8} /* (24, 29, 29) {real, imag} */,
  {32'hbe66caf7, 32'h3d86c01e} /* (24, 29, 28) {real, imag} */,
  {32'h3db88df0, 32'hbe107f8a} /* (24, 29, 27) {real, imag} */,
  {32'h3e103b84, 32'hbcaf3726} /* (24, 29, 26) {real, imag} */,
  {32'h3e0e0da0, 32'h3cd7b064} /* (24, 29, 25) {real, imag} */,
  {32'h3dd0c745, 32'h3bb220b8} /* (24, 29, 24) {real, imag} */,
  {32'hbd5e33f3, 32'hbc9917b5} /* (24, 29, 23) {real, imag} */,
  {32'hbd2b9519, 32'h3c3e5978} /* (24, 29, 22) {real, imag} */,
  {32'h3d543325, 32'h3c531621} /* (24, 29, 21) {real, imag} */,
  {32'hbdb71993, 32'hbcb577e5} /* (24, 29, 20) {real, imag} */,
  {32'hbd984f11, 32'hbd2ed8b4} /* (24, 29, 19) {real, imag} */,
  {32'hbcfd19d8, 32'hbd1bc49d} /* (24, 29, 18) {real, imag} */,
  {32'hbc5335f2, 32'hbd45adba} /* (24, 29, 17) {real, imag} */,
  {32'h3de0d8df, 32'h00000000} /* (24, 29, 16) {real, imag} */,
  {32'hbc5335f2, 32'h3d45adba} /* (24, 29, 15) {real, imag} */,
  {32'hbcfd19d8, 32'h3d1bc49d} /* (24, 29, 14) {real, imag} */,
  {32'hbd984f11, 32'h3d2ed8b4} /* (24, 29, 13) {real, imag} */,
  {32'hbdb71993, 32'h3cb577e5} /* (24, 29, 12) {real, imag} */,
  {32'h3d543325, 32'hbc531621} /* (24, 29, 11) {real, imag} */,
  {32'hbd2b9519, 32'hbc3e5978} /* (24, 29, 10) {real, imag} */,
  {32'hbd5e33f3, 32'h3c9917b5} /* (24, 29, 9) {real, imag} */,
  {32'h3dd0c745, 32'hbbb220b8} /* (24, 29, 8) {real, imag} */,
  {32'h3e0e0da0, 32'hbcd7b064} /* (24, 29, 7) {real, imag} */,
  {32'h3e103b84, 32'h3caf3726} /* (24, 29, 6) {real, imag} */,
  {32'h3db88df0, 32'h3e107f8a} /* (24, 29, 5) {real, imag} */,
  {32'hbe66caf7, 32'hbd86c01e} /* (24, 29, 4) {real, imag} */,
  {32'h3d384fc8, 32'hbc2a08f8} /* (24, 29, 3) {real, imag} */,
  {32'h3f80848d, 32'h3dfa18dc} /* (24, 29, 2) {real, imag} */,
  {32'hc06818bc, 32'hbf9ceaea} /* (24, 29, 1) {real, imag} */,
  {32'hc0888115, 32'h00000000} /* (24, 29, 0) {real, imag} */,
  {32'hc075f335, 32'h3f8a97c2} /* (24, 28, 31) {real, imag} */,
  {32'h3f9414e1, 32'hbe2e60a8} /* (24, 28, 30) {real, imag} */,
  {32'hbde7b16e, 32'hbd29454c} /* (24, 28, 29) {real, imag} */,
  {32'hbe10fe04, 32'h3dc53e8a} /* (24, 28, 28) {real, imag} */,
  {32'h3e1b55f1, 32'hbe5d9435} /* (24, 28, 27) {real, imag} */,
  {32'h3da0f53e, 32'h3d1aca98} /* (24, 28, 26) {real, imag} */,
  {32'hbcf76e2e, 32'h3e04b31c} /* (24, 28, 25) {real, imag} */,
  {32'h3df963b2, 32'hbde7850e} /* (24, 28, 24) {real, imag} */,
  {32'hbd1bd78e, 32'h3b8a9b64} /* (24, 28, 23) {real, imag} */,
  {32'hbd8be113, 32'hbdcc70f8} /* (24, 28, 22) {real, imag} */,
  {32'hbd92c13a, 32'hbe02b109} /* (24, 28, 21) {real, imag} */,
  {32'h3c7fc4b2, 32'h3d0a3f8b} /* (24, 28, 20) {real, imag} */,
  {32'h3c59c22c, 32'h3d56ab72} /* (24, 28, 19) {real, imag} */,
  {32'h3c9f5099, 32'hbd9ca680} /* (24, 28, 18) {real, imag} */,
  {32'h3c00fbe0, 32'hbc578f62} /* (24, 28, 17) {real, imag} */,
  {32'hbd37bea6, 32'h00000000} /* (24, 28, 16) {real, imag} */,
  {32'h3c00fbe0, 32'h3c578f62} /* (24, 28, 15) {real, imag} */,
  {32'h3c9f5099, 32'h3d9ca680} /* (24, 28, 14) {real, imag} */,
  {32'h3c59c22c, 32'hbd56ab72} /* (24, 28, 13) {real, imag} */,
  {32'h3c7fc4b2, 32'hbd0a3f8b} /* (24, 28, 12) {real, imag} */,
  {32'hbd92c13a, 32'h3e02b109} /* (24, 28, 11) {real, imag} */,
  {32'hbd8be113, 32'h3dcc70f8} /* (24, 28, 10) {real, imag} */,
  {32'hbd1bd78e, 32'hbb8a9b64} /* (24, 28, 9) {real, imag} */,
  {32'h3df963b2, 32'h3de7850e} /* (24, 28, 8) {real, imag} */,
  {32'hbcf76e2e, 32'hbe04b31c} /* (24, 28, 7) {real, imag} */,
  {32'h3da0f53e, 32'hbd1aca98} /* (24, 28, 6) {real, imag} */,
  {32'h3e1b55f1, 32'h3e5d9435} /* (24, 28, 5) {real, imag} */,
  {32'hbe10fe04, 32'hbdc53e8a} /* (24, 28, 4) {real, imag} */,
  {32'hbde7b16e, 32'h3d29454c} /* (24, 28, 3) {real, imag} */,
  {32'h3f9414e1, 32'h3e2e60a8} /* (24, 28, 2) {real, imag} */,
  {32'hc075f335, 32'hbf8a97c2} /* (24, 28, 1) {real, imag} */,
  {32'hc08ec3c9, 32'h00000000} /* (24, 28, 0) {real, imag} */,
  {32'hc070f256, 32'h3f7a9168} /* (24, 27, 31) {real, imag} */,
  {32'h3f9e3028, 32'hbe494f11} /* (24, 27, 30) {real, imag} */,
  {32'h3d2c2614, 32'hbe527e47} /* (24, 27, 29) {real, imag} */,
  {32'hbe2955a0, 32'hbb39b320} /* (24, 27, 28) {real, imag} */,
  {32'h3e1d3f60, 32'hbe3f122e} /* (24, 27, 27) {real, imag} */,
  {32'h3d07023b, 32'h3e8ac11e} /* (24, 27, 26) {real, imag} */,
  {32'h3c3d6f8e, 32'h3d483658} /* (24, 27, 25) {real, imag} */,
  {32'h3da1fa50, 32'hbe0040ca} /* (24, 27, 24) {real, imag} */,
  {32'h3d83b3c7, 32'hbcaf78a2} /* (24, 27, 23) {real, imag} */,
  {32'hbd9b919e, 32'hbd8337ea} /* (24, 27, 22) {real, imag} */,
  {32'hbd9d701d, 32'h3cf5c960} /* (24, 27, 21) {real, imag} */,
  {32'h3d4093be, 32'h3d4d49ca} /* (24, 27, 20) {real, imag} */,
  {32'h3d81bb18, 32'h3cdc12de} /* (24, 27, 19) {real, imag} */,
  {32'h3d833435, 32'hbd90782c} /* (24, 27, 18) {real, imag} */,
  {32'h3c619245, 32'h3d2a39e6} /* (24, 27, 17) {real, imag} */,
  {32'hbd587241, 32'h00000000} /* (24, 27, 16) {real, imag} */,
  {32'h3c619245, 32'hbd2a39e6} /* (24, 27, 15) {real, imag} */,
  {32'h3d833435, 32'h3d90782c} /* (24, 27, 14) {real, imag} */,
  {32'h3d81bb18, 32'hbcdc12de} /* (24, 27, 13) {real, imag} */,
  {32'h3d4093be, 32'hbd4d49ca} /* (24, 27, 12) {real, imag} */,
  {32'hbd9d701d, 32'hbcf5c960} /* (24, 27, 11) {real, imag} */,
  {32'hbd9b919e, 32'h3d8337ea} /* (24, 27, 10) {real, imag} */,
  {32'h3d83b3c7, 32'h3caf78a2} /* (24, 27, 9) {real, imag} */,
  {32'h3da1fa50, 32'h3e0040ca} /* (24, 27, 8) {real, imag} */,
  {32'h3c3d6f8e, 32'hbd483658} /* (24, 27, 7) {real, imag} */,
  {32'h3d07023b, 32'hbe8ac11e} /* (24, 27, 6) {real, imag} */,
  {32'h3e1d3f60, 32'h3e3f122e} /* (24, 27, 5) {real, imag} */,
  {32'hbe2955a0, 32'h3b39b320} /* (24, 27, 4) {real, imag} */,
  {32'h3d2c2614, 32'h3e527e47} /* (24, 27, 3) {real, imag} */,
  {32'h3f9e3028, 32'h3e494f11} /* (24, 27, 2) {real, imag} */,
  {32'hc070f256, 32'hbf7a9168} /* (24, 27, 1) {real, imag} */,
  {32'hc08ad12b, 32'h00000000} /* (24, 27, 0) {real, imag} */,
  {32'hc065d2ab, 32'h3f4b37fc} /* (24, 26, 31) {real, imag} */,
  {32'h3fa78be2, 32'hbd0d8770} /* (24, 26, 30) {real, imag} */,
  {32'h3ce2609e, 32'hbde22750} /* (24, 26, 29) {real, imag} */,
  {32'hbd8aea6c, 32'hbd7fa1a5} /* (24, 26, 28) {real, imag} */,
  {32'h3e12ae7c, 32'hbda70042} /* (24, 26, 27) {real, imag} */,
  {32'hbd6f4ca4, 32'h3e2a4e00} /* (24, 26, 26) {real, imag} */,
  {32'h3d7560c2, 32'h3d23e65f} /* (24, 26, 25) {real, imag} */,
  {32'h3df82334, 32'hbd4865fe} /* (24, 26, 24) {real, imag} */,
  {32'hbc4ced4a, 32'h3d503c18} /* (24, 26, 23) {real, imag} */,
  {32'hbd26f18c, 32'hbd67ae35} /* (24, 26, 22) {real, imag} */,
  {32'hbd14faa2, 32'hbd30b932} /* (24, 26, 21) {real, imag} */,
  {32'hbd2e0034, 32'h3d27fabe} /* (24, 26, 20) {real, imag} */,
  {32'h3c4ed562, 32'hbce1103b} /* (24, 26, 19) {real, imag} */,
  {32'hbb33fe40, 32'hbcdeb6a6} /* (24, 26, 18) {real, imag} */,
  {32'hbd595fb2, 32'hbccb814c} /* (24, 26, 17) {real, imag} */,
  {32'h3da8c0d6, 32'h00000000} /* (24, 26, 16) {real, imag} */,
  {32'hbd595fb2, 32'h3ccb814c} /* (24, 26, 15) {real, imag} */,
  {32'hbb33fe40, 32'h3cdeb6a6} /* (24, 26, 14) {real, imag} */,
  {32'h3c4ed562, 32'h3ce1103b} /* (24, 26, 13) {real, imag} */,
  {32'hbd2e0034, 32'hbd27fabe} /* (24, 26, 12) {real, imag} */,
  {32'hbd14faa2, 32'h3d30b932} /* (24, 26, 11) {real, imag} */,
  {32'hbd26f18c, 32'h3d67ae35} /* (24, 26, 10) {real, imag} */,
  {32'hbc4ced4a, 32'hbd503c18} /* (24, 26, 9) {real, imag} */,
  {32'h3df82334, 32'h3d4865fe} /* (24, 26, 8) {real, imag} */,
  {32'h3d7560c2, 32'hbd23e65f} /* (24, 26, 7) {real, imag} */,
  {32'hbd6f4ca4, 32'hbe2a4e00} /* (24, 26, 6) {real, imag} */,
  {32'h3e12ae7c, 32'h3da70042} /* (24, 26, 5) {real, imag} */,
  {32'hbd8aea6c, 32'h3d7fa1a5} /* (24, 26, 4) {real, imag} */,
  {32'h3ce2609e, 32'h3de22750} /* (24, 26, 3) {real, imag} */,
  {32'h3fa78be2, 32'h3d0d8770} /* (24, 26, 2) {real, imag} */,
  {32'hc065d2ab, 32'hbf4b37fc} /* (24, 26, 1) {real, imag} */,
  {32'hc0830d28, 32'h00000000} /* (24, 26, 0) {real, imag} */,
  {32'hc0619377, 32'h3f014af7} /* (24, 25, 31) {real, imag} */,
  {32'h3f9cd62f, 32'h3dab27b7} /* (24, 25, 30) {real, imag} */,
  {32'h3cec7d36, 32'h3b94e804} /* (24, 25, 29) {real, imag} */,
  {32'hbdac581b, 32'hbc07c196} /* (24, 25, 28) {real, imag} */,
  {32'h3e762912, 32'hbc3f8434} /* (24, 25, 27) {real, imag} */,
  {32'h3c8370ae, 32'h3d924c66} /* (24, 25, 26) {real, imag} */,
  {32'h3d2db566, 32'h3d022314} /* (24, 25, 25) {real, imag} */,
  {32'hbdb59be1, 32'hbd272bd2} /* (24, 25, 24) {real, imag} */,
  {32'hbd99ccbc, 32'hbe310993} /* (24, 25, 23) {real, imag} */,
  {32'hbd7e2189, 32'hbb897450} /* (24, 25, 22) {real, imag} */,
  {32'h3cbc76bc, 32'hbdbfd223} /* (24, 25, 21) {real, imag} */,
  {32'hbd8f6c66, 32'h3cbd69c9} /* (24, 25, 20) {real, imag} */,
  {32'hbcdce381, 32'hbce3bcd6} /* (24, 25, 19) {real, imag} */,
  {32'hbdafbcd8, 32'h3db7c5a2} /* (24, 25, 18) {real, imag} */,
  {32'h3cd5f269, 32'h3cf203f0} /* (24, 25, 17) {real, imag} */,
  {32'h3ca8ac09, 32'h00000000} /* (24, 25, 16) {real, imag} */,
  {32'h3cd5f269, 32'hbcf203f0} /* (24, 25, 15) {real, imag} */,
  {32'hbdafbcd8, 32'hbdb7c5a2} /* (24, 25, 14) {real, imag} */,
  {32'hbcdce381, 32'h3ce3bcd6} /* (24, 25, 13) {real, imag} */,
  {32'hbd8f6c66, 32'hbcbd69c9} /* (24, 25, 12) {real, imag} */,
  {32'h3cbc76bc, 32'h3dbfd223} /* (24, 25, 11) {real, imag} */,
  {32'hbd7e2189, 32'h3b897450} /* (24, 25, 10) {real, imag} */,
  {32'hbd99ccbc, 32'h3e310993} /* (24, 25, 9) {real, imag} */,
  {32'hbdb59be1, 32'h3d272bd2} /* (24, 25, 8) {real, imag} */,
  {32'h3d2db566, 32'hbd022314} /* (24, 25, 7) {real, imag} */,
  {32'h3c8370ae, 32'hbd924c66} /* (24, 25, 6) {real, imag} */,
  {32'h3e762912, 32'h3c3f8434} /* (24, 25, 5) {real, imag} */,
  {32'hbdac581b, 32'h3c07c196} /* (24, 25, 4) {real, imag} */,
  {32'h3cec7d36, 32'hbb94e804} /* (24, 25, 3) {real, imag} */,
  {32'h3f9cd62f, 32'hbdab27b7} /* (24, 25, 2) {real, imag} */,
  {32'hc0619377, 32'hbf014af7} /* (24, 25, 1) {real, imag} */,
  {32'hc076c0c2, 32'h00000000} /* (24, 25, 0) {real, imag} */,
  {32'hc044b1d2, 32'h3ee29bf4} /* (24, 24, 31) {real, imag} */,
  {32'h3f939cad, 32'hbdaf7668} /* (24, 24, 30) {real, imag} */,
  {32'hbdf8eaaa, 32'hbc9ccfc6} /* (24, 24, 29) {real, imag} */,
  {32'hbdc7cebe, 32'hbda1da5e} /* (24, 24, 28) {real, imag} */,
  {32'h3e318e06, 32'hbd32fa8c} /* (24, 24, 27) {real, imag} */,
  {32'h3df1fd46, 32'h3c07fb18} /* (24, 24, 26) {real, imag} */,
  {32'h3d344734, 32'h3d3a8796} /* (24, 24, 25) {real, imag} */,
  {32'hbd42d02a, 32'hbceebf8f} /* (24, 24, 24) {real, imag} */,
  {32'hbd68a302, 32'h3a9e36e8} /* (24, 24, 23) {real, imag} */,
  {32'hbcc85b3a, 32'h3da856ee} /* (24, 24, 22) {real, imag} */,
  {32'hbd769ddf, 32'hbd20c7ea} /* (24, 24, 21) {real, imag} */,
  {32'hbc7dbb54, 32'h3d6022c7} /* (24, 24, 20) {real, imag} */,
  {32'hb98bd160, 32'hbd826fdd} /* (24, 24, 19) {real, imag} */,
  {32'h3a8a8980, 32'hbe08281c} /* (24, 24, 18) {real, imag} */,
  {32'hbc6b7b3c, 32'h3ca6e456} /* (24, 24, 17) {real, imag} */,
  {32'hbc8ad264, 32'h00000000} /* (24, 24, 16) {real, imag} */,
  {32'hbc6b7b3c, 32'hbca6e456} /* (24, 24, 15) {real, imag} */,
  {32'h3a8a8980, 32'h3e08281c} /* (24, 24, 14) {real, imag} */,
  {32'hb98bd160, 32'h3d826fdd} /* (24, 24, 13) {real, imag} */,
  {32'hbc7dbb54, 32'hbd6022c7} /* (24, 24, 12) {real, imag} */,
  {32'hbd769ddf, 32'h3d20c7ea} /* (24, 24, 11) {real, imag} */,
  {32'hbcc85b3a, 32'hbda856ee} /* (24, 24, 10) {real, imag} */,
  {32'hbd68a302, 32'hba9e36e8} /* (24, 24, 9) {real, imag} */,
  {32'hbd42d02a, 32'h3ceebf8f} /* (24, 24, 8) {real, imag} */,
  {32'h3d344734, 32'hbd3a8796} /* (24, 24, 7) {real, imag} */,
  {32'h3df1fd46, 32'hbc07fb18} /* (24, 24, 6) {real, imag} */,
  {32'h3e318e06, 32'h3d32fa8c} /* (24, 24, 5) {real, imag} */,
  {32'hbdc7cebe, 32'h3da1da5e} /* (24, 24, 4) {real, imag} */,
  {32'hbdf8eaaa, 32'h3c9ccfc6} /* (24, 24, 3) {real, imag} */,
  {32'h3f939cad, 32'h3daf7668} /* (24, 24, 2) {real, imag} */,
  {32'hc044b1d2, 32'hbee29bf4} /* (24, 24, 1) {real, imag} */,
  {32'hc054edb6, 32'h00000000} /* (24, 24, 0) {real, imag} */,
  {32'hc029e172, 32'h3ebbc3f2} /* (24, 23, 31) {real, imag} */,
  {32'h3f850fde, 32'hbe418478} /* (24, 23, 30) {real, imag} */,
  {32'hbdbb865c, 32'h3c9b8ca6} /* (24, 23, 29) {real, imag} */,
  {32'hbe26d0c5, 32'h3cce6c5a} /* (24, 23, 28) {real, imag} */,
  {32'h3e04d756, 32'hbdc1fc15} /* (24, 23, 27) {real, imag} */,
  {32'hbdd13736, 32'hbe04b6c8} /* (24, 23, 26) {real, imag} */,
  {32'hbc4afbc0, 32'hbcaac09f} /* (24, 23, 25) {real, imag} */,
  {32'h3cffc040, 32'hbd8f4603} /* (24, 23, 24) {real, imag} */,
  {32'h3ddcf3c2, 32'hbe063a6d} /* (24, 23, 23) {real, imag} */,
  {32'hbc88e122, 32'hbd2fee56} /* (24, 23, 22) {real, imag} */,
  {32'h3ddb27f0, 32'hbce240f0} /* (24, 23, 21) {real, imag} */,
  {32'hbd5445f5, 32'h3d6ee038} /* (24, 23, 20) {real, imag} */,
  {32'hbd5c12f1, 32'h3cb8c9f4} /* (24, 23, 19) {real, imag} */,
  {32'h3d0dfab8, 32'hbca81064} /* (24, 23, 18) {real, imag} */,
  {32'h3b50eeae, 32'hbcb181b3} /* (24, 23, 17) {real, imag} */,
  {32'h3d63895d, 32'h00000000} /* (24, 23, 16) {real, imag} */,
  {32'h3b50eeae, 32'h3cb181b3} /* (24, 23, 15) {real, imag} */,
  {32'h3d0dfab8, 32'h3ca81064} /* (24, 23, 14) {real, imag} */,
  {32'hbd5c12f1, 32'hbcb8c9f4} /* (24, 23, 13) {real, imag} */,
  {32'hbd5445f5, 32'hbd6ee038} /* (24, 23, 12) {real, imag} */,
  {32'h3ddb27f0, 32'h3ce240f0} /* (24, 23, 11) {real, imag} */,
  {32'hbc88e122, 32'h3d2fee56} /* (24, 23, 10) {real, imag} */,
  {32'h3ddcf3c2, 32'h3e063a6d} /* (24, 23, 9) {real, imag} */,
  {32'h3cffc040, 32'h3d8f4603} /* (24, 23, 8) {real, imag} */,
  {32'hbc4afbc0, 32'h3caac09f} /* (24, 23, 7) {real, imag} */,
  {32'hbdd13736, 32'h3e04b6c8} /* (24, 23, 6) {real, imag} */,
  {32'h3e04d756, 32'h3dc1fc15} /* (24, 23, 5) {real, imag} */,
  {32'hbe26d0c5, 32'hbcce6c5a} /* (24, 23, 4) {real, imag} */,
  {32'hbdbb865c, 32'hbc9b8ca6} /* (24, 23, 3) {real, imag} */,
  {32'h3f850fde, 32'h3e418478} /* (24, 23, 2) {real, imag} */,
  {32'hc029e172, 32'hbebbc3f2} /* (24, 23, 1) {real, imag} */,
  {32'hc029c570, 32'h00000000} /* (24, 23, 0) {real, imag} */,
  {32'hc00a861b, 32'h3e8405c5} /* (24, 22, 31) {real, imag} */,
  {32'h3f5cede4, 32'hbd7331d8} /* (24, 22, 30) {real, imag} */,
  {32'hbbc0cc30, 32'h3d894662} /* (24, 22, 29) {real, imag} */,
  {32'hbe6fd172, 32'h3e091f6b} /* (24, 22, 28) {real, imag} */,
  {32'h3e89f72d, 32'hbdd9748a} /* (24, 22, 27) {real, imag} */,
  {32'hbe03ea2a, 32'hbdc3df77} /* (24, 22, 26) {real, imag} */,
  {32'hbd07b0f8, 32'h3cf425aa} /* (24, 22, 25) {real, imag} */,
  {32'h3cdd57d2, 32'hbcda7a41} /* (24, 22, 24) {real, imag} */,
  {32'hbc5b5f50, 32'hbd17fc99} /* (24, 22, 23) {real, imag} */,
  {32'hbd0bf15e, 32'hbb8954c4} /* (24, 22, 22) {real, imag} */,
  {32'hbd151428, 32'hbc45ee96} /* (24, 22, 21) {real, imag} */,
  {32'h3cc8e124, 32'h3cdfc524} /* (24, 22, 20) {real, imag} */,
  {32'hbcdec561, 32'h3d169040} /* (24, 22, 19) {real, imag} */,
  {32'h3c6acc5c, 32'h3d4c679c} /* (24, 22, 18) {real, imag} */,
  {32'h3d88f0a1, 32'hbd8a1499} /* (24, 22, 17) {real, imag} */,
  {32'hbcc364a4, 32'h00000000} /* (24, 22, 16) {real, imag} */,
  {32'h3d88f0a1, 32'h3d8a1499} /* (24, 22, 15) {real, imag} */,
  {32'h3c6acc5c, 32'hbd4c679c} /* (24, 22, 14) {real, imag} */,
  {32'hbcdec561, 32'hbd169040} /* (24, 22, 13) {real, imag} */,
  {32'h3cc8e124, 32'hbcdfc524} /* (24, 22, 12) {real, imag} */,
  {32'hbd151428, 32'h3c45ee96} /* (24, 22, 11) {real, imag} */,
  {32'hbd0bf15e, 32'h3b8954c4} /* (24, 22, 10) {real, imag} */,
  {32'hbc5b5f50, 32'h3d17fc99} /* (24, 22, 9) {real, imag} */,
  {32'h3cdd57d2, 32'h3cda7a41} /* (24, 22, 8) {real, imag} */,
  {32'hbd07b0f8, 32'hbcf425aa} /* (24, 22, 7) {real, imag} */,
  {32'hbe03ea2a, 32'h3dc3df77} /* (24, 22, 6) {real, imag} */,
  {32'h3e89f72d, 32'h3dd9748a} /* (24, 22, 5) {real, imag} */,
  {32'hbe6fd172, 32'hbe091f6b} /* (24, 22, 4) {real, imag} */,
  {32'hbbc0cc30, 32'hbd894662} /* (24, 22, 3) {real, imag} */,
  {32'h3f5cede4, 32'h3d7331d8} /* (24, 22, 2) {real, imag} */,
  {32'hc00a861b, 32'hbe8405c5} /* (24, 22, 1) {real, imag} */,
  {32'hbff34d36, 32'h00000000} /* (24, 22, 0) {real, imag} */,
  {32'hbf6602f0, 32'h3dd62940} /* (24, 21, 31) {real, imag} */,
  {32'h3ec5ebe7, 32'hbdd151ee} /* (24, 21, 30) {real, imag} */,
  {32'h3d2e1d4d, 32'h3dbadc45} /* (24, 21, 29) {real, imag} */,
  {32'h3d37dce8, 32'h3ac9c200} /* (24, 21, 28) {real, imag} */,
  {32'h3e261baa, 32'h3d83890d} /* (24, 21, 27) {real, imag} */,
  {32'h3c24fc9d, 32'h3de880a4} /* (24, 21, 26) {real, imag} */,
  {32'h3d358709, 32'hbda56231} /* (24, 21, 25) {real, imag} */,
  {32'hbcbc2b36, 32'h3d219f17} /* (24, 21, 24) {real, imag} */,
  {32'hbe1ca07c, 32'h3cb14c08} /* (24, 21, 23) {real, imag} */,
  {32'h3aad8b68, 32'hbd813ebd} /* (24, 21, 22) {real, imag} */,
  {32'hbdfd67de, 32'h3c54964f} /* (24, 21, 21) {real, imag} */,
  {32'h3cea8528, 32'h3b933610} /* (24, 21, 20) {real, imag} */,
  {32'hbb69d1e4, 32'hbc2f6052} /* (24, 21, 19) {real, imag} */,
  {32'h3d2ed539, 32'h3d2fbe7c} /* (24, 21, 18) {real, imag} */,
  {32'hbcad782e, 32'h3c1f1eec} /* (24, 21, 17) {real, imag} */,
  {32'h3d216a5f, 32'h00000000} /* (24, 21, 16) {real, imag} */,
  {32'hbcad782e, 32'hbc1f1eec} /* (24, 21, 15) {real, imag} */,
  {32'h3d2ed539, 32'hbd2fbe7c} /* (24, 21, 14) {real, imag} */,
  {32'hbb69d1e4, 32'h3c2f6052} /* (24, 21, 13) {real, imag} */,
  {32'h3cea8528, 32'hbb933610} /* (24, 21, 12) {real, imag} */,
  {32'hbdfd67de, 32'hbc54964f} /* (24, 21, 11) {real, imag} */,
  {32'h3aad8b68, 32'h3d813ebd} /* (24, 21, 10) {real, imag} */,
  {32'hbe1ca07c, 32'hbcb14c08} /* (24, 21, 9) {real, imag} */,
  {32'hbcbc2b36, 32'hbd219f17} /* (24, 21, 8) {real, imag} */,
  {32'h3d358709, 32'h3da56231} /* (24, 21, 7) {real, imag} */,
  {32'h3c24fc9d, 32'hbde880a4} /* (24, 21, 6) {real, imag} */,
  {32'h3e261baa, 32'hbd83890d} /* (24, 21, 5) {real, imag} */,
  {32'h3d37dce8, 32'hbac9c200} /* (24, 21, 4) {real, imag} */,
  {32'h3d2e1d4d, 32'hbdbadc45} /* (24, 21, 3) {real, imag} */,
  {32'h3ec5ebe7, 32'h3dd151ee} /* (24, 21, 2) {real, imag} */,
  {32'hbf6602f0, 32'hbdd62940} /* (24, 21, 1) {real, imag} */,
  {32'hbf471abb, 32'h00000000} /* (24, 21, 0) {real, imag} */,
  {32'h3f311f59, 32'hbe537cdc} /* (24, 20, 31) {real, imag} */,
  {32'hbec8b2ec, 32'h3d790f2c} /* (24, 20, 30) {real, imag} */,
  {32'h3d98a550, 32'h3e168d43} /* (24, 20, 29) {real, imag} */,
  {32'h3e16e454, 32'hbe12695d} /* (24, 20, 28) {real, imag} */,
  {32'hbda02581, 32'h3db1cd76} /* (24, 20, 27) {real, imag} */,
  {32'h3d8bbc48, 32'h3d27e60e} /* (24, 20, 26) {real, imag} */,
  {32'h3dbf0696, 32'hbe20b502} /* (24, 20, 25) {real, imag} */,
  {32'hbddd47d9, 32'h3d4b33c6} /* (24, 20, 24) {real, imag} */,
  {32'hbdab7ba0, 32'h3e0b400b} /* (24, 20, 23) {real, imag} */,
  {32'h3d597ffc, 32'hbd3bf132} /* (24, 20, 22) {real, imag} */,
  {32'h3d69f585, 32'h3db0ae92} /* (24, 20, 21) {real, imag} */,
  {32'hbd36782f, 32'hbd20b746} /* (24, 20, 20) {real, imag} */,
  {32'hbdcf2f3e, 32'hbda043f6} /* (24, 20, 19) {real, imag} */,
  {32'h3d8f0c92, 32'h3c8f2650} /* (24, 20, 18) {real, imag} */,
  {32'hbccb7218, 32'h3bd2e570} /* (24, 20, 17) {real, imag} */,
  {32'h3ce3ad3e, 32'h00000000} /* (24, 20, 16) {real, imag} */,
  {32'hbccb7218, 32'hbbd2e570} /* (24, 20, 15) {real, imag} */,
  {32'h3d8f0c92, 32'hbc8f2650} /* (24, 20, 14) {real, imag} */,
  {32'hbdcf2f3e, 32'h3da043f6} /* (24, 20, 13) {real, imag} */,
  {32'hbd36782f, 32'h3d20b746} /* (24, 20, 12) {real, imag} */,
  {32'h3d69f585, 32'hbdb0ae92} /* (24, 20, 11) {real, imag} */,
  {32'h3d597ffc, 32'h3d3bf132} /* (24, 20, 10) {real, imag} */,
  {32'hbdab7ba0, 32'hbe0b400b} /* (24, 20, 9) {real, imag} */,
  {32'hbddd47d9, 32'hbd4b33c6} /* (24, 20, 8) {real, imag} */,
  {32'h3dbf0696, 32'h3e20b502} /* (24, 20, 7) {real, imag} */,
  {32'h3d8bbc48, 32'hbd27e60e} /* (24, 20, 6) {real, imag} */,
  {32'hbda02581, 32'hbdb1cd76} /* (24, 20, 5) {real, imag} */,
  {32'h3e16e454, 32'h3e12695d} /* (24, 20, 4) {real, imag} */,
  {32'h3d98a550, 32'hbe168d43} /* (24, 20, 3) {real, imag} */,
  {32'hbec8b2ec, 32'hbd790f2c} /* (24, 20, 2) {real, imag} */,
  {32'h3f311f59, 32'h3e537cdc} /* (24, 20, 1) {real, imag} */,
  {32'h3eb768c6, 32'h00000000} /* (24, 20, 0) {real, imag} */,
  {32'h3fc5b83a, 32'hbe4443f8} /* (24, 19, 31) {real, imag} */,
  {32'hbf4a3ac8, 32'h3dca1658} /* (24, 19, 30) {real, imag} */,
  {32'h3d13ec54, 32'h3d847107} /* (24, 19, 29) {real, imag} */,
  {32'h3e436692, 32'hbe381637} /* (24, 19, 28) {real, imag} */,
  {32'hbe0f7817, 32'h3df70c11} /* (24, 19, 27) {real, imag} */,
  {32'h3d952ba0, 32'hbd165d93} /* (24, 19, 26) {real, imag} */,
  {32'h3d541370, 32'h3c1d7637} /* (24, 19, 25) {real, imag} */,
  {32'hbe34a3f4, 32'h3db94183} /* (24, 19, 24) {real, imag} */,
  {32'hbd3fcb9b, 32'h3aeb5310} /* (24, 19, 23) {real, imag} */,
  {32'h3a96b580, 32'h3d7f9728} /* (24, 19, 22) {real, imag} */,
  {32'h3c5e6653, 32'h3d29ffdb} /* (24, 19, 21) {real, imag} */,
  {32'h3c8897c8, 32'hbcd50525} /* (24, 19, 20) {real, imag} */,
  {32'hbd48dd06, 32'hbd0ea6ea} /* (24, 19, 19) {real, imag} */,
  {32'hbd0548aa, 32'h3d371039} /* (24, 19, 18) {real, imag} */,
  {32'h3d043c4c, 32'hbd595b1e} /* (24, 19, 17) {real, imag} */,
  {32'h3be9ef48, 32'h00000000} /* (24, 19, 16) {real, imag} */,
  {32'h3d043c4c, 32'h3d595b1e} /* (24, 19, 15) {real, imag} */,
  {32'hbd0548aa, 32'hbd371039} /* (24, 19, 14) {real, imag} */,
  {32'hbd48dd06, 32'h3d0ea6ea} /* (24, 19, 13) {real, imag} */,
  {32'h3c8897c8, 32'h3cd50525} /* (24, 19, 12) {real, imag} */,
  {32'h3c5e6653, 32'hbd29ffdb} /* (24, 19, 11) {real, imag} */,
  {32'h3a96b580, 32'hbd7f9728} /* (24, 19, 10) {real, imag} */,
  {32'hbd3fcb9b, 32'hbaeb5310} /* (24, 19, 9) {real, imag} */,
  {32'hbe34a3f4, 32'hbdb94183} /* (24, 19, 8) {real, imag} */,
  {32'h3d541370, 32'hbc1d7637} /* (24, 19, 7) {real, imag} */,
  {32'h3d952ba0, 32'h3d165d93} /* (24, 19, 6) {real, imag} */,
  {32'hbe0f7817, 32'hbdf70c11} /* (24, 19, 5) {real, imag} */,
  {32'h3e436692, 32'h3e381637} /* (24, 19, 4) {real, imag} */,
  {32'h3d13ec54, 32'hbd847107} /* (24, 19, 3) {real, imag} */,
  {32'hbf4a3ac8, 32'hbdca1658} /* (24, 19, 2) {real, imag} */,
  {32'h3fc5b83a, 32'h3e4443f8} /* (24, 19, 1) {real, imag} */,
  {32'h3f8972b3, 32'h00000000} /* (24, 19, 0) {real, imag} */,
  {32'h40084958, 32'hbe7c266c} /* (24, 18, 31) {real, imag} */,
  {32'hbf514738, 32'h3d4d3806} /* (24, 18, 30) {real, imag} */,
  {32'h3e15ccfe, 32'h3bc8c1c0} /* (24, 18, 29) {real, imag} */,
  {32'h3e778412, 32'hbe54fc58} /* (24, 18, 28) {real, imag} */,
  {32'hbe43802c, 32'h3da8c7dc} /* (24, 18, 27) {real, imag} */,
  {32'h3db88ff4, 32'hbd82dc49} /* (24, 18, 26) {real, imag} */,
  {32'hbd916d1c, 32'h3c6c6e60} /* (24, 18, 25) {real, imag} */,
  {32'hbd62e040, 32'h3e2838bc} /* (24, 18, 24) {real, imag} */,
  {32'h3d3cfc90, 32'hbcbdb7e8} /* (24, 18, 23) {real, imag} */,
  {32'h3d51a4c6, 32'hbe0aa28e} /* (24, 18, 22) {real, imag} */,
  {32'hbe04c81d, 32'h3e135481} /* (24, 18, 21) {real, imag} */,
  {32'h3da06a4a, 32'hbd60ddd4} /* (24, 18, 20) {real, imag} */,
  {32'hbcee9876, 32'h3d00a9e4} /* (24, 18, 19) {real, imag} */,
  {32'h3c2fa871, 32'h3d8e3306} /* (24, 18, 18) {real, imag} */,
  {32'hbd5d9e18, 32'hbc46462f} /* (24, 18, 17) {real, imag} */,
  {32'hbc558a50, 32'h00000000} /* (24, 18, 16) {real, imag} */,
  {32'hbd5d9e18, 32'h3c46462f} /* (24, 18, 15) {real, imag} */,
  {32'h3c2fa871, 32'hbd8e3306} /* (24, 18, 14) {real, imag} */,
  {32'hbcee9876, 32'hbd00a9e4} /* (24, 18, 13) {real, imag} */,
  {32'h3da06a4a, 32'h3d60ddd4} /* (24, 18, 12) {real, imag} */,
  {32'hbe04c81d, 32'hbe135481} /* (24, 18, 11) {real, imag} */,
  {32'h3d51a4c6, 32'h3e0aa28e} /* (24, 18, 10) {real, imag} */,
  {32'h3d3cfc90, 32'h3cbdb7e8} /* (24, 18, 9) {real, imag} */,
  {32'hbd62e040, 32'hbe2838bc} /* (24, 18, 8) {real, imag} */,
  {32'hbd916d1c, 32'hbc6c6e60} /* (24, 18, 7) {real, imag} */,
  {32'h3db88ff4, 32'h3d82dc49} /* (24, 18, 6) {real, imag} */,
  {32'hbe43802c, 32'hbda8c7dc} /* (24, 18, 5) {real, imag} */,
  {32'h3e778412, 32'h3e54fc58} /* (24, 18, 4) {real, imag} */,
  {32'h3e15ccfe, 32'hbbc8c1c0} /* (24, 18, 3) {real, imag} */,
  {32'hbf514738, 32'hbd4d3806} /* (24, 18, 2) {real, imag} */,
  {32'h40084958, 32'h3e7c266c} /* (24, 18, 1) {real, imag} */,
  {32'h3fcb0dd9, 32'h00000000} /* (24, 18, 0) {real, imag} */,
  {32'h40286346, 32'hbeba94a6} /* (24, 17, 31) {real, imag} */,
  {32'hbf576bb6, 32'h3e4d8d3d} /* (24, 17, 30) {real, imag} */,
  {32'h3db2093e, 32'h3d3a8210} /* (24, 17, 29) {real, imag} */,
  {32'h3e716fce, 32'hbdd031b2} /* (24, 17, 28) {real, imag} */,
  {32'hbde32c00, 32'h3d01fd6e} /* (24, 17, 27) {real, imag} */,
  {32'h3d98fa0a, 32'h3d5bea1c} /* (24, 17, 26) {real, imag} */,
  {32'h3da29936, 32'hbb8abce4} /* (24, 17, 25) {real, imag} */,
  {32'h3d24e1a6, 32'h3cc2604c} /* (24, 17, 24) {real, imag} */,
  {32'h3bad7e2c, 32'hbd03c173} /* (24, 17, 23) {real, imag} */,
  {32'h3cdd90a8, 32'h3bb1270c} /* (24, 17, 22) {real, imag} */,
  {32'h3ce0dc80, 32'h3df6a1b5} /* (24, 17, 21) {real, imag} */,
  {32'h3c889737, 32'h3ce0bf06} /* (24, 17, 20) {real, imag} */,
  {32'hbb84539c, 32'h3d1ab4cd} /* (24, 17, 19) {real, imag} */,
  {32'h3dbe4488, 32'hbc8b63d0} /* (24, 17, 18) {real, imag} */,
  {32'hbc7aded4, 32'hbc3b5bbe} /* (24, 17, 17) {real, imag} */,
  {32'hbcf14771, 32'h00000000} /* (24, 17, 16) {real, imag} */,
  {32'hbc7aded4, 32'h3c3b5bbe} /* (24, 17, 15) {real, imag} */,
  {32'h3dbe4488, 32'h3c8b63d0} /* (24, 17, 14) {real, imag} */,
  {32'hbb84539c, 32'hbd1ab4cd} /* (24, 17, 13) {real, imag} */,
  {32'h3c889737, 32'hbce0bf06} /* (24, 17, 12) {real, imag} */,
  {32'h3ce0dc80, 32'hbdf6a1b5} /* (24, 17, 11) {real, imag} */,
  {32'h3cdd90a8, 32'hbbb1270c} /* (24, 17, 10) {real, imag} */,
  {32'h3bad7e2c, 32'h3d03c173} /* (24, 17, 9) {real, imag} */,
  {32'h3d24e1a6, 32'hbcc2604c} /* (24, 17, 8) {real, imag} */,
  {32'h3da29936, 32'h3b8abce4} /* (24, 17, 7) {real, imag} */,
  {32'h3d98fa0a, 32'hbd5bea1c} /* (24, 17, 6) {real, imag} */,
  {32'hbde32c00, 32'hbd01fd6e} /* (24, 17, 5) {real, imag} */,
  {32'h3e716fce, 32'h3dd031b2} /* (24, 17, 4) {real, imag} */,
  {32'h3db2093e, 32'hbd3a8210} /* (24, 17, 3) {real, imag} */,
  {32'hbf576bb6, 32'hbe4d8d3d} /* (24, 17, 2) {real, imag} */,
  {32'h40286346, 32'h3eba94a6} /* (24, 17, 1) {real, imag} */,
  {32'h3fe402eb, 32'h00000000} /* (24, 17, 0) {real, imag} */,
  {32'h40389e85, 32'hbe6b8300} /* (24, 16, 31) {real, imag} */,
  {32'hbf68f100, 32'h3eb2bd8a} /* (24, 16, 30) {real, imag} */,
  {32'hbc8323f8, 32'h3d4b1b94} /* (24, 16, 29) {real, imag} */,
  {32'h3ea77233, 32'hbe3ce9a2} /* (24, 16, 28) {real, imag} */,
  {32'hbe85d903, 32'hbce33589} /* (24, 16, 27) {real, imag} */,
  {32'h3d27c0e8, 32'h3d2d9848} /* (24, 16, 26) {real, imag} */,
  {32'h3db00872, 32'hbbcf771c} /* (24, 16, 25) {real, imag} */,
  {32'hbde8cd90, 32'h3dd26a5d} /* (24, 16, 24) {real, imag} */,
  {32'h3d7b71d3, 32'hb687d800} /* (24, 16, 23) {real, imag} */,
  {32'hbd9ac810, 32'h3d54c88d} /* (24, 16, 22) {real, imag} */,
  {32'hbc938fc6, 32'h3dd59cae} /* (24, 16, 21) {real, imag} */,
  {32'h3be1b30b, 32'hbcf48737} /* (24, 16, 20) {real, imag} */,
  {32'h3c995e28, 32'hbc9e2a2e} /* (24, 16, 19) {real, imag} */,
  {32'h3cbbcf1a, 32'hbc42011b} /* (24, 16, 18) {real, imag} */,
  {32'h3d26b8a3, 32'h3d4e5148} /* (24, 16, 17) {real, imag} */,
  {32'hbd0d51b8, 32'h00000000} /* (24, 16, 16) {real, imag} */,
  {32'h3d26b8a3, 32'hbd4e5148} /* (24, 16, 15) {real, imag} */,
  {32'h3cbbcf1a, 32'h3c42011b} /* (24, 16, 14) {real, imag} */,
  {32'h3c995e28, 32'h3c9e2a2e} /* (24, 16, 13) {real, imag} */,
  {32'h3be1b30b, 32'h3cf48737} /* (24, 16, 12) {real, imag} */,
  {32'hbc938fc6, 32'hbdd59cae} /* (24, 16, 11) {real, imag} */,
  {32'hbd9ac810, 32'hbd54c88d} /* (24, 16, 10) {real, imag} */,
  {32'h3d7b71d3, 32'h3687d800} /* (24, 16, 9) {real, imag} */,
  {32'hbde8cd90, 32'hbdd26a5d} /* (24, 16, 8) {real, imag} */,
  {32'h3db00872, 32'h3bcf771c} /* (24, 16, 7) {real, imag} */,
  {32'h3d27c0e8, 32'hbd2d9848} /* (24, 16, 6) {real, imag} */,
  {32'hbe85d903, 32'h3ce33589} /* (24, 16, 5) {real, imag} */,
  {32'h3ea77233, 32'h3e3ce9a2} /* (24, 16, 4) {real, imag} */,
  {32'hbc8323f8, 32'hbd4b1b94} /* (24, 16, 3) {real, imag} */,
  {32'hbf68f100, 32'hbeb2bd8a} /* (24, 16, 2) {real, imag} */,
  {32'h40389e85, 32'h3e6b8300} /* (24, 16, 1) {real, imag} */,
  {32'h3ff7c388, 32'h00000000} /* (24, 16, 0) {real, imag} */,
  {32'h403350f2, 32'hbe2f4e15} /* (24, 15, 31) {real, imag} */,
  {32'hbf65b0ca, 32'h3e8776fe} /* (24, 15, 30) {real, imag} */,
  {32'hbd6cc200, 32'h3be2cf40} /* (24, 15, 29) {real, imag} */,
  {32'h3e311eca, 32'hbd60824c} /* (24, 15, 28) {real, imag} */,
  {32'hbe5db7f2, 32'h3cd1e001} /* (24, 15, 27) {real, imag} */,
  {32'hbbba61f8, 32'h3d8d7187} /* (24, 15, 26) {real, imag} */,
  {32'h3c346ddc, 32'hba97c870} /* (24, 15, 25) {real, imag} */,
  {32'hbdb27213, 32'h3c0540c1} /* (24, 15, 24) {real, imag} */,
  {32'hbb4aa878, 32'hbd86716a} /* (24, 15, 23) {real, imag} */,
  {32'hbc994240, 32'h3c8c96e5} /* (24, 15, 22) {real, imag} */,
  {32'h3cf89af0, 32'h3d108b5a} /* (24, 15, 21) {real, imag} */,
  {32'hbc6fcdda, 32'hbd945a88} /* (24, 15, 20) {real, imag} */,
  {32'h3d3edc34, 32'h3de3a962} /* (24, 15, 19) {real, imag} */,
  {32'h3b0035e0, 32'h3c32447b} /* (24, 15, 18) {real, imag} */,
  {32'h3c97887a, 32'h3c25e40e} /* (24, 15, 17) {real, imag} */,
  {32'hbce7f9f3, 32'h00000000} /* (24, 15, 16) {real, imag} */,
  {32'h3c97887a, 32'hbc25e40e} /* (24, 15, 15) {real, imag} */,
  {32'h3b0035e0, 32'hbc32447b} /* (24, 15, 14) {real, imag} */,
  {32'h3d3edc34, 32'hbde3a962} /* (24, 15, 13) {real, imag} */,
  {32'hbc6fcdda, 32'h3d945a88} /* (24, 15, 12) {real, imag} */,
  {32'h3cf89af0, 32'hbd108b5a} /* (24, 15, 11) {real, imag} */,
  {32'hbc994240, 32'hbc8c96e5} /* (24, 15, 10) {real, imag} */,
  {32'hbb4aa878, 32'h3d86716a} /* (24, 15, 9) {real, imag} */,
  {32'hbdb27213, 32'hbc0540c1} /* (24, 15, 8) {real, imag} */,
  {32'h3c346ddc, 32'h3a97c870} /* (24, 15, 7) {real, imag} */,
  {32'hbbba61f8, 32'hbd8d7187} /* (24, 15, 6) {real, imag} */,
  {32'hbe5db7f2, 32'hbcd1e001} /* (24, 15, 5) {real, imag} */,
  {32'h3e311eca, 32'h3d60824c} /* (24, 15, 4) {real, imag} */,
  {32'hbd6cc200, 32'hbbe2cf40} /* (24, 15, 3) {real, imag} */,
  {32'hbf65b0ca, 32'hbe8776fe} /* (24, 15, 2) {real, imag} */,
  {32'h403350f2, 32'h3e2f4e15} /* (24, 15, 1) {real, imag} */,
  {32'h3fede86d, 32'h00000000} /* (24, 15, 0) {real, imag} */,
  {32'h402b539c, 32'hbdf0d248} /* (24, 14, 31) {real, imag} */,
  {32'hbf8ffb0f, 32'h3e83294c} /* (24, 14, 30) {real, imag} */,
  {32'hbd2b835a, 32'h3dcd469e} /* (24, 14, 29) {real, imag} */,
  {32'h3e25c904, 32'hbe3b8e86} /* (24, 14, 28) {real, imag} */,
  {32'hbe367528, 32'h3d40efc0} /* (24, 14, 27) {real, imag} */,
  {32'hbc1b06a4, 32'h3adf43f0} /* (24, 14, 26) {real, imag} */,
  {32'h3e1049e4, 32'hbd8b63a8} /* (24, 14, 25) {real, imag} */,
  {32'hbce13b08, 32'hbc7fc818} /* (24, 14, 24) {real, imag} */,
  {32'hbcc3528f, 32'h3d86a725} /* (24, 14, 23) {real, imag} */,
  {32'hbd2614c6, 32'h3a066800} /* (24, 14, 22) {real, imag} */,
  {32'h3d5a7ba3, 32'hbcfa3a08} /* (24, 14, 21) {real, imag} */,
  {32'hbd5e6298, 32'hbd49aade} /* (24, 14, 20) {real, imag} */,
  {32'hbbd1d1b8, 32'h3d4ec6f6} /* (24, 14, 19) {real, imag} */,
  {32'h3c548331, 32'h3bca9028} /* (24, 14, 18) {real, imag} */,
  {32'hbcbd1ce9, 32'hbb98adee} /* (24, 14, 17) {real, imag} */,
  {32'h3d6cd196, 32'h00000000} /* (24, 14, 16) {real, imag} */,
  {32'hbcbd1ce9, 32'h3b98adee} /* (24, 14, 15) {real, imag} */,
  {32'h3c548331, 32'hbbca9028} /* (24, 14, 14) {real, imag} */,
  {32'hbbd1d1b8, 32'hbd4ec6f6} /* (24, 14, 13) {real, imag} */,
  {32'hbd5e6298, 32'h3d49aade} /* (24, 14, 12) {real, imag} */,
  {32'h3d5a7ba3, 32'h3cfa3a08} /* (24, 14, 11) {real, imag} */,
  {32'hbd2614c6, 32'hba066800} /* (24, 14, 10) {real, imag} */,
  {32'hbcc3528f, 32'hbd86a725} /* (24, 14, 9) {real, imag} */,
  {32'hbce13b08, 32'h3c7fc818} /* (24, 14, 8) {real, imag} */,
  {32'h3e1049e4, 32'h3d8b63a8} /* (24, 14, 7) {real, imag} */,
  {32'hbc1b06a4, 32'hbadf43f0} /* (24, 14, 6) {real, imag} */,
  {32'hbe367528, 32'hbd40efc0} /* (24, 14, 5) {real, imag} */,
  {32'h3e25c904, 32'h3e3b8e86} /* (24, 14, 4) {real, imag} */,
  {32'hbd2b835a, 32'hbdcd469e} /* (24, 14, 3) {real, imag} */,
  {32'hbf8ffb0f, 32'hbe83294c} /* (24, 14, 2) {real, imag} */,
  {32'h402b539c, 32'h3df0d248} /* (24, 14, 1) {real, imag} */,
  {32'h3fef6213, 32'h00000000} /* (24, 14, 0) {real, imag} */,
  {32'h401829df, 32'h3b6ea200} /* (24, 13, 31) {real, imag} */,
  {32'hbf8e5552, 32'h3e2e2050} /* (24, 13, 30) {real, imag} */,
  {32'hbe2b7ed3, 32'h3d523cbe} /* (24, 13, 29) {real, imag} */,
  {32'h3e1db460, 32'hbe79cf2b} /* (24, 13, 28) {real, imag} */,
  {32'hbe6eac33, 32'h3d587a6a} /* (24, 13, 27) {real, imag} */,
  {32'h3d480351, 32'h3baeefe8} /* (24, 13, 26) {real, imag} */,
  {32'h3df0eaf8, 32'hbc70e155} /* (24, 13, 25) {real, imag} */,
  {32'h3dcae87b, 32'h3afc01c0} /* (24, 13, 24) {real, imag} */,
  {32'hbdb3667a, 32'hbd578ee4} /* (24, 13, 23) {real, imag} */,
  {32'hbc159908, 32'h3d4969ca} /* (24, 13, 22) {real, imag} */,
  {32'h3c84385a, 32'hbc4dc259} /* (24, 13, 21) {real, imag} */,
  {32'hbbe48ec0, 32'hbd7e5bbe} /* (24, 13, 20) {real, imag} */,
  {32'hbba7f430, 32'h3cfb87cc} /* (24, 13, 19) {real, imag} */,
  {32'h3b423038, 32'h3dd9e124} /* (24, 13, 18) {real, imag} */,
  {32'hbc3da112, 32'hbcbbfae0} /* (24, 13, 17) {real, imag} */,
  {32'hbc808992, 32'h00000000} /* (24, 13, 16) {real, imag} */,
  {32'hbc3da112, 32'h3cbbfae0} /* (24, 13, 15) {real, imag} */,
  {32'h3b423038, 32'hbdd9e124} /* (24, 13, 14) {real, imag} */,
  {32'hbba7f430, 32'hbcfb87cc} /* (24, 13, 13) {real, imag} */,
  {32'hbbe48ec0, 32'h3d7e5bbe} /* (24, 13, 12) {real, imag} */,
  {32'h3c84385a, 32'h3c4dc259} /* (24, 13, 11) {real, imag} */,
  {32'hbc159908, 32'hbd4969ca} /* (24, 13, 10) {real, imag} */,
  {32'hbdb3667a, 32'h3d578ee4} /* (24, 13, 9) {real, imag} */,
  {32'h3dcae87b, 32'hbafc01c0} /* (24, 13, 8) {real, imag} */,
  {32'h3df0eaf8, 32'h3c70e155} /* (24, 13, 7) {real, imag} */,
  {32'h3d480351, 32'hbbaeefe8} /* (24, 13, 6) {real, imag} */,
  {32'hbe6eac33, 32'hbd587a6a} /* (24, 13, 5) {real, imag} */,
  {32'h3e1db460, 32'h3e79cf2b} /* (24, 13, 4) {real, imag} */,
  {32'hbe2b7ed3, 32'hbd523cbe} /* (24, 13, 3) {real, imag} */,
  {32'hbf8e5552, 32'hbe2e2050} /* (24, 13, 2) {real, imag} */,
  {32'h401829df, 32'hbb6ea200} /* (24, 13, 1) {real, imag} */,
  {32'h3fd69d05, 32'h00000000} /* (24, 13, 0) {real, imag} */,
  {32'h3ff8daea, 32'h3e580884} /* (24, 12, 31) {real, imag} */,
  {32'hbf83e80d, 32'hbc228a70} /* (24, 12, 30) {real, imag} */,
  {32'hbd38ac65, 32'h3db79bbc} /* (24, 12, 29) {real, imag} */,
  {32'h3e3f00c0, 32'hbdc159c6} /* (24, 12, 28) {real, imag} */,
  {32'hbdd14cd7, 32'h3e36f08b} /* (24, 12, 27) {real, imag} */,
  {32'h3c993c3a, 32'hbd43bbd0} /* (24, 12, 26) {real, imag} */,
  {32'h3ddbc6d6, 32'h3d0c69ad} /* (24, 12, 25) {real, imag} */,
  {32'hbaa31700, 32'h3dccd9f5} /* (24, 12, 24) {real, imag} */,
  {32'hbd825024, 32'hbdd3b99a} /* (24, 12, 23) {real, imag} */,
  {32'hbb1530e8, 32'h3daecf3b} /* (24, 12, 22) {real, imag} */,
  {32'hbbc2a158, 32'h3c9d4822} /* (24, 12, 21) {real, imag} */,
  {32'h3d68cf65, 32'h3d0ac2f2} /* (24, 12, 20) {real, imag} */,
  {32'h3ccc7a48, 32'h3d9af994} /* (24, 12, 19) {real, imag} */,
  {32'hbd442b76, 32'h3de2d434} /* (24, 12, 18) {real, imag} */,
  {32'hbd8e52de, 32'hbdb25341} /* (24, 12, 17) {real, imag} */,
  {32'h3dc6112e, 32'h00000000} /* (24, 12, 16) {real, imag} */,
  {32'hbd8e52de, 32'h3db25341} /* (24, 12, 15) {real, imag} */,
  {32'hbd442b76, 32'hbde2d434} /* (24, 12, 14) {real, imag} */,
  {32'h3ccc7a48, 32'hbd9af994} /* (24, 12, 13) {real, imag} */,
  {32'h3d68cf65, 32'hbd0ac2f2} /* (24, 12, 12) {real, imag} */,
  {32'hbbc2a158, 32'hbc9d4822} /* (24, 12, 11) {real, imag} */,
  {32'hbb1530e8, 32'hbdaecf3b} /* (24, 12, 10) {real, imag} */,
  {32'hbd825024, 32'h3dd3b99a} /* (24, 12, 9) {real, imag} */,
  {32'hbaa31700, 32'hbdccd9f5} /* (24, 12, 8) {real, imag} */,
  {32'h3ddbc6d6, 32'hbd0c69ad} /* (24, 12, 7) {real, imag} */,
  {32'h3c993c3a, 32'h3d43bbd0} /* (24, 12, 6) {real, imag} */,
  {32'hbdd14cd7, 32'hbe36f08b} /* (24, 12, 5) {real, imag} */,
  {32'h3e3f00c0, 32'h3dc159c6} /* (24, 12, 4) {real, imag} */,
  {32'hbd38ac65, 32'hbdb79bbc} /* (24, 12, 3) {real, imag} */,
  {32'hbf83e80d, 32'h3c228a70} /* (24, 12, 2) {real, imag} */,
  {32'h3ff8daea, 32'hbe580884} /* (24, 12, 1) {real, imag} */,
  {32'h3f91b764, 32'h00000000} /* (24, 12, 0) {real, imag} */,
  {32'h3f737814, 32'h3eafe7f0} /* (24, 11, 31) {real, imag} */,
  {32'hbf4caa70, 32'hbd4a9644} /* (24, 11, 30) {real, imag} */,
  {32'hbd1fe157, 32'h3d95eaab} /* (24, 11, 29) {real, imag} */,
  {32'h3e9dc889, 32'hbe698aec} /* (24, 11, 28) {real, imag} */,
  {32'h3b1a3d60, 32'h3d25620e} /* (24, 11, 27) {real, imag} */,
  {32'hbbe6c92a, 32'h3dbf33d4} /* (24, 11, 26) {real, imag} */,
  {32'hbd742053, 32'hbd809547} /* (24, 11, 25) {real, imag} */,
  {32'hbe164b53, 32'h3c23c733} /* (24, 11, 24) {real, imag} */,
  {32'hbda59b85, 32'h3cd1af34} /* (24, 11, 23) {real, imag} */,
  {32'h3cfc0c84, 32'hbc1d2a86} /* (24, 11, 22) {real, imag} */,
  {32'hbc5672e0, 32'h3cccd2d0} /* (24, 11, 21) {real, imag} */,
  {32'h3ca26636, 32'h3dc90a4a} /* (24, 11, 20) {real, imag} */,
  {32'hbd063211, 32'hbcdc5dcb} /* (24, 11, 19) {real, imag} */,
  {32'h3d9854f8, 32'hbb568c68} /* (24, 11, 18) {real, imag} */,
  {32'h3c592489, 32'h3db31826} /* (24, 11, 17) {real, imag} */,
  {32'h3dd2aadc, 32'h00000000} /* (24, 11, 16) {real, imag} */,
  {32'h3c592489, 32'hbdb31826} /* (24, 11, 15) {real, imag} */,
  {32'h3d9854f8, 32'h3b568c68} /* (24, 11, 14) {real, imag} */,
  {32'hbd063211, 32'h3cdc5dcb} /* (24, 11, 13) {real, imag} */,
  {32'h3ca26636, 32'hbdc90a4a} /* (24, 11, 12) {real, imag} */,
  {32'hbc5672e0, 32'hbcccd2d0} /* (24, 11, 11) {real, imag} */,
  {32'h3cfc0c84, 32'h3c1d2a86} /* (24, 11, 10) {real, imag} */,
  {32'hbda59b85, 32'hbcd1af34} /* (24, 11, 9) {real, imag} */,
  {32'hbe164b53, 32'hbc23c733} /* (24, 11, 8) {real, imag} */,
  {32'hbd742053, 32'h3d809547} /* (24, 11, 7) {real, imag} */,
  {32'hbbe6c92a, 32'hbdbf33d4} /* (24, 11, 6) {real, imag} */,
  {32'h3b1a3d60, 32'hbd25620e} /* (24, 11, 5) {real, imag} */,
  {32'h3e9dc889, 32'h3e698aec} /* (24, 11, 4) {real, imag} */,
  {32'hbd1fe157, 32'hbd95eaab} /* (24, 11, 3) {real, imag} */,
  {32'hbf4caa70, 32'h3d4a9644} /* (24, 11, 2) {real, imag} */,
  {32'h3f737814, 32'hbeafe7f0} /* (24, 11, 1) {real, imag} */,
  {32'h3f12fe9f, 32'h00000000} /* (24, 11, 0) {real, imag} */,
  {32'hbf20177b, 32'h3f1a0276} /* (24, 10, 31) {real, imag} */,
  {32'h3b118a80, 32'hbe2c4fe0} /* (24, 10, 30) {real, imag} */,
  {32'hbe0aefaa, 32'h3c636344} /* (24, 10, 29) {real, imag} */,
  {32'h3de5405c, 32'hbdf6b5aa} /* (24, 10, 28) {real, imag} */,
  {32'h3ddca0d3, 32'hbd0645fc} /* (24, 10, 27) {real, imag} */,
  {32'h3d3a0403, 32'h3cc34ff4} /* (24, 10, 26) {real, imag} */,
  {32'h3cfafd5f, 32'h3dfa5e26} /* (24, 10, 25) {real, imag} */,
  {32'h3c9b721e, 32'hbcd186a5} /* (24, 10, 24) {real, imag} */,
  {32'hbd9ff736, 32'h3d01595f} /* (24, 10, 23) {real, imag} */,
  {32'hbcd61b65, 32'hbcb04525} /* (24, 10, 22) {real, imag} */,
  {32'hbd2fe0e4, 32'hbd97c74f} /* (24, 10, 21) {real, imag} */,
  {32'hbdb82a04, 32'hbdbc3c9f} /* (24, 10, 20) {real, imag} */,
  {32'h3ced3bd1, 32'hbe01e6fc} /* (24, 10, 19) {real, imag} */,
  {32'hbc1a3e00, 32'hbd03afe8} /* (24, 10, 18) {real, imag} */,
  {32'hbc282b4a, 32'h3c15f546} /* (24, 10, 17) {real, imag} */,
  {32'hbd7c5456, 32'h00000000} /* (24, 10, 16) {real, imag} */,
  {32'hbc282b4a, 32'hbc15f546} /* (24, 10, 15) {real, imag} */,
  {32'hbc1a3e00, 32'h3d03afe8} /* (24, 10, 14) {real, imag} */,
  {32'h3ced3bd1, 32'h3e01e6fc} /* (24, 10, 13) {real, imag} */,
  {32'hbdb82a04, 32'h3dbc3c9f} /* (24, 10, 12) {real, imag} */,
  {32'hbd2fe0e4, 32'h3d97c74f} /* (24, 10, 11) {real, imag} */,
  {32'hbcd61b65, 32'h3cb04525} /* (24, 10, 10) {real, imag} */,
  {32'hbd9ff736, 32'hbd01595f} /* (24, 10, 9) {real, imag} */,
  {32'h3c9b721e, 32'h3cd186a5} /* (24, 10, 8) {real, imag} */,
  {32'h3cfafd5f, 32'hbdfa5e26} /* (24, 10, 7) {real, imag} */,
  {32'h3d3a0403, 32'hbcc34ff4} /* (24, 10, 6) {real, imag} */,
  {32'h3ddca0d3, 32'h3d0645fc} /* (24, 10, 5) {real, imag} */,
  {32'h3de5405c, 32'h3df6b5aa} /* (24, 10, 4) {real, imag} */,
  {32'hbe0aefaa, 32'hbc636344} /* (24, 10, 3) {real, imag} */,
  {32'h3b118a80, 32'h3e2c4fe0} /* (24, 10, 2) {real, imag} */,
  {32'hbf20177b, 32'hbf1a0276} /* (24, 10, 1) {real, imag} */,
  {32'hbf2c5009, 32'h00000000} /* (24, 10, 0) {real, imag} */,
  {32'hbfda16e0, 32'h3f6db447} /* (24, 9, 31) {real, imag} */,
  {32'h3efa7478, 32'hbe664fb0} /* (24, 9, 30) {real, imag} */,
  {32'hbb4fd310, 32'hbc545974} /* (24, 9, 29) {real, imag} */,
  {32'hbd096680, 32'hbda8f86c} /* (24, 9, 28) {real, imag} */,
  {32'h3dc48646, 32'hbdc9259b} /* (24, 9, 27) {real, imag} */,
  {32'h3d69a4e3, 32'hbc3dba00} /* (24, 9, 26) {real, imag} */,
  {32'h3ca28680, 32'h3c8dc55f} /* (24, 9, 25) {real, imag} */,
  {32'h3d43753c, 32'h3d0b3c6e} /* (24, 9, 24) {real, imag} */,
  {32'h3d959758, 32'h3d9a5656} /* (24, 9, 23) {real, imag} */,
  {32'h3d0e4db9, 32'hbcc55b13} /* (24, 9, 22) {real, imag} */,
  {32'hbdd927e0, 32'hbd8afc1a} /* (24, 9, 21) {real, imag} */,
  {32'hbd3e5ae1, 32'h3d1f27ac} /* (24, 9, 20) {real, imag} */,
  {32'h3cd62d26, 32'hbda06cf2} /* (24, 9, 19) {real, imag} */,
  {32'h3db5f3ed, 32'h39e0b820} /* (24, 9, 18) {real, imag} */,
  {32'hbc910b40, 32'hbcdd3b35} /* (24, 9, 17) {real, imag} */,
  {32'h3d5f535b, 32'h00000000} /* (24, 9, 16) {real, imag} */,
  {32'hbc910b40, 32'h3cdd3b35} /* (24, 9, 15) {real, imag} */,
  {32'h3db5f3ed, 32'hb9e0b820} /* (24, 9, 14) {real, imag} */,
  {32'h3cd62d26, 32'h3da06cf2} /* (24, 9, 13) {real, imag} */,
  {32'hbd3e5ae1, 32'hbd1f27ac} /* (24, 9, 12) {real, imag} */,
  {32'hbdd927e0, 32'h3d8afc1a} /* (24, 9, 11) {real, imag} */,
  {32'h3d0e4db9, 32'h3cc55b13} /* (24, 9, 10) {real, imag} */,
  {32'h3d959758, 32'hbd9a5656} /* (24, 9, 9) {real, imag} */,
  {32'h3d43753c, 32'hbd0b3c6e} /* (24, 9, 8) {real, imag} */,
  {32'h3ca28680, 32'hbc8dc55f} /* (24, 9, 7) {real, imag} */,
  {32'h3d69a4e3, 32'h3c3dba00} /* (24, 9, 6) {real, imag} */,
  {32'h3dc48646, 32'h3dc9259b} /* (24, 9, 5) {real, imag} */,
  {32'hbd096680, 32'h3da8f86c} /* (24, 9, 4) {real, imag} */,
  {32'hbb4fd310, 32'h3c545974} /* (24, 9, 3) {real, imag} */,
  {32'h3efa7478, 32'h3e664fb0} /* (24, 9, 2) {real, imag} */,
  {32'hbfda16e0, 32'hbf6db447} /* (24, 9, 1) {real, imag} */,
  {32'hbfe9481b, 32'h00000000} /* (24, 9, 0) {real, imag} */,
  {32'hc0120b28, 32'h3f94d9d1} /* (24, 8, 31) {real, imag} */,
  {32'h3f358c36, 32'hbeb9d678} /* (24, 8, 30) {real, imag} */,
  {32'h3e057e3d, 32'h3db31102} /* (24, 8, 29) {real, imag} */,
  {32'hbe172f33, 32'h3d2293fd} /* (24, 8, 28) {real, imag} */,
  {32'h3c4930e8, 32'hbe401e0b} /* (24, 8, 27) {real, imag} */,
  {32'h3d9d4416, 32'hbe09385a} /* (24, 8, 26) {real, imag} */,
  {32'h3d7bb1c4, 32'hbde3f329} /* (24, 8, 25) {real, imag} */,
  {32'h3dec11df, 32'hbd413328} /* (24, 8, 24) {real, imag} */,
  {32'hbdcc06ff, 32'h3cf6c6a2} /* (24, 8, 23) {real, imag} */,
  {32'h3cc62402, 32'h3c011420} /* (24, 8, 22) {real, imag} */,
  {32'h3d8af28d, 32'h3d5d1ac0} /* (24, 8, 21) {real, imag} */,
  {32'h3d699ed9, 32'h3cd14e1a} /* (24, 8, 20) {real, imag} */,
  {32'h3c50f1d9, 32'h3d8fc793} /* (24, 8, 19) {real, imag} */,
  {32'h3d63903c, 32'h3c1ccfe8} /* (24, 8, 18) {real, imag} */,
  {32'h3d4e1ea9, 32'h3d40c937} /* (24, 8, 17) {real, imag} */,
  {32'h3bc1ffb0, 32'h00000000} /* (24, 8, 16) {real, imag} */,
  {32'h3d4e1ea9, 32'hbd40c937} /* (24, 8, 15) {real, imag} */,
  {32'h3d63903c, 32'hbc1ccfe8} /* (24, 8, 14) {real, imag} */,
  {32'h3c50f1d9, 32'hbd8fc793} /* (24, 8, 13) {real, imag} */,
  {32'h3d699ed9, 32'hbcd14e1a} /* (24, 8, 12) {real, imag} */,
  {32'h3d8af28d, 32'hbd5d1ac0} /* (24, 8, 11) {real, imag} */,
  {32'h3cc62402, 32'hbc011420} /* (24, 8, 10) {real, imag} */,
  {32'hbdcc06ff, 32'hbcf6c6a2} /* (24, 8, 9) {real, imag} */,
  {32'h3dec11df, 32'h3d413328} /* (24, 8, 8) {real, imag} */,
  {32'h3d7bb1c4, 32'h3de3f329} /* (24, 8, 7) {real, imag} */,
  {32'h3d9d4416, 32'h3e09385a} /* (24, 8, 6) {real, imag} */,
  {32'h3c4930e8, 32'h3e401e0b} /* (24, 8, 5) {real, imag} */,
  {32'hbe172f33, 32'hbd2293fd} /* (24, 8, 4) {real, imag} */,
  {32'h3e057e3d, 32'hbdb31102} /* (24, 8, 3) {real, imag} */,
  {32'h3f358c36, 32'h3eb9d678} /* (24, 8, 2) {real, imag} */,
  {32'hc0120b28, 32'hbf94d9d1} /* (24, 8, 1) {real, imag} */,
  {32'hc021628e, 32'h00000000} /* (24, 8, 0) {real, imag} */,
  {32'hc025ab9f, 32'h3fb5c158} /* (24, 7, 31) {real, imag} */,
  {32'h3f27217a, 32'hbe9e61da} /* (24, 7, 30) {real, imag} */,
  {32'h3dd9cb72, 32'hbce7881b} /* (24, 7, 29) {real, imag} */,
  {32'hbe63e172, 32'h3ca9675f} /* (24, 7, 28) {real, imag} */,
  {32'h3e2783c2, 32'hbd0f7239} /* (24, 7, 27) {real, imag} */,
  {32'h3daaa0a8, 32'hbd48f723} /* (24, 7, 26) {real, imag} */,
  {32'hbe03b5e0, 32'hbc8b736e} /* (24, 7, 25) {real, imag} */,
  {32'h3ddb72c5, 32'hbd5ee4e6} /* (24, 7, 24) {real, imag} */,
  {32'hbd301335, 32'hbd41aa24} /* (24, 7, 23) {real, imag} */,
  {32'h3dcc6190, 32'h3da2e487} /* (24, 7, 22) {real, imag} */,
  {32'h3c383a18, 32'hbdb0168f} /* (24, 7, 21) {real, imag} */,
  {32'hbde2ad8a, 32'hbd4480e8} /* (24, 7, 20) {real, imag} */,
  {32'h3d286b2c, 32'hbc376a54} /* (24, 7, 19) {real, imag} */,
  {32'h3b1d7f90, 32'hbce69474} /* (24, 7, 18) {real, imag} */,
  {32'hbcd378e9, 32'hbc41af1d} /* (24, 7, 17) {real, imag} */,
  {32'h3b96d75c, 32'h00000000} /* (24, 7, 16) {real, imag} */,
  {32'hbcd378e9, 32'h3c41af1d} /* (24, 7, 15) {real, imag} */,
  {32'h3b1d7f90, 32'h3ce69474} /* (24, 7, 14) {real, imag} */,
  {32'h3d286b2c, 32'h3c376a54} /* (24, 7, 13) {real, imag} */,
  {32'hbde2ad8a, 32'h3d4480e8} /* (24, 7, 12) {real, imag} */,
  {32'h3c383a18, 32'h3db0168f} /* (24, 7, 11) {real, imag} */,
  {32'h3dcc6190, 32'hbda2e487} /* (24, 7, 10) {real, imag} */,
  {32'hbd301335, 32'h3d41aa24} /* (24, 7, 9) {real, imag} */,
  {32'h3ddb72c5, 32'h3d5ee4e6} /* (24, 7, 8) {real, imag} */,
  {32'hbe03b5e0, 32'h3c8b736e} /* (24, 7, 7) {real, imag} */,
  {32'h3daaa0a8, 32'h3d48f723} /* (24, 7, 6) {real, imag} */,
  {32'h3e2783c2, 32'h3d0f7239} /* (24, 7, 5) {real, imag} */,
  {32'hbe63e172, 32'hbca9675f} /* (24, 7, 4) {real, imag} */,
  {32'h3dd9cb72, 32'h3ce7881b} /* (24, 7, 3) {real, imag} */,
  {32'h3f27217a, 32'h3e9e61da} /* (24, 7, 2) {real, imag} */,
  {32'hc025ab9f, 32'hbfb5c158} /* (24, 7, 1) {real, imag} */,
  {32'hc0483cf8, 32'h00000000} /* (24, 7, 0) {real, imag} */,
  {32'hc02d7c4b, 32'h3fe36498} /* (24, 6, 31) {real, imag} */,
  {32'h3f297ff7, 32'hbed00429} /* (24, 6, 30) {real, imag} */,
  {32'hbcdf437e, 32'hbcbe778e} /* (24, 6, 29) {real, imag} */,
  {32'hbe3e3cb6, 32'hbc774d84} /* (24, 6, 28) {real, imag} */,
  {32'h3e53fbe0, 32'hbe05979f} /* (24, 6, 27) {real, imag} */,
  {32'h3acc3b30, 32'hbe15ff8a} /* (24, 6, 26) {real, imag} */,
  {32'h3cb7afa4, 32'hbda095a8} /* (24, 6, 25) {real, imag} */,
  {32'h3bd961c8, 32'hbb891d64} /* (24, 6, 24) {real, imag} */,
  {32'hbd108e16, 32'hbd37cbd8} /* (24, 6, 23) {real, imag} */,
  {32'hbd0604dc, 32'hbc6bfcec} /* (24, 6, 22) {real, imag} */,
  {32'h3c032135, 32'h3cf6fa0d} /* (24, 6, 21) {real, imag} */,
  {32'hbd1de002, 32'h3d0bfa8a} /* (24, 6, 20) {real, imag} */,
  {32'h3d0b5fc0, 32'hbc0b0ad6} /* (24, 6, 19) {real, imag} */,
  {32'h3d599a0b, 32'hbd52eac3} /* (24, 6, 18) {real, imag} */,
  {32'hbcbf6214, 32'h3bca4ef8} /* (24, 6, 17) {real, imag} */,
  {32'hba9f3380, 32'h00000000} /* (24, 6, 16) {real, imag} */,
  {32'hbcbf6214, 32'hbbca4ef8} /* (24, 6, 15) {real, imag} */,
  {32'h3d599a0b, 32'h3d52eac3} /* (24, 6, 14) {real, imag} */,
  {32'h3d0b5fc0, 32'h3c0b0ad6} /* (24, 6, 13) {real, imag} */,
  {32'hbd1de002, 32'hbd0bfa8a} /* (24, 6, 12) {real, imag} */,
  {32'h3c032135, 32'hbcf6fa0d} /* (24, 6, 11) {real, imag} */,
  {32'hbd0604dc, 32'h3c6bfcec} /* (24, 6, 10) {real, imag} */,
  {32'hbd108e16, 32'h3d37cbd8} /* (24, 6, 9) {real, imag} */,
  {32'h3bd961c8, 32'h3b891d64} /* (24, 6, 8) {real, imag} */,
  {32'h3cb7afa4, 32'h3da095a8} /* (24, 6, 7) {real, imag} */,
  {32'h3acc3b30, 32'h3e15ff8a} /* (24, 6, 6) {real, imag} */,
  {32'h3e53fbe0, 32'h3e05979f} /* (24, 6, 5) {real, imag} */,
  {32'hbe3e3cb6, 32'h3c774d84} /* (24, 6, 4) {real, imag} */,
  {32'hbcdf437e, 32'h3cbe778e} /* (24, 6, 3) {real, imag} */,
  {32'h3f297ff7, 32'h3ed00429} /* (24, 6, 2) {real, imag} */,
  {32'hc02d7c4b, 32'hbfe36498} /* (24, 6, 1) {real, imag} */,
  {32'hc068ad58, 32'h00000000} /* (24, 6, 0) {real, imag} */,
  {32'hc029762e, 32'h4018d1a0} /* (24, 5, 31) {real, imag} */,
  {32'h3e44db00, 32'hbf0e0164} /* (24, 5, 30) {real, imag} */,
  {32'h3d83a1b9, 32'h3dddfcda} /* (24, 5, 29) {real, imag} */,
  {32'h3d482ec3, 32'hbde16640} /* (24, 5, 28) {real, imag} */,
  {32'h3dc92f2f, 32'h3d0600aa} /* (24, 5, 27) {real, imag} */,
  {32'h3d2cdf03, 32'hbdab1632} /* (24, 5, 26) {real, imag} */,
  {32'h3ce08bed, 32'h3dc41014} /* (24, 5, 25) {real, imag} */,
  {32'hbccc6c56, 32'hbdcf58b9} /* (24, 5, 24) {real, imag} */,
  {32'hbda57ef7, 32'h3d4cb4b9} /* (24, 5, 23) {real, imag} */,
  {32'h3b4efe90, 32'hbc2c5682} /* (24, 5, 22) {real, imag} */,
  {32'hbd906629, 32'h3bd06462} /* (24, 5, 21) {real, imag} */,
  {32'hbc3fc0f6, 32'hbd36d0b0} /* (24, 5, 20) {real, imag} */,
  {32'h3cd56f9a, 32'hbc80284e} /* (24, 5, 19) {real, imag} */,
  {32'hbd5eda3c, 32'hbd4df555} /* (24, 5, 18) {real, imag} */,
  {32'h3c65a7e9, 32'h3c369d0e} /* (24, 5, 17) {real, imag} */,
  {32'h3dc549e4, 32'h00000000} /* (24, 5, 16) {real, imag} */,
  {32'h3c65a7e9, 32'hbc369d0e} /* (24, 5, 15) {real, imag} */,
  {32'hbd5eda3c, 32'h3d4df555} /* (24, 5, 14) {real, imag} */,
  {32'h3cd56f9a, 32'h3c80284e} /* (24, 5, 13) {real, imag} */,
  {32'hbc3fc0f6, 32'h3d36d0b0} /* (24, 5, 12) {real, imag} */,
  {32'hbd906629, 32'hbbd06462} /* (24, 5, 11) {real, imag} */,
  {32'h3b4efe90, 32'h3c2c5682} /* (24, 5, 10) {real, imag} */,
  {32'hbda57ef7, 32'hbd4cb4b9} /* (24, 5, 9) {real, imag} */,
  {32'hbccc6c56, 32'h3dcf58b9} /* (24, 5, 8) {real, imag} */,
  {32'h3ce08bed, 32'hbdc41014} /* (24, 5, 7) {real, imag} */,
  {32'h3d2cdf03, 32'h3dab1632} /* (24, 5, 6) {real, imag} */,
  {32'h3dc92f2f, 32'hbd0600aa} /* (24, 5, 5) {real, imag} */,
  {32'h3d482ec3, 32'h3de16640} /* (24, 5, 4) {real, imag} */,
  {32'h3d83a1b9, 32'hbdddfcda} /* (24, 5, 3) {real, imag} */,
  {32'h3e44db00, 32'h3f0e0164} /* (24, 5, 2) {real, imag} */,
  {32'hc029762e, 32'hc018d1a0} /* (24, 5, 1) {real, imag} */,
  {32'hc074b4a2, 32'h00000000} /* (24, 5, 0) {real, imag} */,
  {32'hc01be12b, 32'h40365fc3} /* (24, 4, 31) {real, imag} */,
  {32'hbe3e7ff2, 32'hbf2f99b4} /* (24, 4, 30) {real, imag} */,
  {32'h3d438419, 32'h3c8f85d0} /* (24, 4, 29) {real, imag} */,
  {32'h3e1a6a40, 32'hbe4a9325} /* (24, 4, 28) {real, imag} */,
  {32'h3dd5d8d2, 32'h3df5190e} /* (24, 4, 27) {real, imag} */,
  {32'h3c9b5f3c, 32'hbd078d0a} /* (24, 4, 26) {real, imag} */,
  {32'h3d8b0a4c, 32'h3d9e76fd} /* (24, 4, 25) {real, imag} */,
  {32'hbba9b418, 32'hbdaed402} /* (24, 4, 24) {real, imag} */,
  {32'h3c821958, 32'h3cc284d5} /* (24, 4, 23) {real, imag} */,
  {32'h3cee1007, 32'hbd9e6c92} /* (24, 4, 22) {real, imag} */,
  {32'h3d5bac2f, 32'h3d240a6f} /* (24, 4, 21) {real, imag} */,
  {32'hbd5f6f48, 32'hbc27c0d8} /* (24, 4, 20) {real, imag} */,
  {32'h3d69104d, 32'hbd0fac2a} /* (24, 4, 19) {real, imag} */,
  {32'hbca6d41b, 32'hbc90e688} /* (24, 4, 18) {real, imag} */,
  {32'h3c7fa104, 32'hbd8946ec} /* (24, 4, 17) {real, imag} */,
  {32'hbc463f2e, 32'h00000000} /* (24, 4, 16) {real, imag} */,
  {32'h3c7fa104, 32'h3d8946ec} /* (24, 4, 15) {real, imag} */,
  {32'hbca6d41b, 32'h3c90e688} /* (24, 4, 14) {real, imag} */,
  {32'h3d69104d, 32'h3d0fac2a} /* (24, 4, 13) {real, imag} */,
  {32'hbd5f6f48, 32'h3c27c0d8} /* (24, 4, 12) {real, imag} */,
  {32'h3d5bac2f, 32'hbd240a6f} /* (24, 4, 11) {real, imag} */,
  {32'h3cee1007, 32'h3d9e6c92} /* (24, 4, 10) {real, imag} */,
  {32'h3c821958, 32'hbcc284d5} /* (24, 4, 9) {real, imag} */,
  {32'hbba9b418, 32'h3daed402} /* (24, 4, 8) {real, imag} */,
  {32'h3d8b0a4c, 32'hbd9e76fd} /* (24, 4, 7) {real, imag} */,
  {32'h3c9b5f3c, 32'h3d078d0a} /* (24, 4, 6) {real, imag} */,
  {32'h3dd5d8d2, 32'hbdf5190e} /* (24, 4, 5) {real, imag} */,
  {32'h3e1a6a40, 32'h3e4a9325} /* (24, 4, 4) {real, imag} */,
  {32'h3d438419, 32'hbc8f85d0} /* (24, 4, 3) {real, imag} */,
  {32'hbe3e7ff2, 32'h3f2f99b4} /* (24, 4, 2) {real, imag} */,
  {32'hc01be12b, 32'hc0365fc3} /* (24, 4, 1) {real, imag} */,
  {32'hc0833a5b, 32'h00000000} /* (24, 4, 0) {real, imag} */,
  {32'hc0238008, 32'h403edb8f} /* (24, 3, 31) {real, imag} */,
  {32'hbe5f5336, 32'hbf387f7e} /* (24, 3, 30) {real, imag} */,
  {32'h3e281676, 32'h3d7b49ba} /* (24, 3, 29) {real, imag} */,
  {32'h3e0217c1, 32'hbe6c8b05} /* (24, 3, 28) {real, imag} */,
  {32'h3e8b292f, 32'h3d346cca} /* (24, 3, 27) {real, imag} */,
  {32'hbe094730, 32'hbd19d18f} /* (24, 3, 26) {real, imag} */,
  {32'hbc8b7cbe, 32'hbda15589} /* (24, 3, 25) {real, imag} */,
  {32'hbda67fa5, 32'hbc7ddcf8} /* (24, 3, 24) {real, imag} */,
  {32'hbd4e08a7, 32'hbc9d3b29} /* (24, 3, 23) {real, imag} */,
  {32'h3dbc324c, 32'hbd7a29f0} /* (24, 3, 22) {real, imag} */,
  {32'h3da5192e, 32'h3c93b07e} /* (24, 3, 21) {real, imag} */,
  {32'hba40d380, 32'hbcc8cecb} /* (24, 3, 20) {real, imag} */,
  {32'h3d418abf, 32'h3dab122c} /* (24, 3, 19) {real, imag} */,
  {32'h3c14f4f8, 32'h3cefb27a} /* (24, 3, 18) {real, imag} */,
  {32'h3c200f5e, 32'hbd06d758} /* (24, 3, 17) {real, imag} */,
  {32'hbd2a9c5a, 32'h00000000} /* (24, 3, 16) {real, imag} */,
  {32'h3c200f5e, 32'h3d06d758} /* (24, 3, 15) {real, imag} */,
  {32'h3c14f4f8, 32'hbcefb27a} /* (24, 3, 14) {real, imag} */,
  {32'h3d418abf, 32'hbdab122c} /* (24, 3, 13) {real, imag} */,
  {32'hba40d380, 32'h3cc8cecb} /* (24, 3, 12) {real, imag} */,
  {32'h3da5192e, 32'hbc93b07e} /* (24, 3, 11) {real, imag} */,
  {32'h3dbc324c, 32'h3d7a29f0} /* (24, 3, 10) {real, imag} */,
  {32'hbd4e08a7, 32'h3c9d3b29} /* (24, 3, 9) {real, imag} */,
  {32'hbda67fa5, 32'h3c7ddcf8} /* (24, 3, 8) {real, imag} */,
  {32'hbc8b7cbe, 32'h3da15589} /* (24, 3, 7) {real, imag} */,
  {32'hbe094730, 32'h3d19d18f} /* (24, 3, 6) {real, imag} */,
  {32'h3e8b292f, 32'hbd346cca} /* (24, 3, 5) {real, imag} */,
  {32'h3e0217c1, 32'h3e6c8b05} /* (24, 3, 4) {real, imag} */,
  {32'h3e281676, 32'hbd7b49ba} /* (24, 3, 3) {real, imag} */,
  {32'hbe5f5336, 32'h3f387f7e} /* (24, 3, 2) {real, imag} */,
  {32'hc0238008, 32'hc03edb8f} /* (24, 3, 1) {real, imag} */,
  {32'hc082a3e5, 32'h00000000} /* (24, 3, 0) {real, imag} */,
  {32'hc01b7da7, 32'h4040b43a} /* (24, 2, 31) {real, imag} */,
  {32'hbeaad732, 32'hbf3c44ed} /* (24, 2, 30) {real, imag} */,
  {32'h3e7366df, 32'h3d4b66f0} /* (24, 2, 29) {real, imag} */,
  {32'h3dd67e20, 32'hbe987288} /* (24, 2, 28) {real, imag} */,
  {32'h3e062c0e, 32'hb9c24480} /* (24, 2, 27) {real, imag} */,
  {32'h3d621a5d, 32'h3d6a50ec} /* (24, 2, 26) {real, imag} */,
  {32'hbc3ed094, 32'h3d2de2ba} /* (24, 2, 25) {real, imag} */,
  {32'h3cb19444, 32'h3d3a73e2} /* (24, 2, 24) {real, imag} */,
  {32'hbd0e006a, 32'hbcf3e03a} /* (24, 2, 23) {real, imag} */,
  {32'h3d823ff8, 32'hbda2f2bc} /* (24, 2, 22) {real, imag} */,
  {32'h3d40bbd9, 32'h3a384200} /* (24, 2, 21) {real, imag} */,
  {32'hbd8c6d56, 32'hbdaa61ed} /* (24, 2, 20) {real, imag} */,
  {32'h3d8c5d05, 32'h3c299172} /* (24, 2, 19) {real, imag} */,
  {32'hbcf5eebe, 32'h3cd49d58} /* (24, 2, 18) {real, imag} */,
  {32'hbd1e84d6, 32'h3cb4dd0c} /* (24, 2, 17) {real, imag} */,
  {32'h3ca0a15c, 32'h00000000} /* (24, 2, 16) {real, imag} */,
  {32'hbd1e84d6, 32'hbcb4dd0c} /* (24, 2, 15) {real, imag} */,
  {32'hbcf5eebe, 32'hbcd49d58} /* (24, 2, 14) {real, imag} */,
  {32'h3d8c5d05, 32'hbc299172} /* (24, 2, 13) {real, imag} */,
  {32'hbd8c6d56, 32'h3daa61ed} /* (24, 2, 12) {real, imag} */,
  {32'h3d40bbd9, 32'hba384200} /* (24, 2, 11) {real, imag} */,
  {32'h3d823ff8, 32'h3da2f2bc} /* (24, 2, 10) {real, imag} */,
  {32'hbd0e006a, 32'h3cf3e03a} /* (24, 2, 9) {real, imag} */,
  {32'h3cb19444, 32'hbd3a73e2} /* (24, 2, 8) {real, imag} */,
  {32'hbc3ed094, 32'hbd2de2ba} /* (24, 2, 7) {real, imag} */,
  {32'h3d621a5d, 32'hbd6a50ec} /* (24, 2, 6) {real, imag} */,
  {32'h3e062c0e, 32'h39c24480} /* (24, 2, 5) {real, imag} */,
  {32'h3dd67e20, 32'h3e987288} /* (24, 2, 4) {real, imag} */,
  {32'h3e7366df, 32'hbd4b66f0} /* (24, 2, 3) {real, imag} */,
  {32'hbeaad732, 32'h3f3c44ed} /* (24, 2, 2) {real, imag} */,
  {32'hc01b7da7, 32'hc040b43a} /* (24, 2, 1) {real, imag} */,
  {32'hc0822409, 32'h00000000} /* (24, 2, 0) {real, imag} */,
  {32'hc0226249, 32'h40307d30} /* (24, 1, 31) {real, imag} */,
  {32'hbe1e8a3a, 32'hbf21ecfd} /* (24, 1, 30) {real, imag} */,
  {32'h3e86286e, 32'hb83cb500} /* (24, 1, 29) {real, imag} */,
  {32'h3e2f59be, 32'hbe8a8ae6} /* (24, 1, 28) {real, imag} */,
  {32'h3dab3f0f, 32'h3c28539e} /* (24, 1, 27) {real, imag} */,
  {32'h3cdcb41e, 32'hbd5cffea} /* (24, 1, 26) {real, imag} */,
  {32'hbd8cf9e0, 32'h3da427ca} /* (24, 1, 25) {real, imag} */,
  {32'h3d1cd6d2, 32'hbd84e8a2} /* (24, 1, 24) {real, imag} */,
  {32'h3d16ece6, 32'hbcc7340f} /* (24, 1, 23) {real, imag} */,
  {32'hbc84cd0a, 32'h3d01762e} /* (24, 1, 22) {real, imag} */,
  {32'h3bf04446, 32'hbd017486} /* (24, 1, 21) {real, imag} */,
  {32'hbd21dec0, 32'h3ce3c560} /* (24, 1, 20) {real, imag} */,
  {32'hbc0541b0, 32'h3d24ac5f} /* (24, 1, 19) {real, imag} */,
  {32'h3c8700c8, 32'hbdaba606} /* (24, 1, 18) {real, imag} */,
  {32'h3ca79a98, 32'h3dba9d8f} /* (24, 1, 17) {real, imag} */,
  {32'h3d14b840, 32'h00000000} /* (24, 1, 16) {real, imag} */,
  {32'h3ca79a98, 32'hbdba9d8f} /* (24, 1, 15) {real, imag} */,
  {32'h3c8700c8, 32'h3daba606} /* (24, 1, 14) {real, imag} */,
  {32'hbc0541b0, 32'hbd24ac5f} /* (24, 1, 13) {real, imag} */,
  {32'hbd21dec0, 32'hbce3c560} /* (24, 1, 12) {real, imag} */,
  {32'h3bf04446, 32'h3d017486} /* (24, 1, 11) {real, imag} */,
  {32'hbc84cd0a, 32'hbd01762e} /* (24, 1, 10) {real, imag} */,
  {32'h3d16ece6, 32'h3cc7340f} /* (24, 1, 9) {real, imag} */,
  {32'h3d1cd6d2, 32'h3d84e8a2} /* (24, 1, 8) {real, imag} */,
  {32'hbd8cf9e0, 32'hbda427ca} /* (24, 1, 7) {real, imag} */,
  {32'h3cdcb41e, 32'h3d5cffea} /* (24, 1, 6) {real, imag} */,
  {32'h3dab3f0f, 32'hbc28539e} /* (24, 1, 5) {real, imag} */,
  {32'h3e2f59be, 32'h3e8a8ae6} /* (24, 1, 4) {real, imag} */,
  {32'h3e86286e, 32'h383cb500} /* (24, 1, 3) {real, imag} */,
  {32'hbe1e8a3a, 32'h3f21ecfd} /* (24, 1, 2) {real, imag} */,
  {32'hc0226249, 32'hc0307d30} /* (24, 1, 1) {real, imag} */,
  {32'hc082bb5c, 32'h00000000} /* (24, 1, 0) {real, imag} */,
  {32'hc02de981, 32'h400b29c4} /* (24, 0, 31) {real, imag} */,
  {32'h3de7727c, 32'hbe9a0146} /* (24, 0, 30) {real, imag} */,
  {32'h3e2e5ae1, 32'hbc6b19f6} /* (24, 0, 29) {real, imag} */,
  {32'h3ddfdf48, 32'hbe18cb4e} /* (24, 0, 28) {real, imag} */,
  {32'h3dbb7a74, 32'h3cb839ad} /* (24, 0, 27) {real, imag} */,
  {32'hbd0d0566, 32'hbc300c6e} /* (24, 0, 26) {real, imag} */,
  {32'hbc835108, 32'hbc149e6e} /* (24, 0, 25) {real, imag} */,
  {32'h3c9f58a8, 32'h3c0c63c8} /* (24, 0, 24) {real, imag} */,
  {32'h3d824eb6, 32'hbcea97bc} /* (24, 0, 23) {real, imag} */,
  {32'hbdc26272, 32'hbc0f9be4} /* (24, 0, 22) {real, imag} */,
  {32'h3bc65739, 32'hbcded516} /* (24, 0, 21) {real, imag} */,
  {32'h3b5bcb92, 32'h3cd630cd} /* (24, 0, 20) {real, imag} */,
  {32'h3bd7a88e, 32'h3d0a2924} /* (24, 0, 19) {real, imag} */,
  {32'hbc4b34b7, 32'hbbc04b2a} /* (24, 0, 18) {real, imag} */,
  {32'hbd1c984d, 32'hbbed79ec} /* (24, 0, 17) {real, imag} */,
  {32'h3d2190b2, 32'h00000000} /* (24, 0, 16) {real, imag} */,
  {32'hbd1c984d, 32'h3bed79ec} /* (24, 0, 15) {real, imag} */,
  {32'hbc4b34b7, 32'h3bc04b2a} /* (24, 0, 14) {real, imag} */,
  {32'h3bd7a88e, 32'hbd0a2924} /* (24, 0, 13) {real, imag} */,
  {32'h3b5bcb92, 32'hbcd630cd} /* (24, 0, 12) {real, imag} */,
  {32'h3bc65739, 32'h3cded516} /* (24, 0, 11) {real, imag} */,
  {32'hbdc26272, 32'h3c0f9be4} /* (24, 0, 10) {real, imag} */,
  {32'h3d824eb6, 32'h3cea97bc} /* (24, 0, 9) {real, imag} */,
  {32'h3c9f58a8, 32'hbc0c63c8} /* (24, 0, 8) {real, imag} */,
  {32'hbc835108, 32'h3c149e6e} /* (24, 0, 7) {real, imag} */,
  {32'hbd0d0566, 32'h3c300c6e} /* (24, 0, 6) {real, imag} */,
  {32'h3dbb7a74, 32'hbcb839ad} /* (24, 0, 5) {real, imag} */,
  {32'h3ddfdf48, 32'h3e18cb4e} /* (24, 0, 4) {real, imag} */,
  {32'h3e2e5ae1, 32'h3c6b19f6} /* (24, 0, 3) {real, imag} */,
  {32'h3de7727c, 32'h3e9a0146} /* (24, 0, 2) {real, imag} */,
  {32'hc02de981, 32'hc00b29c4} /* (24, 0, 1) {real, imag} */,
  {32'hc080ece3, 32'h00000000} /* (24, 0, 0) {real, imag} */,
  {32'hc067ece0, 32'h40048bc6} /* (23, 31, 31) {real, imag} */,
  {32'h3f34a48c, 32'hbea15588} /* (23, 31, 30) {real, imag} */,
  {32'h3d85f1cd, 32'h3c2b7f4a} /* (23, 31, 29) {real, imag} */,
  {32'hbdde2430, 32'hbc8e2e40} /* (23, 31, 28) {real, imag} */,
  {32'h3dfb60a4, 32'h3c0f0c06} /* (23, 31, 27) {real, imag} */,
  {32'h3b4cc460, 32'h3d251112} /* (23, 31, 26) {real, imag} */,
  {32'hbd220f2c, 32'h3d8f8000} /* (23, 31, 25) {real, imag} */,
  {32'h3dbefa4f, 32'hbd36c5ca} /* (23, 31, 24) {real, imag} */,
  {32'hbb1e2440, 32'hbdf13846} /* (23, 31, 23) {real, imag} */,
  {32'hbd34127e, 32'h3d896780} /* (23, 31, 22) {real, imag} */,
  {32'h3d393498, 32'h3bfde72c} /* (23, 31, 21) {real, imag} */,
  {32'hbd5ffae4, 32'hbcda5f19} /* (23, 31, 20) {real, imag} */,
  {32'h3d192f2e, 32'hbc597fb1} /* (23, 31, 19) {real, imag} */,
  {32'h3d1d7fb8, 32'hbd61bdc7} /* (23, 31, 18) {real, imag} */,
  {32'hbc2a9538, 32'h3bb7dd0c} /* (23, 31, 17) {real, imag} */,
  {32'hbd8bf111, 32'h00000000} /* (23, 31, 16) {real, imag} */,
  {32'hbc2a9538, 32'hbbb7dd0c} /* (23, 31, 15) {real, imag} */,
  {32'h3d1d7fb8, 32'h3d61bdc7} /* (23, 31, 14) {real, imag} */,
  {32'h3d192f2e, 32'h3c597fb1} /* (23, 31, 13) {real, imag} */,
  {32'hbd5ffae4, 32'h3cda5f19} /* (23, 31, 12) {real, imag} */,
  {32'h3d393498, 32'hbbfde72c} /* (23, 31, 11) {real, imag} */,
  {32'hbd34127e, 32'hbd896780} /* (23, 31, 10) {real, imag} */,
  {32'hbb1e2440, 32'h3df13846} /* (23, 31, 9) {real, imag} */,
  {32'h3dbefa4f, 32'h3d36c5ca} /* (23, 31, 8) {real, imag} */,
  {32'hbd220f2c, 32'hbd8f8000} /* (23, 31, 7) {real, imag} */,
  {32'h3b4cc460, 32'hbd251112} /* (23, 31, 6) {real, imag} */,
  {32'h3dfb60a4, 32'hbc0f0c06} /* (23, 31, 5) {real, imag} */,
  {32'hbdde2430, 32'h3c8e2e40} /* (23, 31, 4) {real, imag} */,
  {32'h3d85f1cd, 32'hbc2b7f4a} /* (23, 31, 3) {real, imag} */,
  {32'h3f34a48c, 32'h3ea15588} /* (23, 31, 2) {real, imag} */,
  {32'hc067ece0, 32'hc0048bc6} /* (23, 31, 1) {real, imag} */,
  {32'hc097c953, 32'h00000000} /* (23, 31, 0) {real, imag} */,
  {32'hc082658f, 32'h3fe7d93c} /* (23, 30, 31) {real, imag} */,
  {32'h3f8ed35d, 32'hbe99c8b5} /* (23, 30, 30) {real, imag} */,
  {32'h3d402462, 32'hbd427d0c} /* (23, 30, 29) {real, imag} */,
  {32'hbe39d63e, 32'h3da0cae8} /* (23, 30, 28) {real, imag} */,
  {32'h3e53f456, 32'hbdb50f5f} /* (23, 30, 27) {real, imag} */,
  {32'h3e227f6b, 32'h3db35a1e} /* (23, 30, 26) {real, imag} */,
  {32'hbe1749aa, 32'h3d79d960} /* (23, 30, 25) {real, imag} */,
  {32'h3d633ca5, 32'hbdd52212} /* (23, 30, 24) {real, imag} */,
  {32'h3d0738fe, 32'h3c27d9cc} /* (23, 30, 23) {real, imag} */,
  {32'hbc42185e, 32'h3d3af091} /* (23, 30, 22) {real, imag} */,
  {32'hbd8b33f3, 32'hbe05b733} /* (23, 30, 21) {real, imag} */,
  {32'hbda32415, 32'hbbdd2c70} /* (23, 30, 20) {real, imag} */,
  {32'hbcdfc1f9, 32'h3d1f08d4} /* (23, 30, 19) {real, imag} */,
  {32'h3da827fc, 32'hbd908115} /* (23, 30, 18) {real, imag} */,
  {32'hbd5f0f05, 32'h3d60ed0c} /* (23, 30, 17) {real, imag} */,
  {32'h3ce3418f, 32'h00000000} /* (23, 30, 16) {real, imag} */,
  {32'hbd5f0f05, 32'hbd60ed0c} /* (23, 30, 15) {real, imag} */,
  {32'h3da827fc, 32'h3d908115} /* (23, 30, 14) {real, imag} */,
  {32'hbcdfc1f9, 32'hbd1f08d4} /* (23, 30, 13) {real, imag} */,
  {32'hbda32415, 32'h3bdd2c70} /* (23, 30, 12) {real, imag} */,
  {32'hbd8b33f3, 32'h3e05b733} /* (23, 30, 11) {real, imag} */,
  {32'hbc42185e, 32'hbd3af091} /* (23, 30, 10) {real, imag} */,
  {32'h3d0738fe, 32'hbc27d9cc} /* (23, 30, 9) {real, imag} */,
  {32'h3d633ca5, 32'h3dd52212} /* (23, 30, 8) {real, imag} */,
  {32'hbe1749aa, 32'hbd79d960} /* (23, 30, 7) {real, imag} */,
  {32'h3e227f6b, 32'hbdb35a1e} /* (23, 30, 6) {real, imag} */,
  {32'h3e53f456, 32'h3db50f5f} /* (23, 30, 5) {real, imag} */,
  {32'hbe39d63e, 32'hbda0cae8} /* (23, 30, 4) {real, imag} */,
  {32'h3d402462, 32'h3d427d0c} /* (23, 30, 3) {real, imag} */,
  {32'h3f8ed35d, 32'h3e99c8b5} /* (23, 30, 2) {real, imag} */,
  {32'hc082658f, 32'hbfe7d93c} /* (23, 30, 1) {real, imag} */,
  {32'hc09d1de8, 32'h00000000} /* (23, 30, 0) {real, imag} */,
  {32'hc08b4758, 32'h3fc3c435} /* (23, 29, 31) {real, imag} */,
  {32'h3fae2864, 32'hbe6bcb24} /* (23, 29, 30) {real, imag} */,
  {32'hbc5ceb8c, 32'hbdc48813} /* (23, 29, 29) {real, imag} */,
  {32'hbe70269a, 32'h3e020bc6} /* (23, 29, 28) {real, imag} */,
  {32'h3d077f44, 32'hbe4601d3} /* (23, 29, 27) {real, imag} */,
  {32'h3da90076, 32'h3d3cf0d5} /* (23, 29, 26) {real, imag} */,
  {32'h3d0ed871, 32'hbc9828d0} /* (23, 29, 25) {real, imag} */,
  {32'hbd073735, 32'hbdc66296} /* (23, 29, 24) {real, imag} */,
  {32'h3ce0c00c, 32'h39d5e4c0} /* (23, 29, 23) {real, imag} */,
  {32'h3d85f6e2, 32'h3a72c780} /* (23, 29, 22) {real, imag} */,
  {32'h3d5cbec2, 32'hbb945920} /* (23, 29, 21) {real, imag} */,
  {32'h3d541214, 32'hbc5a93ed} /* (23, 29, 20) {real, imag} */,
  {32'h3cb4c05c, 32'hbc793432} /* (23, 29, 19) {real, imag} */,
  {32'hbd8d70b6, 32'h3c118948} /* (23, 29, 18) {real, imag} */,
  {32'hbcacc649, 32'h3b8e2e8c} /* (23, 29, 17) {real, imag} */,
  {32'h3ccfb844, 32'h00000000} /* (23, 29, 16) {real, imag} */,
  {32'hbcacc649, 32'hbb8e2e8c} /* (23, 29, 15) {real, imag} */,
  {32'hbd8d70b6, 32'hbc118948} /* (23, 29, 14) {real, imag} */,
  {32'h3cb4c05c, 32'h3c793432} /* (23, 29, 13) {real, imag} */,
  {32'h3d541214, 32'h3c5a93ed} /* (23, 29, 12) {real, imag} */,
  {32'h3d5cbec2, 32'h3b945920} /* (23, 29, 11) {real, imag} */,
  {32'h3d85f6e2, 32'hba72c780} /* (23, 29, 10) {real, imag} */,
  {32'h3ce0c00c, 32'hb9d5e4c0} /* (23, 29, 9) {real, imag} */,
  {32'hbd073735, 32'h3dc66296} /* (23, 29, 8) {real, imag} */,
  {32'h3d0ed871, 32'h3c9828d0} /* (23, 29, 7) {real, imag} */,
  {32'h3da90076, 32'hbd3cf0d5} /* (23, 29, 6) {real, imag} */,
  {32'h3d077f44, 32'h3e4601d3} /* (23, 29, 5) {real, imag} */,
  {32'hbe70269a, 32'hbe020bc6} /* (23, 29, 4) {real, imag} */,
  {32'hbc5ceb8c, 32'h3dc48813} /* (23, 29, 3) {real, imag} */,
  {32'h3fae2864, 32'h3e6bcb24} /* (23, 29, 2) {real, imag} */,
  {32'hc08b4758, 32'hbfc3c435} /* (23, 29, 1) {real, imag} */,
  {32'hc0a06884, 32'h00000000} /* (23, 29, 0) {real, imag} */,
  {32'hc093ead0, 32'h3f98881e} /* (23, 28, 31) {real, imag} */,
  {32'h3fc15bd9, 32'hbe9826e8} /* (23, 28, 30) {real, imag} */,
  {32'hbd44152e, 32'hbcf9c5b8} /* (23, 28, 29) {real, imag} */,
  {32'hbe79b573, 32'h3d9ac417} /* (23, 28, 28) {real, imag} */,
  {32'h3dbb3438, 32'hbddc065b} /* (23, 28, 27) {real, imag} */,
  {32'h3e0e3a69, 32'hbb906d18} /* (23, 28, 26) {real, imag} */,
  {32'h3da80e50, 32'h3dbeb484} /* (23, 28, 25) {real, imag} */,
  {32'h3d54379a, 32'hbd7a47aa} /* (23, 28, 24) {real, imag} */,
  {32'hbbb037f8, 32'h3d9ad6ee} /* (23, 28, 23) {real, imag} */,
  {32'h3d9a02c5, 32'h3d467cf0} /* (23, 28, 22) {real, imag} */,
  {32'h3db84883, 32'h3d030d86} /* (23, 28, 21) {real, imag} */,
  {32'hbccf41de, 32'h3cbf1776} /* (23, 28, 20) {real, imag} */,
  {32'h3c319dff, 32'hbd0306a8} /* (23, 28, 19) {real, imag} */,
  {32'h3d3d9de1, 32'h3cc9b820} /* (23, 28, 18) {real, imag} */,
  {32'h3d30faa5, 32'h3d361330} /* (23, 28, 17) {real, imag} */,
  {32'h3d63a37a, 32'h00000000} /* (23, 28, 16) {real, imag} */,
  {32'h3d30faa5, 32'hbd361330} /* (23, 28, 15) {real, imag} */,
  {32'h3d3d9de1, 32'hbcc9b820} /* (23, 28, 14) {real, imag} */,
  {32'h3c319dff, 32'h3d0306a8} /* (23, 28, 13) {real, imag} */,
  {32'hbccf41de, 32'hbcbf1776} /* (23, 28, 12) {real, imag} */,
  {32'h3db84883, 32'hbd030d86} /* (23, 28, 11) {real, imag} */,
  {32'h3d9a02c5, 32'hbd467cf0} /* (23, 28, 10) {real, imag} */,
  {32'hbbb037f8, 32'hbd9ad6ee} /* (23, 28, 9) {real, imag} */,
  {32'h3d54379a, 32'h3d7a47aa} /* (23, 28, 8) {real, imag} */,
  {32'h3da80e50, 32'hbdbeb484} /* (23, 28, 7) {real, imag} */,
  {32'h3e0e3a69, 32'h3b906d18} /* (23, 28, 6) {real, imag} */,
  {32'h3dbb3438, 32'h3ddc065b} /* (23, 28, 5) {real, imag} */,
  {32'hbe79b573, 32'hbd9ac417} /* (23, 28, 4) {real, imag} */,
  {32'hbd44152e, 32'h3cf9c5b8} /* (23, 28, 3) {real, imag} */,
  {32'h3fc15bd9, 32'h3e9826e8} /* (23, 28, 2) {real, imag} */,
  {32'hc093ead0, 32'hbf98881e} /* (23, 28, 1) {real, imag} */,
  {32'hc0a223d2, 32'h00000000} /* (23, 28, 0) {real, imag} */,
  {32'hc093c2ba, 32'h3f801ee0} /* (23, 27, 31) {real, imag} */,
  {32'h3fc514ae, 32'hbe7ffa10} /* (23, 27, 30) {real, imag} */,
  {32'h3de5aeb6, 32'hbd64a0ac} /* (23, 27, 29) {real, imag} */,
  {32'hbd9290e6, 32'h3cd47ace} /* (23, 27, 28) {real, imag} */,
  {32'h3e674efc, 32'hbe30a882} /* (23, 27, 27) {real, imag} */,
  {32'h3d80a7b7, 32'h3e152c42} /* (23, 27, 26) {real, imag} */,
  {32'h3d4591ec, 32'h3d851dc6} /* (23, 27, 25) {real, imag} */,
  {32'h3d8337e6, 32'h3c18944d} /* (23, 27, 24) {real, imag} */,
  {32'h3d9a67cc, 32'h3dafe520} /* (23, 27, 23) {real, imag} */,
  {32'h3c1820c4, 32'h3b761420} /* (23, 27, 22) {real, imag} */,
  {32'hbd383d02, 32'hbd8f7858} /* (23, 27, 21) {real, imag} */,
  {32'hbc241407, 32'hbd2c238b} /* (23, 27, 20) {real, imag} */,
  {32'hbdf11411, 32'h3caf8864} /* (23, 27, 19) {real, imag} */,
  {32'hbd3557c8, 32'hbd5a7a38} /* (23, 27, 18) {real, imag} */,
  {32'hbd04e68e, 32'hbb8fc420} /* (23, 27, 17) {real, imag} */,
  {32'hbc549e34, 32'h00000000} /* (23, 27, 16) {real, imag} */,
  {32'hbd04e68e, 32'h3b8fc420} /* (23, 27, 15) {real, imag} */,
  {32'hbd3557c8, 32'h3d5a7a38} /* (23, 27, 14) {real, imag} */,
  {32'hbdf11411, 32'hbcaf8864} /* (23, 27, 13) {real, imag} */,
  {32'hbc241407, 32'h3d2c238b} /* (23, 27, 12) {real, imag} */,
  {32'hbd383d02, 32'h3d8f7858} /* (23, 27, 11) {real, imag} */,
  {32'h3c1820c4, 32'hbb761420} /* (23, 27, 10) {real, imag} */,
  {32'h3d9a67cc, 32'hbdafe520} /* (23, 27, 9) {real, imag} */,
  {32'h3d8337e6, 32'hbc18944d} /* (23, 27, 8) {real, imag} */,
  {32'h3d4591ec, 32'hbd851dc6} /* (23, 27, 7) {real, imag} */,
  {32'h3d80a7b7, 32'hbe152c42} /* (23, 27, 6) {real, imag} */,
  {32'h3e674efc, 32'h3e30a882} /* (23, 27, 5) {real, imag} */,
  {32'hbd9290e6, 32'hbcd47ace} /* (23, 27, 4) {real, imag} */,
  {32'h3de5aeb6, 32'h3d64a0ac} /* (23, 27, 3) {real, imag} */,
  {32'h3fc514ae, 32'h3e7ffa10} /* (23, 27, 2) {real, imag} */,
  {32'hc093c2ba, 32'hbf801ee0} /* (23, 27, 1) {real, imag} */,
  {32'hc0a3565d, 32'h00000000} /* (23, 27, 0) {real, imag} */,
  {32'hc08d02b3, 32'h3f7407d1} /* (23, 26, 31) {real, imag} */,
  {32'h3fcaa5ec, 32'hbd99891c} /* (23, 26, 30) {real, imag} */,
  {32'h3d8f5127, 32'hbdbe0df0} /* (23, 26, 29) {real, imag} */,
  {32'hbdfbc75e, 32'hbb6a5130} /* (23, 26, 28) {real, imag} */,
  {32'h3e1a5345, 32'hbe3612aa} /* (23, 26, 27) {real, imag} */,
  {32'hbc919a36, 32'hbb2015f8} /* (23, 26, 26) {real, imag} */,
  {32'hbc147398, 32'h3d85d61f} /* (23, 26, 25) {real, imag} */,
  {32'h3cd2995a, 32'h3cd7d419} /* (23, 26, 24) {real, imag} */,
  {32'h3dba969c, 32'hbcc39fa1} /* (23, 26, 23) {real, imag} */,
  {32'hbe0a5c64, 32'hbd57c656} /* (23, 26, 22) {real, imag} */,
  {32'h3cd549ae, 32'h3c891b1e} /* (23, 26, 21) {real, imag} */,
  {32'h3c43a2cc, 32'h3c922d72} /* (23, 26, 20) {real, imag} */,
  {32'h3d40a0a0, 32'h3d09a8b0} /* (23, 26, 19) {real, imag} */,
  {32'hbd06fb68, 32'h3cd08419} /* (23, 26, 18) {real, imag} */,
  {32'h3c1f49e2, 32'hbc87b1e4} /* (23, 26, 17) {real, imag} */,
  {32'hbdb57969, 32'h00000000} /* (23, 26, 16) {real, imag} */,
  {32'h3c1f49e2, 32'h3c87b1e4} /* (23, 26, 15) {real, imag} */,
  {32'hbd06fb68, 32'hbcd08419} /* (23, 26, 14) {real, imag} */,
  {32'h3d40a0a0, 32'hbd09a8b0} /* (23, 26, 13) {real, imag} */,
  {32'h3c43a2cc, 32'hbc922d72} /* (23, 26, 12) {real, imag} */,
  {32'h3cd549ae, 32'hbc891b1e} /* (23, 26, 11) {real, imag} */,
  {32'hbe0a5c64, 32'h3d57c656} /* (23, 26, 10) {real, imag} */,
  {32'h3dba969c, 32'h3cc39fa1} /* (23, 26, 9) {real, imag} */,
  {32'h3cd2995a, 32'hbcd7d419} /* (23, 26, 8) {real, imag} */,
  {32'hbc147398, 32'hbd85d61f} /* (23, 26, 7) {real, imag} */,
  {32'hbc919a36, 32'h3b2015f8} /* (23, 26, 6) {real, imag} */,
  {32'h3e1a5345, 32'h3e3612aa} /* (23, 26, 5) {real, imag} */,
  {32'hbdfbc75e, 32'h3b6a5130} /* (23, 26, 4) {real, imag} */,
  {32'h3d8f5127, 32'h3dbe0df0} /* (23, 26, 3) {real, imag} */,
  {32'h3fcaa5ec, 32'h3d99891c} /* (23, 26, 2) {real, imag} */,
  {32'hc08d02b3, 32'hbf7407d1} /* (23, 26, 1) {real, imag} */,
  {32'hc09cf28f, 32'h00000000} /* (23, 26, 0) {real, imag} */,
  {32'hc086d72f, 32'h3f338da9} /* (23, 25, 31) {real, imag} */,
  {32'h3fcdbaf4, 32'hbe0bafb0} /* (23, 25, 30) {real, imag} */,
  {32'hbd27de3c, 32'h3b649950} /* (23, 25, 29) {real, imag} */,
  {32'hbe0fe36c, 32'hbcde198a} /* (23, 25, 28) {real, imag} */,
  {32'h3eaf554b, 32'h3b70a6c0} /* (23, 25, 27) {real, imag} */,
  {32'h3cda70c3, 32'h3d9bbeb6} /* (23, 25, 26) {real, imag} */,
  {32'h3dcd90f2, 32'hbb99606c} /* (23, 25, 25) {real, imag} */,
  {32'h3e0d2452, 32'hbcbe49e8} /* (23, 25, 24) {real, imag} */,
  {32'h3c758f0c, 32'h3d97837a} /* (23, 25, 23) {real, imag} */,
  {32'hbbf0ce6a, 32'h3d09d626} /* (23, 25, 22) {real, imag} */,
  {32'h3d1b6bdd, 32'hbd8a201f} /* (23, 25, 21) {real, imag} */,
  {32'h3d62def9, 32'h3ce98330} /* (23, 25, 20) {real, imag} */,
  {32'hbc1a8f74, 32'h3b8e0b38} /* (23, 25, 19) {real, imag} */,
  {32'hbc01fbc0, 32'hbd258fa9} /* (23, 25, 18) {real, imag} */,
  {32'hbc36457e, 32'h3d7fa26d} /* (23, 25, 17) {real, imag} */,
  {32'hbcf9214d, 32'h00000000} /* (23, 25, 16) {real, imag} */,
  {32'hbc36457e, 32'hbd7fa26d} /* (23, 25, 15) {real, imag} */,
  {32'hbc01fbc0, 32'h3d258fa9} /* (23, 25, 14) {real, imag} */,
  {32'hbc1a8f74, 32'hbb8e0b38} /* (23, 25, 13) {real, imag} */,
  {32'h3d62def9, 32'hbce98330} /* (23, 25, 12) {real, imag} */,
  {32'h3d1b6bdd, 32'h3d8a201f} /* (23, 25, 11) {real, imag} */,
  {32'hbbf0ce6a, 32'hbd09d626} /* (23, 25, 10) {real, imag} */,
  {32'h3c758f0c, 32'hbd97837a} /* (23, 25, 9) {real, imag} */,
  {32'h3e0d2452, 32'h3cbe49e8} /* (23, 25, 8) {real, imag} */,
  {32'h3dcd90f2, 32'h3b99606c} /* (23, 25, 7) {real, imag} */,
  {32'h3cda70c3, 32'hbd9bbeb6} /* (23, 25, 6) {real, imag} */,
  {32'h3eaf554b, 32'hbb70a6c0} /* (23, 25, 5) {real, imag} */,
  {32'hbe0fe36c, 32'h3cde198a} /* (23, 25, 4) {real, imag} */,
  {32'hbd27de3c, 32'hbb649950} /* (23, 25, 3) {real, imag} */,
  {32'h3fcdbaf4, 32'h3e0bafb0} /* (23, 25, 2) {real, imag} */,
  {32'hc086d72f, 32'hbf338da9} /* (23, 25, 1) {real, imag} */,
  {32'hc08faa32, 32'h00000000} /* (23, 25, 0) {real, imag} */,
  {32'hc07400dc, 32'h3f02142f} /* (23, 24, 31) {real, imag} */,
  {32'h3fc3bc78, 32'hbe55a464} /* (23, 24, 30) {real, imag} */,
  {32'hbdb62828, 32'h3dcbbfa6} /* (23, 24, 29) {real, imag} */,
  {32'hbcf6c75a, 32'h3d054718} /* (23, 24, 28) {real, imag} */,
  {32'h3e707912, 32'hbe1c2b1a} /* (23, 24, 27) {real, imag} */,
  {32'h3c041bc4, 32'hbdad373c} /* (23, 24, 26) {real, imag} */,
  {32'h3d41c535, 32'h3c709520} /* (23, 24, 25) {real, imag} */,
  {32'h3d4e1bc0, 32'h3dc99814} /* (23, 24, 24) {real, imag} */,
  {32'h3ce2445a, 32'hbc50d438} /* (23, 24, 23) {real, imag} */,
  {32'hbc8f8319, 32'h3da44ce2} /* (23, 24, 22) {real, imag} */,
  {32'h3d461941, 32'hbd9aec9b} /* (23, 24, 21) {real, imag} */,
  {32'hbc5b9a30, 32'h3cb5308c} /* (23, 24, 20) {real, imag} */,
  {32'hbd8b682c, 32'hbd25e327} /* (23, 24, 19) {real, imag} */,
  {32'h3c234bd4, 32'h3d2f62fb} /* (23, 24, 18) {real, imag} */,
  {32'hbca3322a, 32'hbcb8abe4} /* (23, 24, 17) {real, imag} */,
  {32'h3e037f4d, 32'h00000000} /* (23, 24, 16) {real, imag} */,
  {32'hbca3322a, 32'h3cb8abe4} /* (23, 24, 15) {real, imag} */,
  {32'h3c234bd4, 32'hbd2f62fb} /* (23, 24, 14) {real, imag} */,
  {32'hbd8b682c, 32'h3d25e327} /* (23, 24, 13) {real, imag} */,
  {32'hbc5b9a30, 32'hbcb5308c} /* (23, 24, 12) {real, imag} */,
  {32'h3d461941, 32'h3d9aec9b} /* (23, 24, 11) {real, imag} */,
  {32'hbc8f8319, 32'hbda44ce2} /* (23, 24, 10) {real, imag} */,
  {32'h3ce2445a, 32'h3c50d438} /* (23, 24, 9) {real, imag} */,
  {32'h3d4e1bc0, 32'hbdc99814} /* (23, 24, 8) {real, imag} */,
  {32'h3d41c535, 32'hbc709520} /* (23, 24, 7) {real, imag} */,
  {32'h3c041bc4, 32'h3dad373c} /* (23, 24, 6) {real, imag} */,
  {32'h3e707912, 32'h3e1c2b1a} /* (23, 24, 5) {real, imag} */,
  {32'hbcf6c75a, 32'hbd054718} /* (23, 24, 4) {real, imag} */,
  {32'hbdb62828, 32'hbdcbbfa6} /* (23, 24, 3) {real, imag} */,
  {32'h3fc3bc78, 32'h3e55a464} /* (23, 24, 2) {real, imag} */,
  {32'hc07400dc, 32'hbf02142f} /* (23, 24, 1) {real, imag} */,
  {32'hc079586c, 32'h00000000} /* (23, 24, 0) {real, imag} */,
  {32'hc04f85b2, 32'h3edbfe52} /* (23, 23, 31) {real, imag} */,
  {32'h3fab9ad8, 32'hbe079ce8} /* (23, 23, 30) {real, imag} */,
  {32'hbd3dbe1c, 32'h3d2801c5} /* (23, 23, 29) {real, imag} */,
  {32'hbdaf5581, 32'h3df89864} /* (23, 23, 28) {real, imag} */,
  {32'h3e126ac2, 32'hbda159ea} /* (23, 23, 27) {real, imag} */,
  {32'hbd84dd79, 32'h3ca259ae} /* (23, 23, 26) {real, imag} */,
  {32'hbce19eb5, 32'h3d5c061a} /* (23, 23, 25) {real, imag} */,
  {32'hbd35c3f2, 32'h3d928923} /* (23, 23, 24) {real, imag} */,
  {32'hbd31b02e, 32'h3c891381} /* (23, 23, 23) {real, imag} */,
  {32'hbd280bc6, 32'h3c7ade8e} /* (23, 23, 22) {real, imag} */,
  {32'h3dd07cc9, 32'hbd55a092} /* (23, 23, 21) {real, imag} */,
  {32'hbb6325b0, 32'h3d3bc5ef} /* (23, 23, 20) {real, imag} */,
  {32'h3c997aec, 32'hbdd19f24} /* (23, 23, 19) {real, imag} */,
  {32'hbd6b033e, 32'h3d0252c9} /* (23, 23, 18) {real, imag} */,
  {32'hbb705148, 32'h3cc58f46} /* (23, 23, 17) {real, imag} */,
  {32'hbc63c82a, 32'h00000000} /* (23, 23, 16) {real, imag} */,
  {32'hbb705148, 32'hbcc58f46} /* (23, 23, 15) {real, imag} */,
  {32'hbd6b033e, 32'hbd0252c9} /* (23, 23, 14) {real, imag} */,
  {32'h3c997aec, 32'h3dd19f24} /* (23, 23, 13) {real, imag} */,
  {32'hbb6325b0, 32'hbd3bc5ef} /* (23, 23, 12) {real, imag} */,
  {32'h3dd07cc9, 32'h3d55a092} /* (23, 23, 11) {real, imag} */,
  {32'hbd280bc6, 32'hbc7ade8e} /* (23, 23, 10) {real, imag} */,
  {32'hbd31b02e, 32'hbc891381} /* (23, 23, 9) {real, imag} */,
  {32'hbd35c3f2, 32'hbd928923} /* (23, 23, 8) {real, imag} */,
  {32'hbce19eb5, 32'hbd5c061a} /* (23, 23, 7) {real, imag} */,
  {32'hbd84dd79, 32'hbca259ae} /* (23, 23, 6) {real, imag} */,
  {32'h3e126ac2, 32'h3da159ea} /* (23, 23, 5) {real, imag} */,
  {32'hbdaf5581, 32'hbdf89864} /* (23, 23, 4) {real, imag} */,
  {32'hbd3dbe1c, 32'hbd2801c5} /* (23, 23, 3) {real, imag} */,
  {32'h3fab9ad8, 32'h3e079ce8} /* (23, 23, 2) {real, imag} */,
  {32'hc04f85b2, 32'hbedbfe52} /* (23, 23, 1) {real, imag} */,
  {32'hc04422d6, 32'h00000000} /* (23, 23, 0) {real, imag} */,
  {32'hc012b5c2, 32'h3e6a84a1} /* (23, 22, 31) {real, imag} */,
  {32'h3f6c861f, 32'hbe04baee} /* (23, 22, 30) {real, imag} */,
  {32'hbd4f8e1a, 32'hbcbf0d6e} /* (23, 22, 29) {real, imag} */,
  {32'hbe0c8ff3, 32'h3e221bb6} /* (23, 22, 28) {real, imag} */,
  {32'h3e54b0c5, 32'hbd8feea9} /* (23, 22, 27) {real, imag} */,
  {32'hbd131dab, 32'h3cdd3fc9} /* (23, 22, 26) {real, imag} */,
  {32'hbd3cf9bc, 32'h3d54d25c} /* (23, 22, 25) {real, imag} */,
  {32'h3ad39be0, 32'hbda2cbca} /* (23, 22, 24) {real, imag} */,
  {32'hbd9e025a, 32'h3cc89ea5} /* (23, 22, 23) {real, imag} */,
  {32'h3c2c35dc, 32'hbc985c66} /* (23, 22, 22) {real, imag} */,
  {32'hbd0914c4, 32'hbb7eb3bc} /* (23, 22, 21) {real, imag} */,
  {32'h3be8f9f8, 32'hbc3c0b60} /* (23, 22, 20) {real, imag} */,
  {32'hbd0de986, 32'h3ad10fd0} /* (23, 22, 19) {real, imag} */,
  {32'h3d83005e, 32'hbccd53e2} /* (23, 22, 18) {real, imag} */,
  {32'hbcc7f47e, 32'hbc8c0710} /* (23, 22, 17) {real, imag} */,
  {32'h3cf23895, 32'h00000000} /* (23, 22, 16) {real, imag} */,
  {32'hbcc7f47e, 32'h3c8c0710} /* (23, 22, 15) {real, imag} */,
  {32'h3d83005e, 32'h3ccd53e2} /* (23, 22, 14) {real, imag} */,
  {32'hbd0de986, 32'hbad10fd0} /* (23, 22, 13) {real, imag} */,
  {32'h3be8f9f8, 32'h3c3c0b60} /* (23, 22, 12) {real, imag} */,
  {32'hbd0914c4, 32'h3b7eb3bc} /* (23, 22, 11) {real, imag} */,
  {32'h3c2c35dc, 32'h3c985c66} /* (23, 22, 10) {real, imag} */,
  {32'hbd9e025a, 32'hbcc89ea5} /* (23, 22, 9) {real, imag} */,
  {32'h3ad39be0, 32'h3da2cbca} /* (23, 22, 8) {real, imag} */,
  {32'hbd3cf9bc, 32'hbd54d25c} /* (23, 22, 7) {real, imag} */,
  {32'hbd131dab, 32'hbcdd3fc9} /* (23, 22, 6) {real, imag} */,
  {32'h3e54b0c5, 32'h3d8feea9} /* (23, 22, 5) {real, imag} */,
  {32'hbe0c8ff3, 32'hbe221bb6} /* (23, 22, 4) {real, imag} */,
  {32'hbd4f8e1a, 32'h3cbf0d6e} /* (23, 22, 3) {real, imag} */,
  {32'h3f6c861f, 32'h3e04baee} /* (23, 22, 2) {real, imag} */,
  {32'hc012b5c2, 32'hbe6a84a1} /* (23, 22, 1) {real, imag} */,
  {32'hc0018be3, 32'h00000000} /* (23, 22, 0) {real, imag} */,
  {32'hbf7c84a0, 32'h3d5e8188} /* (23, 21, 31) {real, imag} */,
  {32'h3eacbe70, 32'hbe114a48} /* (23, 21, 30) {real, imag} */,
  {32'hbd8c9901, 32'h3de97b94} /* (23, 21, 29) {real, imag} */,
  {32'h3d388cff, 32'h3df373b8} /* (23, 21, 28) {real, imag} */,
  {32'h3e28f298, 32'hbda13113} /* (23, 21, 27) {real, imag} */,
  {32'hbd95fc8f, 32'hbce93855} /* (23, 21, 26) {real, imag} */,
  {32'h3de0c03a, 32'hbdd38f5c} /* (23, 21, 25) {real, imag} */,
  {32'hbe16279e, 32'hbb6f357c} /* (23, 21, 24) {real, imag} */,
  {32'hbd8781e5, 32'hbd46932e} /* (23, 21, 23) {real, imag} */,
  {32'hbd09b5b6, 32'h3d544839} /* (23, 21, 22) {real, imag} */,
  {32'h3dc29761, 32'hbd0425e6} /* (23, 21, 21) {real, imag} */,
  {32'hbd3d7327, 32'hbc9ee67b} /* (23, 21, 20) {real, imag} */,
  {32'hbdc731a1, 32'hbcaaf31c} /* (23, 21, 19) {real, imag} */,
  {32'h3d9d52ca, 32'hbbf43488} /* (23, 21, 18) {real, imag} */,
  {32'hbd557074, 32'h3d272a58} /* (23, 21, 17) {real, imag} */,
  {32'hbb3a8d00, 32'h00000000} /* (23, 21, 16) {real, imag} */,
  {32'hbd557074, 32'hbd272a58} /* (23, 21, 15) {real, imag} */,
  {32'h3d9d52ca, 32'h3bf43488} /* (23, 21, 14) {real, imag} */,
  {32'hbdc731a1, 32'h3caaf31c} /* (23, 21, 13) {real, imag} */,
  {32'hbd3d7327, 32'h3c9ee67b} /* (23, 21, 12) {real, imag} */,
  {32'h3dc29761, 32'h3d0425e6} /* (23, 21, 11) {real, imag} */,
  {32'hbd09b5b6, 32'hbd544839} /* (23, 21, 10) {real, imag} */,
  {32'hbd8781e5, 32'h3d46932e} /* (23, 21, 9) {real, imag} */,
  {32'hbe16279e, 32'h3b6f357c} /* (23, 21, 8) {real, imag} */,
  {32'h3de0c03a, 32'h3dd38f5c} /* (23, 21, 7) {real, imag} */,
  {32'hbd95fc8f, 32'h3ce93855} /* (23, 21, 6) {real, imag} */,
  {32'h3e28f298, 32'h3da13113} /* (23, 21, 5) {real, imag} */,
  {32'h3d388cff, 32'hbdf373b8} /* (23, 21, 4) {real, imag} */,
  {32'hbd8c9901, 32'hbde97b94} /* (23, 21, 3) {real, imag} */,
  {32'h3eacbe70, 32'h3e114a48} /* (23, 21, 2) {real, imag} */,
  {32'hbf7c84a0, 32'hbd5e8188} /* (23, 21, 1) {real, imag} */,
  {32'hbf876531, 32'h00000000} /* (23, 21, 0) {real, imag} */,
  {32'h3f651645, 32'hbe204fa8} /* (23, 20, 31) {real, imag} */,
  {32'hbf0a611c, 32'hbe05eeff} /* (23, 20, 30) {real, imag} */,
  {32'hbc3c41a0, 32'h3e2b06ee} /* (23, 20, 29) {real, imag} */,
  {32'h3e1d06e9, 32'hbe125ad9} /* (23, 20, 28) {real, imag} */,
  {32'hbcb12e40, 32'h3d01dc90} /* (23, 20, 27) {real, imag} */,
  {32'hbe054b88, 32'hbdc0fc80} /* (23, 20, 26) {real, imag} */,
  {32'h3d5856a4, 32'hbdadb74a} /* (23, 20, 25) {real, imag} */,
  {32'hbe2b4174, 32'h3d391b56} /* (23, 20, 24) {real, imag} */,
  {32'h3d4e3659, 32'h3c43497c} /* (23, 20, 23) {real, imag} */,
  {32'hbd721796, 32'hbc8c020c} /* (23, 20, 22) {real, imag} */,
  {32'h3e0fa820, 32'h3dce54a7} /* (23, 20, 21) {real, imag} */,
  {32'hbd6ebb44, 32'h3bca4a7c} /* (23, 20, 20) {real, imag} */,
  {32'hbd6a2854, 32'h3e029f96} /* (23, 20, 19) {real, imag} */,
  {32'h3945fa00, 32'h3d6f83aa} /* (23, 20, 18) {real, imag} */,
  {32'hbcdcc77b, 32'hbbb3cd6c} /* (23, 20, 17) {real, imag} */,
  {32'hbccc0d3c, 32'h00000000} /* (23, 20, 16) {real, imag} */,
  {32'hbcdcc77b, 32'h3bb3cd6c} /* (23, 20, 15) {real, imag} */,
  {32'h3945fa00, 32'hbd6f83aa} /* (23, 20, 14) {real, imag} */,
  {32'hbd6a2854, 32'hbe029f96} /* (23, 20, 13) {real, imag} */,
  {32'hbd6ebb44, 32'hbbca4a7c} /* (23, 20, 12) {real, imag} */,
  {32'h3e0fa820, 32'hbdce54a7} /* (23, 20, 11) {real, imag} */,
  {32'hbd721796, 32'h3c8c020c} /* (23, 20, 10) {real, imag} */,
  {32'h3d4e3659, 32'hbc43497c} /* (23, 20, 9) {real, imag} */,
  {32'hbe2b4174, 32'hbd391b56} /* (23, 20, 8) {real, imag} */,
  {32'h3d5856a4, 32'h3dadb74a} /* (23, 20, 7) {real, imag} */,
  {32'hbe054b88, 32'h3dc0fc80} /* (23, 20, 6) {real, imag} */,
  {32'hbcb12e40, 32'hbd01dc90} /* (23, 20, 5) {real, imag} */,
  {32'h3e1d06e9, 32'h3e125ad9} /* (23, 20, 4) {real, imag} */,
  {32'hbc3c41a0, 32'hbe2b06ee} /* (23, 20, 3) {real, imag} */,
  {32'hbf0a611c, 32'h3e05eeff} /* (23, 20, 2) {real, imag} */,
  {32'h3f651645, 32'h3e204fa8} /* (23, 20, 1) {real, imag} */,
  {32'h3eef80ce, 32'h00000000} /* (23, 20, 0) {real, imag} */,
  {32'h4004e26f, 32'hbea85f2d} /* (23, 19, 31) {real, imag} */,
  {32'hbf46084e, 32'h3e636225} /* (23, 19, 30) {real, imag} */,
  {32'hbca62422, 32'h3dd118ac} /* (23, 19, 29) {real, imag} */,
  {32'h3e34c0a7, 32'hbe93ab46} /* (23, 19, 28) {real, imag} */,
  {32'hbde91676, 32'h3cc68324} /* (23, 19, 27) {real, imag} */,
  {32'h3c3e65b8, 32'hbc9cf768} /* (23, 19, 26) {real, imag} */,
  {32'h3d62307f, 32'hbd1b97dc} /* (23, 19, 25) {real, imag} */,
  {32'hbd0c2a7a, 32'h3c88fe91} /* (23, 19, 24) {real, imag} */,
  {32'hbdab8f30, 32'h3db2c6aa} /* (23, 19, 23) {real, imag} */,
  {32'hbd81fadd, 32'hbd017ac7} /* (23, 19, 22) {real, imag} */,
  {32'hbcbf95c0, 32'h3ce391b2} /* (23, 19, 21) {real, imag} */,
  {32'hbdef4c8b, 32'h3d79a28e} /* (23, 19, 20) {real, imag} */,
  {32'h3ca6d912, 32'hbcca9216} /* (23, 19, 19) {real, imag} */,
  {32'h3b81b1e8, 32'hbbbdaf78} /* (23, 19, 18) {real, imag} */,
  {32'h3cd417bd, 32'h3ca87aa1} /* (23, 19, 17) {real, imag} */,
  {32'hbc0b3b36, 32'h00000000} /* (23, 19, 16) {real, imag} */,
  {32'h3cd417bd, 32'hbca87aa1} /* (23, 19, 15) {real, imag} */,
  {32'h3b81b1e8, 32'h3bbdaf78} /* (23, 19, 14) {real, imag} */,
  {32'h3ca6d912, 32'h3cca9216} /* (23, 19, 13) {real, imag} */,
  {32'hbdef4c8b, 32'hbd79a28e} /* (23, 19, 12) {real, imag} */,
  {32'hbcbf95c0, 32'hbce391b2} /* (23, 19, 11) {real, imag} */,
  {32'hbd81fadd, 32'h3d017ac7} /* (23, 19, 10) {real, imag} */,
  {32'hbdab8f30, 32'hbdb2c6aa} /* (23, 19, 9) {real, imag} */,
  {32'hbd0c2a7a, 32'hbc88fe91} /* (23, 19, 8) {real, imag} */,
  {32'h3d62307f, 32'h3d1b97dc} /* (23, 19, 7) {real, imag} */,
  {32'h3c3e65b8, 32'h3c9cf768} /* (23, 19, 6) {real, imag} */,
  {32'hbde91676, 32'hbcc68324} /* (23, 19, 5) {real, imag} */,
  {32'h3e34c0a7, 32'h3e93ab46} /* (23, 19, 4) {real, imag} */,
  {32'hbca62422, 32'hbdd118ac} /* (23, 19, 3) {real, imag} */,
  {32'hbf46084e, 32'hbe636225} /* (23, 19, 2) {real, imag} */,
  {32'h4004e26f, 32'h3ea85f2d} /* (23, 19, 1) {real, imag} */,
  {32'h3faf93c8, 32'h00000000} /* (23, 19, 0) {real, imag} */,
  {32'h403a755a, 32'hbe8aeb90} /* (23, 18, 31) {real, imag} */,
  {32'hbf85029c, 32'h3e83646e} /* (23, 18, 30) {real, imag} */,
  {32'h3bdebb10, 32'h3cb1a6f9} /* (23, 18, 29) {real, imag} */,
  {32'h3e9fca81, 32'hbe772bf6} /* (23, 18, 28) {real, imag} */,
  {32'hbe9e73d8, 32'h3d86bbb2} /* (23, 18, 27) {real, imag} */,
  {32'h3d956017, 32'h3d8ae5a3} /* (23, 18, 26) {real, imag} */,
  {32'hbd3cba30, 32'h3cdef434} /* (23, 18, 25) {real, imag} */,
  {32'h3be91978, 32'h3e19c1db} /* (23, 18, 24) {real, imag} */,
  {32'hbbf12f1f, 32'h3c9dd4fb} /* (23, 18, 23) {real, imag} */,
  {32'hbd0db31c, 32'h3dd25e9e} /* (23, 18, 22) {real, imag} */,
  {32'h3b745818, 32'h3dc4e476} /* (23, 18, 21) {real, imag} */,
  {32'hbc65d736, 32'hbce0aa8a} /* (23, 18, 20) {real, imag} */,
  {32'h3d687e9c, 32'h3c515586} /* (23, 18, 19) {real, imag} */,
  {32'hbcaa285d, 32'h3cdfcd9b} /* (23, 18, 18) {real, imag} */,
  {32'hbced5694, 32'hbd51e129} /* (23, 18, 17) {real, imag} */,
  {32'hbcdc6df0, 32'h00000000} /* (23, 18, 16) {real, imag} */,
  {32'hbced5694, 32'h3d51e129} /* (23, 18, 15) {real, imag} */,
  {32'hbcaa285d, 32'hbcdfcd9b} /* (23, 18, 14) {real, imag} */,
  {32'h3d687e9c, 32'hbc515586} /* (23, 18, 13) {real, imag} */,
  {32'hbc65d736, 32'h3ce0aa8a} /* (23, 18, 12) {real, imag} */,
  {32'h3b745818, 32'hbdc4e476} /* (23, 18, 11) {real, imag} */,
  {32'hbd0db31c, 32'hbdd25e9e} /* (23, 18, 10) {real, imag} */,
  {32'hbbf12f1f, 32'hbc9dd4fb} /* (23, 18, 9) {real, imag} */,
  {32'h3be91978, 32'hbe19c1db} /* (23, 18, 8) {real, imag} */,
  {32'hbd3cba30, 32'hbcdef434} /* (23, 18, 7) {real, imag} */,
  {32'h3d956017, 32'hbd8ae5a3} /* (23, 18, 6) {real, imag} */,
  {32'hbe9e73d8, 32'hbd86bbb2} /* (23, 18, 5) {real, imag} */,
  {32'h3e9fca81, 32'h3e772bf6} /* (23, 18, 4) {real, imag} */,
  {32'h3bdebb10, 32'hbcb1a6f9} /* (23, 18, 3) {real, imag} */,
  {32'hbf85029c, 32'hbe83646e} /* (23, 18, 2) {real, imag} */,
  {32'h403a755a, 32'h3e8aeb90} /* (23, 18, 1) {real, imag} */,
  {32'h3ff075c4, 32'h00000000} /* (23, 18, 0) {real, imag} */,
  {32'h405eef41, 32'hbeb4a511} /* (23, 17, 31) {real, imag} */,
  {32'hbf9534c8, 32'h3e9be5d7} /* (23, 17, 30) {real, imag} */,
  {32'h3d16ce4e, 32'hbc2499c8} /* (23, 17, 29) {real, imag} */,
  {32'h3ebf64e7, 32'hbe83b61b} /* (23, 17, 28) {real, imag} */,
  {32'hbe3b185a, 32'h3db8cb2f} /* (23, 17, 27) {real, imag} */,
  {32'hbd89bcd7, 32'h3d254944} /* (23, 17, 26) {real, imag} */,
  {32'h3d22e8d4, 32'hbcff5356} /* (23, 17, 25) {real, imag} */,
  {32'h3d38b8a7, 32'h3dd2e44c} /* (23, 17, 24) {real, imag} */,
  {32'hbcdf9222, 32'hbd1999f0} /* (23, 17, 23) {real, imag} */,
  {32'h3ccdcefe, 32'hbe09e442} /* (23, 17, 22) {real, imag} */,
  {32'hbd979034, 32'h3c387891} /* (23, 17, 21) {real, imag} */,
  {32'h3a2a52c0, 32'h3c91f8bb} /* (23, 17, 20) {real, imag} */,
  {32'hbdc0142a, 32'h3d2694ae} /* (23, 17, 19) {real, imag} */,
  {32'hbc94509b, 32'h3da1e943} /* (23, 17, 18) {real, imag} */,
  {32'h3ca48631, 32'hbbc23ab4} /* (23, 17, 17) {real, imag} */,
  {32'hbc6607fa, 32'h00000000} /* (23, 17, 16) {real, imag} */,
  {32'h3ca48631, 32'h3bc23ab4} /* (23, 17, 15) {real, imag} */,
  {32'hbc94509b, 32'hbda1e943} /* (23, 17, 14) {real, imag} */,
  {32'hbdc0142a, 32'hbd2694ae} /* (23, 17, 13) {real, imag} */,
  {32'h3a2a52c0, 32'hbc91f8bb} /* (23, 17, 12) {real, imag} */,
  {32'hbd979034, 32'hbc387891} /* (23, 17, 11) {real, imag} */,
  {32'h3ccdcefe, 32'h3e09e442} /* (23, 17, 10) {real, imag} */,
  {32'hbcdf9222, 32'h3d1999f0} /* (23, 17, 9) {real, imag} */,
  {32'h3d38b8a7, 32'hbdd2e44c} /* (23, 17, 8) {real, imag} */,
  {32'h3d22e8d4, 32'h3cff5356} /* (23, 17, 7) {real, imag} */,
  {32'hbd89bcd7, 32'hbd254944} /* (23, 17, 6) {real, imag} */,
  {32'hbe3b185a, 32'hbdb8cb2f} /* (23, 17, 5) {real, imag} */,
  {32'h3ebf64e7, 32'h3e83b61b} /* (23, 17, 4) {real, imag} */,
  {32'h3d16ce4e, 32'h3c2499c8} /* (23, 17, 3) {real, imag} */,
  {32'hbf9534c8, 32'hbe9be5d7} /* (23, 17, 2) {real, imag} */,
  {32'h405eef41, 32'h3eb4a511} /* (23, 17, 1) {real, imag} */,
  {32'h4005a853, 32'h00000000} /* (23, 17, 0) {real, imag} */,
  {32'h4068c5ee, 32'hbecbf708} /* (23, 16, 31) {real, imag} */,
  {32'hbfa0c1dd, 32'h3ea30785} /* (23, 16, 30) {real, imag} */,
  {32'h3ccc402a, 32'h3dd67ffc} /* (23, 16, 29) {real, imag} */,
  {32'h3ea548a6, 32'hbe0d8802} /* (23, 16, 28) {real, imag} */,
  {32'hbe8288d2, 32'h3da30f6d} /* (23, 16, 27) {real, imag} */,
  {32'hbe0a9bd1, 32'hbb834470} /* (23, 16, 26) {real, imag} */,
  {32'h3dd1c41a, 32'hbb894d78} /* (23, 16, 25) {real, imag} */,
  {32'hbd9b74a6, 32'h3dc32716} /* (23, 16, 24) {real, imag} */,
  {32'hbd85db8c, 32'h3dc31e25} /* (23, 16, 23) {real, imag} */,
  {32'hbbc31545, 32'hbc92d176} /* (23, 16, 22) {real, imag} */,
  {32'hbd5e0010, 32'h3c577865} /* (23, 16, 21) {real, imag} */,
  {32'hbd12de2b, 32'h3c835090} /* (23, 16, 20) {real, imag} */,
  {32'h3c856ba4, 32'hbd861b2e} /* (23, 16, 19) {real, imag} */,
  {32'h3d516b20, 32'hbda38b0c} /* (23, 16, 18) {real, imag} */,
  {32'h3c71304a, 32'hbc202802} /* (23, 16, 17) {real, imag} */,
  {32'hbdc573be, 32'h00000000} /* (23, 16, 16) {real, imag} */,
  {32'h3c71304a, 32'h3c202802} /* (23, 16, 15) {real, imag} */,
  {32'h3d516b20, 32'h3da38b0c} /* (23, 16, 14) {real, imag} */,
  {32'h3c856ba4, 32'h3d861b2e} /* (23, 16, 13) {real, imag} */,
  {32'hbd12de2b, 32'hbc835090} /* (23, 16, 12) {real, imag} */,
  {32'hbd5e0010, 32'hbc577865} /* (23, 16, 11) {real, imag} */,
  {32'hbbc31545, 32'h3c92d176} /* (23, 16, 10) {real, imag} */,
  {32'hbd85db8c, 32'hbdc31e25} /* (23, 16, 9) {real, imag} */,
  {32'hbd9b74a6, 32'hbdc32716} /* (23, 16, 8) {real, imag} */,
  {32'h3dd1c41a, 32'h3b894d78} /* (23, 16, 7) {real, imag} */,
  {32'hbe0a9bd1, 32'h3b834470} /* (23, 16, 6) {real, imag} */,
  {32'hbe8288d2, 32'hbda30f6d} /* (23, 16, 5) {real, imag} */,
  {32'h3ea548a6, 32'h3e0d8802} /* (23, 16, 4) {real, imag} */,
  {32'h3ccc402a, 32'hbdd67ffc} /* (23, 16, 3) {real, imag} */,
  {32'hbfa0c1dd, 32'hbea30785} /* (23, 16, 2) {real, imag} */,
  {32'h4068c5ee, 32'h3ecbf708} /* (23, 16, 1) {real, imag} */,
  {32'h401d55d4, 32'h00000000} /* (23, 16, 0) {real, imag} */,
  {32'h406cff65, 32'hbe977057} /* (23, 15, 31) {real, imag} */,
  {32'hbfa2f2c0, 32'h3e5407aa} /* (23, 15, 30) {real, imag} */,
  {32'hbe2d85fe, 32'h3de1fa41} /* (23, 15, 29) {real, imag} */,
  {32'h3e8c12b1, 32'hbdc3f174} /* (23, 15, 28) {real, imag} */,
  {32'hbe72dc1a, 32'h3de1f2f5} /* (23, 15, 27) {real, imag} */,
  {32'hbc137ca8, 32'hbd1a7ba8} /* (23, 15, 26) {real, imag} */,
  {32'h3daab047, 32'hbc770f9c} /* (23, 15, 25) {real, imag} */,
  {32'hbe1a1afa, 32'hbdb76228} /* (23, 15, 24) {real, imag} */,
  {32'h3c2155f4, 32'h3dbc7f02} /* (23, 15, 23) {real, imag} */,
  {32'h3b887aa2, 32'h3d782916} /* (23, 15, 22) {real, imag} */,
  {32'h3d3dbf5c, 32'hbcb5e8ee} /* (23, 15, 21) {real, imag} */,
  {32'h3dd59b6c, 32'h3d2de9a4} /* (23, 15, 20) {real, imag} */,
  {32'hbcfe3850, 32'hbdea3941} /* (23, 15, 19) {real, imag} */,
  {32'h388e0100, 32'h3cdc77c0} /* (23, 15, 18) {real, imag} */,
  {32'h3cc6bea9, 32'hbd448a00} /* (23, 15, 17) {real, imag} */,
  {32'hbd8929a9, 32'h00000000} /* (23, 15, 16) {real, imag} */,
  {32'h3cc6bea9, 32'h3d448a00} /* (23, 15, 15) {real, imag} */,
  {32'h388e0100, 32'hbcdc77c0} /* (23, 15, 14) {real, imag} */,
  {32'hbcfe3850, 32'h3dea3941} /* (23, 15, 13) {real, imag} */,
  {32'h3dd59b6c, 32'hbd2de9a4} /* (23, 15, 12) {real, imag} */,
  {32'h3d3dbf5c, 32'h3cb5e8ee} /* (23, 15, 11) {real, imag} */,
  {32'h3b887aa2, 32'hbd782916} /* (23, 15, 10) {real, imag} */,
  {32'h3c2155f4, 32'hbdbc7f02} /* (23, 15, 9) {real, imag} */,
  {32'hbe1a1afa, 32'h3db76228} /* (23, 15, 8) {real, imag} */,
  {32'h3daab047, 32'h3c770f9c} /* (23, 15, 7) {real, imag} */,
  {32'hbc137ca8, 32'h3d1a7ba8} /* (23, 15, 6) {real, imag} */,
  {32'hbe72dc1a, 32'hbde1f2f5} /* (23, 15, 5) {real, imag} */,
  {32'h3e8c12b1, 32'h3dc3f174} /* (23, 15, 4) {real, imag} */,
  {32'hbe2d85fe, 32'hbde1fa41} /* (23, 15, 3) {real, imag} */,
  {32'hbfa2f2c0, 32'hbe5407aa} /* (23, 15, 2) {real, imag} */,
  {32'h406cff65, 32'h3e977057} /* (23, 15, 1) {real, imag} */,
  {32'h40205b67, 32'h00000000} /* (23, 15, 0) {real, imag} */,
  {32'h4055db62, 32'hbddb9320} /* (23, 14, 31) {real, imag} */,
  {32'hbfab1dd8, 32'h3e629c5f} /* (23, 14, 30) {real, imag} */,
  {32'hbdafe72d, 32'h3d37febc} /* (23, 14, 29) {real, imag} */,
  {32'h3eb2d9d7, 32'hbe5834be} /* (23, 14, 28) {real, imag} */,
  {32'hbe756034, 32'h3d7dd9d3} /* (23, 14, 27) {real, imag} */,
  {32'hbdd2bfed, 32'h3b1ed460} /* (23, 14, 26) {real, imag} */,
  {32'h3df1d47e, 32'hbd3114da} /* (23, 14, 25) {real, imag} */,
  {32'h3dc390a8, 32'hbd2825c5} /* (23, 14, 24) {real, imag} */,
  {32'h3c457e68, 32'hbc314e62} /* (23, 14, 23) {real, imag} */,
  {32'h3b67b1f8, 32'h3d210ef7} /* (23, 14, 22) {real, imag} */,
  {32'hbc895fdd, 32'h3da2021e} /* (23, 14, 21) {real, imag} */,
  {32'h3d0e2170, 32'hbd64afc7} /* (23, 14, 20) {real, imag} */,
  {32'h3d09c000, 32'h3d3c0f12} /* (23, 14, 19) {real, imag} */,
  {32'hbcff85ff, 32'h3d2e5ca2} /* (23, 14, 18) {real, imag} */,
  {32'h3c278d9b, 32'h3cddb7d2} /* (23, 14, 17) {real, imag} */,
  {32'h3d082dcb, 32'h00000000} /* (23, 14, 16) {real, imag} */,
  {32'h3c278d9b, 32'hbcddb7d2} /* (23, 14, 15) {real, imag} */,
  {32'hbcff85ff, 32'hbd2e5ca2} /* (23, 14, 14) {real, imag} */,
  {32'h3d09c000, 32'hbd3c0f12} /* (23, 14, 13) {real, imag} */,
  {32'h3d0e2170, 32'h3d64afc7} /* (23, 14, 12) {real, imag} */,
  {32'hbc895fdd, 32'hbda2021e} /* (23, 14, 11) {real, imag} */,
  {32'h3b67b1f8, 32'hbd210ef7} /* (23, 14, 10) {real, imag} */,
  {32'h3c457e68, 32'h3c314e62} /* (23, 14, 9) {real, imag} */,
  {32'h3dc390a8, 32'h3d2825c5} /* (23, 14, 8) {real, imag} */,
  {32'h3df1d47e, 32'h3d3114da} /* (23, 14, 7) {real, imag} */,
  {32'hbdd2bfed, 32'hbb1ed460} /* (23, 14, 6) {real, imag} */,
  {32'hbe756034, 32'hbd7dd9d3} /* (23, 14, 5) {real, imag} */,
  {32'h3eb2d9d7, 32'h3e5834be} /* (23, 14, 4) {real, imag} */,
  {32'hbdafe72d, 32'hbd37febc} /* (23, 14, 3) {real, imag} */,
  {32'hbfab1dd8, 32'hbe629c5f} /* (23, 14, 2) {real, imag} */,
  {32'h4055db62, 32'h3ddb9320} /* (23, 14, 1) {real, imag} */,
  {32'h4022e7e0, 32'h00000000} /* (23, 14, 0) {real, imag} */,
  {32'h40351305, 32'hbd58ea98} /* (23, 13, 31) {real, imag} */,
  {32'hbfad1131, 32'h3e231c1f} /* (23, 13, 30) {real, imag} */,
  {32'hbdae87e8, 32'hbc1f4f90} /* (23, 13, 29) {real, imag} */,
  {32'h3ea13e0c, 32'hbe98083c} /* (23, 13, 28) {real, imag} */,
  {32'hbe91c26a, 32'h3e02a688} /* (23, 13, 27) {real, imag} */,
  {32'h3da787e3, 32'h3ca2a9a4} /* (23, 13, 26) {real, imag} */,
  {32'h3e3569e3, 32'h3d50d1d2} /* (23, 13, 25) {real, imag} */,
  {32'hbb05e9a0, 32'hbc536cf2} /* (23, 13, 24) {real, imag} */,
  {32'h3da7fdac, 32'h3c0a7d60} /* (23, 13, 23) {real, imag} */,
  {32'h3bc835bc, 32'h3bb486f8} /* (23, 13, 22) {real, imag} */,
  {32'h3d882d14, 32'h3db50654} /* (23, 13, 21) {real, imag} */,
  {32'h3bbb4c50, 32'h3c87b8f4} /* (23, 13, 20) {real, imag} */,
  {32'hbd93d4cc, 32'hbce11a60} /* (23, 13, 19) {real, imag} */,
  {32'h3d19298d, 32'hbd22c123} /* (23, 13, 18) {real, imag} */,
  {32'hbd895245, 32'h3c7e8f42} /* (23, 13, 17) {real, imag} */,
  {32'hbd434c56, 32'h00000000} /* (23, 13, 16) {real, imag} */,
  {32'hbd895245, 32'hbc7e8f42} /* (23, 13, 15) {real, imag} */,
  {32'h3d19298d, 32'h3d22c123} /* (23, 13, 14) {real, imag} */,
  {32'hbd93d4cc, 32'h3ce11a60} /* (23, 13, 13) {real, imag} */,
  {32'h3bbb4c50, 32'hbc87b8f4} /* (23, 13, 12) {real, imag} */,
  {32'h3d882d14, 32'hbdb50654} /* (23, 13, 11) {real, imag} */,
  {32'h3bc835bc, 32'hbbb486f8} /* (23, 13, 10) {real, imag} */,
  {32'h3da7fdac, 32'hbc0a7d60} /* (23, 13, 9) {real, imag} */,
  {32'hbb05e9a0, 32'h3c536cf2} /* (23, 13, 8) {real, imag} */,
  {32'h3e3569e3, 32'hbd50d1d2} /* (23, 13, 7) {real, imag} */,
  {32'h3da787e3, 32'hbca2a9a4} /* (23, 13, 6) {real, imag} */,
  {32'hbe91c26a, 32'hbe02a688} /* (23, 13, 5) {real, imag} */,
  {32'h3ea13e0c, 32'h3e98083c} /* (23, 13, 4) {real, imag} */,
  {32'hbdae87e8, 32'h3c1f4f90} /* (23, 13, 3) {real, imag} */,
  {32'hbfad1131, 32'hbe231c1f} /* (23, 13, 2) {real, imag} */,
  {32'h40351305, 32'h3d58ea98} /* (23, 13, 1) {real, imag} */,
  {32'h4008f8be, 32'h00000000} /* (23, 13, 0) {real, imag} */,
  {32'h40147b31, 32'h3e34fe98} /* (23, 12, 31) {real, imag} */,
  {32'hbf928008, 32'h3dd2b5d2} /* (23, 12, 30) {real, imag} */,
  {32'hbd842e50, 32'h3c1fd7e0} /* (23, 12, 29) {real, imag} */,
  {32'h3e8712dc, 32'hbe737d13} /* (23, 12, 28) {real, imag} */,
  {32'hbe49c80e, 32'h3e98aea4} /* (23, 12, 27) {real, imag} */,
  {32'h3c6fc3a4, 32'hbd9a73a0} /* (23, 12, 26) {real, imag} */,
  {32'h3dec5088, 32'hbcb4305c} /* (23, 12, 25) {real, imag} */,
  {32'hbe053afc, 32'h3caae8f0} /* (23, 12, 24) {real, imag} */,
  {32'hbd0bd3f9, 32'h3d933e2e} /* (23, 12, 23) {real, imag} */,
  {32'h3d26b924, 32'hbd8bf754} /* (23, 12, 22) {real, imag} */,
  {32'hbcd5b642, 32'hbd0fa8a2} /* (23, 12, 21) {real, imag} */,
  {32'hbb947760, 32'hbcd34e53} /* (23, 12, 20) {real, imag} */,
  {32'hbb1f2dd8, 32'hbd1a4232} /* (23, 12, 19) {real, imag} */,
  {32'hbd168159, 32'h3db133f3} /* (23, 12, 18) {real, imag} */,
  {32'hbcd4c067, 32'h3d02f98e} /* (23, 12, 17) {real, imag} */,
  {32'h3dc64e15, 32'h00000000} /* (23, 12, 16) {real, imag} */,
  {32'hbcd4c067, 32'hbd02f98e} /* (23, 12, 15) {real, imag} */,
  {32'hbd168159, 32'hbdb133f3} /* (23, 12, 14) {real, imag} */,
  {32'hbb1f2dd8, 32'h3d1a4232} /* (23, 12, 13) {real, imag} */,
  {32'hbb947760, 32'h3cd34e53} /* (23, 12, 12) {real, imag} */,
  {32'hbcd5b642, 32'h3d0fa8a2} /* (23, 12, 11) {real, imag} */,
  {32'h3d26b924, 32'h3d8bf754} /* (23, 12, 10) {real, imag} */,
  {32'hbd0bd3f9, 32'hbd933e2e} /* (23, 12, 9) {real, imag} */,
  {32'hbe053afc, 32'hbcaae8f0} /* (23, 12, 8) {real, imag} */,
  {32'h3dec5088, 32'h3cb4305c} /* (23, 12, 7) {real, imag} */,
  {32'h3c6fc3a4, 32'h3d9a73a0} /* (23, 12, 6) {real, imag} */,
  {32'hbe49c80e, 32'hbe98aea4} /* (23, 12, 5) {real, imag} */,
  {32'h3e8712dc, 32'h3e737d13} /* (23, 12, 4) {real, imag} */,
  {32'hbd842e50, 32'hbc1fd7e0} /* (23, 12, 3) {real, imag} */,
  {32'hbf928008, 32'hbdd2b5d2} /* (23, 12, 2) {real, imag} */,
  {32'h40147b31, 32'hbe34fe98} /* (23, 12, 1) {real, imag} */,
  {32'h3fbd5ca4, 32'h00000000} /* (23, 12, 0) {real, imag} */,
  {32'h3f95d2fc, 32'h3e59ea6e} /* (23, 11, 31) {real, imag} */,
  {32'hbf38e32a, 32'hbdb4b46f} /* (23, 11, 30) {real, imag} */,
  {32'hbe3a60c0, 32'hbc797c24} /* (23, 11, 29) {real, imag} */,
  {32'h3e2a69bc, 32'hbd7d1f68} /* (23, 11, 28) {real, imag} */,
  {32'hbe38138c, 32'h3df3a763} /* (23, 11, 27) {real, imag} */,
  {32'hbd6c0231, 32'h3cab3da3} /* (23, 11, 26) {real, imag} */,
  {32'h3d95a0a8, 32'hbb3f1f00} /* (23, 11, 25) {real, imag} */,
  {32'hbd99af60, 32'h3bde940a} /* (23, 11, 24) {real, imag} */,
  {32'h3cf6e655, 32'hbd8ed31f} /* (23, 11, 23) {real, imag} */,
  {32'hbc40605a, 32'hbceb3b8e} /* (23, 11, 22) {real, imag} */,
  {32'hbd350716, 32'h3d5f210a} /* (23, 11, 21) {real, imag} */,
  {32'hbd42bc65, 32'hbb30ac08} /* (23, 11, 20) {real, imag} */,
  {32'hbd6f1ba2, 32'h3d06d379} /* (23, 11, 19) {real, imag} */,
  {32'h3cd482e4, 32'hbd875c1e} /* (23, 11, 18) {real, imag} */,
  {32'h3cafc5c0, 32'h3c46e1ac} /* (23, 11, 17) {real, imag} */,
  {32'h3db7f5b3, 32'h00000000} /* (23, 11, 16) {real, imag} */,
  {32'h3cafc5c0, 32'hbc46e1ac} /* (23, 11, 15) {real, imag} */,
  {32'h3cd482e4, 32'h3d875c1e} /* (23, 11, 14) {real, imag} */,
  {32'hbd6f1ba2, 32'hbd06d379} /* (23, 11, 13) {real, imag} */,
  {32'hbd42bc65, 32'h3b30ac08} /* (23, 11, 12) {real, imag} */,
  {32'hbd350716, 32'hbd5f210a} /* (23, 11, 11) {real, imag} */,
  {32'hbc40605a, 32'h3ceb3b8e} /* (23, 11, 10) {real, imag} */,
  {32'h3cf6e655, 32'h3d8ed31f} /* (23, 11, 9) {real, imag} */,
  {32'hbd99af60, 32'hbbde940a} /* (23, 11, 8) {real, imag} */,
  {32'h3d95a0a8, 32'h3b3f1f00} /* (23, 11, 7) {real, imag} */,
  {32'hbd6c0231, 32'hbcab3da3} /* (23, 11, 6) {real, imag} */,
  {32'hbe38138c, 32'hbdf3a763} /* (23, 11, 5) {real, imag} */,
  {32'h3e2a69bc, 32'h3d7d1f68} /* (23, 11, 4) {real, imag} */,
  {32'hbe3a60c0, 32'h3c797c24} /* (23, 11, 3) {real, imag} */,
  {32'hbf38e32a, 32'h3db4b46f} /* (23, 11, 2) {real, imag} */,
  {32'h3f95d2fc, 32'hbe59ea6e} /* (23, 11, 1) {real, imag} */,
  {32'h3f08ef3a, 32'h00000000} /* (23, 11, 0) {real, imag} */,
  {32'hbf24b28f, 32'h3f15887a} /* (23, 10, 31) {real, imag} */,
  {32'h3b80fa80, 32'hbeaff770} /* (23, 10, 30) {real, imag} */,
  {32'hbe2e0572, 32'hbd5c8e4b} /* (23, 10, 29) {real, imag} */,
  {32'h3e4e6633, 32'h3db3b628} /* (23, 10, 28) {real, imag} */,
  {32'h3e09e1d7, 32'hbd9a4a7b} /* (23, 10, 27) {real, imag} */,
  {32'hbb9e4086, 32'hbc3bfdde} /* (23, 10, 26) {real, imag} */,
  {32'hbd9d417a, 32'h3ce02c60} /* (23, 10, 25) {real, imag} */,
  {32'h3dced292, 32'h3e0e4823} /* (23, 10, 24) {real, imag} */,
  {32'h3d236099, 32'h3d0faa44} /* (23, 10, 23) {real, imag} */,
  {32'hbda2a876, 32'hbda0bc42} /* (23, 10, 22) {real, imag} */,
  {32'hbd6cfc7e, 32'hbbac7abe} /* (23, 10, 21) {real, imag} */,
  {32'h3d3646c0, 32'hbc4c46a4} /* (23, 10, 20) {real, imag} */,
  {32'h3d14af44, 32'hbd59fff6} /* (23, 10, 19) {real, imag} */,
  {32'h3cce8a88, 32'hbd1d99a7} /* (23, 10, 18) {real, imag} */,
  {32'h3cded882, 32'h3da55c2e} /* (23, 10, 17) {real, imag} */,
  {32'h3d94b030, 32'h00000000} /* (23, 10, 16) {real, imag} */,
  {32'h3cded882, 32'hbda55c2e} /* (23, 10, 15) {real, imag} */,
  {32'h3cce8a88, 32'h3d1d99a7} /* (23, 10, 14) {real, imag} */,
  {32'h3d14af44, 32'h3d59fff6} /* (23, 10, 13) {real, imag} */,
  {32'h3d3646c0, 32'h3c4c46a4} /* (23, 10, 12) {real, imag} */,
  {32'hbd6cfc7e, 32'h3bac7abe} /* (23, 10, 11) {real, imag} */,
  {32'hbda2a876, 32'h3da0bc42} /* (23, 10, 10) {real, imag} */,
  {32'h3d236099, 32'hbd0faa44} /* (23, 10, 9) {real, imag} */,
  {32'h3dced292, 32'hbe0e4823} /* (23, 10, 8) {real, imag} */,
  {32'hbd9d417a, 32'hbce02c60} /* (23, 10, 7) {real, imag} */,
  {32'hbb9e4086, 32'h3c3bfdde} /* (23, 10, 6) {real, imag} */,
  {32'h3e09e1d7, 32'h3d9a4a7b} /* (23, 10, 5) {real, imag} */,
  {32'h3e4e6633, 32'hbdb3b628} /* (23, 10, 4) {real, imag} */,
  {32'hbe2e0572, 32'h3d5c8e4b} /* (23, 10, 3) {real, imag} */,
  {32'h3b80fa80, 32'h3eaff770} /* (23, 10, 2) {real, imag} */,
  {32'hbf24b28f, 32'hbf15887a} /* (23, 10, 1) {real, imag} */,
  {32'hbf625ccf, 32'h00000000} /* (23, 10, 0) {real, imag} */,
  {32'hbff6a76c, 32'h3f84d124} /* (23, 9, 31) {real, imag} */,
  {32'h3f2e194f, 32'hbe96a720} /* (23, 9, 30) {real, imag} */,
  {32'hbd9d620e, 32'h3dcbbb5c} /* (23, 9, 29) {real, imag} */,
  {32'hbc8bc84c, 32'h3d896fda} /* (23, 9, 28) {real, imag} */,
  {32'h3e69171c, 32'hbd624dc8} /* (23, 9, 27) {real, imag} */,
  {32'h3d4c3a56, 32'hbb82ac46} /* (23, 9, 26) {real, imag} */,
  {32'h3d042977, 32'hbcc935ac} /* (23, 9, 25) {real, imag} */,
  {32'h3da55689, 32'hbd526ea6} /* (23, 9, 24) {real, imag} */,
  {32'h3cd45627, 32'h3ceccbcf} /* (23, 9, 23) {real, imag} */,
  {32'hbc803ebe, 32'h3d3f9ce4} /* (23, 9, 22) {real, imag} */,
  {32'h3d9a8f13, 32'h3ca898f8} /* (23, 9, 21) {real, imag} */,
  {32'hbd9dd556, 32'h3d2c81b9} /* (23, 9, 20) {real, imag} */,
  {32'hbd4a722e, 32'hbc0b63f4} /* (23, 9, 19) {real, imag} */,
  {32'hbc8900bd, 32'hbb8d71aa} /* (23, 9, 18) {real, imag} */,
  {32'h3d1fe26a, 32'h3cd2ae6e} /* (23, 9, 17) {real, imag} */,
  {32'hbd756e60, 32'h00000000} /* (23, 9, 16) {real, imag} */,
  {32'h3d1fe26a, 32'hbcd2ae6e} /* (23, 9, 15) {real, imag} */,
  {32'hbc8900bd, 32'h3b8d71aa} /* (23, 9, 14) {real, imag} */,
  {32'hbd4a722e, 32'h3c0b63f4} /* (23, 9, 13) {real, imag} */,
  {32'hbd9dd556, 32'hbd2c81b9} /* (23, 9, 12) {real, imag} */,
  {32'h3d9a8f13, 32'hbca898f8} /* (23, 9, 11) {real, imag} */,
  {32'hbc803ebe, 32'hbd3f9ce4} /* (23, 9, 10) {real, imag} */,
  {32'h3cd45627, 32'hbceccbcf} /* (23, 9, 9) {real, imag} */,
  {32'h3da55689, 32'h3d526ea6} /* (23, 9, 8) {real, imag} */,
  {32'h3d042977, 32'h3cc935ac} /* (23, 9, 7) {real, imag} */,
  {32'h3d4c3a56, 32'h3b82ac46} /* (23, 9, 6) {real, imag} */,
  {32'h3e69171c, 32'h3d624dc8} /* (23, 9, 5) {real, imag} */,
  {32'hbc8bc84c, 32'hbd896fda} /* (23, 9, 4) {real, imag} */,
  {32'hbd9d620e, 32'hbdcbbb5c} /* (23, 9, 3) {real, imag} */,
  {32'h3f2e194f, 32'h3e96a720} /* (23, 9, 2) {real, imag} */,
  {32'hbff6a76c, 32'hbf84d124} /* (23, 9, 1) {real, imag} */,
  {32'hc00b7d1a, 32'h00000000} /* (23, 9, 0) {real, imag} */,
  {32'hc030b814, 32'h3fb8ab3e} /* (23, 8, 31) {real, imag} */,
  {32'h3f6316c7, 32'hbee5fbc0} /* (23, 8, 30) {real, imag} */,
  {32'h3e18f415, 32'h3db5d76a} /* (23, 8, 29) {real, imag} */,
  {32'hbe0eedc1, 32'h3db2339f} /* (23, 8, 28) {real, imag} */,
  {32'h3e3c80c4, 32'hbdfe296b} /* (23, 8, 27) {real, imag} */,
  {32'h3dfa7be8, 32'hbca6c0f6} /* (23, 8, 26) {real, imag} */,
  {32'hbd885378, 32'h3d9fe3e0} /* (23, 8, 25) {real, imag} */,
  {32'h3d7ade62, 32'h3c500b94} /* (23, 8, 24) {real, imag} */,
  {32'hbde21a72, 32'h3d877aa7} /* (23, 8, 23) {real, imag} */,
  {32'h3d034a9d, 32'hbe044ffd} /* (23, 8, 22) {real, imag} */,
  {32'h3d3fd98b, 32'h3d15ef3a} /* (23, 8, 21) {real, imag} */,
  {32'hbe24ce81, 32'hbd6ccff8} /* (23, 8, 20) {real, imag} */,
  {32'h3d0c7552, 32'h3d4483bd} /* (23, 8, 19) {real, imag} */,
  {32'h3c24a210, 32'hbd451633} /* (23, 8, 18) {real, imag} */,
  {32'h3ca92d00, 32'hbd3a8a0a} /* (23, 8, 17) {real, imag} */,
  {32'h3d0b68c1, 32'h00000000} /* (23, 8, 16) {real, imag} */,
  {32'h3ca92d00, 32'h3d3a8a0a} /* (23, 8, 15) {real, imag} */,
  {32'h3c24a210, 32'h3d451633} /* (23, 8, 14) {real, imag} */,
  {32'h3d0c7552, 32'hbd4483bd} /* (23, 8, 13) {real, imag} */,
  {32'hbe24ce81, 32'h3d6ccff8} /* (23, 8, 12) {real, imag} */,
  {32'h3d3fd98b, 32'hbd15ef3a} /* (23, 8, 11) {real, imag} */,
  {32'h3d034a9d, 32'h3e044ffd} /* (23, 8, 10) {real, imag} */,
  {32'hbde21a72, 32'hbd877aa7} /* (23, 8, 9) {real, imag} */,
  {32'h3d7ade62, 32'hbc500b94} /* (23, 8, 8) {real, imag} */,
  {32'hbd885378, 32'hbd9fe3e0} /* (23, 8, 7) {real, imag} */,
  {32'h3dfa7be8, 32'h3ca6c0f6} /* (23, 8, 6) {real, imag} */,
  {32'h3e3c80c4, 32'h3dfe296b} /* (23, 8, 5) {real, imag} */,
  {32'hbe0eedc1, 32'hbdb2339f} /* (23, 8, 4) {real, imag} */,
  {32'h3e18f415, 32'hbdb5d76a} /* (23, 8, 3) {real, imag} */,
  {32'h3f6316c7, 32'h3ee5fbc0} /* (23, 8, 2) {real, imag} */,
  {32'hc030b814, 32'hbfb8ab3e} /* (23, 8, 1) {real, imag} */,
  {32'hc0446c44, 32'h00000000} /* (23, 8, 0) {real, imag} */,
  {32'hc0485fc9, 32'h3fdb29a6} /* (23, 7, 31) {real, imag} */,
  {32'h3f6f3921, 32'hbecb0544} /* (23, 7, 30) {real, imag} */,
  {32'h3dc91dbe, 32'hbdbbfd38} /* (23, 7, 29) {real, imag} */,
  {32'hbdf16274, 32'hbcd75dce} /* (23, 7, 28) {real, imag} */,
  {32'h3e09a334, 32'hbde46984} /* (23, 7, 27) {real, imag} */,
  {32'h3d702da6, 32'hbdcc1636} /* (23, 7, 26) {real, imag} */,
  {32'hbdcb581e, 32'h3cdb7b2d} /* (23, 7, 25) {real, imag} */,
  {32'h3dedb8ec, 32'h3c8f2c16} /* (23, 7, 24) {real, imag} */,
  {32'h3db17c80, 32'hbad53080} /* (23, 7, 23) {real, imag} */,
  {32'h3c24d5e1, 32'h3d8b2079} /* (23, 7, 22) {real, imag} */,
  {32'hbd2d6217, 32'h3b35a340} /* (23, 7, 21) {real, imag} */,
  {32'h3dad6600, 32'h3c8f8e1a} /* (23, 7, 20) {real, imag} */,
  {32'h3c3f0f7c, 32'hbd815748} /* (23, 7, 19) {real, imag} */,
  {32'h3d1c745f, 32'h3caca27e} /* (23, 7, 18) {real, imag} */,
  {32'h3b89d364, 32'h3d9b9c26} /* (23, 7, 17) {real, imag} */,
  {32'hbd2adc6c, 32'h00000000} /* (23, 7, 16) {real, imag} */,
  {32'h3b89d364, 32'hbd9b9c26} /* (23, 7, 15) {real, imag} */,
  {32'h3d1c745f, 32'hbcaca27e} /* (23, 7, 14) {real, imag} */,
  {32'h3c3f0f7c, 32'h3d815748} /* (23, 7, 13) {real, imag} */,
  {32'h3dad6600, 32'hbc8f8e1a} /* (23, 7, 12) {real, imag} */,
  {32'hbd2d6217, 32'hbb35a340} /* (23, 7, 11) {real, imag} */,
  {32'h3c24d5e1, 32'hbd8b2079} /* (23, 7, 10) {real, imag} */,
  {32'h3db17c80, 32'h3ad53080} /* (23, 7, 9) {real, imag} */,
  {32'h3dedb8ec, 32'hbc8f2c16} /* (23, 7, 8) {real, imag} */,
  {32'hbdcb581e, 32'hbcdb7b2d} /* (23, 7, 7) {real, imag} */,
  {32'h3d702da6, 32'h3dcc1636} /* (23, 7, 6) {real, imag} */,
  {32'h3e09a334, 32'h3de46984} /* (23, 7, 5) {real, imag} */,
  {32'hbdf16274, 32'h3cd75dce} /* (23, 7, 4) {real, imag} */,
  {32'h3dc91dbe, 32'h3dbbfd38} /* (23, 7, 3) {real, imag} */,
  {32'h3f6f3921, 32'h3ecb0544} /* (23, 7, 2) {real, imag} */,
  {32'hc0485fc9, 32'hbfdb29a6} /* (23, 7, 1) {real, imag} */,
  {32'hc06df3f4, 32'h00000000} /* (23, 7, 0) {real, imag} */,
  {32'hc0543844, 32'h400b3ef6} /* (23, 6, 31) {real, imag} */,
  {32'h3f3ea0fb, 32'hbf17c97a} /* (23, 6, 30) {real, imag} */,
  {32'h3d38c9a2, 32'h3d5cbc2d} /* (23, 6, 29) {real, imag} */,
  {32'hbdfc44c2, 32'h3cdf9b3a} /* (23, 6, 28) {real, imag} */,
  {32'h3dfa863e, 32'hbdd403cb} /* (23, 6, 27) {real, imag} */,
  {32'hbc36d3a3, 32'hbc69003e} /* (23, 6, 26) {real, imag} */,
  {32'hbd979839, 32'hbc7ad7b8} /* (23, 6, 25) {real, imag} */,
  {32'h3d631a81, 32'hbd75a252} /* (23, 6, 24) {real, imag} */,
  {32'hbbd4d838, 32'h3bb27d24} /* (23, 6, 23) {real, imag} */,
  {32'hbd7f8c48, 32'h3d0d22a0} /* (23, 6, 22) {real, imag} */,
  {32'hbd264d45, 32'hbd684e89} /* (23, 6, 21) {real, imag} */,
  {32'h3c878788, 32'hbbb21ba0} /* (23, 6, 20) {real, imag} */,
  {32'hbd14f676, 32'hbbdbc55c} /* (23, 6, 19) {real, imag} */,
  {32'h3d0a10ac, 32'hbc024066} /* (23, 6, 18) {real, imag} */,
  {32'hbcc702fb, 32'h3cf44754} /* (23, 6, 17) {real, imag} */,
  {32'hbcf430c7, 32'h00000000} /* (23, 6, 16) {real, imag} */,
  {32'hbcc702fb, 32'hbcf44754} /* (23, 6, 15) {real, imag} */,
  {32'h3d0a10ac, 32'h3c024066} /* (23, 6, 14) {real, imag} */,
  {32'hbd14f676, 32'h3bdbc55c} /* (23, 6, 13) {real, imag} */,
  {32'h3c878788, 32'h3bb21ba0} /* (23, 6, 12) {real, imag} */,
  {32'hbd264d45, 32'h3d684e89} /* (23, 6, 11) {real, imag} */,
  {32'hbd7f8c48, 32'hbd0d22a0} /* (23, 6, 10) {real, imag} */,
  {32'hbbd4d838, 32'hbbb27d24} /* (23, 6, 9) {real, imag} */,
  {32'h3d631a81, 32'h3d75a252} /* (23, 6, 8) {real, imag} */,
  {32'hbd979839, 32'h3c7ad7b8} /* (23, 6, 7) {real, imag} */,
  {32'hbc36d3a3, 32'h3c69003e} /* (23, 6, 6) {real, imag} */,
  {32'h3dfa863e, 32'h3dd403cb} /* (23, 6, 5) {real, imag} */,
  {32'hbdfc44c2, 32'hbcdf9b3a} /* (23, 6, 4) {real, imag} */,
  {32'h3d38c9a2, 32'hbd5cbc2d} /* (23, 6, 3) {real, imag} */,
  {32'h3f3ea0fb, 32'h3f17c97a} /* (23, 6, 2) {real, imag} */,
  {32'hc0543844, 32'hc00b3ef6} /* (23, 6, 1) {real, imag} */,
  {32'hc0810825, 32'h00000000} /* (23, 6, 0) {real, imag} */,
  {32'hc04c8eeb, 32'h4038d601} /* (23, 5, 31) {real, imag} */,
  {32'h3e675b68, 32'hbf2c2312} /* (23, 5, 30) {real, imag} */,
  {32'h3dd822fa, 32'hbcbc0a9c} /* (23, 5, 29) {real, imag} */,
  {32'h3cb17936, 32'hbd68171f} /* (23, 5, 28) {real, imag} */,
  {32'h3e08380c, 32'h3cab0a38} /* (23, 5, 27) {real, imag} */,
  {32'hbc6f22c2, 32'hbce6a824} /* (23, 5, 26) {real, imag} */,
  {32'h3c87a3a0, 32'h3a312500} /* (23, 5, 25) {real, imag} */,
  {32'hbd8ff56a, 32'h3c261c8d} /* (23, 5, 24) {real, imag} */,
  {32'h3cc56b88, 32'hbd075910} /* (23, 5, 23) {real, imag} */,
  {32'hbdbf54e2, 32'hbd08eafa} /* (23, 5, 22) {real, imag} */,
  {32'h3d1af306, 32'hbceea3c9} /* (23, 5, 21) {real, imag} */,
  {32'h3b2be9ec, 32'h3d9894ee} /* (23, 5, 20) {real, imag} */,
  {32'hbcc303b4, 32'h3d0dd1ab} /* (23, 5, 19) {real, imag} */,
  {32'h3c033a78, 32'hbd0aea1c} /* (23, 5, 18) {real, imag} */,
  {32'h3d62489e, 32'hbd502641} /* (23, 5, 17) {real, imag} */,
  {32'h3b840208, 32'h00000000} /* (23, 5, 16) {real, imag} */,
  {32'h3d62489e, 32'h3d502641} /* (23, 5, 15) {real, imag} */,
  {32'h3c033a78, 32'h3d0aea1c} /* (23, 5, 14) {real, imag} */,
  {32'hbcc303b4, 32'hbd0dd1ab} /* (23, 5, 13) {real, imag} */,
  {32'h3b2be9ec, 32'hbd9894ee} /* (23, 5, 12) {real, imag} */,
  {32'h3d1af306, 32'h3ceea3c9} /* (23, 5, 11) {real, imag} */,
  {32'hbdbf54e2, 32'h3d08eafa} /* (23, 5, 10) {real, imag} */,
  {32'h3cc56b88, 32'h3d075910} /* (23, 5, 9) {real, imag} */,
  {32'hbd8ff56a, 32'hbc261c8d} /* (23, 5, 8) {real, imag} */,
  {32'h3c87a3a0, 32'hba312500} /* (23, 5, 7) {real, imag} */,
  {32'hbc6f22c2, 32'h3ce6a824} /* (23, 5, 6) {real, imag} */,
  {32'h3e08380c, 32'hbcab0a38} /* (23, 5, 5) {real, imag} */,
  {32'h3cb17936, 32'h3d68171f} /* (23, 5, 4) {real, imag} */,
  {32'h3dd822fa, 32'h3cbc0a9c} /* (23, 5, 3) {real, imag} */,
  {32'h3e675b68, 32'h3f2c2312} /* (23, 5, 2) {real, imag} */,
  {32'hc04c8eeb, 32'hc038d601} /* (23, 5, 1) {real, imag} */,
  {32'hc0914ed7, 32'h00000000} /* (23, 5, 0) {real, imag} */,
  {32'hc0463803, 32'h405c3d95} /* (23, 4, 31) {real, imag} */,
  {32'hbd8c95f0, 32'hbf2ffb0e} /* (23, 4, 30) {real, imag} */,
  {32'h3e116c9c, 32'hbe02d2ef} /* (23, 4, 29) {real, imag} */,
  {32'h3e08d1ef, 32'hbe5328a2} /* (23, 4, 28) {real, imag} */,
  {32'h3e3fb7a6, 32'h3e19233e} /* (23, 4, 27) {real, imag} */,
  {32'h3de380a6, 32'h3e03b274} /* (23, 4, 26) {real, imag} */,
  {32'h3dc2e41e, 32'hba465280} /* (23, 4, 25) {real, imag} */,
  {32'hbdb2ffbf, 32'h3c8484b0} /* (23, 4, 24) {real, imag} */,
  {32'h3d213677, 32'hbd856a3e} /* (23, 4, 23) {real, imag} */,
  {32'h3d2c2ee0, 32'hbd76975a} /* (23, 4, 22) {real, imag} */,
  {32'h3cc64808, 32'h3d85cd83} /* (23, 4, 21) {real, imag} */,
  {32'h3bc01d66, 32'hbddc4ff0} /* (23, 4, 20) {real, imag} */,
  {32'hbd0cb715, 32'h3cad930a} /* (23, 4, 19) {real, imag} */,
  {32'h3b6d05a0, 32'hbd1f2f5c} /* (23, 4, 18) {real, imag} */,
  {32'h3cd7f242, 32'hbd599b9c} /* (23, 4, 17) {real, imag} */,
  {32'hbc47e9f8, 32'h00000000} /* (23, 4, 16) {real, imag} */,
  {32'h3cd7f242, 32'h3d599b9c} /* (23, 4, 15) {real, imag} */,
  {32'h3b6d05a0, 32'h3d1f2f5c} /* (23, 4, 14) {real, imag} */,
  {32'hbd0cb715, 32'hbcad930a} /* (23, 4, 13) {real, imag} */,
  {32'h3bc01d66, 32'h3ddc4ff0} /* (23, 4, 12) {real, imag} */,
  {32'h3cc64808, 32'hbd85cd83} /* (23, 4, 11) {real, imag} */,
  {32'h3d2c2ee0, 32'h3d76975a} /* (23, 4, 10) {real, imag} */,
  {32'h3d213677, 32'h3d856a3e} /* (23, 4, 9) {real, imag} */,
  {32'hbdb2ffbf, 32'hbc8484b0} /* (23, 4, 8) {real, imag} */,
  {32'h3dc2e41e, 32'h3a465280} /* (23, 4, 7) {real, imag} */,
  {32'h3de380a6, 32'hbe03b274} /* (23, 4, 6) {real, imag} */,
  {32'h3e3fb7a6, 32'hbe19233e} /* (23, 4, 5) {real, imag} */,
  {32'h3e08d1ef, 32'h3e5328a2} /* (23, 4, 4) {real, imag} */,
  {32'h3e116c9c, 32'h3e02d2ef} /* (23, 4, 3) {real, imag} */,
  {32'hbd8c95f0, 32'h3f2ffb0e} /* (23, 4, 2) {real, imag} */,
  {32'hc0463803, 32'hc05c3d95} /* (23, 4, 1) {real, imag} */,
  {32'hc09cc802, 32'h00000000} /* (23, 4, 0) {real, imag} */,
  {32'hc04b27fd, 32'h40631154} /* (23, 3, 31) {real, imag} */,
  {32'hbebab94a, 32'hbf5c0adf} /* (23, 3, 30) {real, imag} */,
  {32'h3df70486, 32'h3c06a898} /* (23, 3, 29) {real, imag} */,
  {32'h3d6929fe, 32'hbe9df64f} /* (23, 3, 28) {real, imag} */,
  {32'h3e6b9ec5, 32'h3e135c7d} /* (23, 3, 27) {real, imag} */,
  {32'h3e0a179a, 32'h3c73140c} /* (23, 3, 26) {real, imag} */,
  {32'h3d337533, 32'h3e05bd04} /* (23, 3, 25) {real, imag} */,
  {32'hbd434851, 32'hbd2c80d8} /* (23, 3, 24) {real, imag} */,
  {32'h3d95c05a, 32'hbcc90673} /* (23, 3, 23) {real, imag} */,
  {32'h3bd39e28, 32'h3b9d1660} /* (23, 3, 22) {real, imag} */,
  {32'h3d23639a, 32'hbcfd7728} /* (23, 3, 21) {real, imag} */,
  {32'hbcd14d57, 32'h3ab72168} /* (23, 3, 20) {real, imag} */,
  {32'h3c3a7390, 32'hbd84ffd2} /* (23, 3, 19) {real, imag} */,
  {32'hbdde51b6, 32'h3d8ef7d4} /* (23, 3, 18) {real, imag} */,
  {32'hbcef2eb1, 32'hbcf5f0d5} /* (23, 3, 17) {real, imag} */,
  {32'hbe1f5d9a, 32'h00000000} /* (23, 3, 16) {real, imag} */,
  {32'hbcef2eb1, 32'h3cf5f0d5} /* (23, 3, 15) {real, imag} */,
  {32'hbdde51b6, 32'hbd8ef7d4} /* (23, 3, 14) {real, imag} */,
  {32'h3c3a7390, 32'h3d84ffd2} /* (23, 3, 13) {real, imag} */,
  {32'hbcd14d57, 32'hbab72168} /* (23, 3, 12) {real, imag} */,
  {32'h3d23639a, 32'h3cfd7728} /* (23, 3, 11) {real, imag} */,
  {32'h3bd39e28, 32'hbb9d1660} /* (23, 3, 10) {real, imag} */,
  {32'h3d95c05a, 32'h3cc90673} /* (23, 3, 9) {real, imag} */,
  {32'hbd434851, 32'h3d2c80d8} /* (23, 3, 8) {real, imag} */,
  {32'h3d337533, 32'hbe05bd04} /* (23, 3, 7) {real, imag} */,
  {32'h3e0a179a, 32'hbc73140c} /* (23, 3, 6) {real, imag} */,
  {32'h3e6b9ec5, 32'hbe135c7d} /* (23, 3, 5) {real, imag} */,
  {32'h3d6929fe, 32'h3e9df64f} /* (23, 3, 4) {real, imag} */,
  {32'h3df70486, 32'hbc06a898} /* (23, 3, 3) {real, imag} */,
  {32'hbebab94a, 32'h3f5c0adf} /* (23, 3, 2) {real, imag} */,
  {32'hc04b27fd, 32'hc0631154} /* (23, 3, 1) {real, imag} */,
  {32'hc09e39b4, 32'h00000000} /* (23, 3, 0) {real, imag} */,
  {32'hc03f4755, 32'h406401f6} /* (23, 2, 31) {real, imag} */,
  {32'hbe84ec55, 32'hbf564150} /* (23, 2, 30) {real, imag} */,
  {32'h3e5e3f74, 32'h3c01f212} /* (23, 2, 29) {real, imag} */,
  {32'h3d238cf8, 32'hbeb2d2a4} /* (23, 2, 28) {real, imag} */,
  {32'h3e9a624b, 32'hbccfb150} /* (23, 2, 27) {real, imag} */,
  {32'hbd002c8c, 32'h3c0e8060} /* (23, 2, 26) {real, imag} */,
  {32'h3d8f230e, 32'h3dce2692} /* (23, 2, 25) {real, imag} */,
  {32'hbdd26c96, 32'h3be14d58} /* (23, 2, 24) {real, imag} */,
  {32'hbc70cb9e, 32'hbde83dfa} /* (23, 2, 23) {real, imag} */,
  {32'hbd892f04, 32'h3daefe5e} /* (23, 2, 22) {real, imag} */,
  {32'h3da488d3, 32'h3d42097c} /* (23, 2, 21) {real, imag} */,
  {32'h3a5ffe80, 32'h3e022782} /* (23, 2, 20) {real, imag} */,
  {32'hbd9812b4, 32'h3dcec2d0} /* (23, 2, 19) {real, imag} */,
  {32'h3acfa1a0, 32'hbd62768a} /* (23, 2, 18) {real, imag} */,
  {32'h3d0f46e7, 32'hbd5f5ade} /* (23, 2, 17) {real, imag} */,
  {32'hbd8452b6, 32'h00000000} /* (23, 2, 16) {real, imag} */,
  {32'h3d0f46e7, 32'h3d5f5ade} /* (23, 2, 15) {real, imag} */,
  {32'h3acfa1a0, 32'h3d62768a} /* (23, 2, 14) {real, imag} */,
  {32'hbd9812b4, 32'hbdcec2d0} /* (23, 2, 13) {real, imag} */,
  {32'h3a5ffe80, 32'hbe022782} /* (23, 2, 12) {real, imag} */,
  {32'h3da488d3, 32'hbd42097c} /* (23, 2, 11) {real, imag} */,
  {32'hbd892f04, 32'hbdaefe5e} /* (23, 2, 10) {real, imag} */,
  {32'hbc70cb9e, 32'h3de83dfa} /* (23, 2, 9) {real, imag} */,
  {32'hbdd26c96, 32'hbbe14d58} /* (23, 2, 8) {real, imag} */,
  {32'h3d8f230e, 32'hbdce2692} /* (23, 2, 7) {real, imag} */,
  {32'hbd002c8c, 32'hbc0e8060} /* (23, 2, 6) {real, imag} */,
  {32'h3e9a624b, 32'h3ccfb150} /* (23, 2, 5) {real, imag} */,
  {32'h3d238cf8, 32'h3eb2d2a4} /* (23, 2, 4) {real, imag} */,
  {32'h3e5e3f74, 32'hbc01f212} /* (23, 2, 3) {real, imag} */,
  {32'hbe84ec55, 32'h3f564150} /* (23, 2, 2) {real, imag} */,
  {32'hc03f4755, 32'hc06401f6} /* (23, 2, 1) {real, imag} */,
  {32'hc0a4b13c, 32'h00000000} /* (23, 2, 0) {real, imag} */,
  {32'hc043445e, 32'h40537ada} /* (23, 1, 31) {real, imag} */,
  {32'hbe17e736, 32'hbf25f07e} /* (23, 1, 30) {real, imag} */,
  {32'h3e9e758e, 32'hbd10d2b2} /* (23, 1, 29) {real, imag} */,
  {32'h3dae3520, 32'hbe9d918e} /* (23, 1, 28) {real, imag} */,
  {32'h3e5f1122, 32'h3d66febe} /* (23, 1, 27) {real, imag} */,
  {32'hbdd617c7, 32'h3d377366} /* (23, 1, 26) {real, imag} */,
  {32'hbcf281fc, 32'hbc14f8d0} /* (23, 1, 25) {real, imag} */,
  {32'h3cc7c2d0, 32'hbb58eff8} /* (23, 1, 24) {real, imag} */,
  {32'h3d43d84e, 32'h3d03f198} /* (23, 1, 23) {real, imag} */,
  {32'hbda02d57, 32'hbdd87cca} /* (23, 1, 22) {real, imag} */,
  {32'h3d74bfdc, 32'hbd34210c} /* (23, 1, 21) {real, imag} */,
  {32'hbd3f925a, 32'h3d1231ec} /* (23, 1, 20) {real, imag} */,
  {32'hbd498c42, 32'h3cf2cb02} /* (23, 1, 19) {real, imag} */,
  {32'hbcbf0533, 32'hbcc4c636} /* (23, 1, 18) {real, imag} */,
  {32'h3d968a65, 32'hbd47b14c} /* (23, 1, 17) {real, imag} */,
  {32'h3d925085, 32'h00000000} /* (23, 1, 16) {real, imag} */,
  {32'h3d968a65, 32'h3d47b14c} /* (23, 1, 15) {real, imag} */,
  {32'hbcbf0533, 32'h3cc4c636} /* (23, 1, 14) {real, imag} */,
  {32'hbd498c42, 32'hbcf2cb02} /* (23, 1, 13) {real, imag} */,
  {32'hbd3f925a, 32'hbd1231ec} /* (23, 1, 12) {real, imag} */,
  {32'h3d74bfdc, 32'h3d34210c} /* (23, 1, 11) {real, imag} */,
  {32'hbda02d57, 32'h3dd87cca} /* (23, 1, 10) {real, imag} */,
  {32'h3d43d84e, 32'hbd03f198} /* (23, 1, 9) {real, imag} */,
  {32'h3cc7c2d0, 32'h3b58eff8} /* (23, 1, 8) {real, imag} */,
  {32'hbcf281fc, 32'h3c14f8d0} /* (23, 1, 7) {real, imag} */,
  {32'hbdd617c7, 32'hbd377366} /* (23, 1, 6) {real, imag} */,
  {32'h3e5f1122, 32'hbd66febe} /* (23, 1, 5) {real, imag} */,
  {32'h3dae3520, 32'h3e9d918e} /* (23, 1, 4) {real, imag} */,
  {32'h3e9e758e, 32'h3d10d2b2} /* (23, 1, 3) {real, imag} */,
  {32'hbe17e736, 32'h3f25f07e} /* (23, 1, 2) {real, imag} */,
  {32'hc043445e, 32'hc0537ada} /* (23, 1, 1) {real, imag} */,
  {32'hc09860d5, 32'h00000000} /* (23, 1, 0) {real, imag} */,
  {32'hc04ce74e, 32'h402c21bf} /* (23, 0, 31) {real, imag} */,
  {32'h3e565a38, 32'hbee30377} /* (23, 0, 30) {real, imag} */,
  {32'h3e0ea3bf, 32'hbc3d9fd4} /* (23, 0, 29) {real, imag} */,
  {32'h3d8bb0c8, 32'hbe65a2cc} /* (23, 0, 28) {real, imag} */,
  {32'h3d33790c, 32'h3db7502b} /* (23, 0, 27) {real, imag} */,
  {32'hbadbf280, 32'hbd185360} /* (23, 0, 26) {real, imag} */,
  {32'h3d003b10, 32'h3ba1d0b8} /* (23, 0, 25) {real, imag} */,
  {32'h3d05e2ed, 32'h3c998b76} /* (23, 0, 24) {real, imag} */,
  {32'h3d92c37c, 32'h3d683f9a} /* (23, 0, 23) {real, imag} */,
  {32'h39bcf6b0, 32'hbdbe6e5a} /* (23, 0, 22) {real, imag} */,
  {32'hbd9cffce, 32'hbd1eff03} /* (23, 0, 21) {real, imag} */,
  {32'h3cb94a76, 32'h3c8832dc} /* (23, 0, 20) {real, imag} */,
  {32'h3b887912, 32'h3d0ca853} /* (23, 0, 19) {real, imag} */,
  {32'hbd3188ea, 32'h3d07139c} /* (23, 0, 18) {real, imag} */,
  {32'h3c89195d, 32'hbd60fc60} /* (23, 0, 17) {real, imag} */,
  {32'h3d6814a8, 32'h00000000} /* (23, 0, 16) {real, imag} */,
  {32'h3c89195d, 32'h3d60fc60} /* (23, 0, 15) {real, imag} */,
  {32'hbd3188ea, 32'hbd07139c} /* (23, 0, 14) {real, imag} */,
  {32'h3b887912, 32'hbd0ca853} /* (23, 0, 13) {real, imag} */,
  {32'h3cb94a76, 32'hbc8832dc} /* (23, 0, 12) {real, imag} */,
  {32'hbd9cffce, 32'h3d1eff03} /* (23, 0, 11) {real, imag} */,
  {32'h39bcf6b0, 32'h3dbe6e5a} /* (23, 0, 10) {real, imag} */,
  {32'h3d92c37c, 32'hbd683f9a} /* (23, 0, 9) {real, imag} */,
  {32'h3d05e2ed, 32'hbc998b76} /* (23, 0, 8) {real, imag} */,
  {32'h3d003b10, 32'hbba1d0b8} /* (23, 0, 7) {real, imag} */,
  {32'hbadbf280, 32'h3d185360} /* (23, 0, 6) {real, imag} */,
  {32'h3d33790c, 32'hbdb7502b} /* (23, 0, 5) {real, imag} */,
  {32'h3d8bb0c8, 32'h3e65a2cc} /* (23, 0, 4) {real, imag} */,
  {32'h3e0ea3bf, 32'h3c3d9fd4} /* (23, 0, 3) {real, imag} */,
  {32'h3e565a38, 32'h3ee30377} /* (23, 0, 2) {real, imag} */,
  {32'hc04ce74e, 32'hc02c21bf} /* (23, 0, 1) {real, imag} */,
  {32'hc0967900, 32'h00000000} /* (23, 0, 0) {real, imag} */,
  {32'hc07d526d, 32'h40153968} /* (22, 31, 31) {real, imag} */,
  {32'h3f3c123b, 32'hbedce955} /* (22, 31, 30) {real, imag} */,
  {32'h3cb07878, 32'h3cbf9e88} /* (22, 31, 29) {real, imag} */,
  {32'hbdefaa3a, 32'hbce035f8} /* (22, 31, 28) {real, imag} */,
  {32'h3dbe0aa6, 32'hbcbc9630} /* (22, 31, 27) {real, imag} */,
  {32'h3d205888, 32'hbc735a26} /* (22, 31, 26) {real, imag} */,
  {32'hbd4fca44, 32'h3cb65660} /* (22, 31, 25) {real, imag} */,
  {32'hbba72e34, 32'hbd592186} /* (22, 31, 24) {real, imag} */,
  {32'h3aebc888, 32'h3cd8b79a} /* (22, 31, 23) {real, imag} */,
  {32'h3dc8b8ac, 32'hbd56b8bc} /* (22, 31, 22) {real, imag} */,
  {32'h3d03bc4c, 32'hba5302e0} /* (22, 31, 21) {real, imag} */,
  {32'hbcfbf2a1, 32'hbd8a1b70} /* (22, 31, 20) {real, imag} */,
  {32'h3d568739, 32'h3d4e8e96} /* (22, 31, 19) {real, imag} */,
  {32'h3d05ee50, 32'h3c38cb36} /* (22, 31, 18) {real, imag} */,
  {32'hbc0e1496, 32'h3bb63462} /* (22, 31, 17) {real, imag} */,
  {32'h3bd557e6, 32'h00000000} /* (22, 31, 16) {real, imag} */,
  {32'hbc0e1496, 32'hbbb63462} /* (22, 31, 15) {real, imag} */,
  {32'h3d05ee50, 32'hbc38cb36} /* (22, 31, 14) {real, imag} */,
  {32'h3d568739, 32'hbd4e8e96} /* (22, 31, 13) {real, imag} */,
  {32'hbcfbf2a1, 32'h3d8a1b70} /* (22, 31, 12) {real, imag} */,
  {32'h3d03bc4c, 32'h3a5302e0} /* (22, 31, 11) {real, imag} */,
  {32'h3dc8b8ac, 32'h3d56b8bc} /* (22, 31, 10) {real, imag} */,
  {32'h3aebc888, 32'hbcd8b79a} /* (22, 31, 9) {real, imag} */,
  {32'hbba72e34, 32'h3d592186} /* (22, 31, 8) {real, imag} */,
  {32'hbd4fca44, 32'hbcb65660} /* (22, 31, 7) {real, imag} */,
  {32'h3d205888, 32'h3c735a26} /* (22, 31, 6) {real, imag} */,
  {32'h3dbe0aa6, 32'h3cbc9630} /* (22, 31, 5) {real, imag} */,
  {32'hbdefaa3a, 32'h3ce035f8} /* (22, 31, 4) {real, imag} */,
  {32'h3cb07878, 32'hbcbf9e88} /* (22, 31, 3) {real, imag} */,
  {32'h3f3c123b, 32'h3edce955} /* (22, 31, 2) {real, imag} */,
  {32'hc07d526d, 32'hc0153968} /* (22, 31, 1) {real, imag} */,
  {32'hc0a381fb, 32'h00000000} /* (22, 31, 0) {real, imag} */,
  {32'hc08fe08b, 32'h3ffb98f6} /* (22, 30, 31) {real, imag} */,
  {32'h3f9c5391, 32'hbec3e39c} /* (22, 30, 30) {real, imag} */,
  {32'hbd0599ea, 32'hbcb83612} /* (22, 30, 29) {real, imag} */,
  {32'hbe9fce2d, 32'h3c881eb0} /* (22, 30, 28) {real, imag} */,
  {32'h3e6c2e92, 32'h3d0d6cbe} /* (22, 30, 27) {real, imag} */,
  {32'h3d1293e1, 32'hbba23d40} /* (22, 30, 26) {real, imag} */,
  {32'hbd744db7, 32'hbd8f8763} /* (22, 30, 25) {real, imag} */,
  {32'h3cf119d0, 32'hbdb0686f} /* (22, 30, 24) {real, imag} */,
  {32'hbe024fcf, 32'hbd0b003c} /* (22, 30, 23) {real, imag} */,
  {32'h3da5f1e2, 32'h3cda5a7e} /* (22, 30, 22) {real, imag} */,
  {32'h3da5e53f, 32'h3ca901f8} /* (22, 30, 21) {real, imag} */,
  {32'hbd8be628, 32'h3c9a224e} /* (22, 30, 20) {real, imag} */,
  {32'h3d13ce5c, 32'h3d77e912} /* (22, 30, 19) {real, imag} */,
  {32'h3ce7bb7f, 32'hbdc9b0da} /* (22, 30, 18) {real, imag} */,
  {32'hbcfd60c9, 32'hbcf7593e} /* (22, 30, 17) {real, imag} */,
  {32'h3d4eac42, 32'h00000000} /* (22, 30, 16) {real, imag} */,
  {32'hbcfd60c9, 32'h3cf7593e} /* (22, 30, 15) {real, imag} */,
  {32'h3ce7bb7f, 32'h3dc9b0da} /* (22, 30, 14) {real, imag} */,
  {32'h3d13ce5c, 32'hbd77e912} /* (22, 30, 13) {real, imag} */,
  {32'hbd8be628, 32'hbc9a224e} /* (22, 30, 12) {real, imag} */,
  {32'h3da5e53f, 32'hbca901f8} /* (22, 30, 11) {real, imag} */,
  {32'h3da5f1e2, 32'hbcda5a7e} /* (22, 30, 10) {real, imag} */,
  {32'hbe024fcf, 32'h3d0b003c} /* (22, 30, 9) {real, imag} */,
  {32'h3cf119d0, 32'h3db0686f} /* (22, 30, 8) {real, imag} */,
  {32'hbd744db7, 32'h3d8f8763} /* (22, 30, 7) {real, imag} */,
  {32'h3d1293e1, 32'h3ba23d40} /* (22, 30, 6) {real, imag} */,
  {32'h3e6c2e92, 32'hbd0d6cbe} /* (22, 30, 5) {real, imag} */,
  {32'hbe9fce2d, 32'hbc881eb0} /* (22, 30, 4) {real, imag} */,
  {32'hbd0599ea, 32'h3cb83612} /* (22, 30, 3) {real, imag} */,
  {32'h3f9c5391, 32'h3ec3e39c} /* (22, 30, 2) {real, imag} */,
  {32'hc08fe08b, 32'hbffb98f6} /* (22, 30, 1) {real, imag} */,
  {32'hc0ab546d, 32'h00000000} /* (22, 30, 0) {real, imag} */,
  {32'hc09db42a, 32'h3fcba777} /* (22, 29, 31) {real, imag} */,
  {32'h3fc401aa, 32'hbeb2acc2} /* (22, 29, 30) {real, imag} */,
  {32'hbdb68426, 32'hbd616c00} /* (22, 29, 29) {real, imag} */,
  {32'hbe85da77, 32'h3dc63643} /* (22, 29, 28) {real, imag} */,
  {32'h3e4ae450, 32'hbe5e9cdf} /* (22, 29, 27) {real, imag} */,
  {32'hbd809994, 32'hbd659a61} /* (22, 29, 26) {real, imag} */,
  {32'hbd60b0bb, 32'hbd27730a} /* (22, 29, 25) {real, imag} */,
  {32'h3d6d6d5c, 32'hbe3012c8} /* (22, 29, 24) {real, imag} */,
  {32'hbd2284e2, 32'hbc3d5c16} /* (22, 29, 23) {real, imag} */,
  {32'h3e0b15ac, 32'hbcdb9f74} /* (22, 29, 22) {real, imag} */,
  {32'h3cebd520, 32'hbd51f742} /* (22, 29, 21) {real, imag} */,
  {32'h3c8248f0, 32'h3d668e88} /* (22, 29, 20) {real, imag} */,
  {32'h3c811a5a, 32'hbdc83984} /* (22, 29, 19) {real, imag} */,
  {32'hbcc9f636, 32'h3d3b3de2} /* (22, 29, 18) {real, imag} */,
  {32'h3cbdefe4, 32'h3cf329a7} /* (22, 29, 17) {real, imag} */,
  {32'hbbf48888, 32'h00000000} /* (22, 29, 16) {real, imag} */,
  {32'h3cbdefe4, 32'hbcf329a7} /* (22, 29, 15) {real, imag} */,
  {32'hbcc9f636, 32'hbd3b3de2} /* (22, 29, 14) {real, imag} */,
  {32'h3c811a5a, 32'h3dc83984} /* (22, 29, 13) {real, imag} */,
  {32'h3c8248f0, 32'hbd668e88} /* (22, 29, 12) {real, imag} */,
  {32'h3cebd520, 32'h3d51f742} /* (22, 29, 11) {real, imag} */,
  {32'h3e0b15ac, 32'h3cdb9f74} /* (22, 29, 10) {real, imag} */,
  {32'hbd2284e2, 32'h3c3d5c16} /* (22, 29, 9) {real, imag} */,
  {32'h3d6d6d5c, 32'h3e3012c8} /* (22, 29, 8) {real, imag} */,
  {32'hbd60b0bb, 32'h3d27730a} /* (22, 29, 7) {real, imag} */,
  {32'hbd809994, 32'h3d659a61} /* (22, 29, 6) {real, imag} */,
  {32'h3e4ae450, 32'h3e5e9cdf} /* (22, 29, 5) {real, imag} */,
  {32'hbe85da77, 32'hbdc63643} /* (22, 29, 4) {real, imag} */,
  {32'hbdb68426, 32'h3d616c00} /* (22, 29, 3) {real, imag} */,
  {32'h3fc401aa, 32'h3eb2acc2} /* (22, 29, 2) {real, imag} */,
  {32'hc09db42a, 32'hbfcba777} /* (22, 29, 1) {real, imag} */,
  {32'hc0abf71c, 32'h00000000} /* (22, 29, 0) {real, imag} */,
  {32'hc0a58dc3, 32'h3faa7dc2} /* (22, 28, 31) {real, imag} */,
  {32'h3fe691e8, 32'hbeb34409} /* (22, 28, 30) {real, imag} */,
  {32'hbd1b0fcc, 32'hbde55dd0} /* (22, 28, 29) {real, imag} */,
  {32'hbe5d97aa, 32'h3e2d0bef} /* (22, 28, 28) {real, imag} */,
  {32'h3e7467eb, 32'hbe05d509} /* (22, 28, 27) {real, imag} */,
  {32'hbb4e51f0, 32'hbd8a947b} /* (22, 28, 26) {real, imag} */,
  {32'hbbb85e8c, 32'h3d87858c} /* (22, 28, 25) {real, imag} */,
  {32'h3d7fc589, 32'hbe49ca06} /* (22, 28, 24) {real, imag} */,
  {32'h3c1b8ea4, 32'h3d8ce0b4} /* (22, 28, 23) {real, imag} */,
  {32'h3c023cde, 32'hbbdff778} /* (22, 28, 22) {real, imag} */,
  {32'h3d4ee2f4, 32'h3d8df3cb} /* (22, 28, 21) {real, imag} */,
  {32'hbcb81076, 32'hbd6d24df} /* (22, 28, 20) {real, imag} */,
  {32'hbcfcd356, 32'h3cfa4876} /* (22, 28, 19) {real, imag} */,
  {32'h3c8161b6, 32'h3d1534ad} /* (22, 28, 18) {real, imag} */,
  {32'h3ca0e8ec, 32'h3cbb54ba} /* (22, 28, 17) {real, imag} */,
  {32'h3bfe0fcc, 32'h00000000} /* (22, 28, 16) {real, imag} */,
  {32'h3ca0e8ec, 32'hbcbb54ba} /* (22, 28, 15) {real, imag} */,
  {32'h3c8161b6, 32'hbd1534ad} /* (22, 28, 14) {real, imag} */,
  {32'hbcfcd356, 32'hbcfa4876} /* (22, 28, 13) {real, imag} */,
  {32'hbcb81076, 32'h3d6d24df} /* (22, 28, 12) {real, imag} */,
  {32'h3d4ee2f4, 32'hbd8df3cb} /* (22, 28, 11) {real, imag} */,
  {32'h3c023cde, 32'h3bdff778} /* (22, 28, 10) {real, imag} */,
  {32'h3c1b8ea4, 32'hbd8ce0b4} /* (22, 28, 9) {real, imag} */,
  {32'h3d7fc589, 32'h3e49ca06} /* (22, 28, 8) {real, imag} */,
  {32'hbbb85e8c, 32'hbd87858c} /* (22, 28, 7) {real, imag} */,
  {32'hbb4e51f0, 32'h3d8a947b} /* (22, 28, 6) {real, imag} */,
  {32'h3e7467eb, 32'h3e05d509} /* (22, 28, 5) {real, imag} */,
  {32'hbe5d97aa, 32'hbe2d0bef} /* (22, 28, 4) {real, imag} */,
  {32'hbd1b0fcc, 32'h3de55dd0} /* (22, 28, 3) {real, imag} */,
  {32'h3fe691e8, 32'h3eb34409} /* (22, 28, 2) {real, imag} */,
  {32'hc0a58dc3, 32'hbfaa7dc2} /* (22, 28, 1) {real, imag} */,
  {32'hc0b0a1ab, 32'h00000000} /* (22, 28, 0) {real, imag} */,
  {32'hc0a5aa94, 32'h3f750a72} /* (22, 27, 31) {real, imag} */,
  {32'h3febd140, 32'hbec66bda} /* (22, 27, 30) {real, imag} */,
  {32'h3da4d861, 32'hbc96337c} /* (22, 27, 29) {real, imag} */,
  {32'hbe59d8e7, 32'hbbe70d20} /* (22, 27, 28) {real, imag} */,
  {32'h3e344539, 32'hbe293df4} /* (22, 27, 27) {real, imag} */,
  {32'hbc888096, 32'h3d94f6ad} /* (22, 27, 26) {real, imag} */,
  {32'hbe1acee0, 32'h3d8b1f80} /* (22, 27, 25) {real, imag} */,
  {32'hbd9374f8, 32'hbd0625a0} /* (22, 27, 24) {real, imag} */,
  {32'h3c58b290, 32'hbd905754} /* (22, 27, 23) {real, imag} */,
  {32'h3db1311d, 32'h3c9ed4c8} /* (22, 27, 22) {real, imag} */,
  {32'h3d3484a8, 32'hbd6659d5} /* (22, 27, 21) {real, imag} */,
  {32'hbd91bed8, 32'hbd5d3d1c} /* (22, 27, 20) {real, imag} */,
  {32'hbcc52a36, 32'h3c0c01c8} /* (22, 27, 19) {real, imag} */,
  {32'hbd4d5d1e, 32'hbd4e7878} /* (22, 27, 18) {real, imag} */,
  {32'h3ccb7e88, 32'hbc73ca80} /* (22, 27, 17) {real, imag} */,
  {32'h3c229631, 32'h00000000} /* (22, 27, 16) {real, imag} */,
  {32'h3ccb7e88, 32'h3c73ca80} /* (22, 27, 15) {real, imag} */,
  {32'hbd4d5d1e, 32'h3d4e7878} /* (22, 27, 14) {real, imag} */,
  {32'hbcc52a36, 32'hbc0c01c8} /* (22, 27, 13) {real, imag} */,
  {32'hbd91bed8, 32'h3d5d3d1c} /* (22, 27, 12) {real, imag} */,
  {32'h3d3484a8, 32'h3d6659d5} /* (22, 27, 11) {real, imag} */,
  {32'h3db1311d, 32'hbc9ed4c8} /* (22, 27, 10) {real, imag} */,
  {32'h3c58b290, 32'h3d905754} /* (22, 27, 9) {real, imag} */,
  {32'hbd9374f8, 32'h3d0625a0} /* (22, 27, 8) {real, imag} */,
  {32'hbe1acee0, 32'hbd8b1f80} /* (22, 27, 7) {real, imag} */,
  {32'hbc888096, 32'hbd94f6ad} /* (22, 27, 6) {real, imag} */,
  {32'h3e344539, 32'h3e293df4} /* (22, 27, 5) {real, imag} */,
  {32'hbe59d8e7, 32'h3be70d20} /* (22, 27, 4) {real, imag} */,
  {32'h3da4d861, 32'h3c96337c} /* (22, 27, 3) {real, imag} */,
  {32'h3febd140, 32'h3ec66bda} /* (22, 27, 2) {real, imag} */,
  {32'hc0a5aa94, 32'hbf750a72} /* (22, 27, 1) {real, imag} */,
  {32'hc0b04050, 32'h00000000} /* (22, 27, 0) {real, imag} */,
  {32'hc09c964c, 32'h3f6ad84a} /* (22, 26, 31) {real, imag} */,
  {32'h3fe6f03a, 32'hbecf5658} /* (22, 26, 30) {real, imag} */,
  {32'hbc0fd04a, 32'hbd5daf91} /* (22, 26, 29) {real, imag} */,
  {32'hbe854caa, 32'hbbec56d8} /* (22, 26, 28) {real, imag} */,
  {32'h3e9a8b5a, 32'hbe5f8dc6} /* (22, 26, 27) {real, imag} */,
  {32'h3c87ff04, 32'h3d8efa38} /* (22, 26, 26) {real, imag} */,
  {32'hbdb10d41, 32'hbd1f6664} /* (22, 26, 25) {real, imag} */,
  {32'h3d0ebdb0, 32'hbd7a4188} /* (22, 26, 24) {real, imag} */,
  {32'h3caecaac, 32'hbccfd6ce} /* (22, 26, 23) {real, imag} */,
  {32'hbd030906, 32'h3dc317a6} /* (22, 26, 22) {real, imag} */,
  {32'hbd0f3682, 32'hbdf1e53c} /* (22, 26, 21) {real, imag} */,
  {32'h3dac5350, 32'hbd4ed240} /* (22, 26, 20) {real, imag} */,
  {32'h3d2b28d8, 32'h3c9d13b3} /* (22, 26, 19) {real, imag} */,
  {32'h3cd8e926, 32'h3cee81e8} /* (22, 26, 18) {real, imag} */,
  {32'h3c8d9736, 32'hbd013faf} /* (22, 26, 17) {real, imag} */,
  {32'hbc7e1372, 32'h00000000} /* (22, 26, 16) {real, imag} */,
  {32'h3c8d9736, 32'h3d013faf} /* (22, 26, 15) {real, imag} */,
  {32'h3cd8e926, 32'hbcee81e8} /* (22, 26, 14) {real, imag} */,
  {32'h3d2b28d8, 32'hbc9d13b3} /* (22, 26, 13) {real, imag} */,
  {32'h3dac5350, 32'h3d4ed240} /* (22, 26, 12) {real, imag} */,
  {32'hbd0f3682, 32'h3df1e53c} /* (22, 26, 11) {real, imag} */,
  {32'hbd030906, 32'hbdc317a6} /* (22, 26, 10) {real, imag} */,
  {32'h3caecaac, 32'h3ccfd6ce} /* (22, 26, 9) {real, imag} */,
  {32'h3d0ebdb0, 32'h3d7a4188} /* (22, 26, 8) {real, imag} */,
  {32'hbdb10d41, 32'h3d1f6664} /* (22, 26, 7) {real, imag} */,
  {32'h3c87ff04, 32'hbd8efa38} /* (22, 26, 6) {real, imag} */,
  {32'h3e9a8b5a, 32'h3e5f8dc6} /* (22, 26, 5) {real, imag} */,
  {32'hbe854caa, 32'h3bec56d8} /* (22, 26, 4) {real, imag} */,
  {32'hbc0fd04a, 32'h3d5daf91} /* (22, 26, 3) {real, imag} */,
  {32'h3fe6f03a, 32'h3ecf5658} /* (22, 26, 2) {real, imag} */,
  {32'hc09c964c, 32'hbf6ad84a} /* (22, 26, 1) {real, imag} */,
  {32'hc0a993f6, 32'h00000000} /* (22, 26, 0) {real, imag} */,
  {32'hc092013c, 32'h3f3af51f} /* (22, 25, 31) {real, imag} */,
  {32'h3fe85ea2, 32'hbea75e27} /* (22, 25, 30) {real, imag} */,
  {32'hbe06334c, 32'hbd8bc1ca} /* (22, 25, 29) {real, imag} */,
  {32'hbe530d8f, 32'h3dc30b82} /* (22, 25, 28) {real, imag} */,
  {32'h3e816ce0, 32'hbdd6e804} /* (22, 25, 27) {real, imag} */,
  {32'h3cd61536, 32'hbc68f132} /* (22, 25, 26) {real, imag} */,
  {32'hbdb3c6ed, 32'hbd44f47e} /* (22, 25, 25) {real, imag} */,
  {32'h3da1ce93, 32'hbd82a0b4} /* (22, 25, 24) {real, imag} */,
  {32'h3d9a5438, 32'hbcdf65e8} /* (22, 25, 23) {real, imag} */,
  {32'hbad32aa0, 32'hbc5588d8} /* (22, 25, 22) {real, imag} */,
  {32'hbd09fad8, 32'hbd36e3fb} /* (22, 25, 21) {real, imag} */,
  {32'hbc66313d, 32'h3d6a5cfd} /* (22, 25, 20) {real, imag} */,
  {32'h3d3e1aae, 32'h3b9dd1f8} /* (22, 25, 19) {real, imag} */,
  {32'h3deee210, 32'hbca0cae3} /* (22, 25, 18) {real, imag} */,
  {32'hbc1f08c6, 32'h3c9f0b70} /* (22, 25, 17) {real, imag} */,
  {32'hbce40055, 32'h00000000} /* (22, 25, 16) {real, imag} */,
  {32'hbc1f08c6, 32'hbc9f0b70} /* (22, 25, 15) {real, imag} */,
  {32'h3deee210, 32'h3ca0cae3} /* (22, 25, 14) {real, imag} */,
  {32'h3d3e1aae, 32'hbb9dd1f8} /* (22, 25, 13) {real, imag} */,
  {32'hbc66313d, 32'hbd6a5cfd} /* (22, 25, 12) {real, imag} */,
  {32'hbd09fad8, 32'h3d36e3fb} /* (22, 25, 11) {real, imag} */,
  {32'hbad32aa0, 32'h3c5588d8} /* (22, 25, 10) {real, imag} */,
  {32'h3d9a5438, 32'h3cdf65e8} /* (22, 25, 9) {real, imag} */,
  {32'h3da1ce93, 32'h3d82a0b4} /* (22, 25, 8) {real, imag} */,
  {32'hbdb3c6ed, 32'h3d44f47e} /* (22, 25, 7) {real, imag} */,
  {32'h3cd61536, 32'h3c68f132} /* (22, 25, 6) {real, imag} */,
  {32'h3e816ce0, 32'h3dd6e804} /* (22, 25, 5) {real, imag} */,
  {32'hbe530d8f, 32'hbdc30b82} /* (22, 25, 4) {real, imag} */,
  {32'hbe06334c, 32'h3d8bc1ca} /* (22, 25, 3) {real, imag} */,
  {32'h3fe85ea2, 32'h3ea75e27} /* (22, 25, 2) {real, imag} */,
  {32'hc092013c, 32'hbf3af51f} /* (22, 25, 1) {real, imag} */,
  {32'hc09bd282, 32'h00000000} /* (22, 25, 0) {real, imag} */,
  {32'hc0848d57, 32'h3f0c892a} /* (22, 24, 31) {real, imag} */,
  {32'h3fdd1d48, 32'hbe428386} /* (22, 24, 30) {real, imag} */,
  {32'hbdf992da, 32'h3d8ca6b5} /* (22, 24, 29) {real, imag} */,
  {32'hbd2e04c8, 32'h3e264515} /* (22, 24, 28) {real, imag} */,
  {32'h3e501d60, 32'hbe00e333} /* (22, 24, 27) {real, imag} */,
  {32'h3d3f7984, 32'hbd0c71c7} /* (22, 24, 26) {real, imag} */,
  {32'h3d3bc214, 32'h3dbbdd4e} /* (22, 24, 25) {real, imag} */,
  {32'h3d8bacf6, 32'hbd3ae646} /* (22, 24, 24) {real, imag} */,
  {32'hbd15830e, 32'h3d2b2d44} /* (22, 24, 23) {real, imag} */,
  {32'h3d496623, 32'hbc77631c} /* (22, 24, 22) {real, imag} */,
  {32'h3da13a3a, 32'h3ca92c68} /* (22, 24, 21) {real, imag} */,
  {32'hbd94ac79, 32'hbd815b64} /* (22, 24, 20) {real, imag} */,
  {32'hbdffc44b, 32'hbd585584} /* (22, 24, 19) {real, imag} */,
  {32'hbba4a69c, 32'h3c9833e3} /* (22, 24, 18) {real, imag} */,
  {32'h3d36a799, 32'h3da677e2} /* (22, 24, 17) {real, imag} */,
  {32'hbdb387b2, 32'h00000000} /* (22, 24, 16) {real, imag} */,
  {32'h3d36a799, 32'hbda677e2} /* (22, 24, 15) {real, imag} */,
  {32'hbba4a69c, 32'hbc9833e3} /* (22, 24, 14) {real, imag} */,
  {32'hbdffc44b, 32'h3d585584} /* (22, 24, 13) {real, imag} */,
  {32'hbd94ac79, 32'h3d815b64} /* (22, 24, 12) {real, imag} */,
  {32'h3da13a3a, 32'hbca92c68} /* (22, 24, 11) {real, imag} */,
  {32'h3d496623, 32'h3c77631c} /* (22, 24, 10) {real, imag} */,
  {32'hbd15830e, 32'hbd2b2d44} /* (22, 24, 9) {real, imag} */,
  {32'h3d8bacf6, 32'h3d3ae646} /* (22, 24, 8) {real, imag} */,
  {32'h3d3bc214, 32'hbdbbdd4e} /* (22, 24, 7) {real, imag} */,
  {32'h3d3f7984, 32'h3d0c71c7} /* (22, 24, 6) {real, imag} */,
  {32'h3e501d60, 32'h3e00e333} /* (22, 24, 5) {real, imag} */,
  {32'hbd2e04c8, 32'hbe264515} /* (22, 24, 4) {real, imag} */,
  {32'hbdf992da, 32'hbd8ca6b5} /* (22, 24, 3) {real, imag} */,
  {32'h3fdd1d48, 32'h3e428386} /* (22, 24, 2) {real, imag} */,
  {32'hc0848d57, 32'hbf0c892a} /* (22, 24, 1) {real, imag} */,
  {32'hc0838923, 32'h00000000} /* (22, 24, 0) {real, imag} */,
  {32'hc05ac0c8, 32'h3ecf228a} /* (22, 23, 31) {real, imag} */,
  {32'h3fa6e68d, 32'hbe966fd9} /* (22, 23, 30) {real, imag} */,
  {32'h3d1dae5f, 32'hbd038af2} /* (22, 23, 29) {real, imag} */,
  {32'hbda6284e, 32'h3e29972b} /* (22, 23, 28) {real, imag} */,
  {32'h3e8065dc, 32'hbda2ccc6} /* (22, 23, 27) {real, imag} */,
  {32'h3cfc17ae, 32'hbe0c4a24} /* (22, 23, 26) {real, imag} */,
  {32'h3c98c467, 32'h3d7a2e46} /* (22, 23, 25) {real, imag} */,
  {32'h3d5b1c22, 32'h3d7d802c} /* (22, 23, 24) {real, imag} */,
  {32'hbd3b0847, 32'hbd34ad73} /* (22, 23, 23) {real, imag} */,
  {32'hbd3204c9, 32'hbd7f9fd0} /* (22, 23, 22) {real, imag} */,
  {32'hbb5c8f28, 32'h3d02dfdf} /* (22, 23, 21) {real, imag} */,
  {32'h3caab9b4, 32'h3c7b61ec} /* (22, 23, 20) {real, imag} */,
  {32'hbd88ea0f, 32'hbd8da21c} /* (22, 23, 19) {real, imag} */,
  {32'hbd292720, 32'h3c1f2a74} /* (22, 23, 18) {real, imag} */,
  {32'h3c53f5aa, 32'hbcb85596} /* (22, 23, 17) {real, imag} */,
  {32'h3d7ff021, 32'h00000000} /* (22, 23, 16) {real, imag} */,
  {32'h3c53f5aa, 32'h3cb85596} /* (22, 23, 15) {real, imag} */,
  {32'hbd292720, 32'hbc1f2a74} /* (22, 23, 14) {real, imag} */,
  {32'hbd88ea0f, 32'h3d8da21c} /* (22, 23, 13) {real, imag} */,
  {32'h3caab9b4, 32'hbc7b61ec} /* (22, 23, 12) {real, imag} */,
  {32'hbb5c8f28, 32'hbd02dfdf} /* (22, 23, 11) {real, imag} */,
  {32'hbd3204c9, 32'h3d7f9fd0} /* (22, 23, 10) {real, imag} */,
  {32'hbd3b0847, 32'h3d34ad73} /* (22, 23, 9) {real, imag} */,
  {32'h3d5b1c22, 32'hbd7d802c} /* (22, 23, 8) {real, imag} */,
  {32'h3c98c467, 32'hbd7a2e46} /* (22, 23, 7) {real, imag} */,
  {32'h3cfc17ae, 32'h3e0c4a24} /* (22, 23, 6) {real, imag} */,
  {32'h3e8065dc, 32'h3da2ccc6} /* (22, 23, 5) {real, imag} */,
  {32'hbda6284e, 32'hbe29972b} /* (22, 23, 4) {real, imag} */,
  {32'h3d1dae5f, 32'h3d038af2} /* (22, 23, 3) {real, imag} */,
  {32'h3fa6e68d, 32'h3e966fd9} /* (22, 23, 2) {real, imag} */,
  {32'hc05ac0c8, 32'hbecf228a} /* (22, 23, 1) {real, imag} */,
  {32'hc05e7834, 32'h00000000} /* (22, 23, 0) {real, imag} */,
  {32'hc0177fbf, 32'h3e8eacca} /* (22, 22, 31) {real, imag} */,
  {32'h3f5734c4, 32'hbe50bd50} /* (22, 22, 30) {real, imag} */,
  {32'h3c97b3de, 32'h3d8e6952} /* (22, 22, 29) {real, imag} */,
  {32'hbe0195f7, 32'h3e374e45} /* (22, 22, 28) {real, imag} */,
  {32'h3e5019b9, 32'hbdca67ae} /* (22, 22, 27) {real, imag} */,
  {32'hbc18fea9, 32'hbda418b2} /* (22, 22, 26) {real, imag} */,
  {32'hbdae1bcc, 32'hbd0ed82e} /* (22, 22, 25) {real, imag} */,
  {32'h3da50014, 32'hbd53c684} /* (22, 22, 24) {real, imag} */,
  {32'h3cb423d0, 32'h3c210f62} /* (22, 22, 23) {real, imag} */,
  {32'hbd40141d, 32'h3ca1727b} /* (22, 22, 22) {real, imag} */,
  {32'h3c7fab36, 32'hbdafb028} /* (22, 22, 21) {real, imag} */,
  {32'h3cb20219, 32'hbdbc7a6b} /* (22, 22, 20) {real, imag} */,
  {32'h3cc7db74, 32'hbc91101b} /* (22, 22, 19) {real, imag} */,
  {32'hbcd73348, 32'hbd7b6f85} /* (22, 22, 18) {real, imag} */,
  {32'hbca371d0, 32'h3c9e9491} /* (22, 22, 17) {real, imag} */,
  {32'h3d796f0b, 32'h00000000} /* (22, 22, 16) {real, imag} */,
  {32'hbca371d0, 32'hbc9e9491} /* (22, 22, 15) {real, imag} */,
  {32'hbcd73348, 32'h3d7b6f85} /* (22, 22, 14) {real, imag} */,
  {32'h3cc7db74, 32'h3c91101b} /* (22, 22, 13) {real, imag} */,
  {32'h3cb20219, 32'h3dbc7a6b} /* (22, 22, 12) {real, imag} */,
  {32'h3c7fab36, 32'h3dafb028} /* (22, 22, 11) {real, imag} */,
  {32'hbd40141d, 32'hbca1727b} /* (22, 22, 10) {real, imag} */,
  {32'h3cb423d0, 32'hbc210f62} /* (22, 22, 9) {real, imag} */,
  {32'h3da50014, 32'h3d53c684} /* (22, 22, 8) {real, imag} */,
  {32'hbdae1bcc, 32'h3d0ed82e} /* (22, 22, 7) {real, imag} */,
  {32'hbc18fea9, 32'h3da418b2} /* (22, 22, 6) {real, imag} */,
  {32'h3e5019b9, 32'h3dca67ae} /* (22, 22, 5) {real, imag} */,
  {32'hbe0195f7, 32'hbe374e45} /* (22, 22, 4) {real, imag} */,
  {32'h3c97b3de, 32'hbd8e6952} /* (22, 22, 3) {real, imag} */,
  {32'h3f5734c4, 32'h3e50bd50} /* (22, 22, 2) {real, imag} */,
  {32'hc0177fbf, 32'hbe8eacca} /* (22, 22, 1) {real, imag} */,
  {32'hc01a84e4, 32'h00000000} /* (22, 22, 0) {real, imag} */,
  {32'hbf6c99e0, 32'h3dc373e4} /* (22, 21, 31) {real, imag} */,
  {32'h3e896fd2, 32'hbe3db3ef} /* (22, 21, 30) {real, imag} */,
  {32'h3cfeee68, 32'h3e1f189d} /* (22, 21, 29) {real, imag} */,
  {32'hbe0bd2d9, 32'h3d448b41} /* (22, 21, 28) {real, imag} */,
  {32'h3e19cabf, 32'hbd9299cc} /* (22, 21, 27) {real, imag} */,
  {32'hbd764f36, 32'h3c05e1be} /* (22, 21, 26) {real, imag} */,
  {32'hbc80c700, 32'hbda84c92} /* (22, 21, 25) {real, imag} */,
  {32'h3df79728, 32'hbd7c182b} /* (22, 21, 24) {real, imag} */,
  {32'hbdd80930, 32'h3d14a110} /* (22, 21, 23) {real, imag} */,
  {32'h3d5068e8, 32'hbd993e68} /* (22, 21, 22) {real, imag} */,
  {32'h3d648517, 32'hbd4d6c45} /* (22, 21, 21) {real, imag} */,
  {32'h3c86b200, 32'h3dae0060} /* (22, 21, 20) {real, imag} */,
  {32'h3d4b35b7, 32'hbd4a81a7} /* (22, 21, 19) {real, imag} */,
  {32'hbd630931, 32'hbd10aecc} /* (22, 21, 18) {real, imag} */,
  {32'h3d0ff327, 32'h3d3bdbdb} /* (22, 21, 17) {real, imag} */,
  {32'hbc76afdb, 32'h00000000} /* (22, 21, 16) {real, imag} */,
  {32'h3d0ff327, 32'hbd3bdbdb} /* (22, 21, 15) {real, imag} */,
  {32'hbd630931, 32'h3d10aecc} /* (22, 21, 14) {real, imag} */,
  {32'h3d4b35b7, 32'h3d4a81a7} /* (22, 21, 13) {real, imag} */,
  {32'h3c86b200, 32'hbdae0060} /* (22, 21, 12) {real, imag} */,
  {32'h3d648517, 32'h3d4d6c45} /* (22, 21, 11) {real, imag} */,
  {32'h3d5068e8, 32'h3d993e68} /* (22, 21, 10) {real, imag} */,
  {32'hbdd80930, 32'hbd14a110} /* (22, 21, 9) {real, imag} */,
  {32'h3df79728, 32'h3d7c182b} /* (22, 21, 8) {real, imag} */,
  {32'hbc80c700, 32'h3da84c92} /* (22, 21, 7) {real, imag} */,
  {32'hbd764f36, 32'hbc05e1be} /* (22, 21, 6) {real, imag} */,
  {32'h3e19cabf, 32'h3d9299cc} /* (22, 21, 5) {real, imag} */,
  {32'hbe0bd2d9, 32'hbd448b41} /* (22, 21, 4) {real, imag} */,
  {32'h3cfeee68, 32'hbe1f189d} /* (22, 21, 3) {real, imag} */,
  {32'h3e896fd2, 32'h3e3db3ef} /* (22, 21, 2) {real, imag} */,
  {32'hbf6c99e0, 32'hbdc373e4} /* (22, 21, 1) {real, imag} */,
  {32'hbf8e074e, 32'h00000000} /* (22, 21, 0) {real, imag} */,
  {32'h3f91d7c4, 32'hbe45bf4c} /* (22, 20, 31) {real, imag} */,
  {32'hbf0f2b29, 32'hbdca2ef5} /* (22, 20, 30) {real, imag} */,
  {32'hbd9ecd36, 32'h3df4d36e} /* (22, 20, 29) {real, imag} */,
  {32'hbc2b5ac0, 32'hbe076504} /* (22, 20, 28) {real, imag} */,
  {32'hbddc4fd4, 32'hbc312f08} /* (22, 20, 27) {real, imag} */,
  {32'hbd8e65b4, 32'hbe072828} /* (22, 20, 26) {real, imag} */,
  {32'h3c0ee10c, 32'h3d738417} /* (22, 20, 25) {real, imag} */,
  {32'hbd0cdcc3, 32'hbc2b71c8} /* (22, 20, 24) {real, imag} */,
  {32'hbd51afbe, 32'h3b67f050} /* (22, 20, 23) {real, imag} */,
  {32'hbd8fc8bf, 32'hbd1d5aca} /* (22, 20, 22) {real, imag} */,
  {32'h3ce270da, 32'h3d9c673c} /* (22, 20, 21) {real, imag} */,
  {32'h3befd668, 32'h3d255a4e} /* (22, 20, 20) {real, imag} */,
  {32'h3b114e94, 32'hbd9f45fe} /* (22, 20, 19) {real, imag} */,
  {32'h3c6b4c2c, 32'h3c93b7f0} /* (22, 20, 18) {real, imag} */,
  {32'h3b248bb0, 32'h3c5aa362} /* (22, 20, 17) {real, imag} */,
  {32'h3a8d8d20, 32'h00000000} /* (22, 20, 16) {real, imag} */,
  {32'h3b248bb0, 32'hbc5aa362} /* (22, 20, 15) {real, imag} */,
  {32'h3c6b4c2c, 32'hbc93b7f0} /* (22, 20, 14) {real, imag} */,
  {32'h3b114e94, 32'h3d9f45fe} /* (22, 20, 13) {real, imag} */,
  {32'h3befd668, 32'hbd255a4e} /* (22, 20, 12) {real, imag} */,
  {32'h3ce270da, 32'hbd9c673c} /* (22, 20, 11) {real, imag} */,
  {32'hbd8fc8bf, 32'h3d1d5aca} /* (22, 20, 10) {real, imag} */,
  {32'hbd51afbe, 32'hbb67f050} /* (22, 20, 9) {real, imag} */,
  {32'hbd0cdcc3, 32'h3c2b71c8} /* (22, 20, 8) {real, imag} */,
  {32'h3c0ee10c, 32'hbd738417} /* (22, 20, 7) {real, imag} */,
  {32'hbd8e65b4, 32'h3e072828} /* (22, 20, 6) {real, imag} */,
  {32'hbddc4fd4, 32'h3c312f08} /* (22, 20, 5) {real, imag} */,
  {32'hbc2b5ac0, 32'h3e076504} /* (22, 20, 4) {real, imag} */,
  {32'hbd9ecd36, 32'hbdf4d36e} /* (22, 20, 3) {real, imag} */,
  {32'hbf0f2b29, 32'h3dca2ef5} /* (22, 20, 2) {real, imag} */,
  {32'h3f91d7c4, 32'h3e45bf4c} /* (22, 20, 1) {real, imag} */,
  {32'h3eea602c, 32'h00000000} /* (22, 20, 0) {real, imag} */,
  {32'h401a822a, 32'hbebe9b41} /* (22, 19, 31) {real, imag} */,
  {32'hbf82e57e, 32'h3e938af9} /* (22, 19, 30) {real, imag} */,
  {32'hbe06263a, 32'h3d64a838} /* (22, 19, 29) {real, imag} */,
  {32'h3db82e0c, 32'hbd9aa04c} /* (22, 19, 28) {real, imag} */,
  {32'hbe3d3235, 32'h3d60f14c} /* (22, 19, 27) {real, imag} */,
  {32'h3d5f4b0d, 32'hbd37d8e5} /* (22, 19, 26) {real, imag} */,
  {32'h3e04613f, 32'h3c1c3858} /* (22, 19, 25) {real, imag} */,
  {32'hbdc26f76, 32'hbdcbddd8} /* (22, 19, 24) {real, imag} */,
  {32'h3d35c4bb, 32'hbd806069} /* (22, 19, 23) {real, imag} */,
  {32'hbc41e782, 32'h3c815699} /* (22, 19, 22) {real, imag} */,
  {32'hbc218631, 32'h3c883441} /* (22, 19, 21) {real, imag} */,
  {32'h3c901da0, 32'h3d409e0b} /* (22, 19, 20) {real, imag} */,
  {32'h3d08641d, 32'hbd199c97} /* (22, 19, 19) {real, imag} */,
  {32'hbbc7f0e8, 32'hbd3765e2} /* (22, 19, 18) {real, imag} */,
  {32'hbafb5fb8, 32'hbbf00bf4} /* (22, 19, 17) {real, imag} */,
  {32'hbd8a1ff9, 32'h00000000} /* (22, 19, 16) {real, imag} */,
  {32'hbafb5fb8, 32'h3bf00bf4} /* (22, 19, 15) {real, imag} */,
  {32'hbbc7f0e8, 32'h3d3765e2} /* (22, 19, 14) {real, imag} */,
  {32'h3d08641d, 32'h3d199c97} /* (22, 19, 13) {real, imag} */,
  {32'h3c901da0, 32'hbd409e0b} /* (22, 19, 12) {real, imag} */,
  {32'hbc218631, 32'hbc883441} /* (22, 19, 11) {real, imag} */,
  {32'hbc41e782, 32'hbc815699} /* (22, 19, 10) {real, imag} */,
  {32'h3d35c4bb, 32'h3d806069} /* (22, 19, 9) {real, imag} */,
  {32'hbdc26f76, 32'h3dcbddd8} /* (22, 19, 8) {real, imag} */,
  {32'h3e04613f, 32'hbc1c3858} /* (22, 19, 7) {real, imag} */,
  {32'h3d5f4b0d, 32'h3d37d8e5} /* (22, 19, 6) {real, imag} */,
  {32'hbe3d3235, 32'hbd60f14c} /* (22, 19, 5) {real, imag} */,
  {32'h3db82e0c, 32'h3d9aa04c} /* (22, 19, 4) {real, imag} */,
  {32'hbe06263a, 32'hbd64a838} /* (22, 19, 3) {real, imag} */,
  {32'hbf82e57e, 32'hbe938af9} /* (22, 19, 2) {real, imag} */,
  {32'h401a822a, 32'h3ebe9b41} /* (22, 19, 1) {real, imag} */,
  {32'h3fa335ac, 32'h00000000} /* (22, 19, 0) {real, imag} */,
  {32'h40588703, 32'hbed48f9a} /* (22, 18, 31) {real, imag} */,
  {32'hbf9f070b, 32'h3e9d94c8} /* (22, 18, 30) {real, imag} */,
  {32'hbd845c88, 32'hbd973c94} /* (22, 18, 29) {real, imag} */,
  {32'h3e80142c, 32'hbe07969e} /* (22, 18, 28) {real, imag} */,
  {32'hbd1029aa, 32'h3e30347c} /* (22, 18, 27) {real, imag} */,
  {32'hbdae5c5d, 32'h3d04155e} /* (22, 18, 26) {real, imag} */,
  {32'hbcc8d3d2, 32'hbd3dffee} /* (22, 18, 25) {real, imag} */,
  {32'hba376280, 32'h3d8b29d7} /* (22, 18, 24) {real, imag} */,
  {32'hbd6ad8df, 32'hbcec3521} /* (22, 18, 23) {real, imag} */,
  {32'hbcd11234, 32'h3c0eca1c} /* (22, 18, 22) {real, imag} */,
  {32'hbd581f18, 32'h3b28a1c4} /* (22, 18, 21) {real, imag} */,
  {32'hbd9132b8, 32'h3d3a4dc9} /* (22, 18, 20) {real, imag} */,
  {32'hbcce8e07, 32'hbcca9110} /* (22, 18, 19) {real, imag} */,
  {32'hbc988602, 32'h3cf08e16} /* (22, 18, 18) {real, imag} */,
  {32'h3d5c2992, 32'h3c1888d5} /* (22, 18, 17) {real, imag} */,
  {32'hbc7bd686, 32'h00000000} /* (22, 18, 16) {real, imag} */,
  {32'h3d5c2992, 32'hbc1888d5} /* (22, 18, 15) {real, imag} */,
  {32'hbc988602, 32'hbcf08e16} /* (22, 18, 14) {real, imag} */,
  {32'hbcce8e07, 32'h3cca9110} /* (22, 18, 13) {real, imag} */,
  {32'hbd9132b8, 32'hbd3a4dc9} /* (22, 18, 12) {real, imag} */,
  {32'hbd581f18, 32'hbb28a1c4} /* (22, 18, 11) {real, imag} */,
  {32'hbcd11234, 32'hbc0eca1c} /* (22, 18, 10) {real, imag} */,
  {32'hbd6ad8df, 32'h3cec3521} /* (22, 18, 9) {real, imag} */,
  {32'hba376280, 32'hbd8b29d7} /* (22, 18, 8) {real, imag} */,
  {32'hbcc8d3d2, 32'h3d3dffee} /* (22, 18, 7) {real, imag} */,
  {32'hbdae5c5d, 32'hbd04155e} /* (22, 18, 6) {real, imag} */,
  {32'hbd1029aa, 32'hbe30347c} /* (22, 18, 5) {real, imag} */,
  {32'h3e80142c, 32'h3e07969e} /* (22, 18, 4) {real, imag} */,
  {32'hbd845c88, 32'h3d973c94} /* (22, 18, 3) {real, imag} */,
  {32'hbf9f070b, 32'hbe9d94c8} /* (22, 18, 2) {real, imag} */,
  {32'h40588703, 32'h3ed48f9a} /* (22, 18, 1) {real, imag} */,
  {32'h3ff3bb48, 32'h00000000} /* (22, 18, 0) {real, imag} */,
  {32'h407e681b, 32'hbecc9794} /* (22, 17, 31) {real, imag} */,
  {32'hbfbb3a38, 32'h3ebcb830} /* (22, 17, 30) {real, imag} */,
  {32'hbc629f20, 32'h3d895059} /* (22, 17, 29) {real, imag} */,
  {32'h3ee31cd0, 32'hbe543ba0} /* (22, 17, 28) {real, imag} */,
  {32'hbe825f20, 32'h3e0ae443} /* (22, 17, 27) {real, imag} */,
  {32'hbd9f2018, 32'hbd2dea1c} /* (22, 17, 26) {real, imag} */,
  {32'h3cd13d78, 32'h3d77203e} /* (22, 17, 25) {real, imag} */,
  {32'h3d9a3f16, 32'h3ddd19e9} /* (22, 17, 24) {real, imag} */,
  {32'hbc92f442, 32'hbd2a47f3} /* (22, 17, 23) {real, imag} */,
  {32'hbb9bf602, 32'h3d9d6906} /* (22, 17, 22) {real, imag} */,
  {32'hbd0083f2, 32'hbdaeeed1} /* (22, 17, 21) {real, imag} */,
  {32'hbd5a2868, 32'h3abf0340} /* (22, 17, 20) {real, imag} */,
  {32'hbd1651ed, 32'h3b4bcaf0} /* (22, 17, 19) {real, imag} */,
  {32'hba5b1700, 32'hbdb0cea1} /* (22, 17, 18) {real, imag} */,
  {32'h3d5b257e, 32'h3c27afe6} /* (22, 17, 17) {real, imag} */,
  {32'hbc8ef04e, 32'h00000000} /* (22, 17, 16) {real, imag} */,
  {32'h3d5b257e, 32'hbc27afe6} /* (22, 17, 15) {real, imag} */,
  {32'hba5b1700, 32'h3db0cea1} /* (22, 17, 14) {real, imag} */,
  {32'hbd1651ed, 32'hbb4bcaf0} /* (22, 17, 13) {real, imag} */,
  {32'hbd5a2868, 32'hbabf0340} /* (22, 17, 12) {real, imag} */,
  {32'hbd0083f2, 32'h3daeeed1} /* (22, 17, 11) {real, imag} */,
  {32'hbb9bf602, 32'hbd9d6906} /* (22, 17, 10) {real, imag} */,
  {32'hbc92f442, 32'h3d2a47f3} /* (22, 17, 9) {real, imag} */,
  {32'h3d9a3f16, 32'hbddd19e9} /* (22, 17, 8) {real, imag} */,
  {32'h3cd13d78, 32'hbd77203e} /* (22, 17, 7) {real, imag} */,
  {32'hbd9f2018, 32'h3d2dea1c} /* (22, 17, 6) {real, imag} */,
  {32'hbe825f20, 32'hbe0ae443} /* (22, 17, 5) {real, imag} */,
  {32'h3ee31cd0, 32'h3e543ba0} /* (22, 17, 4) {real, imag} */,
  {32'hbc629f20, 32'hbd895059} /* (22, 17, 3) {real, imag} */,
  {32'hbfbb3a38, 32'hbebcb830} /* (22, 17, 2) {real, imag} */,
  {32'h407e681b, 32'h3ecc9794} /* (22, 17, 1) {real, imag} */,
  {32'h401eee1c, 32'h00000000} /* (22, 17, 0) {real, imag} */,
  {32'h4085459a, 32'hbedf07ac} /* (22, 16, 31) {real, imag} */,
  {32'hbfbf009f, 32'h3e8e3925} /* (22, 16, 30) {real, imag} */,
  {32'hbd9feb8a, 32'h3e7211a0} /* (22, 16, 29) {real, imag} */,
  {32'h3eccfc3c, 32'hbe8e6fc8} /* (22, 16, 28) {real, imag} */,
  {32'hbe848297, 32'h3d92aae2} /* (22, 16, 27) {real, imag} */,
  {32'hbd7508e4, 32'hbda42723} /* (22, 16, 26) {real, imag} */,
  {32'h3d5901bf, 32'hbd5f649a} /* (22, 16, 25) {real, imag} */,
  {32'hbd6ffaa8, 32'h3d57deec} /* (22, 16, 24) {real, imag} */,
  {32'hbd1528b6, 32'h3c4e8f50} /* (22, 16, 23) {real, imag} */,
  {32'h3dc77f0d, 32'h3c555a54} /* (22, 16, 22) {real, imag} */,
  {32'h3ca2ebd4, 32'hbd03a66d} /* (22, 16, 21) {real, imag} */,
  {32'hbd9f4127, 32'h3e21e6de} /* (22, 16, 20) {real, imag} */,
  {32'hbc9e19c4, 32'hbcfd21a0} /* (22, 16, 19) {real, imag} */,
  {32'h3b3c47d8, 32'h3d239db5} /* (22, 16, 18) {real, imag} */,
  {32'hbcb8f861, 32'hbc277320} /* (22, 16, 17) {real, imag} */,
  {32'hbd4c7e3f, 32'h00000000} /* (22, 16, 16) {real, imag} */,
  {32'hbcb8f861, 32'h3c277320} /* (22, 16, 15) {real, imag} */,
  {32'h3b3c47d8, 32'hbd239db5} /* (22, 16, 14) {real, imag} */,
  {32'hbc9e19c4, 32'h3cfd21a0} /* (22, 16, 13) {real, imag} */,
  {32'hbd9f4127, 32'hbe21e6de} /* (22, 16, 12) {real, imag} */,
  {32'h3ca2ebd4, 32'h3d03a66d} /* (22, 16, 11) {real, imag} */,
  {32'h3dc77f0d, 32'hbc555a54} /* (22, 16, 10) {real, imag} */,
  {32'hbd1528b6, 32'hbc4e8f50} /* (22, 16, 9) {real, imag} */,
  {32'hbd6ffaa8, 32'hbd57deec} /* (22, 16, 8) {real, imag} */,
  {32'h3d5901bf, 32'h3d5f649a} /* (22, 16, 7) {real, imag} */,
  {32'hbd7508e4, 32'h3da42723} /* (22, 16, 6) {real, imag} */,
  {32'hbe848297, 32'hbd92aae2} /* (22, 16, 5) {real, imag} */,
  {32'h3eccfc3c, 32'h3e8e6fc8} /* (22, 16, 4) {real, imag} */,
  {32'hbd9feb8a, 32'hbe7211a0} /* (22, 16, 3) {real, imag} */,
  {32'hbfbf009f, 32'hbe8e3925} /* (22, 16, 2) {real, imag} */,
  {32'h4085459a, 32'h3edf07ac} /* (22, 16, 1) {real, imag} */,
  {32'h402e8e02, 32'h00000000} /* (22, 16, 0) {real, imag} */,
  {32'h4085a3e2, 32'hbebc6b64} /* (22, 15, 31) {real, imag} */,
  {32'hbfb37df4, 32'h3e965eec} /* (22, 15, 30) {real, imag} */,
  {32'hbe5fdf80, 32'h3e0c902e} /* (22, 15, 29) {real, imag} */,
  {32'h3e949784, 32'hbe588df6} /* (22, 15, 28) {real, imag} */,
  {32'hbe86155e, 32'h3e237639} /* (22, 15, 27) {real, imag} */,
  {32'hbe59468c, 32'hbc92702c} /* (22, 15, 26) {real, imag} */,
  {32'h3dd48c7a, 32'hbd9af241} /* (22, 15, 25) {real, imag} */,
  {32'hbcc46bd6, 32'h3d5a84f6} /* (22, 15, 24) {real, imag} */,
  {32'h3c1d40db, 32'h3b0785b0} /* (22, 15, 23) {real, imag} */,
  {32'hbc1d0301, 32'hbc5e68d0} /* (22, 15, 22) {real, imag} */,
  {32'hbade4638, 32'h3dcaffdf} /* (22, 15, 21) {real, imag} */,
  {32'hbcf07297, 32'hbd096012} /* (22, 15, 20) {real, imag} */,
  {32'h3c27b4b5, 32'h3d924a64} /* (22, 15, 19) {real, imag} */,
  {32'hbd2f5846, 32'h3b6e3020} /* (22, 15, 18) {real, imag} */,
  {32'h38b92900, 32'h3b8e1011} /* (22, 15, 17) {real, imag} */,
  {32'h3cc69d24, 32'h00000000} /* (22, 15, 16) {real, imag} */,
  {32'h38b92900, 32'hbb8e1011} /* (22, 15, 15) {real, imag} */,
  {32'hbd2f5846, 32'hbb6e3020} /* (22, 15, 14) {real, imag} */,
  {32'h3c27b4b5, 32'hbd924a64} /* (22, 15, 13) {real, imag} */,
  {32'hbcf07297, 32'h3d096012} /* (22, 15, 12) {real, imag} */,
  {32'hbade4638, 32'hbdcaffdf} /* (22, 15, 11) {real, imag} */,
  {32'hbc1d0301, 32'h3c5e68d0} /* (22, 15, 10) {real, imag} */,
  {32'h3c1d40db, 32'hbb0785b0} /* (22, 15, 9) {real, imag} */,
  {32'hbcc46bd6, 32'hbd5a84f6} /* (22, 15, 8) {real, imag} */,
  {32'h3dd48c7a, 32'h3d9af241} /* (22, 15, 7) {real, imag} */,
  {32'hbe59468c, 32'h3c92702c} /* (22, 15, 6) {real, imag} */,
  {32'hbe86155e, 32'hbe237639} /* (22, 15, 5) {real, imag} */,
  {32'h3e949784, 32'h3e588df6} /* (22, 15, 4) {real, imag} */,
  {32'hbe5fdf80, 32'hbe0c902e} /* (22, 15, 3) {real, imag} */,
  {32'hbfb37df4, 32'hbe965eec} /* (22, 15, 2) {real, imag} */,
  {32'h4085a3e2, 32'h3ebc6b64} /* (22, 15, 1) {real, imag} */,
  {32'h40332340, 32'h00000000} /* (22, 15, 0) {real, imag} */,
  {32'h407535e5, 32'hbeb214fe} /* (22, 14, 31) {real, imag} */,
  {32'hbfbb22f3, 32'h3e7af3b4} /* (22, 14, 30) {real, imag} */,
  {32'hbd82fcce, 32'h3d4ba4ad} /* (22, 14, 29) {real, imag} */,
  {32'h3eca1be0, 32'hbe0cce7a} /* (22, 14, 28) {real, imag} */,
  {32'hbe52edf0, 32'h3dad9a28} /* (22, 14, 27) {real, imag} */,
  {32'hbdb5b4d7, 32'hbc30fe20} /* (22, 14, 26) {real, imag} */,
  {32'h3dfc3540, 32'hbd5f2742} /* (22, 14, 25) {real, imag} */,
  {32'hbdeb611f, 32'h3b8d32d0} /* (22, 14, 24) {real, imag} */,
  {32'h3d54ea1b, 32'h3db24681} /* (22, 14, 23) {real, imag} */,
  {32'h3e0a64a0, 32'h3dfbb162} /* (22, 14, 22) {real, imag} */,
  {32'hbc8e4317, 32'hbca3428e} /* (22, 14, 21) {real, imag} */,
  {32'h3c4fe964, 32'h3da80758} /* (22, 14, 20) {real, imag} */,
  {32'h3b4612b8, 32'hbd0144d7} /* (22, 14, 19) {real, imag} */,
  {32'h3d3d59fb, 32'h3d5f7fc9} /* (22, 14, 18) {real, imag} */,
  {32'h3d3a286c, 32'hbc03804f} /* (22, 14, 17) {real, imag} */,
  {32'h3d1f13ee, 32'h00000000} /* (22, 14, 16) {real, imag} */,
  {32'h3d3a286c, 32'h3c03804f} /* (22, 14, 15) {real, imag} */,
  {32'h3d3d59fb, 32'hbd5f7fc9} /* (22, 14, 14) {real, imag} */,
  {32'h3b4612b8, 32'h3d0144d7} /* (22, 14, 13) {real, imag} */,
  {32'h3c4fe964, 32'hbda80758} /* (22, 14, 12) {real, imag} */,
  {32'hbc8e4317, 32'h3ca3428e} /* (22, 14, 11) {real, imag} */,
  {32'h3e0a64a0, 32'hbdfbb162} /* (22, 14, 10) {real, imag} */,
  {32'h3d54ea1b, 32'hbdb24681} /* (22, 14, 9) {real, imag} */,
  {32'hbdeb611f, 32'hbb8d32d0} /* (22, 14, 8) {real, imag} */,
  {32'h3dfc3540, 32'h3d5f2742} /* (22, 14, 7) {real, imag} */,
  {32'hbdb5b4d7, 32'h3c30fe20} /* (22, 14, 6) {real, imag} */,
  {32'hbe52edf0, 32'hbdad9a28} /* (22, 14, 5) {real, imag} */,
  {32'h3eca1be0, 32'h3e0cce7a} /* (22, 14, 4) {real, imag} */,
  {32'hbd82fcce, 32'hbd4ba4ad} /* (22, 14, 3) {real, imag} */,
  {32'hbfbb22f3, 32'hbe7af3b4} /* (22, 14, 2) {real, imag} */,
  {32'h407535e5, 32'h3eb214fe} /* (22, 14, 1) {real, imag} */,
  {32'h40379dc4, 32'h00000000} /* (22, 14, 0) {real, imag} */,
  {32'h404f5b7c, 32'hb861e000} /* (22, 13, 31) {real, imag} */,
  {32'hbfb24bbe, 32'h3e113430} /* (22, 13, 30) {real, imag} */,
  {32'hbcd5bfce, 32'hbce30ee8} /* (22, 13, 29) {real, imag} */,
  {32'h3e9ccdaf, 32'hbe7bfd6e} /* (22, 13, 28) {real, imag} */,
  {32'hbe3f1d3f, 32'h3e641c5b} /* (22, 13, 27) {real, imag} */,
  {32'h3b1a4550, 32'hbd7816cb} /* (22, 13, 26) {real, imag} */,
  {32'h3d830034, 32'hbdec17b9} /* (22, 13, 25) {real, imag} */,
  {32'hbdcec5b8, 32'h3e22c8aa} /* (22, 13, 24) {real, imag} */,
  {32'h3d549231, 32'h3d931285} /* (22, 13, 23) {real, imag} */,
  {32'h3d198dcc, 32'hbc96586b} /* (22, 13, 22) {real, imag} */,
  {32'hbc01c7fb, 32'h3d152e54} /* (22, 13, 21) {real, imag} */,
  {32'hbd38baa6, 32'hbc92c62a} /* (22, 13, 20) {real, imag} */,
  {32'h3d99fe02, 32'h3c9ba1e2} /* (22, 13, 19) {real, imag} */,
  {32'hbc0ca0ac, 32'h3d888e0f} /* (22, 13, 18) {real, imag} */,
  {32'hbaa3c488, 32'h3d1c2f54} /* (22, 13, 17) {real, imag} */,
  {32'h3d2d8bca, 32'h00000000} /* (22, 13, 16) {real, imag} */,
  {32'hbaa3c488, 32'hbd1c2f54} /* (22, 13, 15) {real, imag} */,
  {32'hbc0ca0ac, 32'hbd888e0f} /* (22, 13, 14) {real, imag} */,
  {32'h3d99fe02, 32'hbc9ba1e2} /* (22, 13, 13) {real, imag} */,
  {32'hbd38baa6, 32'h3c92c62a} /* (22, 13, 12) {real, imag} */,
  {32'hbc01c7fb, 32'hbd152e54} /* (22, 13, 11) {real, imag} */,
  {32'h3d198dcc, 32'h3c96586b} /* (22, 13, 10) {real, imag} */,
  {32'h3d549231, 32'hbd931285} /* (22, 13, 9) {real, imag} */,
  {32'hbdcec5b8, 32'hbe22c8aa} /* (22, 13, 8) {real, imag} */,
  {32'h3d830034, 32'h3dec17b9} /* (22, 13, 7) {real, imag} */,
  {32'h3b1a4550, 32'h3d7816cb} /* (22, 13, 6) {real, imag} */,
  {32'hbe3f1d3f, 32'hbe641c5b} /* (22, 13, 5) {real, imag} */,
  {32'h3e9ccdaf, 32'h3e7bfd6e} /* (22, 13, 4) {real, imag} */,
  {32'hbcd5bfce, 32'h3ce30ee8} /* (22, 13, 3) {real, imag} */,
  {32'hbfb24bbe, 32'hbe113430} /* (22, 13, 2) {real, imag} */,
  {32'h404f5b7c, 32'h3861e000} /* (22, 13, 1) {real, imag} */,
  {32'h401e6b6e, 32'h00000000} /* (22, 13, 0) {real, imag} */,
  {32'h40174166, 32'h3e2a20fc} /* (22, 12, 31) {real, imag} */,
  {32'hbf9de9e2, 32'h3d9464c5} /* (22, 12, 30) {real, imag} */,
  {32'hbdb82142, 32'h3dcdfd56} /* (22, 12, 29) {real, imag} */,
  {32'h3e7ef67a, 32'hbe907bc6} /* (22, 12, 28) {real, imag} */,
  {32'hbe97aac2, 32'h3e29036e} /* (22, 12, 27) {real, imag} */,
  {32'h3deed624, 32'h3dc48754} /* (22, 12, 26) {real, imag} */,
  {32'h3dc30bce, 32'h3cc7f6ea} /* (22, 12, 25) {real, imag} */,
  {32'hbdb5a86e, 32'h3b269420} /* (22, 12, 24) {real, imag} */,
  {32'hbc44de50, 32'hbddefcfe} /* (22, 12, 23) {real, imag} */,
  {32'hbd5b3c23, 32'h3d40bc3c} /* (22, 12, 22) {real, imag} */,
  {32'hbd88ce3c, 32'hbd1fc3d9} /* (22, 12, 21) {real, imag} */,
  {32'hbd89676a, 32'hbdbd97b7} /* (22, 12, 20) {real, imag} */,
  {32'h3d08c0b4, 32'h3dd3846c} /* (22, 12, 19) {real, imag} */,
  {32'hbd46f879, 32'h3c2b6d9b} /* (22, 12, 18) {real, imag} */,
  {32'hbd2a7cbd, 32'h3b61bb48} /* (22, 12, 17) {real, imag} */,
  {32'hbd93d100, 32'h00000000} /* (22, 12, 16) {real, imag} */,
  {32'hbd2a7cbd, 32'hbb61bb48} /* (22, 12, 15) {real, imag} */,
  {32'hbd46f879, 32'hbc2b6d9b} /* (22, 12, 14) {real, imag} */,
  {32'h3d08c0b4, 32'hbdd3846c} /* (22, 12, 13) {real, imag} */,
  {32'hbd89676a, 32'h3dbd97b7} /* (22, 12, 12) {real, imag} */,
  {32'hbd88ce3c, 32'h3d1fc3d9} /* (22, 12, 11) {real, imag} */,
  {32'hbd5b3c23, 32'hbd40bc3c} /* (22, 12, 10) {real, imag} */,
  {32'hbc44de50, 32'h3ddefcfe} /* (22, 12, 9) {real, imag} */,
  {32'hbdb5a86e, 32'hbb269420} /* (22, 12, 8) {real, imag} */,
  {32'h3dc30bce, 32'hbcc7f6ea} /* (22, 12, 7) {real, imag} */,
  {32'h3deed624, 32'hbdc48754} /* (22, 12, 6) {real, imag} */,
  {32'hbe97aac2, 32'hbe29036e} /* (22, 12, 5) {real, imag} */,
  {32'h3e7ef67a, 32'h3e907bc6} /* (22, 12, 4) {real, imag} */,
  {32'hbdb82142, 32'hbdcdfd56} /* (22, 12, 3) {real, imag} */,
  {32'hbf9de9e2, 32'hbd9464c5} /* (22, 12, 2) {real, imag} */,
  {32'h40174166, 32'hbe2a20fc} /* (22, 12, 1) {real, imag} */,
  {32'h3fd7b7e9, 32'h00000000} /* (22, 12, 0) {real, imag} */,
  {32'h3f93a188, 32'h3ee0f843} /* (22, 11, 31) {real, imag} */,
  {32'hbf4bca6d, 32'h396e2c00} /* (22, 11, 30) {real, imag} */,
  {32'hbdbe43f8, 32'h3cb0bf08} /* (22, 11, 29) {real, imag} */,
  {32'h3ea03258, 32'hbd5b1e2d} /* (22, 11, 28) {real, imag} */,
  {32'hbe11afb7, 32'h3def338e} /* (22, 11, 27) {real, imag} */,
  {32'hbcd84e01, 32'h3d4c07aa} /* (22, 11, 26) {real, imag} */,
  {32'h3dd60a3d, 32'hbdd7ab96} /* (22, 11, 25) {real, imag} */,
  {32'hbd0e2b49, 32'hbd446b51} /* (22, 11, 24) {real, imag} */,
  {32'h3d96219e, 32'h3d80b86a} /* (22, 11, 23) {real, imag} */,
  {32'hbc6815e0, 32'h3df71efa} /* (22, 11, 22) {real, imag} */,
  {32'hbd7ea41b, 32'hbb864eb8} /* (22, 11, 21) {real, imag} */,
  {32'h3da22e0b, 32'hbdc500f4} /* (22, 11, 20) {real, imag} */,
  {32'h3ca0694e, 32'h3c5c1aec} /* (22, 11, 19) {real, imag} */,
  {32'hbd8093d8, 32'h3d843e1c} /* (22, 11, 18) {real, imag} */,
  {32'hbc3fbfb4, 32'h3c892642} /* (22, 11, 17) {real, imag} */,
  {32'h3c63b1e1, 32'h00000000} /* (22, 11, 16) {real, imag} */,
  {32'hbc3fbfb4, 32'hbc892642} /* (22, 11, 15) {real, imag} */,
  {32'hbd8093d8, 32'hbd843e1c} /* (22, 11, 14) {real, imag} */,
  {32'h3ca0694e, 32'hbc5c1aec} /* (22, 11, 13) {real, imag} */,
  {32'h3da22e0b, 32'h3dc500f4} /* (22, 11, 12) {real, imag} */,
  {32'hbd7ea41b, 32'h3b864eb8} /* (22, 11, 11) {real, imag} */,
  {32'hbc6815e0, 32'hbdf71efa} /* (22, 11, 10) {real, imag} */,
  {32'h3d96219e, 32'hbd80b86a} /* (22, 11, 9) {real, imag} */,
  {32'hbd0e2b49, 32'h3d446b51} /* (22, 11, 8) {real, imag} */,
  {32'h3dd60a3d, 32'h3dd7ab96} /* (22, 11, 7) {real, imag} */,
  {32'hbcd84e01, 32'hbd4c07aa} /* (22, 11, 6) {real, imag} */,
  {32'hbe11afb7, 32'hbdef338e} /* (22, 11, 5) {real, imag} */,
  {32'h3ea03258, 32'h3d5b1e2d} /* (22, 11, 4) {real, imag} */,
  {32'hbdbe43f8, 32'hbcb0bf08} /* (22, 11, 3) {real, imag} */,
  {32'hbf4bca6d, 32'hb96e2c00} /* (22, 11, 2) {real, imag} */,
  {32'h3f93a188, 32'hbee0f843} /* (22, 11, 1) {real, imag} */,
  {32'h3f10fdac, 32'h00000000} /* (22, 11, 0) {real, imag} */,
  {32'hbf22cd29, 32'h3f4e4ca1} /* (22, 10, 31) {real, imag} */,
  {32'h3d020f38, 32'hbe2a2f4a} /* (22, 10, 30) {real, imag} */,
  {32'hbc94993a, 32'hbd5745de} /* (22, 10, 29) {real, imag} */,
  {32'h3dc2892e, 32'h3e1c3181} /* (22, 10, 28) {real, imag} */,
  {32'h3e0c48af, 32'hba8ea1e0} /* (22, 10, 27) {real, imag} */,
  {32'h3d0199d2, 32'h3d94bd64} /* (22, 10, 26) {real, imag} */,
  {32'h3cf8d75a, 32'h3c549fda} /* (22, 10, 25) {real, imag} */,
  {32'h3d28e334, 32'hbdca73c2} /* (22, 10, 24) {real, imag} */,
  {32'hbc92ef78, 32'h3d83fe5c} /* (22, 10, 23) {real, imag} */,
  {32'h3d79d0ab, 32'h3d3bc410} /* (22, 10, 22) {real, imag} */,
  {32'hbd452bae, 32'hbda9a566} /* (22, 10, 21) {real, imag} */,
  {32'h3cf56347, 32'h3d9df69d} /* (22, 10, 20) {real, imag} */,
  {32'h3d3ddd0a, 32'h3ba9e8a4} /* (22, 10, 19) {real, imag} */,
  {32'hbd97dc7f, 32'h3ced061e} /* (22, 10, 18) {real, imag} */,
  {32'hbcecd81c, 32'h3d320b6c} /* (22, 10, 17) {real, imag} */,
  {32'h3cb5124a, 32'h00000000} /* (22, 10, 16) {real, imag} */,
  {32'hbcecd81c, 32'hbd320b6c} /* (22, 10, 15) {real, imag} */,
  {32'hbd97dc7f, 32'hbced061e} /* (22, 10, 14) {real, imag} */,
  {32'h3d3ddd0a, 32'hbba9e8a4} /* (22, 10, 13) {real, imag} */,
  {32'h3cf56347, 32'hbd9df69d} /* (22, 10, 12) {real, imag} */,
  {32'hbd452bae, 32'h3da9a566} /* (22, 10, 11) {real, imag} */,
  {32'h3d79d0ab, 32'hbd3bc410} /* (22, 10, 10) {real, imag} */,
  {32'hbc92ef78, 32'hbd83fe5c} /* (22, 10, 9) {real, imag} */,
  {32'h3d28e334, 32'h3dca73c2} /* (22, 10, 8) {real, imag} */,
  {32'h3cf8d75a, 32'hbc549fda} /* (22, 10, 7) {real, imag} */,
  {32'h3d0199d2, 32'hbd94bd64} /* (22, 10, 6) {real, imag} */,
  {32'h3e0c48af, 32'h3a8ea1e0} /* (22, 10, 5) {real, imag} */,
  {32'h3dc2892e, 32'hbe1c3181} /* (22, 10, 4) {real, imag} */,
  {32'hbc94993a, 32'h3d5745de} /* (22, 10, 3) {real, imag} */,
  {32'h3d020f38, 32'h3e2a2f4a} /* (22, 10, 2) {real, imag} */,
  {32'hbf22cd29, 32'hbf4e4ca1} /* (22, 10, 1) {real, imag} */,
  {32'hbf655a96, 32'h00000000} /* (22, 10, 0) {real, imag} */,
  {32'hc00a79b4, 32'h3f8a5f02} /* (22, 9, 31) {real, imag} */,
  {32'h3f09ec0a, 32'hbedd6491} /* (22, 9, 30) {real, imag} */,
  {32'hbd2b697d, 32'hbcf3c9a8} /* (22, 9, 29) {real, imag} */,
  {32'h3c31f444, 32'h3e0a3d75} /* (22, 9, 28) {real, imag} */,
  {32'h3e09a9d6, 32'hbe2bf506} /* (22, 9, 27) {real, imag} */,
  {32'h3d0f079b, 32'h3cef48e4} /* (22, 9, 26) {real, imag} */,
  {32'h3ad3da70, 32'h3c83aadc} /* (22, 9, 25) {real, imag} */,
  {32'h3c916e77, 32'hbc2e7772} /* (22, 9, 24) {real, imag} */,
  {32'hbd6523e3, 32'h3ccfc89a} /* (22, 9, 23) {real, imag} */,
  {32'hbd378787, 32'hbdcb04da} /* (22, 9, 22) {real, imag} */,
  {32'hbd7924b4, 32'hbdef4fb6} /* (22, 9, 21) {real, imag} */,
  {32'h3c8316f0, 32'hbdd25d62} /* (22, 9, 20) {real, imag} */,
  {32'h3c853b1f, 32'h3d11f21b} /* (22, 9, 19) {real, imag} */,
  {32'h3caef6d0, 32'hbdee20c6} /* (22, 9, 18) {real, imag} */,
  {32'h3a89d904, 32'h3c830c62} /* (22, 9, 17) {real, imag} */,
  {32'h3d4ee867, 32'h00000000} /* (22, 9, 16) {real, imag} */,
  {32'h3a89d904, 32'hbc830c62} /* (22, 9, 15) {real, imag} */,
  {32'h3caef6d0, 32'h3dee20c6} /* (22, 9, 14) {real, imag} */,
  {32'h3c853b1f, 32'hbd11f21b} /* (22, 9, 13) {real, imag} */,
  {32'h3c8316f0, 32'h3dd25d62} /* (22, 9, 12) {real, imag} */,
  {32'hbd7924b4, 32'h3def4fb6} /* (22, 9, 11) {real, imag} */,
  {32'hbd378787, 32'h3dcb04da} /* (22, 9, 10) {real, imag} */,
  {32'hbd6523e3, 32'hbccfc89a} /* (22, 9, 9) {real, imag} */,
  {32'h3c916e77, 32'h3c2e7772} /* (22, 9, 8) {real, imag} */,
  {32'h3ad3da70, 32'hbc83aadc} /* (22, 9, 7) {real, imag} */,
  {32'h3d0f079b, 32'hbcef48e4} /* (22, 9, 6) {real, imag} */,
  {32'h3e09a9d6, 32'h3e2bf506} /* (22, 9, 5) {real, imag} */,
  {32'h3c31f444, 32'hbe0a3d75} /* (22, 9, 4) {real, imag} */,
  {32'hbd2b697d, 32'h3cf3c9a8} /* (22, 9, 3) {real, imag} */,
  {32'h3f09ec0a, 32'h3edd6491} /* (22, 9, 2) {real, imag} */,
  {32'hc00a79b4, 32'hbf8a5f02} /* (22, 9, 1) {real, imag} */,
  {32'hc00f16cc, 32'h00000000} /* (22, 9, 0) {real, imag} */,
  {32'hc03c90a8, 32'h3fc0451d} /* (22, 8, 31) {real, imag} */,
  {32'h3f7b90c0, 32'hbede17eb} /* (22, 8, 30) {real, imag} */,
  {32'h3b4b5e50, 32'hbdb671df} /* (22, 8, 29) {real, imag} */,
  {32'hbe00afa6, 32'h3dc18d66} /* (22, 8, 28) {real, imag} */,
  {32'h3e5b6dec, 32'hbd28092c} /* (22, 8, 27) {real, imag} */,
  {32'h3d80a381, 32'h3c800b74} /* (22, 8, 26) {real, imag} */,
  {32'h3d8d2883, 32'hbcdd83e8} /* (22, 8, 25) {real, imag} */,
  {32'hbd12ed6a, 32'hbd3d62ca} /* (22, 8, 24) {real, imag} */,
  {32'h3e2d155e, 32'hbd0d9aa0} /* (22, 8, 23) {real, imag} */,
  {32'h3cb23d3a, 32'h3c0b7894} /* (22, 8, 22) {real, imag} */,
  {32'h3d65130b, 32'hbdce0b47} /* (22, 8, 21) {real, imag} */,
  {32'hbc5893d6, 32'h3d756c40} /* (22, 8, 20) {real, imag} */,
  {32'h3de3ff75, 32'h3ccacf65} /* (22, 8, 19) {real, imag} */,
  {32'h3d0fc338, 32'h3c75d9f2} /* (22, 8, 18) {real, imag} */,
  {32'hbd3001a7, 32'hbbeca2e0} /* (22, 8, 17) {real, imag} */,
  {32'h3bbd0d80, 32'h00000000} /* (22, 8, 16) {real, imag} */,
  {32'hbd3001a7, 32'h3beca2e0} /* (22, 8, 15) {real, imag} */,
  {32'h3d0fc338, 32'hbc75d9f2} /* (22, 8, 14) {real, imag} */,
  {32'h3de3ff75, 32'hbccacf65} /* (22, 8, 13) {real, imag} */,
  {32'hbc5893d6, 32'hbd756c40} /* (22, 8, 12) {real, imag} */,
  {32'h3d65130b, 32'h3dce0b47} /* (22, 8, 11) {real, imag} */,
  {32'h3cb23d3a, 32'hbc0b7894} /* (22, 8, 10) {real, imag} */,
  {32'h3e2d155e, 32'h3d0d9aa0} /* (22, 8, 9) {real, imag} */,
  {32'hbd12ed6a, 32'h3d3d62ca} /* (22, 8, 8) {real, imag} */,
  {32'h3d8d2883, 32'h3cdd83e8} /* (22, 8, 7) {real, imag} */,
  {32'h3d80a381, 32'hbc800b74} /* (22, 8, 6) {real, imag} */,
  {32'h3e5b6dec, 32'h3d28092c} /* (22, 8, 5) {real, imag} */,
  {32'hbe00afa6, 32'hbdc18d66} /* (22, 8, 4) {real, imag} */,
  {32'h3b4b5e50, 32'h3db671df} /* (22, 8, 3) {real, imag} */,
  {32'h3f7b90c0, 32'h3ede17eb} /* (22, 8, 2) {real, imag} */,
  {32'hc03c90a8, 32'hbfc0451d} /* (22, 8, 1) {real, imag} */,
  {32'hc04d750e, 32'h00000000} /* (22, 8, 0) {real, imag} */,
  {32'hc05e4f94, 32'h3ffa7ee8} /* (22, 7, 31) {real, imag} */,
  {32'h3f76ef49, 32'hbf0f5ad1} /* (22, 7, 30) {real, imag} */,
  {32'h3da49e49, 32'hbdf24126} /* (22, 7, 29) {real, imag} */,
  {32'hbd9b4202, 32'h3d6aa824} /* (22, 7, 28) {real, imag} */,
  {32'h3e61f3b1, 32'hbca5ce06} /* (22, 7, 27) {real, imag} */,
  {32'h3bc77848, 32'h3d0c9220} /* (22, 7, 26) {real, imag} */,
  {32'h3db1029b, 32'hbd4802f6} /* (22, 7, 25) {real, imag} */,
  {32'h3dc0651d, 32'hbde0589c} /* (22, 7, 24) {real, imag} */,
  {32'h3cf1b2da, 32'hbd4f70de} /* (22, 7, 23) {real, imag} */,
  {32'h3d7874ad, 32'h3dfc4cd1} /* (22, 7, 22) {real, imag} */,
  {32'h3d8b93e0, 32'h3cf8a262} /* (22, 7, 21) {real, imag} */,
  {32'hbd359623, 32'h3da4e6c4} /* (22, 7, 20) {real, imag} */,
  {32'hbdb4a979, 32'hbdaa1128} /* (22, 7, 19) {real, imag} */,
  {32'hbdcbe024, 32'hbd629c28} /* (22, 7, 18) {real, imag} */,
  {32'h3ca6bbd4, 32'h3c790e09} /* (22, 7, 17) {real, imag} */,
  {32'hbcb5f9cb, 32'h00000000} /* (22, 7, 16) {real, imag} */,
  {32'h3ca6bbd4, 32'hbc790e09} /* (22, 7, 15) {real, imag} */,
  {32'hbdcbe024, 32'h3d629c28} /* (22, 7, 14) {real, imag} */,
  {32'hbdb4a979, 32'h3daa1128} /* (22, 7, 13) {real, imag} */,
  {32'hbd359623, 32'hbda4e6c4} /* (22, 7, 12) {real, imag} */,
  {32'h3d8b93e0, 32'hbcf8a262} /* (22, 7, 11) {real, imag} */,
  {32'h3d7874ad, 32'hbdfc4cd1} /* (22, 7, 10) {real, imag} */,
  {32'h3cf1b2da, 32'h3d4f70de} /* (22, 7, 9) {real, imag} */,
  {32'h3dc0651d, 32'h3de0589c} /* (22, 7, 8) {real, imag} */,
  {32'h3db1029b, 32'h3d4802f6} /* (22, 7, 7) {real, imag} */,
  {32'h3bc77848, 32'hbd0c9220} /* (22, 7, 6) {real, imag} */,
  {32'h3e61f3b1, 32'h3ca5ce06} /* (22, 7, 5) {real, imag} */,
  {32'hbd9b4202, 32'hbd6aa824} /* (22, 7, 4) {real, imag} */,
  {32'h3da49e49, 32'h3df24126} /* (22, 7, 3) {real, imag} */,
  {32'h3f76ef49, 32'h3f0f5ad1} /* (22, 7, 2) {real, imag} */,
  {32'hc05e4f94, 32'hbffa7ee8} /* (22, 7, 1) {real, imag} */,
  {32'hc07dfa91, 32'h00000000} /* (22, 7, 0) {real, imag} */,
  {32'hc0690f08, 32'h401c4712} /* (22, 6, 31) {real, imag} */,
  {32'h3f476cb4, 32'hbf184eec} /* (22, 6, 30) {real, imag} */,
  {32'h3d8e0fea, 32'hbc55220c} /* (22, 6, 29) {real, imag} */,
  {32'hbd437b90, 32'hbda04fae} /* (22, 6, 28) {real, imag} */,
  {32'h3e041655, 32'hbd9f6f6f} /* (22, 6, 27) {real, imag} */,
  {32'hbd2f0106, 32'hbcfbb888} /* (22, 6, 26) {real, imag} */,
  {32'hbd8fb56f, 32'h3d2c2084} /* (22, 6, 25) {real, imag} */,
  {32'h3db3236c, 32'hbd8a06ac} /* (22, 6, 24) {real, imag} */,
  {32'hbd4f3d2e, 32'h3c9f19ec} /* (22, 6, 23) {real, imag} */,
  {32'hbda81e30, 32'h3d1f150c} /* (22, 6, 22) {real, imag} */,
  {32'h3a1a51c0, 32'h3b2c2fb0} /* (22, 6, 21) {real, imag} */,
  {32'hbd1bd3c8, 32'hbdb9742a} /* (22, 6, 20) {real, imag} */,
  {32'h3dd697ce, 32'hbce7fc09} /* (22, 6, 19) {real, imag} */,
  {32'hbaae0818, 32'hbb84ee60} /* (22, 6, 18) {real, imag} */,
  {32'h3a495b90, 32'h3d8006e0} /* (22, 6, 17) {real, imag} */,
  {32'hbd2c40c6, 32'h00000000} /* (22, 6, 16) {real, imag} */,
  {32'h3a495b90, 32'hbd8006e0} /* (22, 6, 15) {real, imag} */,
  {32'hbaae0818, 32'h3b84ee60} /* (22, 6, 14) {real, imag} */,
  {32'h3dd697ce, 32'h3ce7fc09} /* (22, 6, 13) {real, imag} */,
  {32'hbd1bd3c8, 32'h3db9742a} /* (22, 6, 12) {real, imag} */,
  {32'h3a1a51c0, 32'hbb2c2fb0} /* (22, 6, 11) {real, imag} */,
  {32'hbda81e30, 32'hbd1f150c} /* (22, 6, 10) {real, imag} */,
  {32'hbd4f3d2e, 32'hbc9f19ec} /* (22, 6, 9) {real, imag} */,
  {32'h3db3236c, 32'h3d8a06ac} /* (22, 6, 8) {real, imag} */,
  {32'hbd8fb56f, 32'hbd2c2084} /* (22, 6, 7) {real, imag} */,
  {32'hbd2f0106, 32'h3cfbb888} /* (22, 6, 6) {real, imag} */,
  {32'h3e041655, 32'h3d9f6f6f} /* (22, 6, 5) {real, imag} */,
  {32'hbd437b90, 32'h3da04fae} /* (22, 6, 4) {real, imag} */,
  {32'h3d8e0fea, 32'h3c55220c} /* (22, 6, 3) {real, imag} */,
  {32'h3f476cb4, 32'h3f184eec} /* (22, 6, 2) {real, imag} */,
  {32'hc0690f08, 32'hc01c4712} /* (22, 6, 1) {real, imag} */,
  {32'hc08a9bea, 32'h00000000} /* (22, 6, 0) {real, imag} */,
  {32'hc0641607, 32'h404ff2a2} /* (22, 5, 31) {real, imag} */,
  {32'h3e50889c, 32'hbf3c7ab3} /* (22, 5, 30) {real, imag} */,
  {32'h3e20625e, 32'hbdb1f501} /* (22, 5, 29) {real, imag} */,
  {32'h3d20f304, 32'hbe3f83c5} /* (22, 5, 28) {real, imag} */,
  {32'h3e73b8a1, 32'h3c9e11d4} /* (22, 5, 27) {real, imag} */,
  {32'h3d90c0e0, 32'h3d388e74} /* (22, 5, 26) {real, imag} */,
  {32'h3d9cc758, 32'h3defc950} /* (22, 5, 25) {real, imag} */,
  {32'hbdaaeb34, 32'hbd9960ba} /* (22, 5, 24) {real, imag} */,
  {32'h3e1250ee, 32'h3c35b392} /* (22, 5, 23) {real, imag} */,
  {32'h3c895784, 32'h3df3ba38} /* (22, 5, 22) {real, imag} */,
  {32'h3a8e3dc0, 32'hbd0c5b53} /* (22, 5, 21) {real, imag} */,
  {32'hbd3ba7d2, 32'hbd80954f} /* (22, 5, 20) {real, imag} */,
  {32'hbd0277f7, 32'hbca0965c} /* (22, 5, 19) {real, imag} */,
  {32'hbdb7f611, 32'hbcf69c17} /* (22, 5, 18) {real, imag} */,
  {32'hbc437558, 32'hbdb1b1bc} /* (22, 5, 17) {real, imag} */,
  {32'h3c502ccd, 32'h00000000} /* (22, 5, 16) {real, imag} */,
  {32'hbc437558, 32'h3db1b1bc} /* (22, 5, 15) {real, imag} */,
  {32'hbdb7f611, 32'h3cf69c17} /* (22, 5, 14) {real, imag} */,
  {32'hbd0277f7, 32'h3ca0965c} /* (22, 5, 13) {real, imag} */,
  {32'hbd3ba7d2, 32'h3d80954f} /* (22, 5, 12) {real, imag} */,
  {32'h3a8e3dc0, 32'h3d0c5b53} /* (22, 5, 11) {real, imag} */,
  {32'h3c895784, 32'hbdf3ba38} /* (22, 5, 10) {real, imag} */,
  {32'h3e1250ee, 32'hbc35b392} /* (22, 5, 9) {real, imag} */,
  {32'hbdaaeb34, 32'h3d9960ba} /* (22, 5, 8) {real, imag} */,
  {32'h3d9cc758, 32'hbdefc950} /* (22, 5, 7) {real, imag} */,
  {32'h3d90c0e0, 32'hbd388e74} /* (22, 5, 6) {real, imag} */,
  {32'h3e73b8a1, 32'hbc9e11d4} /* (22, 5, 5) {real, imag} */,
  {32'h3d20f304, 32'h3e3f83c5} /* (22, 5, 4) {real, imag} */,
  {32'h3e20625e, 32'h3db1f501} /* (22, 5, 3) {real, imag} */,
  {32'h3e50889c, 32'h3f3c7ab3} /* (22, 5, 2) {real, imag} */,
  {32'hc0641607, 32'hc04ff2a2} /* (22, 5, 1) {real, imag} */,
  {32'hc09abef4, 32'h00000000} /* (22, 5, 0) {real, imag} */,
  {32'hc05f1e4f, 32'h4073dcd3} /* (22, 4, 31) {real, imag} */,
  {32'hbe54e340, 32'hbf55939c} /* (22, 4, 30) {real, imag} */,
  {32'h3e692c63, 32'hbe09acce} /* (22, 4, 29) {real, imag} */,
  {32'h3e4732d8, 32'hbe7193f9} /* (22, 4, 28) {real, imag} */,
  {32'h3e198a63, 32'h3df78426} /* (22, 4, 27) {real, imag} */,
  {32'hbd18841d, 32'h3c95afd0} /* (22, 4, 26) {real, imag} */,
  {32'h3d357918, 32'h3bd175e0} /* (22, 4, 25) {real, imag} */,
  {32'hbd898764, 32'h3c93b1e4} /* (22, 4, 24) {real, imag} */,
  {32'h3d768cdd, 32'h3c95d0a6} /* (22, 4, 23) {real, imag} */,
  {32'hbd585294, 32'hbd670a99} /* (22, 4, 22) {real, imag} */,
  {32'h3d8a7e1d, 32'hbd95ee79} /* (22, 4, 21) {real, imag} */,
  {32'hbd1ba5e9, 32'h3cec7026} /* (22, 4, 20) {real, imag} */,
  {32'hbd73481d, 32'h3d7595bb} /* (22, 4, 19) {real, imag} */,
  {32'hbd31713d, 32'hbc99e9b4} /* (22, 4, 18) {real, imag} */,
  {32'h3d3025be, 32'hbac12a80} /* (22, 4, 17) {real, imag} */,
  {32'h3b9a08bc, 32'h00000000} /* (22, 4, 16) {real, imag} */,
  {32'h3d3025be, 32'h3ac12a80} /* (22, 4, 15) {real, imag} */,
  {32'hbd31713d, 32'h3c99e9b4} /* (22, 4, 14) {real, imag} */,
  {32'hbd73481d, 32'hbd7595bb} /* (22, 4, 13) {real, imag} */,
  {32'hbd1ba5e9, 32'hbcec7026} /* (22, 4, 12) {real, imag} */,
  {32'h3d8a7e1d, 32'h3d95ee79} /* (22, 4, 11) {real, imag} */,
  {32'hbd585294, 32'h3d670a99} /* (22, 4, 10) {real, imag} */,
  {32'h3d768cdd, 32'hbc95d0a6} /* (22, 4, 9) {real, imag} */,
  {32'hbd898764, 32'hbc93b1e4} /* (22, 4, 8) {real, imag} */,
  {32'h3d357918, 32'hbbd175e0} /* (22, 4, 7) {real, imag} */,
  {32'hbd18841d, 32'hbc95afd0} /* (22, 4, 6) {real, imag} */,
  {32'h3e198a63, 32'hbdf78426} /* (22, 4, 5) {real, imag} */,
  {32'h3e4732d8, 32'h3e7193f9} /* (22, 4, 4) {real, imag} */,
  {32'h3e692c63, 32'h3e09acce} /* (22, 4, 3) {real, imag} */,
  {32'hbe54e340, 32'h3f55939c} /* (22, 4, 2) {real, imag} */,
  {32'hc05f1e4f, 32'hc073dcd3} /* (22, 4, 1) {real, imag} */,
  {32'hc0a1a571, 32'h00000000} /* (22, 4, 0) {real, imag} */,
  {32'hc063230c, 32'h407d6a7c} /* (22, 3, 31) {real, imag} */,
  {32'hbe8b77ca, 32'hbf80e984} /* (22, 3, 30) {real, imag} */,
  {32'h3e71119b, 32'hbe60de58} /* (22, 3, 29) {real, imag} */,
  {32'h3e1c62e2, 32'hbead30fd} /* (22, 3, 28) {real, imag} */,
  {32'h3e9c4fc4, 32'h3ccc30d8} /* (22, 3, 27) {real, imag} */,
  {32'hbc921fec, 32'hbd54e9c7} /* (22, 3, 26) {real, imag} */,
  {32'h3d56bf5f, 32'h3e0af6fa} /* (22, 3, 25) {real, imag} */,
  {32'hbdae6820, 32'hbd087a4a} /* (22, 3, 24) {real, imag} */,
  {32'h3dd13f5f, 32'hbd0dd242} /* (22, 3, 23) {real, imag} */,
  {32'h3d8c982c, 32'hbc48e0f3} /* (22, 3, 22) {real, imag} */,
  {32'hbcdfb67c, 32'h3d0c29da} /* (22, 3, 21) {real, imag} */,
  {32'h3dab828f, 32'h3cd3d21d} /* (22, 3, 20) {real, imag} */,
  {32'hbd98c91a, 32'hbd8d8388} /* (22, 3, 19) {real, imag} */,
  {32'hbdf75136, 32'h3d28d112} /* (22, 3, 18) {real, imag} */,
  {32'hbcd2f124, 32'h3d4ae9a0} /* (22, 3, 17) {real, imag} */,
  {32'h3da1c122, 32'h00000000} /* (22, 3, 16) {real, imag} */,
  {32'hbcd2f124, 32'hbd4ae9a0} /* (22, 3, 15) {real, imag} */,
  {32'hbdf75136, 32'hbd28d112} /* (22, 3, 14) {real, imag} */,
  {32'hbd98c91a, 32'h3d8d8388} /* (22, 3, 13) {real, imag} */,
  {32'h3dab828f, 32'hbcd3d21d} /* (22, 3, 12) {real, imag} */,
  {32'hbcdfb67c, 32'hbd0c29da} /* (22, 3, 11) {real, imag} */,
  {32'h3d8c982c, 32'h3c48e0f3} /* (22, 3, 10) {real, imag} */,
  {32'h3dd13f5f, 32'h3d0dd242} /* (22, 3, 9) {real, imag} */,
  {32'hbdae6820, 32'h3d087a4a} /* (22, 3, 8) {real, imag} */,
  {32'h3d56bf5f, 32'hbe0af6fa} /* (22, 3, 7) {real, imag} */,
  {32'hbc921fec, 32'h3d54e9c7} /* (22, 3, 6) {real, imag} */,
  {32'h3e9c4fc4, 32'hbccc30d8} /* (22, 3, 5) {real, imag} */,
  {32'h3e1c62e2, 32'h3ead30fd} /* (22, 3, 4) {real, imag} */,
  {32'h3e71119b, 32'h3e60de58} /* (22, 3, 3) {real, imag} */,
  {32'hbe8b77ca, 32'h3f80e984} /* (22, 3, 2) {real, imag} */,
  {32'hc063230c, 32'hc07d6a7c} /* (22, 3, 1) {real, imag} */,
  {32'hc0ad2dd0, 32'h00000000} /* (22, 3, 0) {real, imag} */,
  {32'hc05e5e92, 32'h40735cd5} /* (22, 2, 31) {real, imag} */,
  {32'hbeab9b2c, 32'hbf601c42} /* (22, 2, 30) {real, imag} */,
  {32'h3d8fb063, 32'hbdc5ffea} /* (22, 2, 29) {real, imag} */,
  {32'h3da2327c, 32'hbe922c77} /* (22, 2, 28) {real, imag} */,
  {32'h3e876cdd, 32'h3ddabcc9} /* (22, 2, 27) {real, imag} */,
  {32'h3d6a5c8d, 32'hbdcef329} /* (22, 2, 26) {real, imag} */,
  {32'h3dda964c, 32'hbd885e51} /* (22, 2, 25) {real, imag} */,
  {32'h3d11654c, 32'hbd6ceb3e} /* (22, 2, 24) {real, imag} */,
  {32'h3e06ab7b, 32'hbd4ddad2} /* (22, 2, 23) {real, imag} */,
  {32'hbb93d148, 32'hbd858c76} /* (22, 2, 22) {real, imag} */,
  {32'h3d4295aa, 32'hbd2c0174} /* (22, 2, 21) {real, imag} */,
  {32'h3d64baa7, 32'h3db06548} /* (22, 2, 20) {real, imag} */,
  {32'hbc1cb1e6, 32'hbc83dfd3} /* (22, 2, 19) {real, imag} */,
  {32'h3b959b94, 32'h39a10b80} /* (22, 2, 18) {real, imag} */,
  {32'hbc2b7dc6, 32'h3d295231} /* (22, 2, 17) {real, imag} */,
  {32'h3da9de29, 32'h00000000} /* (22, 2, 16) {real, imag} */,
  {32'hbc2b7dc6, 32'hbd295231} /* (22, 2, 15) {real, imag} */,
  {32'h3b959b94, 32'hb9a10b80} /* (22, 2, 14) {real, imag} */,
  {32'hbc1cb1e6, 32'h3c83dfd3} /* (22, 2, 13) {real, imag} */,
  {32'h3d64baa7, 32'hbdb06548} /* (22, 2, 12) {real, imag} */,
  {32'h3d4295aa, 32'h3d2c0174} /* (22, 2, 11) {real, imag} */,
  {32'hbb93d148, 32'h3d858c76} /* (22, 2, 10) {real, imag} */,
  {32'h3e06ab7b, 32'h3d4ddad2} /* (22, 2, 9) {real, imag} */,
  {32'h3d11654c, 32'h3d6ceb3e} /* (22, 2, 8) {real, imag} */,
  {32'h3dda964c, 32'h3d885e51} /* (22, 2, 7) {real, imag} */,
  {32'h3d6a5c8d, 32'h3dcef329} /* (22, 2, 6) {real, imag} */,
  {32'h3e876cdd, 32'hbddabcc9} /* (22, 2, 5) {real, imag} */,
  {32'h3da2327c, 32'h3e922c77} /* (22, 2, 4) {real, imag} */,
  {32'h3d8fb063, 32'h3dc5ffea} /* (22, 2, 3) {real, imag} */,
  {32'hbeab9b2c, 32'h3f601c42} /* (22, 2, 2) {real, imag} */,
  {32'hc05e5e92, 32'hc0735cd5} /* (22, 2, 1) {real, imag} */,
  {32'hc0ae534f, 32'h00000000} /* (22, 2, 0) {real, imag} */,
  {32'hc0578861, 32'h4064a5ac} /* (22, 1, 31) {real, imag} */,
  {32'hbe0d3774, 32'hbf55ec82} /* (22, 1, 30) {real, imag} */,
  {32'h3e1abde9, 32'hbe01e0da} /* (22, 1, 29) {real, imag} */,
  {32'h3c721e50, 32'hbeb6c2ae} /* (22, 1, 28) {real, imag} */,
  {32'h3e45f4b9, 32'h3e1b846f} /* (22, 1, 27) {real, imag} */,
  {32'hbd5d97bc, 32'hbd203372} /* (22, 1, 26) {real, imag} */,
  {32'h3de10d4a, 32'h3d27f504} /* (22, 1, 25) {real, imag} */,
  {32'h3c505c9a, 32'hbd42a7f2} /* (22, 1, 24) {real, imag} */,
  {32'h3c8b5d4e, 32'hbc55949d} /* (22, 1, 23) {real, imag} */,
  {32'hbda4b6a0, 32'hbc63ca42} /* (22, 1, 22) {real, imag} */,
  {32'h3c240409, 32'h3d54fa5c} /* (22, 1, 21) {real, imag} */,
  {32'h3d91a950, 32'hbb88e200} /* (22, 1, 20) {real, imag} */,
  {32'hbc92821e, 32'h3cb993a7} /* (22, 1, 19) {real, imag} */,
  {32'h3ca809dc, 32'h3b5a7bb8} /* (22, 1, 18) {real, imag} */,
  {32'hbd664644, 32'h3aa11d8e} /* (22, 1, 17) {real, imag} */,
  {32'h3ba2981e, 32'h00000000} /* (22, 1, 16) {real, imag} */,
  {32'hbd664644, 32'hbaa11d8e} /* (22, 1, 15) {real, imag} */,
  {32'h3ca809dc, 32'hbb5a7bb8} /* (22, 1, 14) {real, imag} */,
  {32'hbc92821e, 32'hbcb993a7} /* (22, 1, 13) {real, imag} */,
  {32'h3d91a950, 32'h3b88e200} /* (22, 1, 12) {real, imag} */,
  {32'h3c240409, 32'hbd54fa5c} /* (22, 1, 11) {real, imag} */,
  {32'hbda4b6a0, 32'h3c63ca42} /* (22, 1, 10) {real, imag} */,
  {32'h3c8b5d4e, 32'h3c55949d} /* (22, 1, 9) {real, imag} */,
  {32'h3c505c9a, 32'h3d42a7f2} /* (22, 1, 8) {real, imag} */,
  {32'h3de10d4a, 32'hbd27f504} /* (22, 1, 7) {real, imag} */,
  {32'hbd5d97bc, 32'h3d203372} /* (22, 1, 6) {real, imag} */,
  {32'h3e45f4b9, 32'hbe1b846f} /* (22, 1, 5) {real, imag} */,
  {32'h3c721e50, 32'h3eb6c2ae} /* (22, 1, 4) {real, imag} */,
  {32'h3e1abde9, 32'h3e01e0da} /* (22, 1, 3) {real, imag} */,
  {32'hbe0d3774, 32'h3f55ec82} /* (22, 1, 2) {real, imag} */,
  {32'hc0578861, 32'hc064a5ac} /* (22, 1, 1) {real, imag} */,
  {32'hc0aaf37d, 32'h00000000} /* (22, 1, 0) {real, imag} */,
  {32'hc063ca4d, 32'h403b8352} /* (22, 0, 31) {real, imag} */,
  {32'h3e67a458, 32'hbf1e11ca} /* (22, 0, 30) {real, imag} */,
  {32'h3e235c11, 32'hbce33c44} /* (22, 0, 29) {real, imag} */,
  {32'hbd60803c, 32'hbe6e554d} /* (22, 0, 28) {real, imag} */,
  {32'h3c7f1aa0, 32'hbccf3cc4} /* (22, 0, 27) {real, imag} */,
  {32'hbdc62a22, 32'h3c5c7758} /* (22, 0, 26) {real, imag} */,
  {32'h3d26340f, 32'h3d30ba3e} /* (22, 0, 25) {real, imag} */,
  {32'h3cdbb023, 32'hbd8d8ca3} /* (22, 0, 24) {real, imag} */,
  {32'h3d873d71, 32'hbda4a704} /* (22, 0, 23) {real, imag} */,
  {32'hbe09fc32, 32'hbda8e122} /* (22, 0, 22) {real, imag} */,
  {32'hbcf979b8, 32'h3cf439de} /* (22, 0, 21) {real, imag} */,
  {32'h3d2f6ada, 32'h3d31f776} /* (22, 0, 20) {real, imag} */,
  {32'hbd51cc98, 32'hbd7628d0} /* (22, 0, 19) {real, imag} */,
  {32'h3d3bb08e, 32'h3c46ba43} /* (22, 0, 18) {real, imag} */,
  {32'hbc04c146, 32'hbd786220} /* (22, 0, 17) {real, imag} */,
  {32'hbd5c3935, 32'h00000000} /* (22, 0, 16) {real, imag} */,
  {32'hbc04c146, 32'h3d786220} /* (22, 0, 15) {real, imag} */,
  {32'h3d3bb08e, 32'hbc46ba43} /* (22, 0, 14) {real, imag} */,
  {32'hbd51cc98, 32'h3d7628d0} /* (22, 0, 13) {real, imag} */,
  {32'h3d2f6ada, 32'hbd31f776} /* (22, 0, 12) {real, imag} */,
  {32'hbcf979b8, 32'hbcf439de} /* (22, 0, 11) {real, imag} */,
  {32'hbe09fc32, 32'h3da8e122} /* (22, 0, 10) {real, imag} */,
  {32'h3d873d71, 32'h3da4a704} /* (22, 0, 9) {real, imag} */,
  {32'h3cdbb023, 32'h3d8d8ca3} /* (22, 0, 8) {real, imag} */,
  {32'h3d26340f, 32'hbd30ba3e} /* (22, 0, 7) {real, imag} */,
  {32'hbdc62a22, 32'hbc5c7758} /* (22, 0, 6) {real, imag} */,
  {32'h3c7f1aa0, 32'h3ccf3cc4} /* (22, 0, 5) {real, imag} */,
  {32'hbd60803c, 32'h3e6e554d} /* (22, 0, 4) {real, imag} */,
  {32'h3e235c11, 32'h3ce33c44} /* (22, 0, 3) {real, imag} */,
  {32'h3e67a458, 32'h3f1e11ca} /* (22, 0, 2) {real, imag} */,
  {32'hc063ca4d, 32'hc03b8352} /* (22, 0, 1) {real, imag} */,
  {32'hc0a5510d, 32'h00000000} /* (22, 0, 0) {real, imag} */,
  {32'hc083f146, 32'h4015235c} /* (21, 31, 31) {real, imag} */,
  {32'h3f47e62b, 32'hbf040067} /* (21, 31, 30) {real, imag} */,
  {32'h3cdd09b8, 32'h3d77b55c} /* (21, 31, 29) {real, imag} */,
  {32'hbdde38ed, 32'hbd0f3da0} /* (21, 31, 28) {real, imag} */,
  {32'h3d410f80, 32'hbca538e6} /* (21, 31, 27) {real, imag} */,
  {32'h3c3d54a8, 32'hbd45a486} /* (21, 31, 26) {real, imag} */,
  {32'h3d98a9fb, 32'h3cb82382} /* (21, 31, 25) {real, imag} */,
  {32'h3d09b68a, 32'h3b074518} /* (21, 31, 24) {real, imag} */,
  {32'hb7a49000, 32'h3d45ba37} /* (21, 31, 23) {real, imag} */,
  {32'h3c5bbbf4, 32'h3ce1a820} /* (21, 31, 22) {real, imag} */,
  {32'h3c779bd8, 32'hbd8f7a23} /* (21, 31, 21) {real, imag} */,
  {32'h3d39f976, 32'hbcc716dc} /* (21, 31, 20) {real, imag} */,
  {32'hbc7d1262, 32'h3c992f46} /* (21, 31, 19) {real, imag} */,
  {32'hbd29faec, 32'hbc8eed1e} /* (21, 31, 18) {real, imag} */,
  {32'hbc1123bb, 32'hbcd32df3} /* (21, 31, 17) {real, imag} */,
  {32'h3d000ee4, 32'h00000000} /* (21, 31, 16) {real, imag} */,
  {32'hbc1123bb, 32'h3cd32df3} /* (21, 31, 15) {real, imag} */,
  {32'hbd29faec, 32'h3c8eed1e} /* (21, 31, 14) {real, imag} */,
  {32'hbc7d1262, 32'hbc992f46} /* (21, 31, 13) {real, imag} */,
  {32'h3d39f976, 32'h3cc716dc} /* (21, 31, 12) {real, imag} */,
  {32'h3c779bd8, 32'h3d8f7a23} /* (21, 31, 11) {real, imag} */,
  {32'h3c5bbbf4, 32'hbce1a820} /* (21, 31, 10) {real, imag} */,
  {32'hb7a49000, 32'hbd45ba37} /* (21, 31, 9) {real, imag} */,
  {32'h3d09b68a, 32'hbb074518} /* (21, 31, 8) {real, imag} */,
  {32'h3d98a9fb, 32'hbcb82382} /* (21, 31, 7) {real, imag} */,
  {32'h3c3d54a8, 32'h3d45a486} /* (21, 31, 6) {real, imag} */,
  {32'h3d410f80, 32'h3ca538e6} /* (21, 31, 5) {real, imag} */,
  {32'hbdde38ed, 32'h3d0f3da0} /* (21, 31, 4) {real, imag} */,
  {32'h3cdd09b8, 32'hbd77b55c} /* (21, 31, 3) {real, imag} */,
  {32'h3f47e62b, 32'h3f040067} /* (21, 31, 2) {real, imag} */,
  {32'hc083f146, 32'hc015235c} /* (21, 31, 1) {real, imag} */,
  {32'hc0a6ed23, 32'h00000000} /* (21, 31, 0) {real, imag} */,
  {32'hc0967bf2, 32'h4001178e} /* (21, 30, 31) {real, imag} */,
  {32'h3f91c5ce, 32'hbefd97cc} /* (21, 30, 30) {real, imag} */,
  {32'hbccf4c4c, 32'h3d3878aa} /* (21, 30, 29) {real, imag} */,
  {32'hbe8abaf4, 32'h3be51d80} /* (21, 30, 28) {real, imag} */,
  {32'h3e522419, 32'hbd8ed907} /* (21, 30, 27) {real, imag} */,
  {32'hbe034682, 32'hbe1f7dfa} /* (21, 30, 26) {real, imag} */,
  {32'h3ca7cabe, 32'h3d0e0754} /* (21, 30, 25) {real, imag} */,
  {32'h3d73ddaa, 32'hbdbd5efa} /* (21, 30, 24) {real, imag} */,
  {32'h3d390803, 32'hbc0d5406} /* (21, 30, 23) {real, imag} */,
  {32'h3cedf2f6, 32'h3d978160} /* (21, 30, 22) {real, imag} */,
  {32'h3cc38786, 32'h3c34aa74} /* (21, 30, 21) {real, imag} */,
  {32'h3df27eee, 32'hbda4b384} /* (21, 30, 20) {real, imag} */,
  {32'hbd2ea698, 32'hbcc2ca76} /* (21, 30, 19) {real, imag} */,
  {32'h3d44169e, 32'h3d23deee} /* (21, 30, 18) {real, imag} */,
  {32'h3ce34f22, 32'hbd0e7902} /* (21, 30, 17) {real, imag} */,
  {32'hbcd44e4b, 32'h00000000} /* (21, 30, 16) {real, imag} */,
  {32'h3ce34f22, 32'h3d0e7902} /* (21, 30, 15) {real, imag} */,
  {32'h3d44169e, 32'hbd23deee} /* (21, 30, 14) {real, imag} */,
  {32'hbd2ea698, 32'h3cc2ca76} /* (21, 30, 13) {real, imag} */,
  {32'h3df27eee, 32'h3da4b384} /* (21, 30, 12) {real, imag} */,
  {32'h3cc38786, 32'hbc34aa74} /* (21, 30, 11) {real, imag} */,
  {32'h3cedf2f6, 32'hbd978160} /* (21, 30, 10) {real, imag} */,
  {32'h3d390803, 32'h3c0d5406} /* (21, 30, 9) {real, imag} */,
  {32'h3d73ddaa, 32'h3dbd5efa} /* (21, 30, 8) {real, imag} */,
  {32'h3ca7cabe, 32'hbd0e0754} /* (21, 30, 7) {real, imag} */,
  {32'hbe034682, 32'h3e1f7dfa} /* (21, 30, 6) {real, imag} */,
  {32'h3e522419, 32'h3d8ed907} /* (21, 30, 5) {real, imag} */,
  {32'hbe8abaf4, 32'hbbe51d80} /* (21, 30, 4) {real, imag} */,
  {32'hbccf4c4c, 32'hbd3878aa} /* (21, 30, 3) {real, imag} */,
  {32'h3f91c5ce, 32'h3efd97cc} /* (21, 30, 2) {real, imag} */,
  {32'hc0967bf2, 32'hc001178e} /* (21, 30, 1) {real, imag} */,
  {32'hc0a8a248, 32'h00000000} /* (21, 30, 0) {real, imag} */,
  {32'hc0a5df93, 32'h3fcada0f} /* (21, 29, 31) {real, imag} */,
  {32'h3fb96039, 32'hbe925047} /* (21, 29, 30) {real, imag} */,
  {32'hbce6ddc8, 32'hbda680f9} /* (21, 29, 29) {real, imag} */,
  {32'hbeada238, 32'h3e16d57a} /* (21, 29, 28) {real, imag} */,
  {32'h3e828922, 32'hbd9af5b4} /* (21, 29, 27) {real, imag} */,
  {32'h3c86600d, 32'h3d503f88} /* (21, 29, 26) {real, imag} */,
  {32'h3b01020c, 32'h3d1b4047} /* (21, 29, 25) {real, imag} */,
  {32'h3da1b061, 32'hbd3dd0a3} /* (21, 29, 24) {real, imag} */,
  {32'h3d69278e, 32'hbbb74d68} /* (21, 29, 23) {real, imag} */,
  {32'h3d5f1bea, 32'h3b595ce4} /* (21, 29, 22) {real, imag} */,
  {32'h3ddafa8b, 32'h3ca64624} /* (21, 29, 21) {real, imag} */,
  {32'h3d5e68f6, 32'hbdf806b7} /* (21, 29, 20) {real, imag} */,
  {32'h3d16a31a, 32'hbc98457a} /* (21, 29, 19) {real, imag} */,
  {32'hb9c4f780, 32'hbd2b247b} /* (21, 29, 18) {real, imag} */,
  {32'hbd04588e, 32'h3caa0f90} /* (21, 29, 17) {real, imag} */,
  {32'h3d8a2aa9, 32'h00000000} /* (21, 29, 16) {real, imag} */,
  {32'hbd04588e, 32'hbcaa0f90} /* (21, 29, 15) {real, imag} */,
  {32'hb9c4f780, 32'h3d2b247b} /* (21, 29, 14) {real, imag} */,
  {32'h3d16a31a, 32'h3c98457a} /* (21, 29, 13) {real, imag} */,
  {32'h3d5e68f6, 32'h3df806b7} /* (21, 29, 12) {real, imag} */,
  {32'h3ddafa8b, 32'hbca64624} /* (21, 29, 11) {real, imag} */,
  {32'h3d5f1bea, 32'hbb595ce4} /* (21, 29, 10) {real, imag} */,
  {32'h3d69278e, 32'h3bb74d68} /* (21, 29, 9) {real, imag} */,
  {32'h3da1b061, 32'h3d3dd0a3} /* (21, 29, 8) {real, imag} */,
  {32'h3b01020c, 32'hbd1b4047} /* (21, 29, 7) {real, imag} */,
  {32'h3c86600d, 32'hbd503f88} /* (21, 29, 6) {real, imag} */,
  {32'h3e828922, 32'h3d9af5b4} /* (21, 29, 5) {real, imag} */,
  {32'hbeada238, 32'hbe16d57a} /* (21, 29, 4) {real, imag} */,
  {32'hbce6ddc8, 32'h3da680f9} /* (21, 29, 3) {real, imag} */,
  {32'h3fb96039, 32'h3e925047} /* (21, 29, 2) {real, imag} */,
  {32'hc0a5df93, 32'hbfcada0f} /* (21, 29, 1) {real, imag} */,
  {32'hc0a9a986, 32'h00000000} /* (21, 29, 0) {real, imag} */,
  {32'hc0ab00b6, 32'h3fa98c96} /* (21, 28, 31) {real, imag} */,
  {32'h3fe4d8ac, 32'hbee9d5b4} /* (21, 28, 30) {real, imag} */,
  {32'hbcffaeb0, 32'hbca5ebbc} /* (21, 28, 29) {real, imag} */,
  {32'hbe8c686e, 32'h3e24dfbe} /* (21, 28, 28) {real, imag} */,
  {32'h3e60a86a, 32'hbe45ca52} /* (21, 28, 27) {real, imag} */,
  {32'hbd05e580, 32'h3d495d4f} /* (21, 28, 26) {real, imag} */,
  {32'hbdea3b88, 32'h3d949646} /* (21, 28, 25) {real, imag} */,
  {32'hbb7d48e0, 32'hbdd7bb48} /* (21, 28, 24) {real, imag} */,
  {32'hbc96e03e, 32'h3dafcc20} /* (21, 28, 23) {real, imag} */,
  {32'hbd849bb5, 32'hbc923150} /* (21, 28, 22) {real, imag} */,
  {32'h3d02242c, 32'hbdc90f1a} /* (21, 28, 21) {real, imag} */,
  {32'h3cf6bc80, 32'hbd9491b3} /* (21, 28, 20) {real, imag} */,
  {32'hbd22912b, 32'hbdc9ee7a} /* (21, 28, 19) {real, imag} */,
  {32'hbdca01b6, 32'h3cf88950} /* (21, 28, 18) {real, imag} */,
  {32'hbd7451c6, 32'hbc63dfb3} /* (21, 28, 17) {real, imag} */,
  {32'h3dc51e36, 32'h00000000} /* (21, 28, 16) {real, imag} */,
  {32'hbd7451c6, 32'h3c63dfb3} /* (21, 28, 15) {real, imag} */,
  {32'hbdca01b6, 32'hbcf88950} /* (21, 28, 14) {real, imag} */,
  {32'hbd22912b, 32'h3dc9ee7a} /* (21, 28, 13) {real, imag} */,
  {32'h3cf6bc80, 32'h3d9491b3} /* (21, 28, 12) {real, imag} */,
  {32'h3d02242c, 32'h3dc90f1a} /* (21, 28, 11) {real, imag} */,
  {32'hbd849bb5, 32'h3c923150} /* (21, 28, 10) {real, imag} */,
  {32'hbc96e03e, 32'hbdafcc20} /* (21, 28, 9) {real, imag} */,
  {32'hbb7d48e0, 32'h3dd7bb48} /* (21, 28, 8) {real, imag} */,
  {32'hbdea3b88, 32'hbd949646} /* (21, 28, 7) {real, imag} */,
  {32'hbd05e580, 32'hbd495d4f} /* (21, 28, 6) {real, imag} */,
  {32'h3e60a86a, 32'h3e45ca52} /* (21, 28, 5) {real, imag} */,
  {32'hbe8c686e, 32'hbe24dfbe} /* (21, 28, 4) {real, imag} */,
  {32'hbcffaeb0, 32'h3ca5ebbc} /* (21, 28, 3) {real, imag} */,
  {32'h3fe4d8ac, 32'h3ee9d5b4} /* (21, 28, 2) {real, imag} */,
  {32'hc0ab00b6, 32'hbfa98c96} /* (21, 28, 1) {real, imag} */,
  {32'hc0b4669b, 32'h00000000} /* (21, 28, 0) {real, imag} */,
  {32'hc0a9521a, 32'h3f929c13} /* (21, 27, 31) {real, imag} */,
  {32'h3feada86, 32'hbf027ef1} /* (21, 27, 30) {real, imag} */,
  {32'hbc0bd296, 32'h3b5e1ca0} /* (21, 27, 29) {real, imag} */,
  {32'hbe70cfe4, 32'h3d894972} /* (21, 27, 28) {real, imag} */,
  {32'h3e45d038, 32'hbe34a808} /* (21, 27, 27) {real, imag} */,
  {32'hbd2cb339, 32'hbe1ddf3f} /* (21, 27, 26) {real, imag} */,
  {32'hbdc0b8bf, 32'hbb661890} /* (21, 27, 25) {real, imag} */,
  {32'h3cb28eaf, 32'hbd3804a9} /* (21, 27, 24) {real, imag} */,
  {32'h3db16636, 32'h3c1f7c4f} /* (21, 27, 23) {real, imag} */,
  {32'hbd013311, 32'h3cc5a20e} /* (21, 27, 22) {real, imag} */,
  {32'h3d669882, 32'h3d811c14} /* (21, 27, 21) {real, imag} */,
  {32'hbd79b1d6, 32'h3ccfd993} /* (21, 27, 20) {real, imag} */,
  {32'h3b9605e0, 32'h3cb10704} /* (21, 27, 19) {real, imag} */,
  {32'h3d35389c, 32'h3c4a2b3c} /* (21, 27, 18) {real, imag} */,
  {32'hbb2fc074, 32'h3d1d9ba4} /* (21, 27, 17) {real, imag} */,
  {32'hbe12b8a9, 32'h00000000} /* (21, 27, 16) {real, imag} */,
  {32'hbb2fc074, 32'hbd1d9ba4} /* (21, 27, 15) {real, imag} */,
  {32'h3d35389c, 32'hbc4a2b3c} /* (21, 27, 14) {real, imag} */,
  {32'h3b9605e0, 32'hbcb10704} /* (21, 27, 13) {real, imag} */,
  {32'hbd79b1d6, 32'hbccfd993} /* (21, 27, 12) {real, imag} */,
  {32'h3d669882, 32'hbd811c14} /* (21, 27, 11) {real, imag} */,
  {32'hbd013311, 32'hbcc5a20e} /* (21, 27, 10) {real, imag} */,
  {32'h3db16636, 32'hbc1f7c4f} /* (21, 27, 9) {real, imag} */,
  {32'h3cb28eaf, 32'h3d3804a9} /* (21, 27, 8) {real, imag} */,
  {32'hbdc0b8bf, 32'h3b661890} /* (21, 27, 7) {real, imag} */,
  {32'hbd2cb339, 32'h3e1ddf3f} /* (21, 27, 6) {real, imag} */,
  {32'h3e45d038, 32'h3e34a808} /* (21, 27, 5) {real, imag} */,
  {32'hbe70cfe4, 32'hbd894972} /* (21, 27, 4) {real, imag} */,
  {32'hbc0bd296, 32'hbb5e1ca0} /* (21, 27, 3) {real, imag} */,
  {32'h3feada86, 32'h3f027ef1} /* (21, 27, 2) {real, imag} */,
  {32'hc0a9521a, 32'hbf929c13} /* (21, 27, 1) {real, imag} */,
  {32'hc0b9eb55, 32'h00000000} /* (21, 27, 0) {real, imag} */,
  {32'hc0a4d6b2, 32'h3f76f4dd} /* (21, 26, 31) {real, imag} */,
  {32'h3ff94024, 32'hbec89274} /* (21, 26, 30) {real, imag} */,
  {32'hbcb1a601, 32'h3c21316a} /* (21, 26, 29) {real, imag} */,
  {32'hbeb6c335, 32'h3bb0acb0} /* (21, 26, 28) {real, imag} */,
  {32'h3e825d06, 32'hbe168607} /* (21, 26, 27) {real, imag} */,
  {32'h3d387ef6, 32'h3d4dfa6c} /* (21, 26, 26) {real, imag} */,
  {32'hbceb1864, 32'hbdbbeee3} /* (21, 26, 25) {real, imag} */,
  {32'h3d7b1879, 32'hbb40e328} /* (21, 26, 24) {real, imag} */,
  {32'h3d73af6a, 32'h3db393fb} /* (21, 26, 23) {real, imag} */,
  {32'h3df23e48, 32'hbde1a068} /* (21, 26, 22) {real, imag} */,
  {32'hbd9d83da, 32'hbe6b4bd6} /* (21, 26, 21) {real, imag} */,
  {32'hbd35e344, 32'hbd1d8eed} /* (21, 26, 20) {real, imag} */,
  {32'hbd045f50, 32'h3cc6134d} /* (21, 26, 19) {real, imag} */,
  {32'h3b26ef00, 32'h3c2b0d42} /* (21, 26, 18) {real, imag} */,
  {32'h3c30285a, 32'hbcdbf87f} /* (21, 26, 17) {real, imag} */,
  {32'hbc95addf, 32'h00000000} /* (21, 26, 16) {real, imag} */,
  {32'h3c30285a, 32'h3cdbf87f} /* (21, 26, 15) {real, imag} */,
  {32'h3b26ef00, 32'hbc2b0d42} /* (21, 26, 14) {real, imag} */,
  {32'hbd045f50, 32'hbcc6134d} /* (21, 26, 13) {real, imag} */,
  {32'hbd35e344, 32'h3d1d8eed} /* (21, 26, 12) {real, imag} */,
  {32'hbd9d83da, 32'h3e6b4bd6} /* (21, 26, 11) {real, imag} */,
  {32'h3df23e48, 32'h3de1a068} /* (21, 26, 10) {real, imag} */,
  {32'h3d73af6a, 32'hbdb393fb} /* (21, 26, 9) {real, imag} */,
  {32'h3d7b1879, 32'h3b40e328} /* (21, 26, 8) {real, imag} */,
  {32'hbceb1864, 32'h3dbbeee3} /* (21, 26, 7) {real, imag} */,
  {32'h3d387ef6, 32'hbd4dfa6c} /* (21, 26, 6) {real, imag} */,
  {32'h3e825d06, 32'h3e168607} /* (21, 26, 5) {real, imag} */,
  {32'hbeb6c335, 32'hbbb0acb0} /* (21, 26, 4) {real, imag} */,
  {32'hbcb1a601, 32'hbc21316a} /* (21, 26, 3) {real, imag} */,
  {32'h3ff94024, 32'h3ec89274} /* (21, 26, 2) {real, imag} */,
  {32'hc0a4d6b2, 32'hbf76f4dd} /* (21, 26, 1) {real, imag} */,
  {32'hc0b00a7f, 32'h00000000} /* (21, 26, 0) {real, imag} */,
  {32'hc09c1ad5, 32'h3f4aa897} /* (21, 25, 31) {real, imag} */,
  {32'h3ff2da24, 32'hbeca8274} /* (21, 25, 30) {real, imag} */,
  {32'hbda13a00, 32'h3c9addfe} /* (21, 25, 29) {real, imag} */,
  {32'hbe395ce1, 32'hbd9986de} /* (21, 25, 28) {real, imag} */,
  {32'h3e8b5af2, 32'hbe6623be} /* (21, 25, 27) {real, imag} */,
  {32'hbd890a7c, 32'h3d34f54d} /* (21, 25, 26) {real, imag} */,
  {32'hbc6d1b28, 32'h3dae1cef} /* (21, 25, 25) {real, imag} */,
  {32'h3ce2923a, 32'hbdbabdee} /* (21, 25, 24) {real, imag} */,
  {32'h3d8807e4, 32'h3db5db92} /* (21, 25, 23) {real, imag} */,
  {32'hbb1c7bf0, 32'h3c2b72be} /* (21, 25, 22) {real, imag} */,
  {32'h3d2d8dac, 32'hbd079a9d} /* (21, 25, 21) {real, imag} */,
  {32'hbd3aea4a, 32'h3d92318e} /* (21, 25, 20) {real, imag} */,
  {32'hbd44da92, 32'h3d6345bb} /* (21, 25, 19) {real, imag} */,
  {32'h3ca8f5aa, 32'h3cdfc91d} /* (21, 25, 18) {real, imag} */,
  {32'hbca0000e, 32'hbd0ca0dc} /* (21, 25, 17) {real, imag} */,
  {32'hbab30e20, 32'h00000000} /* (21, 25, 16) {real, imag} */,
  {32'hbca0000e, 32'h3d0ca0dc} /* (21, 25, 15) {real, imag} */,
  {32'h3ca8f5aa, 32'hbcdfc91d} /* (21, 25, 14) {real, imag} */,
  {32'hbd44da92, 32'hbd6345bb} /* (21, 25, 13) {real, imag} */,
  {32'hbd3aea4a, 32'hbd92318e} /* (21, 25, 12) {real, imag} */,
  {32'h3d2d8dac, 32'h3d079a9d} /* (21, 25, 11) {real, imag} */,
  {32'hbb1c7bf0, 32'hbc2b72be} /* (21, 25, 10) {real, imag} */,
  {32'h3d8807e4, 32'hbdb5db92} /* (21, 25, 9) {real, imag} */,
  {32'h3ce2923a, 32'h3dbabdee} /* (21, 25, 8) {real, imag} */,
  {32'hbc6d1b28, 32'hbdae1cef} /* (21, 25, 7) {real, imag} */,
  {32'hbd890a7c, 32'hbd34f54d} /* (21, 25, 6) {real, imag} */,
  {32'h3e8b5af2, 32'h3e6623be} /* (21, 25, 5) {real, imag} */,
  {32'hbe395ce1, 32'h3d9986de} /* (21, 25, 4) {real, imag} */,
  {32'hbda13a00, 32'hbc9addfe} /* (21, 25, 3) {real, imag} */,
  {32'h3ff2da24, 32'h3eca8274} /* (21, 25, 2) {real, imag} */,
  {32'hc09c1ad5, 32'hbf4aa897} /* (21, 25, 1) {real, imag} */,
  {32'hc09f28fd, 32'h00000000} /* (21, 25, 0) {real, imag} */,
  {32'hc088f257, 32'h3f016d16} /* (21, 24, 31) {real, imag} */,
  {32'h3fd5b090, 32'hbef1ba10} /* (21, 24, 30) {real, imag} */,
  {32'hbd8fdbc3, 32'hbd68d4e2} /* (21, 24, 29) {real, imag} */,
  {32'hbe64e92e, 32'h3de7391f} /* (21, 24, 28) {real, imag} */,
  {32'h3e7ae9b2, 32'hbe47afd9} /* (21, 24, 27) {real, imag} */,
  {32'hbd8bdd4a, 32'hbdb1db42} /* (21, 24, 26) {real, imag} */,
  {32'hbab792d0, 32'h3d301d35} /* (21, 24, 25) {real, imag} */,
  {32'h3ddd34f4, 32'hbdeb958c} /* (21, 24, 24) {real, imag} */,
  {32'h3d7ea4d9, 32'h3e00b2aa} /* (21, 24, 23) {real, imag} */,
  {32'h3c788123, 32'hbd8787a1} /* (21, 24, 22) {real, imag} */,
  {32'hbd370dde, 32'h3c52f2f6} /* (21, 24, 21) {real, imag} */,
  {32'h3d67fbc4, 32'hbc9fac0c} /* (21, 24, 20) {real, imag} */,
  {32'h3b129070, 32'h3db295ed} /* (21, 24, 19) {real, imag} */,
  {32'h3dc91d7f, 32'hbd0940c1} /* (21, 24, 18) {real, imag} */,
  {32'hbd6b6418, 32'hbcf1e73e} /* (21, 24, 17) {real, imag} */,
  {32'h3af0a298, 32'h00000000} /* (21, 24, 16) {real, imag} */,
  {32'hbd6b6418, 32'h3cf1e73e} /* (21, 24, 15) {real, imag} */,
  {32'h3dc91d7f, 32'h3d0940c1} /* (21, 24, 14) {real, imag} */,
  {32'h3b129070, 32'hbdb295ed} /* (21, 24, 13) {real, imag} */,
  {32'h3d67fbc4, 32'h3c9fac0c} /* (21, 24, 12) {real, imag} */,
  {32'hbd370dde, 32'hbc52f2f6} /* (21, 24, 11) {real, imag} */,
  {32'h3c788123, 32'h3d8787a1} /* (21, 24, 10) {real, imag} */,
  {32'h3d7ea4d9, 32'hbe00b2aa} /* (21, 24, 9) {real, imag} */,
  {32'h3ddd34f4, 32'h3deb958c} /* (21, 24, 8) {real, imag} */,
  {32'hbab792d0, 32'hbd301d35} /* (21, 24, 7) {real, imag} */,
  {32'hbd8bdd4a, 32'h3db1db42} /* (21, 24, 6) {real, imag} */,
  {32'h3e7ae9b2, 32'h3e47afd9} /* (21, 24, 5) {real, imag} */,
  {32'hbe64e92e, 32'hbde7391f} /* (21, 24, 4) {real, imag} */,
  {32'hbd8fdbc3, 32'h3d68d4e2} /* (21, 24, 3) {real, imag} */,
  {32'h3fd5b090, 32'h3ef1ba10} /* (21, 24, 2) {real, imag} */,
  {32'hc088f257, 32'hbf016d16} /* (21, 24, 1) {real, imag} */,
  {32'hc082342c, 32'h00000000} /* (21, 24, 0) {real, imag} */,
  {32'hc05fa34c, 32'h3ec07232} /* (21, 23, 31) {real, imag} */,
  {32'h3fa8bf49, 32'hbebc09aa} /* (21, 23, 30) {real, imag} */,
  {32'hbc9ace06, 32'hb9cff360} /* (21, 23, 29) {real, imag} */,
  {32'hbdc6c4f6, 32'h3df0af06} /* (21, 23, 28) {real, imag} */,
  {32'h3e82f420, 32'hbcf94652} /* (21, 23, 27) {real, imag} */,
  {32'h3cde1909, 32'hbc7bc308} /* (21, 23, 26) {real, imag} */,
  {32'hbdd6be16, 32'hbc3033cc} /* (21, 23, 25) {real, imag} */,
  {32'h3e02bf7b, 32'hbd6a6573} /* (21, 23, 24) {real, imag} */,
  {32'hbdbbd81a, 32'hbd5aa690} /* (21, 23, 23) {real, imag} */,
  {32'hbcbce542, 32'hbd677b78} /* (21, 23, 22) {real, imag} */,
  {32'h3c91f4b4, 32'hbd365814} /* (21, 23, 21) {real, imag} */,
  {32'hbca25cb6, 32'h3c66cba2} /* (21, 23, 20) {real, imag} */,
  {32'hbc0cf480, 32'h3d22950e} /* (21, 23, 19) {real, imag} */,
  {32'hbadd8a28, 32'hbdd8a56b} /* (21, 23, 18) {real, imag} */,
  {32'hbcfa1334, 32'hbc154af0} /* (21, 23, 17) {real, imag} */,
  {32'h3d905d3e, 32'h00000000} /* (21, 23, 16) {real, imag} */,
  {32'hbcfa1334, 32'h3c154af0} /* (21, 23, 15) {real, imag} */,
  {32'hbadd8a28, 32'h3dd8a56b} /* (21, 23, 14) {real, imag} */,
  {32'hbc0cf480, 32'hbd22950e} /* (21, 23, 13) {real, imag} */,
  {32'hbca25cb6, 32'hbc66cba2} /* (21, 23, 12) {real, imag} */,
  {32'h3c91f4b4, 32'h3d365814} /* (21, 23, 11) {real, imag} */,
  {32'hbcbce542, 32'h3d677b78} /* (21, 23, 10) {real, imag} */,
  {32'hbdbbd81a, 32'h3d5aa690} /* (21, 23, 9) {real, imag} */,
  {32'h3e02bf7b, 32'h3d6a6573} /* (21, 23, 8) {real, imag} */,
  {32'hbdd6be16, 32'h3c3033cc} /* (21, 23, 7) {real, imag} */,
  {32'h3cde1909, 32'h3c7bc308} /* (21, 23, 6) {real, imag} */,
  {32'h3e82f420, 32'h3cf94652} /* (21, 23, 5) {real, imag} */,
  {32'hbdc6c4f6, 32'hbdf0af06} /* (21, 23, 4) {real, imag} */,
  {32'hbc9ace06, 32'h39cff360} /* (21, 23, 3) {real, imag} */,
  {32'h3fa8bf49, 32'h3ebc09aa} /* (21, 23, 2) {real, imag} */,
  {32'hc05fa34c, 32'hbec07232} /* (21, 23, 1) {real, imag} */,
  {32'hc0603cea, 32'h00000000} /* (21, 23, 0) {real, imag} */,
  {32'hc021986b, 32'h3e32bf70} /* (21, 22, 31) {real, imag} */,
  {32'h3f54bd0d, 32'hbebd62ea} /* (21, 22, 30) {real, imag} */,
  {32'hbd213f66, 32'hbc2b728c} /* (21, 22, 29) {real, imag} */,
  {32'hbdebd888, 32'h3d79c787} /* (21, 22, 28) {real, imag} */,
  {32'h3e8e062e, 32'hbd274f77} /* (21, 22, 27) {real, imag} */,
  {32'hbc37fe78, 32'hbd9028c9} /* (21, 22, 26) {real, imag} */,
  {32'hbceeb084, 32'h3cf51c09} /* (21, 22, 25) {real, imag} */,
  {32'h3d5a231b, 32'h3cb262f0} /* (21, 22, 24) {real, imag} */,
  {32'hbda9fdaf, 32'h3ad16cb0} /* (21, 22, 23) {real, imag} */,
  {32'h3d510c2e, 32'hbde84e8a} /* (21, 22, 22) {real, imag} */,
  {32'h3be3cc74, 32'hbd01def7} /* (21, 22, 21) {real, imag} */,
  {32'hbd1f2c52, 32'hbd811056} /* (21, 22, 20) {real, imag} */,
  {32'h3ca609f8, 32'hbb73976e} /* (21, 22, 19) {real, imag} */,
  {32'h3d35380a, 32'hbded7952} /* (21, 22, 18) {real, imag} */,
  {32'h3a8d9328, 32'h3d6302cc} /* (21, 22, 17) {real, imag} */,
  {32'h3d26e010, 32'h00000000} /* (21, 22, 16) {real, imag} */,
  {32'h3a8d9328, 32'hbd6302cc} /* (21, 22, 15) {real, imag} */,
  {32'h3d35380a, 32'h3ded7952} /* (21, 22, 14) {real, imag} */,
  {32'h3ca609f8, 32'h3b73976e} /* (21, 22, 13) {real, imag} */,
  {32'hbd1f2c52, 32'h3d811056} /* (21, 22, 12) {real, imag} */,
  {32'h3be3cc74, 32'h3d01def7} /* (21, 22, 11) {real, imag} */,
  {32'h3d510c2e, 32'h3de84e8a} /* (21, 22, 10) {real, imag} */,
  {32'hbda9fdaf, 32'hbad16cb0} /* (21, 22, 9) {real, imag} */,
  {32'h3d5a231b, 32'hbcb262f0} /* (21, 22, 8) {real, imag} */,
  {32'hbceeb084, 32'hbcf51c09} /* (21, 22, 7) {real, imag} */,
  {32'hbc37fe78, 32'h3d9028c9} /* (21, 22, 6) {real, imag} */,
  {32'h3e8e062e, 32'h3d274f77} /* (21, 22, 5) {real, imag} */,
  {32'hbdebd888, 32'hbd79c787} /* (21, 22, 4) {real, imag} */,
  {32'hbd213f66, 32'h3c2b728c} /* (21, 22, 3) {real, imag} */,
  {32'h3f54bd0d, 32'h3ebd62ea} /* (21, 22, 2) {real, imag} */,
  {32'hc021986b, 32'hbe32bf70} /* (21, 22, 1) {real, imag} */,
  {32'hc01fbb0d, 32'h00000000} /* (21, 22, 0) {real, imag} */,
  {32'hbf49cc11, 32'h3d175ae0} /* (21, 21, 31) {real, imag} */,
  {32'h3e018d42, 32'hbe4f30ae} /* (21, 21, 30) {real, imag} */,
  {32'hbd4f86e2, 32'h3d6e68c5} /* (21, 21, 29) {real, imag} */,
  {32'hbe12aeb5, 32'hbd6b3c08} /* (21, 21, 28) {real, imag} */,
  {32'h3d469014, 32'hbd39ff65} /* (21, 21, 27) {real, imag} */,
  {32'hbda32c65, 32'hbca7e82c} /* (21, 21, 26) {real, imag} */,
  {32'hbb8a5a1c, 32'hbc272703} /* (21, 21, 25) {real, imag} */,
  {32'h3c699070, 32'hbd54a416} /* (21, 21, 24) {real, imag} */,
  {32'hbc66659f, 32'h3c55b8b9} /* (21, 21, 23) {real, imag} */,
  {32'hbd046bc3, 32'hbdc9f851} /* (21, 21, 22) {real, imag} */,
  {32'h3b4e5020, 32'h3b4b7420} /* (21, 21, 21) {real, imag} */,
  {32'h3d0e4eb8, 32'hbc8d94f3} /* (21, 21, 20) {real, imag} */,
  {32'hbb42d340, 32'hbd075237} /* (21, 21, 19) {real, imag} */,
  {32'h3d18f72b, 32'hbd964e39} /* (21, 21, 18) {real, imag} */,
  {32'h3db3962e, 32'hbae35a68} /* (21, 21, 17) {real, imag} */,
  {32'hbc9aa541, 32'h00000000} /* (21, 21, 16) {real, imag} */,
  {32'h3db3962e, 32'h3ae35a68} /* (21, 21, 15) {real, imag} */,
  {32'h3d18f72b, 32'h3d964e39} /* (21, 21, 14) {real, imag} */,
  {32'hbb42d340, 32'h3d075237} /* (21, 21, 13) {real, imag} */,
  {32'h3d0e4eb8, 32'h3c8d94f3} /* (21, 21, 12) {real, imag} */,
  {32'h3b4e5020, 32'hbb4b7420} /* (21, 21, 11) {real, imag} */,
  {32'hbd046bc3, 32'h3dc9f851} /* (21, 21, 10) {real, imag} */,
  {32'hbc66659f, 32'hbc55b8b9} /* (21, 21, 9) {real, imag} */,
  {32'h3c699070, 32'h3d54a416} /* (21, 21, 8) {real, imag} */,
  {32'hbb8a5a1c, 32'h3c272703} /* (21, 21, 7) {real, imag} */,
  {32'hbda32c65, 32'h3ca7e82c} /* (21, 21, 6) {real, imag} */,
  {32'h3d469014, 32'h3d39ff65} /* (21, 21, 5) {real, imag} */,
  {32'hbe12aeb5, 32'h3d6b3c08} /* (21, 21, 4) {real, imag} */,
  {32'hbd4f86e2, 32'hbd6e68c5} /* (21, 21, 3) {real, imag} */,
  {32'h3e018d42, 32'h3e4f30ae} /* (21, 21, 2) {real, imag} */,
  {32'hbf49cc11, 32'hbd175ae0} /* (21, 21, 1) {real, imag} */,
  {32'hbf862669, 32'h00000000} /* (21, 21, 0) {real, imag} */,
  {32'h3fa00c5f, 32'hbe3a804c} /* (21, 20, 31) {real, imag} */,
  {32'hbf245fbb, 32'h3d846104} /* (21, 20, 30) {real, imag} */,
  {32'hbda03e4c, 32'h3e276568} /* (21, 20, 29) {real, imag} */,
  {32'hbdba0f3e, 32'hbdaabf02} /* (21, 20, 28) {real, imag} */,
  {32'hbdd8dcea, 32'h3d84b96e} /* (21, 20, 27) {real, imag} */,
  {32'hbe020b5f, 32'hbe024399} /* (21, 20, 26) {real, imag} */,
  {32'h3d33831a, 32'h3d0d953c} /* (21, 20, 25) {real, imag} */,
  {32'h3d388039, 32'hbd09b3cb} /* (21, 20, 24) {real, imag} */,
  {32'hbcc576ce, 32'h3d82d49a} /* (21, 20, 23) {real, imag} */,
  {32'h3b40ad78, 32'hbe0e4bf0} /* (21, 20, 22) {real, imag} */,
  {32'h3d291083, 32'h3e1cd1e4} /* (21, 20, 21) {real, imag} */,
  {32'h3c97fcf8, 32'h3cce09ae} /* (21, 20, 20) {real, imag} */,
  {32'h3c111380, 32'hbd8abb72} /* (21, 20, 19) {real, imag} */,
  {32'h3d2b7d18, 32'hbd7fbe00} /* (21, 20, 18) {real, imag} */,
  {32'hbdcace22, 32'hbd1aa9f0} /* (21, 20, 17) {real, imag} */,
  {32'h3d8bdfdc, 32'h00000000} /* (21, 20, 16) {real, imag} */,
  {32'hbdcace22, 32'h3d1aa9f0} /* (21, 20, 15) {real, imag} */,
  {32'h3d2b7d18, 32'h3d7fbe00} /* (21, 20, 14) {real, imag} */,
  {32'h3c111380, 32'h3d8abb72} /* (21, 20, 13) {real, imag} */,
  {32'h3c97fcf8, 32'hbcce09ae} /* (21, 20, 12) {real, imag} */,
  {32'h3d291083, 32'hbe1cd1e4} /* (21, 20, 11) {real, imag} */,
  {32'h3b40ad78, 32'h3e0e4bf0} /* (21, 20, 10) {real, imag} */,
  {32'hbcc576ce, 32'hbd82d49a} /* (21, 20, 9) {real, imag} */,
  {32'h3d388039, 32'h3d09b3cb} /* (21, 20, 8) {real, imag} */,
  {32'h3d33831a, 32'hbd0d953c} /* (21, 20, 7) {real, imag} */,
  {32'hbe020b5f, 32'h3e024399} /* (21, 20, 6) {real, imag} */,
  {32'hbdd8dcea, 32'hbd84b96e} /* (21, 20, 5) {real, imag} */,
  {32'hbdba0f3e, 32'h3daabf02} /* (21, 20, 4) {real, imag} */,
  {32'hbda03e4c, 32'hbe276568} /* (21, 20, 3) {real, imag} */,
  {32'hbf245fbb, 32'hbd846104} /* (21, 20, 2) {real, imag} */,
  {32'h3fa00c5f, 32'h3e3a804c} /* (21, 20, 1) {real, imag} */,
  {32'h3e92d1c4, 32'h00000000} /* (21, 20, 0) {real, imag} */,
  {32'h402a3934, 32'hbef09bb4} /* (21, 19, 31) {real, imag} */,
  {32'hbf88cf5e, 32'h3e490f6c} /* (21, 19, 30) {real, imag} */,
  {32'h3b62fbe0, 32'h3d5aa2b1} /* (21, 19, 29) {real, imag} */,
  {32'h3d7307fc, 32'hbd1b379c} /* (21, 19, 28) {real, imag} */,
  {32'hbe35bb87, 32'h3dabece8} /* (21, 19, 27) {real, imag} */,
  {32'hbdbbcfca, 32'h3cbc44fc} /* (21, 19, 26) {real, imag} */,
  {32'hbcc34476, 32'h3dd38008} /* (21, 19, 25) {real, imag} */,
  {32'hbe184ac5, 32'h3ca2238a} /* (21, 19, 24) {real, imag} */,
  {32'hbd5dd2e1, 32'hbcc7035c} /* (21, 19, 23) {real, imag} */,
  {32'hbbd0709c, 32'hbdd79260} /* (21, 19, 22) {real, imag} */,
  {32'h3cc63d5a, 32'hbcbdd0d6} /* (21, 19, 21) {real, imag} */,
  {32'h3db03115, 32'hbd7397ac} /* (21, 19, 20) {real, imag} */,
  {32'hbd8b42bf, 32'hbcdc2efc} /* (21, 19, 19) {real, imag} */,
  {32'hbb945098, 32'h3cccb82e} /* (21, 19, 18) {real, imag} */,
  {32'h3ce11d90, 32'hbcffc02d} /* (21, 19, 17) {real, imag} */,
  {32'h3d223d52, 32'h00000000} /* (21, 19, 16) {real, imag} */,
  {32'h3ce11d90, 32'h3cffc02d} /* (21, 19, 15) {real, imag} */,
  {32'hbb945098, 32'hbcccb82e} /* (21, 19, 14) {real, imag} */,
  {32'hbd8b42bf, 32'h3cdc2efc} /* (21, 19, 13) {real, imag} */,
  {32'h3db03115, 32'h3d7397ac} /* (21, 19, 12) {real, imag} */,
  {32'h3cc63d5a, 32'h3cbdd0d6} /* (21, 19, 11) {real, imag} */,
  {32'hbbd0709c, 32'h3dd79260} /* (21, 19, 10) {real, imag} */,
  {32'hbd5dd2e1, 32'h3cc7035c} /* (21, 19, 9) {real, imag} */,
  {32'hbe184ac5, 32'hbca2238a} /* (21, 19, 8) {real, imag} */,
  {32'hbcc34476, 32'hbdd38008} /* (21, 19, 7) {real, imag} */,
  {32'hbdbbcfca, 32'hbcbc44fc} /* (21, 19, 6) {real, imag} */,
  {32'hbe35bb87, 32'hbdabece8} /* (21, 19, 5) {real, imag} */,
  {32'h3d7307fc, 32'h3d1b379c} /* (21, 19, 4) {real, imag} */,
  {32'h3b62fbe0, 32'hbd5aa2b1} /* (21, 19, 3) {real, imag} */,
  {32'hbf88cf5e, 32'hbe490f6c} /* (21, 19, 2) {real, imag} */,
  {32'h402a3934, 32'h3ef09bb4} /* (21, 19, 1) {real, imag} */,
  {32'h3f9d0f4c, 32'h00000000} /* (21, 19, 0) {real, imag} */,
  {32'h40659d8b, 32'hbef30184} /* (21, 18, 31) {real, imag} */,
  {32'hbfb13d7c, 32'h3e6ec7e5} /* (21, 18, 30) {real, imag} */,
  {32'h3b86e3b0, 32'h3de82fc7} /* (21, 18, 29) {real, imag} */,
  {32'h3ddf42ca, 32'hbdef717e} /* (21, 18, 28) {real, imag} */,
  {32'hbd55de0a, 32'h3dd01456} /* (21, 18, 27) {real, imag} */,
  {32'hbdc55101, 32'h3da0d55e} /* (21, 18, 26) {real, imag} */,
  {32'h3d080322, 32'h3dc8aaa5} /* (21, 18, 25) {real, imag} */,
  {32'hbc153340, 32'h3d040dc4} /* (21, 18, 24) {real, imag} */,
  {32'hbd63dc25, 32'hbb70cee0} /* (21, 18, 23) {real, imag} */,
  {32'h3c7c3268, 32'h3d9911e9} /* (21, 18, 22) {real, imag} */,
  {32'hbd1ee4ca, 32'hbe4020f2} /* (21, 18, 21) {real, imag} */,
  {32'hbd58eed0, 32'h3d8b51e6} /* (21, 18, 20) {real, imag} */,
  {32'h3b8b165a, 32'hbc7fa339} /* (21, 18, 19) {real, imag} */,
  {32'hbcaf1606, 32'hbd205bda} /* (21, 18, 18) {real, imag} */,
  {32'hbd618b59, 32'hbcad794f} /* (21, 18, 17) {real, imag} */,
  {32'hbd1a9c73, 32'h00000000} /* (21, 18, 16) {real, imag} */,
  {32'hbd618b59, 32'h3cad794f} /* (21, 18, 15) {real, imag} */,
  {32'hbcaf1606, 32'h3d205bda} /* (21, 18, 14) {real, imag} */,
  {32'h3b8b165a, 32'h3c7fa339} /* (21, 18, 13) {real, imag} */,
  {32'hbd58eed0, 32'hbd8b51e6} /* (21, 18, 12) {real, imag} */,
  {32'hbd1ee4ca, 32'h3e4020f2} /* (21, 18, 11) {real, imag} */,
  {32'h3c7c3268, 32'hbd9911e9} /* (21, 18, 10) {real, imag} */,
  {32'hbd63dc25, 32'h3b70cee0} /* (21, 18, 9) {real, imag} */,
  {32'hbc153340, 32'hbd040dc4} /* (21, 18, 8) {real, imag} */,
  {32'h3d080322, 32'hbdc8aaa5} /* (21, 18, 7) {real, imag} */,
  {32'hbdc55101, 32'hbda0d55e} /* (21, 18, 6) {real, imag} */,
  {32'hbd55de0a, 32'hbdd01456} /* (21, 18, 5) {real, imag} */,
  {32'h3ddf42ca, 32'h3def717e} /* (21, 18, 4) {real, imag} */,
  {32'h3b86e3b0, 32'hbde82fc7} /* (21, 18, 3) {real, imag} */,
  {32'hbfb13d7c, 32'hbe6ec7e5} /* (21, 18, 2) {real, imag} */,
  {32'h40659d8b, 32'h3ef30184} /* (21, 18, 1) {real, imag} */,
  {32'h400b3ad0, 32'h00000000} /* (21, 18, 0) {real, imag} */,
  {32'h408742d6, 32'hbf076aae} /* (21, 17, 31) {real, imag} */,
  {32'hbfc1a9f6, 32'h3ea84092} /* (21, 17, 30) {real, imag} */,
  {32'hbcd96478, 32'h3e913159} /* (21, 17, 29) {real, imag} */,
  {32'h3e08d176, 32'hbe0461aa} /* (21, 17, 28) {real, imag} */,
  {32'hbe0f9474, 32'h3e6b872a} /* (21, 17, 27) {real, imag} */,
  {32'h3c149c94, 32'h3d264f72} /* (21, 17, 26) {real, imag} */,
  {32'h3d0d65ff, 32'h3e26187f} /* (21, 17, 25) {real, imag} */,
  {32'h3d31da78, 32'h3d880235} /* (21, 17, 24) {real, imag} */,
  {32'hbdab447f, 32'h3d977de6} /* (21, 17, 23) {real, imag} */,
  {32'hbd905778, 32'h3d14042c} /* (21, 17, 22) {real, imag} */,
  {32'hbd2bd5a9, 32'h3d2f032a} /* (21, 17, 21) {real, imag} */,
  {32'hbc6563ec, 32'hbd66ac94} /* (21, 17, 20) {real, imag} */,
  {32'h3d18538b, 32'h3c82ecb8} /* (21, 17, 19) {real, imag} */,
  {32'h3d3ef4e1, 32'h3d086004} /* (21, 17, 18) {real, imag} */,
  {32'hbd93485e, 32'hbccf0331} /* (21, 17, 17) {real, imag} */,
  {32'hbd6b2c4e, 32'h00000000} /* (21, 17, 16) {real, imag} */,
  {32'hbd93485e, 32'h3ccf0331} /* (21, 17, 15) {real, imag} */,
  {32'h3d3ef4e1, 32'hbd086004} /* (21, 17, 14) {real, imag} */,
  {32'h3d18538b, 32'hbc82ecb8} /* (21, 17, 13) {real, imag} */,
  {32'hbc6563ec, 32'h3d66ac94} /* (21, 17, 12) {real, imag} */,
  {32'hbd2bd5a9, 32'hbd2f032a} /* (21, 17, 11) {real, imag} */,
  {32'hbd905778, 32'hbd14042c} /* (21, 17, 10) {real, imag} */,
  {32'hbdab447f, 32'hbd977de6} /* (21, 17, 9) {real, imag} */,
  {32'h3d31da78, 32'hbd880235} /* (21, 17, 8) {real, imag} */,
  {32'h3d0d65ff, 32'hbe26187f} /* (21, 17, 7) {real, imag} */,
  {32'h3c149c94, 32'hbd264f72} /* (21, 17, 6) {real, imag} */,
  {32'hbe0f9474, 32'hbe6b872a} /* (21, 17, 5) {real, imag} */,
  {32'h3e08d176, 32'h3e0461aa} /* (21, 17, 4) {real, imag} */,
  {32'hbcd96478, 32'hbe913159} /* (21, 17, 3) {real, imag} */,
  {32'hbfc1a9f6, 32'hbea84092} /* (21, 17, 2) {real, imag} */,
  {32'h408742d6, 32'h3f076aae} /* (21, 17, 1) {real, imag} */,
  {32'h402e1f78, 32'h00000000} /* (21, 17, 0) {real, imag} */,
  {32'h408df644, 32'hbee09fb8} /* (21, 16, 31) {real, imag} */,
  {32'hbfbb78ba, 32'h3eb74fe6} /* (21, 16, 30) {real, imag} */,
  {32'hbdd02b58, 32'h3e0561a4} /* (21, 16, 29) {real, imag} */,
  {32'h3e9ba107, 32'hbd57bc85} /* (21, 16, 28) {real, imag} */,
  {32'hbea2e972, 32'h3d3ca48e} /* (21, 16, 27) {real, imag} */,
  {32'h3de08d46, 32'h3d52cb64} /* (21, 16, 26) {real, imag} */,
  {32'hbcf45928, 32'hbd226e04} /* (21, 16, 25) {real, imag} */,
  {32'hbcfec6bb, 32'h3e06d587} /* (21, 16, 24) {real, imag} */,
  {32'hbd9c2c15, 32'h3d4f4668} /* (21, 16, 23) {real, imag} */,
  {32'hbc60a30d, 32'hbd32c03a} /* (21, 16, 22) {real, imag} */,
  {32'h3b491c70, 32'h3d8e7421} /* (21, 16, 21) {real, imag} */,
  {32'h3d036c4b, 32'hbd649694} /* (21, 16, 20) {real, imag} */,
  {32'hbd41ac1c, 32'h3c3cd702} /* (21, 16, 19) {real, imag} */,
  {32'h3bd96b18, 32'h3dd30eda} /* (21, 16, 18) {real, imag} */,
  {32'hbbe14900, 32'h3d584c0a} /* (21, 16, 17) {real, imag} */,
  {32'h3d421127, 32'h00000000} /* (21, 16, 16) {real, imag} */,
  {32'hbbe14900, 32'hbd584c0a} /* (21, 16, 15) {real, imag} */,
  {32'h3bd96b18, 32'hbdd30eda} /* (21, 16, 14) {real, imag} */,
  {32'hbd41ac1c, 32'hbc3cd702} /* (21, 16, 13) {real, imag} */,
  {32'h3d036c4b, 32'h3d649694} /* (21, 16, 12) {real, imag} */,
  {32'h3b491c70, 32'hbd8e7421} /* (21, 16, 11) {real, imag} */,
  {32'hbc60a30d, 32'h3d32c03a} /* (21, 16, 10) {real, imag} */,
  {32'hbd9c2c15, 32'hbd4f4668} /* (21, 16, 9) {real, imag} */,
  {32'hbcfec6bb, 32'hbe06d587} /* (21, 16, 8) {real, imag} */,
  {32'hbcf45928, 32'h3d226e04} /* (21, 16, 7) {real, imag} */,
  {32'h3de08d46, 32'hbd52cb64} /* (21, 16, 6) {real, imag} */,
  {32'hbea2e972, 32'hbd3ca48e} /* (21, 16, 5) {real, imag} */,
  {32'h3e9ba107, 32'h3d57bc85} /* (21, 16, 4) {real, imag} */,
  {32'hbdd02b58, 32'hbe0561a4} /* (21, 16, 3) {real, imag} */,
  {32'hbfbb78ba, 32'hbeb74fe6} /* (21, 16, 2) {real, imag} */,
  {32'h408df644, 32'h3ee09fb8} /* (21, 16, 1) {real, imag} */,
  {32'h403dd41c, 32'h00000000} /* (21, 16, 0) {real, imag} */,
  {32'h408c83f8, 32'hbedef6a3} /* (21, 15, 31) {real, imag} */,
  {32'hbfb8fafa, 32'h3ea2473a} /* (21, 15, 30) {real, imag} */,
  {32'hbe1a74d4, 32'h3de3fb40} /* (21, 15, 29) {real, imag} */,
  {32'h3e915360, 32'hbd0051c8} /* (21, 15, 28) {real, imag} */,
  {32'hbe8481ee, 32'h3ceb8d30} /* (21, 15, 27) {real, imag} */,
  {32'hbd2e7d67, 32'hbde1879b} /* (21, 15, 26) {real, imag} */,
  {32'h3ce3fcfb, 32'hbd9b54b6} /* (21, 15, 25) {real, imag} */,
  {32'hbd5628e0, 32'h3df842b7} /* (21, 15, 24) {real, imag} */,
  {32'h3d2dd25a, 32'h3d9bf45c} /* (21, 15, 23) {real, imag} */,
  {32'h3da2e3c8, 32'h3ca13da9} /* (21, 15, 22) {real, imag} */,
  {32'hbdec07c0, 32'h3d54a8e6} /* (21, 15, 21) {real, imag} */,
  {32'hbdb5ca42, 32'h3daea814} /* (21, 15, 20) {real, imag} */,
  {32'hbdb35130, 32'h3d4fc49a} /* (21, 15, 19) {real, imag} */,
  {32'h3d0a7559, 32'h3dcc45b6} /* (21, 15, 18) {real, imag} */,
  {32'h3d000267, 32'hbd95dcc8} /* (21, 15, 17) {real, imag} */,
  {32'hbdd04af9, 32'h00000000} /* (21, 15, 16) {real, imag} */,
  {32'h3d000267, 32'h3d95dcc8} /* (21, 15, 15) {real, imag} */,
  {32'h3d0a7559, 32'hbdcc45b6} /* (21, 15, 14) {real, imag} */,
  {32'hbdb35130, 32'hbd4fc49a} /* (21, 15, 13) {real, imag} */,
  {32'hbdb5ca42, 32'hbdaea814} /* (21, 15, 12) {real, imag} */,
  {32'hbdec07c0, 32'hbd54a8e6} /* (21, 15, 11) {real, imag} */,
  {32'h3da2e3c8, 32'hbca13da9} /* (21, 15, 10) {real, imag} */,
  {32'h3d2dd25a, 32'hbd9bf45c} /* (21, 15, 9) {real, imag} */,
  {32'hbd5628e0, 32'hbdf842b7} /* (21, 15, 8) {real, imag} */,
  {32'h3ce3fcfb, 32'h3d9b54b6} /* (21, 15, 7) {real, imag} */,
  {32'hbd2e7d67, 32'h3de1879b} /* (21, 15, 6) {real, imag} */,
  {32'hbe8481ee, 32'hbceb8d30} /* (21, 15, 5) {real, imag} */,
  {32'h3e915360, 32'h3d0051c8} /* (21, 15, 4) {real, imag} */,
  {32'hbe1a74d4, 32'hbde3fb40} /* (21, 15, 3) {real, imag} */,
  {32'hbfb8fafa, 32'hbea2473a} /* (21, 15, 2) {real, imag} */,
  {32'h408c83f8, 32'h3edef6a3} /* (21, 15, 1) {real, imag} */,
  {32'h40443f04, 32'h00000000} /* (21, 15, 0) {real, imag} */,
  {32'h4083eb43, 32'hbeafa7cc} /* (21, 14, 31) {real, imag} */,
  {32'hbfb2f544, 32'h3eadeee0} /* (21, 14, 30) {real, imag} */,
  {32'hbe21ba46, 32'hbd2a896a} /* (21, 14, 29) {real, imag} */,
  {32'h3e5f4beb, 32'hbdd06362} /* (21, 14, 28) {real, imag} */,
  {32'hbde9a825, 32'h3e43e649} /* (21, 14, 27) {real, imag} */,
  {32'hbdc3043b, 32'h3b5827c0} /* (21, 14, 26) {real, imag} */,
  {32'h3c9e2faf, 32'h3bfa0c10} /* (21, 14, 25) {real, imag} */,
  {32'hbd965bc0, 32'h3e41f98b} /* (21, 14, 24) {real, imag} */,
  {32'h3c6004fc, 32'h3df0d96b} /* (21, 14, 23) {real, imag} */,
  {32'hbd21516c, 32'h3d4e16ae} /* (21, 14, 22) {real, imag} */,
  {32'hbde57e93, 32'h3d710196} /* (21, 14, 21) {real, imag} */,
  {32'hbb6a7fa8, 32'hbd0751e3} /* (21, 14, 20) {real, imag} */,
  {32'hbb3f7e2c, 32'hbc2f7d2d} /* (21, 14, 19) {real, imag} */,
  {32'h3d34021d, 32'h3c0d37c6} /* (21, 14, 18) {real, imag} */,
  {32'hbd7a5239, 32'hbd33f338} /* (21, 14, 17) {real, imag} */,
  {32'hbc6a0abb, 32'h00000000} /* (21, 14, 16) {real, imag} */,
  {32'hbd7a5239, 32'h3d33f338} /* (21, 14, 15) {real, imag} */,
  {32'h3d34021d, 32'hbc0d37c6} /* (21, 14, 14) {real, imag} */,
  {32'hbb3f7e2c, 32'h3c2f7d2d} /* (21, 14, 13) {real, imag} */,
  {32'hbb6a7fa8, 32'h3d0751e3} /* (21, 14, 12) {real, imag} */,
  {32'hbde57e93, 32'hbd710196} /* (21, 14, 11) {real, imag} */,
  {32'hbd21516c, 32'hbd4e16ae} /* (21, 14, 10) {real, imag} */,
  {32'h3c6004fc, 32'hbdf0d96b} /* (21, 14, 9) {real, imag} */,
  {32'hbd965bc0, 32'hbe41f98b} /* (21, 14, 8) {real, imag} */,
  {32'h3c9e2faf, 32'hbbfa0c10} /* (21, 14, 7) {real, imag} */,
  {32'hbdc3043b, 32'hbb5827c0} /* (21, 14, 6) {real, imag} */,
  {32'hbde9a825, 32'hbe43e649} /* (21, 14, 5) {real, imag} */,
  {32'h3e5f4beb, 32'h3dd06362} /* (21, 14, 4) {real, imag} */,
  {32'hbe21ba46, 32'h3d2a896a} /* (21, 14, 3) {real, imag} */,
  {32'hbfb2f544, 32'hbeadeee0} /* (21, 14, 2) {real, imag} */,
  {32'h4083eb43, 32'h3eafa7cc} /* (21, 14, 1) {real, imag} */,
  {32'h403e096c, 32'h00000000} /* (21, 14, 0) {real, imag} */,
  {32'h405c4a74, 32'hbe2227f8} /* (21, 13, 31) {real, imag} */,
  {32'hbfacf42c, 32'h3e8c0d5c} /* (21, 13, 30) {real, imag} */,
  {32'hbdf49d88, 32'hbd6a8d1b} /* (21, 13, 29) {real, imag} */,
  {32'h3e93dace, 32'hbe1c67c2} /* (21, 13, 28) {real, imag} */,
  {32'hbe5b0e8d, 32'h3e8814bc} /* (21, 13, 27) {real, imag} */,
  {32'h3d9ceb22, 32'h3dce97e3} /* (21, 13, 26) {real, imag} */,
  {32'h3da80a24, 32'hbe101fde} /* (21, 13, 25) {real, imag} */,
  {32'hbcd4b408, 32'h3ded77d6} /* (21, 13, 24) {real, imag} */,
  {32'hbd2633e1, 32'h3e0002e2} /* (21, 13, 23) {real, imag} */,
  {32'hbd15d3d4, 32'h3dc3139c} /* (21, 13, 22) {real, imag} */,
  {32'hbc9a5efa, 32'h3ca72ea2} /* (21, 13, 21) {real, imag} */,
  {32'hbc8ad9d4, 32'h3c4bb518} /* (21, 13, 20) {real, imag} */,
  {32'h3dfba83d, 32'hbd47397a} /* (21, 13, 19) {real, imag} */,
  {32'hbdc88c52, 32'hbcb02a9e} /* (21, 13, 18) {real, imag} */,
  {32'hbd83d1a5, 32'h3d2a59da} /* (21, 13, 17) {real, imag} */,
  {32'h3dae0cdb, 32'h00000000} /* (21, 13, 16) {real, imag} */,
  {32'hbd83d1a5, 32'hbd2a59da} /* (21, 13, 15) {real, imag} */,
  {32'hbdc88c52, 32'h3cb02a9e} /* (21, 13, 14) {real, imag} */,
  {32'h3dfba83d, 32'h3d47397a} /* (21, 13, 13) {real, imag} */,
  {32'hbc8ad9d4, 32'hbc4bb518} /* (21, 13, 12) {real, imag} */,
  {32'hbc9a5efa, 32'hbca72ea2} /* (21, 13, 11) {real, imag} */,
  {32'hbd15d3d4, 32'hbdc3139c} /* (21, 13, 10) {real, imag} */,
  {32'hbd2633e1, 32'hbe0002e2} /* (21, 13, 9) {real, imag} */,
  {32'hbcd4b408, 32'hbded77d6} /* (21, 13, 8) {real, imag} */,
  {32'h3da80a24, 32'h3e101fde} /* (21, 13, 7) {real, imag} */,
  {32'h3d9ceb22, 32'hbdce97e3} /* (21, 13, 6) {real, imag} */,
  {32'hbe5b0e8d, 32'hbe8814bc} /* (21, 13, 5) {real, imag} */,
  {32'h3e93dace, 32'h3e1c67c2} /* (21, 13, 4) {real, imag} */,
  {32'hbdf49d88, 32'h3d6a8d1b} /* (21, 13, 3) {real, imag} */,
  {32'hbfacf42c, 32'hbe8c0d5c} /* (21, 13, 2) {real, imag} */,
  {32'h405c4a74, 32'h3e2227f8} /* (21, 13, 1) {real, imag} */,
  {32'h40212bfe, 32'h00000000} /* (21, 13, 0) {real, imag} */,
  {32'h4016322a, 32'h3dddfdf8} /* (21, 12, 31) {real, imag} */,
  {32'hbfa02b56, 32'h3e1a2562} /* (21, 12, 30) {real, imag} */,
  {32'h3d966f70, 32'hbcfd26f4} /* (21, 12, 29) {real, imag} */,
  {32'h3e7bee09, 32'hbdfd1eee} /* (21, 12, 28) {real, imag} */,
  {32'hbe8e3018, 32'h3dfcf446} /* (21, 12, 27) {real, imag} */,
  {32'h3e1ccc85, 32'h3d2329d4} /* (21, 12, 26) {real, imag} */,
  {32'h3de6fcb7, 32'hbd035440} /* (21, 12, 25) {real, imag} */,
  {32'h3cfbac76, 32'hbcd9a826} /* (21, 12, 24) {real, imag} */,
  {32'hbdb102a4, 32'h3d9fa958} /* (21, 12, 23) {real, imag} */,
  {32'h3d14dd68, 32'hbc4f9358} /* (21, 12, 22) {real, imag} */,
  {32'hbdfa336a, 32'h3e088000} /* (21, 12, 21) {real, imag} */,
  {32'hbd5588ae, 32'h3c0e395c} /* (21, 12, 20) {real, imag} */,
  {32'h3d8d1ebd, 32'hbc9b743a} /* (21, 12, 19) {real, imag} */,
  {32'hbd7c1500, 32'h3bd86350} /* (21, 12, 18) {real, imag} */,
  {32'h3bafac10, 32'hbcec5667} /* (21, 12, 17) {real, imag} */,
  {32'h3adc6ea0, 32'h00000000} /* (21, 12, 16) {real, imag} */,
  {32'h3bafac10, 32'h3cec5667} /* (21, 12, 15) {real, imag} */,
  {32'hbd7c1500, 32'hbbd86350} /* (21, 12, 14) {real, imag} */,
  {32'h3d8d1ebd, 32'h3c9b743a} /* (21, 12, 13) {real, imag} */,
  {32'hbd5588ae, 32'hbc0e395c} /* (21, 12, 12) {real, imag} */,
  {32'hbdfa336a, 32'hbe088000} /* (21, 12, 11) {real, imag} */,
  {32'h3d14dd68, 32'h3c4f9358} /* (21, 12, 10) {real, imag} */,
  {32'hbdb102a4, 32'hbd9fa958} /* (21, 12, 9) {real, imag} */,
  {32'h3cfbac76, 32'h3cd9a826} /* (21, 12, 8) {real, imag} */,
  {32'h3de6fcb7, 32'h3d035440} /* (21, 12, 7) {real, imag} */,
  {32'h3e1ccc85, 32'hbd2329d4} /* (21, 12, 6) {real, imag} */,
  {32'hbe8e3018, 32'hbdfcf446} /* (21, 12, 5) {real, imag} */,
  {32'h3e7bee09, 32'h3dfd1eee} /* (21, 12, 4) {real, imag} */,
  {32'h3d966f70, 32'h3cfd26f4} /* (21, 12, 3) {real, imag} */,
  {32'hbfa02b56, 32'hbe1a2562} /* (21, 12, 2) {real, imag} */,
  {32'h4016322a, 32'hbdddfdf8} /* (21, 12, 1) {real, imag} */,
  {32'h3fcfd0db, 32'h00000000} /* (21, 12, 0) {real, imag} */,
  {32'h3f8ba3c0, 32'h3ef2d3e4} /* (21, 11, 31) {real, imag} */,
  {32'hbf33bf26, 32'h3b69b680} /* (21, 11, 30) {real, imag} */,
  {32'h3d5e8b76, 32'hbd04a1ed} /* (21, 11, 29) {real, imag} */,
  {32'h3e38ae39, 32'hbde035a4} /* (21, 11, 28) {real, imag} */,
  {32'hbd85fc80, 32'hbd223be3} /* (21, 11, 27) {real, imag} */,
  {32'h3d8119ef, 32'h3d76e31a} /* (21, 11, 26) {real, imag} */,
  {32'h3d461438, 32'h3d29190a} /* (21, 11, 25) {real, imag} */,
  {32'hbe03770d, 32'h3d993211} /* (21, 11, 24) {real, imag} */,
  {32'h3b25939c, 32'h3ce7dcf8} /* (21, 11, 23) {real, imag} */,
  {32'h3d85166a, 32'hbd80bc29} /* (21, 11, 22) {real, imag} */,
  {32'hbe0da14e, 32'h3da3a9db} /* (21, 11, 21) {real, imag} */,
  {32'hbd8ebcff, 32'h3d1fed08} /* (21, 11, 20) {real, imag} */,
  {32'h3dba3854, 32'hbd457f95} /* (21, 11, 19) {real, imag} */,
  {32'hbd098e61, 32'hbcb9c84d} /* (21, 11, 18) {real, imag} */,
  {32'hbcb198b4, 32'h3cc901ca} /* (21, 11, 17) {real, imag} */,
  {32'h3d8ead12, 32'h00000000} /* (21, 11, 16) {real, imag} */,
  {32'hbcb198b4, 32'hbcc901ca} /* (21, 11, 15) {real, imag} */,
  {32'hbd098e61, 32'h3cb9c84d} /* (21, 11, 14) {real, imag} */,
  {32'h3dba3854, 32'h3d457f95} /* (21, 11, 13) {real, imag} */,
  {32'hbd8ebcff, 32'hbd1fed08} /* (21, 11, 12) {real, imag} */,
  {32'hbe0da14e, 32'hbda3a9db} /* (21, 11, 11) {real, imag} */,
  {32'h3d85166a, 32'h3d80bc29} /* (21, 11, 10) {real, imag} */,
  {32'h3b25939c, 32'hbce7dcf8} /* (21, 11, 9) {real, imag} */,
  {32'hbe03770d, 32'hbd993211} /* (21, 11, 8) {real, imag} */,
  {32'h3d461438, 32'hbd29190a} /* (21, 11, 7) {real, imag} */,
  {32'h3d8119ef, 32'hbd76e31a} /* (21, 11, 6) {real, imag} */,
  {32'hbd85fc80, 32'h3d223be3} /* (21, 11, 5) {real, imag} */,
  {32'h3e38ae39, 32'h3de035a4} /* (21, 11, 4) {real, imag} */,
  {32'h3d5e8b76, 32'h3d04a1ed} /* (21, 11, 3) {real, imag} */,
  {32'hbf33bf26, 32'hbb69b680} /* (21, 11, 2) {real, imag} */,
  {32'h3f8ba3c0, 32'hbef2d3e4} /* (21, 11, 1) {real, imag} */,
  {32'h3f598ba2, 32'h00000000} /* (21, 11, 0) {real, imag} */,
  {32'hbf2b7b08, 32'h3f4d888e} /* (21, 10, 31) {real, imag} */,
  {32'h3e1ac18c, 32'hbe2c0cbc} /* (21, 10, 30) {real, imag} */,
  {32'h3c1bddf2, 32'hbc95bea8} /* (21, 10, 29) {real, imag} */,
  {32'h3d79bf3c, 32'hbd7df095} /* (21, 10, 28) {real, imag} */,
  {32'h3dfc9e82, 32'hbd819b9c} /* (21, 10, 27) {real, imag} */,
  {32'hbd98eb1d, 32'h3ae612c0} /* (21, 10, 26) {real, imag} */,
  {32'hbe1de222, 32'h3dac6f1c} /* (21, 10, 25) {real, imag} */,
  {32'h3d368831, 32'hbd8e2060} /* (21, 10, 24) {real, imag} */,
  {32'hbd7f9a2e, 32'hbcc73b5f} /* (21, 10, 23) {real, imag} */,
  {32'hbc0ecce6, 32'h3cd0a34a} /* (21, 10, 22) {real, imag} */,
  {32'h3c7d7ad2, 32'hbdb93112} /* (21, 10, 21) {real, imag} */,
  {32'hbdb022cf, 32'hbd5d82f4} /* (21, 10, 20) {real, imag} */,
  {32'hbd17829e, 32'hbb4facf2} /* (21, 10, 19) {real, imag} */,
  {32'h3d14e448, 32'h3c225e50} /* (21, 10, 18) {real, imag} */,
  {32'h3ca74f9a, 32'hbcd7f507} /* (21, 10, 17) {real, imag} */,
  {32'h3e019d02, 32'h00000000} /* (21, 10, 16) {real, imag} */,
  {32'h3ca74f9a, 32'h3cd7f507} /* (21, 10, 15) {real, imag} */,
  {32'h3d14e448, 32'hbc225e50} /* (21, 10, 14) {real, imag} */,
  {32'hbd17829e, 32'h3b4facf2} /* (21, 10, 13) {real, imag} */,
  {32'hbdb022cf, 32'h3d5d82f4} /* (21, 10, 12) {real, imag} */,
  {32'h3c7d7ad2, 32'h3db93112} /* (21, 10, 11) {real, imag} */,
  {32'hbc0ecce6, 32'hbcd0a34a} /* (21, 10, 10) {real, imag} */,
  {32'hbd7f9a2e, 32'h3cc73b5f} /* (21, 10, 9) {real, imag} */,
  {32'h3d368831, 32'h3d8e2060} /* (21, 10, 8) {real, imag} */,
  {32'hbe1de222, 32'hbdac6f1c} /* (21, 10, 7) {real, imag} */,
  {32'hbd98eb1d, 32'hbae612c0} /* (21, 10, 6) {real, imag} */,
  {32'h3dfc9e82, 32'h3d819b9c} /* (21, 10, 5) {real, imag} */,
  {32'h3d79bf3c, 32'h3d7df095} /* (21, 10, 4) {real, imag} */,
  {32'h3c1bddf2, 32'h3c95bea8} /* (21, 10, 3) {real, imag} */,
  {32'h3e1ac18c, 32'h3e2c0cbc} /* (21, 10, 2) {real, imag} */,
  {32'hbf2b7b08, 32'hbf4d888e} /* (21, 10, 1) {real, imag} */,
  {32'hbf53598d, 32'h00000000} /* (21, 10, 0) {real, imag} */,
  {32'hc008dd34, 32'h3f829d78} /* (21, 9, 31) {real, imag} */,
  {32'h3f4794c2, 32'hbebe49e0} /* (21, 9, 30) {real, imag} */,
  {32'h3dd4b6a6, 32'hb9384740} /* (21, 9, 29) {real, imag} */,
  {32'h3a673000, 32'h3de0e58a} /* (21, 9, 28) {real, imag} */,
  {32'h3e1ad770, 32'hbd247cf3} /* (21, 9, 27) {real, imag} */,
  {32'h3d74c9d0, 32'hbd9a57e2} /* (21, 9, 26) {real, imag} */,
  {32'hbdaaf224, 32'h3deae69c} /* (21, 9, 25) {real, imag} */,
  {32'h3d9dd0a6, 32'hbdef4344} /* (21, 9, 24) {real, imag} */,
  {32'hbd8b1c76, 32'hbd5937cc} /* (21, 9, 23) {real, imag} */,
  {32'hbca02f1e, 32'h3d23d408} /* (21, 9, 22) {real, imag} */,
  {32'hbde1c88f, 32'hbd9bf294} /* (21, 9, 21) {real, imag} */,
  {32'h3b95a7ca, 32'h3d3926e4} /* (21, 9, 20) {real, imag} */,
  {32'h3d6bd6f8, 32'h3dad1369} /* (21, 9, 19) {real, imag} */,
  {32'h398284a0, 32'h3d0e2e12} /* (21, 9, 18) {real, imag} */,
  {32'hbd6161ca, 32'h3de6de0b} /* (21, 9, 17) {real, imag} */,
  {32'h3d1dc04a, 32'h00000000} /* (21, 9, 16) {real, imag} */,
  {32'hbd6161ca, 32'hbde6de0b} /* (21, 9, 15) {real, imag} */,
  {32'h398284a0, 32'hbd0e2e12} /* (21, 9, 14) {real, imag} */,
  {32'h3d6bd6f8, 32'hbdad1369} /* (21, 9, 13) {real, imag} */,
  {32'h3b95a7ca, 32'hbd3926e4} /* (21, 9, 12) {real, imag} */,
  {32'hbde1c88f, 32'h3d9bf294} /* (21, 9, 11) {real, imag} */,
  {32'hbca02f1e, 32'hbd23d408} /* (21, 9, 10) {real, imag} */,
  {32'hbd8b1c76, 32'h3d5937cc} /* (21, 9, 9) {real, imag} */,
  {32'h3d9dd0a6, 32'h3def4344} /* (21, 9, 8) {real, imag} */,
  {32'hbdaaf224, 32'hbdeae69c} /* (21, 9, 7) {real, imag} */,
  {32'h3d74c9d0, 32'h3d9a57e2} /* (21, 9, 6) {real, imag} */,
  {32'h3e1ad770, 32'h3d247cf3} /* (21, 9, 5) {real, imag} */,
  {32'h3a673000, 32'hbde0e58a} /* (21, 9, 4) {real, imag} */,
  {32'h3dd4b6a6, 32'h39384740} /* (21, 9, 3) {real, imag} */,
  {32'h3f4794c2, 32'h3ebe49e0} /* (21, 9, 2) {real, imag} */,
  {32'hc008dd34, 32'hbf829d78} /* (21, 9, 1) {real, imag} */,
  {32'hc0120600, 32'h00000000} /* (21, 9, 0) {real, imag} */,
  {32'hc043a334, 32'h3fc99c3f} /* (21, 8, 31) {real, imag} */,
  {32'h3f763c20, 32'hbedc0184} /* (21, 8, 30) {real, imag} */,
  {32'h39fc6f00, 32'hbc0ee248} /* (21, 8, 29) {real, imag} */,
  {32'h3bf9e030, 32'h3e0daf44} /* (21, 8, 28) {real, imag} */,
  {32'h3e53707c, 32'hbde0095a} /* (21, 8, 27) {real, imag} */,
  {32'h3d54343b, 32'hbd949cea} /* (21, 8, 26) {real, imag} */,
  {32'h3d5fd8a0, 32'h3d82cf5a} /* (21, 8, 25) {real, imag} */,
  {32'h3d785540, 32'hbe4315d6} /* (21, 8, 24) {real, imag} */,
  {32'h3d801cb0, 32'hbb31a840} /* (21, 8, 23) {real, imag} */,
  {32'hbcb7947c, 32'h3ddf2ecf} /* (21, 8, 22) {real, imag} */,
  {32'h3d530d72, 32'hbb8ab524} /* (21, 8, 21) {real, imag} */,
  {32'h3c9acc70, 32'h3d1ebf94} /* (21, 8, 20) {real, imag} */,
  {32'h3d3aa243, 32'hbcdfba44} /* (21, 8, 19) {real, imag} */,
  {32'hbcdf15ac, 32'hbd5c0b15} /* (21, 8, 18) {real, imag} */,
  {32'h3da1dc0c, 32'h3d36f1b5} /* (21, 8, 17) {real, imag} */,
  {32'hbd04586f, 32'h00000000} /* (21, 8, 16) {real, imag} */,
  {32'h3da1dc0c, 32'hbd36f1b5} /* (21, 8, 15) {real, imag} */,
  {32'hbcdf15ac, 32'h3d5c0b15} /* (21, 8, 14) {real, imag} */,
  {32'h3d3aa243, 32'h3cdfba44} /* (21, 8, 13) {real, imag} */,
  {32'h3c9acc70, 32'hbd1ebf94} /* (21, 8, 12) {real, imag} */,
  {32'h3d530d72, 32'h3b8ab524} /* (21, 8, 11) {real, imag} */,
  {32'hbcb7947c, 32'hbddf2ecf} /* (21, 8, 10) {real, imag} */,
  {32'h3d801cb0, 32'h3b31a840} /* (21, 8, 9) {real, imag} */,
  {32'h3d785540, 32'h3e4315d6} /* (21, 8, 8) {real, imag} */,
  {32'h3d5fd8a0, 32'hbd82cf5a} /* (21, 8, 7) {real, imag} */,
  {32'h3d54343b, 32'h3d949cea} /* (21, 8, 6) {real, imag} */,
  {32'h3e53707c, 32'h3de0095a} /* (21, 8, 5) {real, imag} */,
  {32'h3bf9e030, 32'hbe0daf44} /* (21, 8, 4) {real, imag} */,
  {32'h39fc6f00, 32'h3c0ee248} /* (21, 8, 3) {real, imag} */,
  {32'h3f763c20, 32'h3edc0184} /* (21, 8, 2) {real, imag} */,
  {32'hc043a334, 32'hbfc99c3f} /* (21, 8, 1) {real, imag} */,
  {32'hc04622dc, 32'h00000000} /* (21, 8, 0) {real, imag} */,
  {32'hc06d0d36, 32'h4001c2b2} /* (21, 7, 31) {real, imag} */,
  {32'h3f745fb4, 32'hbf0b5481} /* (21, 7, 30) {real, imag} */,
  {32'h3b9a4008, 32'hbd0d6621} /* (21, 7, 29) {real, imag} */,
  {32'hbc678d80, 32'h3d48b68a} /* (21, 7, 28) {real, imag} */,
  {32'h3e1adf34, 32'h3ce48fa4} /* (21, 7, 27) {real, imag} */,
  {32'h3ca429d7, 32'h3c7efe24} /* (21, 7, 26) {real, imag} */,
  {32'h3dd14ab7, 32'h3d35c01e} /* (21, 7, 25) {real, imag} */,
  {32'h3db60a26, 32'hbe238f41} /* (21, 7, 24) {real, imag} */,
  {32'hbbffc658, 32'hbd6d988c} /* (21, 7, 23) {real, imag} */,
  {32'h3d0ccb1f, 32'hbd2c27c0} /* (21, 7, 22) {real, imag} */,
  {32'h3c514f90, 32'h3c4425d4} /* (21, 7, 21) {real, imag} */,
  {32'hbc233b08, 32'h3ba3aa40} /* (21, 7, 20) {real, imag} */,
  {32'h3bd29acc, 32'h3d4b00a5} /* (21, 7, 19) {real, imag} */,
  {32'h3d78d97f, 32'h3d3958ce} /* (21, 7, 18) {real, imag} */,
  {32'hbd6e8f09, 32'h3c95a63c} /* (21, 7, 17) {real, imag} */,
  {32'h3dad2248, 32'h00000000} /* (21, 7, 16) {real, imag} */,
  {32'hbd6e8f09, 32'hbc95a63c} /* (21, 7, 15) {real, imag} */,
  {32'h3d78d97f, 32'hbd3958ce} /* (21, 7, 14) {real, imag} */,
  {32'h3bd29acc, 32'hbd4b00a5} /* (21, 7, 13) {real, imag} */,
  {32'hbc233b08, 32'hbba3aa40} /* (21, 7, 12) {real, imag} */,
  {32'h3c514f90, 32'hbc4425d4} /* (21, 7, 11) {real, imag} */,
  {32'h3d0ccb1f, 32'h3d2c27c0} /* (21, 7, 10) {real, imag} */,
  {32'hbbffc658, 32'h3d6d988c} /* (21, 7, 9) {real, imag} */,
  {32'h3db60a26, 32'h3e238f41} /* (21, 7, 8) {real, imag} */,
  {32'h3dd14ab7, 32'hbd35c01e} /* (21, 7, 7) {real, imag} */,
  {32'h3ca429d7, 32'hbc7efe24} /* (21, 7, 6) {real, imag} */,
  {32'h3e1adf34, 32'hbce48fa4} /* (21, 7, 5) {real, imag} */,
  {32'hbc678d80, 32'hbd48b68a} /* (21, 7, 4) {real, imag} */,
  {32'h3b9a4008, 32'h3d0d6621} /* (21, 7, 3) {real, imag} */,
  {32'h3f745fb4, 32'h3f0b5481} /* (21, 7, 2) {real, imag} */,
  {32'hc06d0d36, 32'hc001c2b2} /* (21, 7, 1) {real, imag} */,
  {32'hc07ca1ee, 32'h00000000} /* (21, 7, 0) {real, imag} */,
  {32'hc078d328, 32'h401b5521} /* (21, 6, 31) {real, imag} */,
  {32'h3f5fa9e1, 32'hbf3594bc} /* (21, 6, 30) {real, imag} */,
  {32'hbcb52e29, 32'hbd8b837f} /* (21, 6, 29) {real, imag} */,
  {32'hbca520f0, 32'hbe2fc0f2} /* (21, 6, 28) {real, imag} */,
  {32'h3e30a375, 32'hbd031fdc} /* (21, 6, 27) {real, imag} */,
  {32'hbda8de43, 32'h3adc24f0} /* (21, 6, 26) {real, imag} */,
  {32'h3ddf826b, 32'h3ccda744} /* (21, 6, 25) {real, imag} */,
  {32'h3c02546c, 32'hbd0e3cb0} /* (21, 6, 24) {real, imag} */,
  {32'h3d4159f2, 32'h3d4d5fca} /* (21, 6, 23) {real, imag} */,
  {32'h3d918206, 32'h3e0311e2} /* (21, 6, 22) {real, imag} */,
  {32'hbc6dc84c, 32'h3d94edf3} /* (21, 6, 21) {real, imag} */,
  {32'hbd3fc808, 32'hbdaf3426} /* (21, 6, 20) {real, imag} */,
  {32'hbc25c5f7, 32'h3be49cc4} /* (21, 6, 19) {real, imag} */,
  {32'h3c482ed0, 32'hbd7730a0} /* (21, 6, 18) {real, imag} */,
  {32'h3ccfc683, 32'h3dab5562} /* (21, 6, 17) {real, imag} */,
  {32'hbb7df608, 32'h00000000} /* (21, 6, 16) {real, imag} */,
  {32'h3ccfc683, 32'hbdab5562} /* (21, 6, 15) {real, imag} */,
  {32'h3c482ed0, 32'h3d7730a0} /* (21, 6, 14) {real, imag} */,
  {32'hbc25c5f7, 32'hbbe49cc4} /* (21, 6, 13) {real, imag} */,
  {32'hbd3fc808, 32'h3daf3426} /* (21, 6, 12) {real, imag} */,
  {32'hbc6dc84c, 32'hbd94edf3} /* (21, 6, 11) {real, imag} */,
  {32'h3d918206, 32'hbe0311e2} /* (21, 6, 10) {real, imag} */,
  {32'h3d4159f2, 32'hbd4d5fca} /* (21, 6, 9) {real, imag} */,
  {32'h3c02546c, 32'h3d0e3cb0} /* (21, 6, 8) {real, imag} */,
  {32'h3ddf826b, 32'hbccda744} /* (21, 6, 7) {real, imag} */,
  {32'hbda8de43, 32'hbadc24f0} /* (21, 6, 6) {real, imag} */,
  {32'h3e30a375, 32'h3d031fdc} /* (21, 6, 5) {real, imag} */,
  {32'hbca520f0, 32'h3e2fc0f2} /* (21, 6, 4) {real, imag} */,
  {32'hbcb52e29, 32'h3d8b837f} /* (21, 6, 3) {real, imag} */,
  {32'h3f5fa9e1, 32'h3f3594bc} /* (21, 6, 2) {real, imag} */,
  {32'hc078d328, 32'hc01b5521} /* (21, 6, 1) {real, imag} */,
  {32'hc089d7f9, 32'h00000000} /* (21, 6, 0) {real, imag} */,
  {32'hc073ca9b, 32'h40525d84} /* (21, 5, 31) {real, imag} */,
  {32'h3e8b6638, 32'hbf67149b} /* (21, 5, 30) {real, imag} */,
  {32'h3d824b19, 32'hbe0b0598} /* (21, 5, 29) {real, imag} */,
  {32'h3e4566fe, 32'hbe49954d} /* (21, 5, 28) {real, imag} */,
  {32'h3e364c48, 32'h3d5f2c92} /* (21, 5, 27) {real, imag} */,
  {32'hbe03d81d, 32'h3d83fd22} /* (21, 5, 26) {real, imag} */,
  {32'h3dbb7793, 32'h3d96d138} /* (21, 5, 25) {real, imag} */,
  {32'hbbcaf9f4, 32'hbdfa352e} /* (21, 5, 24) {real, imag} */,
  {32'h3d1dedf3, 32'h3cf64eb4} /* (21, 5, 23) {real, imag} */,
  {32'hbcad34d2, 32'h3c3f0654} /* (21, 5, 22) {real, imag} */,
  {32'hbdcc5b91, 32'hbd1d90f4} /* (21, 5, 21) {real, imag} */,
  {32'hbb67f3c0, 32'hbd9f186a} /* (21, 5, 20) {real, imag} */,
  {32'h3d13ef41, 32'h3cd04104} /* (21, 5, 19) {real, imag} */,
  {32'hbbde88b0, 32'hbc895cbc} /* (21, 5, 18) {real, imag} */,
  {32'hbc5bd6c5, 32'h3cd0599f} /* (21, 5, 17) {real, imag} */,
  {32'h3c19ec80, 32'h00000000} /* (21, 5, 16) {real, imag} */,
  {32'hbc5bd6c5, 32'hbcd0599f} /* (21, 5, 15) {real, imag} */,
  {32'hbbde88b0, 32'h3c895cbc} /* (21, 5, 14) {real, imag} */,
  {32'h3d13ef41, 32'hbcd04104} /* (21, 5, 13) {real, imag} */,
  {32'hbb67f3c0, 32'h3d9f186a} /* (21, 5, 12) {real, imag} */,
  {32'hbdcc5b91, 32'h3d1d90f4} /* (21, 5, 11) {real, imag} */,
  {32'hbcad34d2, 32'hbc3f0654} /* (21, 5, 10) {real, imag} */,
  {32'h3d1dedf3, 32'hbcf64eb4} /* (21, 5, 9) {real, imag} */,
  {32'hbbcaf9f4, 32'h3dfa352e} /* (21, 5, 8) {real, imag} */,
  {32'h3dbb7793, 32'hbd96d138} /* (21, 5, 7) {real, imag} */,
  {32'hbe03d81d, 32'hbd83fd22} /* (21, 5, 6) {real, imag} */,
  {32'h3e364c48, 32'hbd5f2c92} /* (21, 5, 5) {real, imag} */,
  {32'h3e4566fe, 32'h3e49954d} /* (21, 5, 4) {real, imag} */,
  {32'h3d824b19, 32'h3e0b0598} /* (21, 5, 3) {real, imag} */,
  {32'h3e8b6638, 32'h3f67149b} /* (21, 5, 2) {real, imag} */,
  {32'hc073ca9b, 32'hc0525d84} /* (21, 5, 1) {real, imag} */,
  {32'hc0955c8b, 32'h00000000} /* (21, 5, 0) {real, imag} */,
  {32'hc05f0c5c, 32'h40749b6d} /* (21, 4, 31) {real, imag} */,
  {32'hbdbec1c8, 32'hbf886e2d} /* (21, 4, 30) {real, imag} */,
  {32'h3decd48c, 32'hbe531bc0} /* (21, 4, 29) {real, imag} */,
  {32'h3dd633fa, 32'hbedddd09} /* (21, 4, 28) {real, imag} */,
  {32'h3dc1b2ac, 32'h3d76aac8} /* (21, 4, 27) {real, imag} */,
  {32'h3da65b7a, 32'h3d59af8d} /* (21, 4, 26) {real, imag} */,
  {32'h3ddbd7c6, 32'hbc597644} /* (21, 4, 25) {real, imag} */,
  {32'hbe214392, 32'h3ce45396} /* (21, 4, 24) {real, imag} */,
  {32'h3df71414, 32'hbd47701c} /* (21, 4, 23) {real, imag} */,
  {32'h3d503f89, 32'h3c985670} /* (21, 4, 22) {real, imag} */,
  {32'hbdb17c22, 32'h3cd954ba} /* (21, 4, 21) {real, imag} */,
  {32'hbdbfea43, 32'h3d9364b5} /* (21, 4, 20) {real, imag} */,
  {32'hbb99ccf8, 32'hbb443030} /* (21, 4, 19) {real, imag} */,
  {32'hbc4ce940, 32'hbb69a564} /* (21, 4, 18) {real, imag} */,
  {32'hbbccd8a0, 32'hbd0b26ba} /* (21, 4, 17) {real, imag} */,
  {32'hbca45942, 32'h00000000} /* (21, 4, 16) {real, imag} */,
  {32'hbbccd8a0, 32'h3d0b26ba} /* (21, 4, 15) {real, imag} */,
  {32'hbc4ce940, 32'h3b69a564} /* (21, 4, 14) {real, imag} */,
  {32'hbb99ccf8, 32'h3b443030} /* (21, 4, 13) {real, imag} */,
  {32'hbdbfea43, 32'hbd9364b5} /* (21, 4, 12) {real, imag} */,
  {32'hbdb17c22, 32'hbcd954ba} /* (21, 4, 11) {real, imag} */,
  {32'h3d503f89, 32'hbc985670} /* (21, 4, 10) {real, imag} */,
  {32'h3df71414, 32'h3d47701c} /* (21, 4, 9) {real, imag} */,
  {32'hbe214392, 32'hbce45396} /* (21, 4, 8) {real, imag} */,
  {32'h3ddbd7c6, 32'h3c597644} /* (21, 4, 7) {real, imag} */,
  {32'h3da65b7a, 32'hbd59af8d} /* (21, 4, 6) {real, imag} */,
  {32'h3dc1b2ac, 32'hbd76aac8} /* (21, 4, 5) {real, imag} */,
  {32'h3dd633fa, 32'h3edddd09} /* (21, 4, 4) {real, imag} */,
  {32'h3decd48c, 32'h3e531bc0} /* (21, 4, 3) {real, imag} */,
  {32'hbdbec1c8, 32'h3f886e2d} /* (21, 4, 2) {real, imag} */,
  {32'hc05f0c5c, 32'hc0749b6d} /* (21, 4, 1) {real, imag} */,
  {32'hc0a4c735, 32'h00000000} /* (21, 4, 0) {real, imag} */,
  {32'hc05f470e, 32'h4080f8e8} /* (21, 3, 31) {real, imag} */,
  {32'hbea63174, 32'hbf81e7fa} /* (21, 3, 30) {real, imag} */,
  {32'h3c111498, 32'hbdc12c13} /* (21, 3, 29) {real, imag} */,
  {32'h3d98c176, 32'hbecba501} /* (21, 3, 28) {real, imag} */,
  {32'h3ea12b3e, 32'h3df8958c} /* (21, 3, 27) {real, imag} */,
  {32'h3c9e9359, 32'hbd8368e8} /* (21, 3, 26) {real, imag} */,
  {32'h3c29f10b, 32'h3d6e7201} /* (21, 3, 25) {real, imag} */,
  {32'hbcbc0ecb, 32'hbdbc427e} /* (21, 3, 24) {real, imag} */,
  {32'h3e0c2208, 32'h3d1a998d} /* (21, 3, 23) {real, imag} */,
  {32'h3d92ddd3, 32'hbce18a78} /* (21, 3, 22) {real, imag} */,
  {32'h3cf4ee34, 32'hbcdaf740} /* (21, 3, 21) {real, imag} */,
  {32'hbd552e86, 32'hbde865fd} /* (21, 3, 20) {real, imag} */,
  {32'h3c465026, 32'hbd5b95e3} /* (21, 3, 19) {real, imag} */,
  {32'h3d83e030, 32'hbdbdf4e4} /* (21, 3, 18) {real, imag} */,
  {32'h3c0bf682, 32'h3c704dcc} /* (21, 3, 17) {real, imag} */,
  {32'h3c982cbb, 32'h00000000} /* (21, 3, 16) {real, imag} */,
  {32'h3c0bf682, 32'hbc704dcc} /* (21, 3, 15) {real, imag} */,
  {32'h3d83e030, 32'h3dbdf4e4} /* (21, 3, 14) {real, imag} */,
  {32'h3c465026, 32'h3d5b95e3} /* (21, 3, 13) {real, imag} */,
  {32'hbd552e86, 32'h3de865fd} /* (21, 3, 12) {real, imag} */,
  {32'h3cf4ee34, 32'h3cdaf740} /* (21, 3, 11) {real, imag} */,
  {32'h3d92ddd3, 32'h3ce18a78} /* (21, 3, 10) {real, imag} */,
  {32'h3e0c2208, 32'hbd1a998d} /* (21, 3, 9) {real, imag} */,
  {32'hbcbc0ecb, 32'h3dbc427e} /* (21, 3, 8) {real, imag} */,
  {32'h3c29f10b, 32'hbd6e7201} /* (21, 3, 7) {real, imag} */,
  {32'h3c9e9359, 32'h3d8368e8} /* (21, 3, 6) {real, imag} */,
  {32'h3ea12b3e, 32'hbdf8958c} /* (21, 3, 5) {real, imag} */,
  {32'h3d98c176, 32'h3ecba501} /* (21, 3, 4) {real, imag} */,
  {32'h3c111498, 32'h3dc12c13} /* (21, 3, 3) {real, imag} */,
  {32'hbea63174, 32'h3f81e7fa} /* (21, 3, 2) {real, imag} */,
  {32'hc05f470e, 32'hc080f8e8} /* (21, 3, 1) {real, imag} */,
  {32'hc0ae27c6, 32'h00000000} /* (21, 3, 0) {real, imag} */,
  {32'hc05ea37c, 32'h407a541a} /* (21, 2, 31) {real, imag} */,
  {32'hbe8a4e0a, 32'hbf75b01e} /* (21, 2, 30) {real, imag} */,
  {32'h3c816884, 32'hbe293158} /* (21, 2, 29) {real, imag} */,
  {32'h3ddc4a03, 32'hbe8a40c2} /* (21, 2, 28) {real, imag} */,
  {32'h3e67f41b, 32'h3d67951a} /* (21, 2, 27) {real, imag} */,
  {32'h3d029a62, 32'hbc7b0748} /* (21, 2, 26) {real, imag} */,
  {32'h3dc854f8, 32'hbc3c4cfe} /* (21, 2, 25) {real, imag} */,
  {32'hbce923cb, 32'hbd83b4fa} /* (21, 2, 24) {real, imag} */,
  {32'h3ca0c256, 32'hbd7d0c4e} /* (21, 2, 23) {real, imag} */,
  {32'h3d7d5037, 32'hbc13b800} /* (21, 2, 22) {real, imag} */,
  {32'h3dc3083e, 32'hbd1d0d67} /* (21, 2, 21) {real, imag} */,
  {32'h3d10c77c, 32'h3cac7390} /* (21, 2, 20) {real, imag} */,
  {32'h3d706eba, 32'h3ca63322} /* (21, 2, 19) {real, imag} */,
  {32'hbc84f474, 32'h3be22bbc} /* (21, 2, 18) {real, imag} */,
  {32'hbc5ed70c, 32'h3d828ea9} /* (21, 2, 17) {real, imag} */,
  {32'h3988f600, 32'h00000000} /* (21, 2, 16) {real, imag} */,
  {32'hbc5ed70c, 32'hbd828ea9} /* (21, 2, 15) {real, imag} */,
  {32'hbc84f474, 32'hbbe22bbc} /* (21, 2, 14) {real, imag} */,
  {32'h3d706eba, 32'hbca63322} /* (21, 2, 13) {real, imag} */,
  {32'h3d10c77c, 32'hbcac7390} /* (21, 2, 12) {real, imag} */,
  {32'h3dc3083e, 32'h3d1d0d67} /* (21, 2, 11) {real, imag} */,
  {32'h3d7d5037, 32'h3c13b800} /* (21, 2, 10) {real, imag} */,
  {32'h3ca0c256, 32'h3d7d0c4e} /* (21, 2, 9) {real, imag} */,
  {32'hbce923cb, 32'h3d83b4fa} /* (21, 2, 8) {real, imag} */,
  {32'h3dc854f8, 32'h3c3c4cfe} /* (21, 2, 7) {real, imag} */,
  {32'h3d029a62, 32'h3c7b0748} /* (21, 2, 6) {real, imag} */,
  {32'h3e67f41b, 32'hbd67951a} /* (21, 2, 5) {real, imag} */,
  {32'h3ddc4a03, 32'h3e8a40c2} /* (21, 2, 4) {real, imag} */,
  {32'h3c816884, 32'h3e293158} /* (21, 2, 3) {real, imag} */,
  {32'hbe8a4e0a, 32'h3f75b01e} /* (21, 2, 2) {real, imag} */,
  {32'hc05ea37c, 32'hc07a541a} /* (21, 2, 1) {real, imag} */,
  {32'hc0ae2d8e, 32'h00000000} /* (21, 2, 0) {real, imag} */,
  {32'hc0631050, 32'h406ec5da} /* (21, 1, 31) {real, imag} */,
  {32'h3bc79180, 32'hbf70b41f} /* (21, 1, 30) {real, imag} */,
  {32'h3e1a3542, 32'hbe0163f5} /* (21, 1, 29) {real, imag} */,
  {32'h3dde13e9, 32'hbe693a30} /* (21, 1, 28) {real, imag} */,
  {32'h3e80d744, 32'hbd51db61} /* (21, 1, 27) {real, imag} */,
  {32'h3d91a8c3, 32'hbd8aa9d3} /* (21, 1, 26) {real, imag} */,
  {32'h3dbca11f, 32'h3c686b7c} /* (21, 1, 25) {real, imag} */,
  {32'hbd8d2ba7, 32'h3d42a8fe} /* (21, 1, 24) {real, imag} */,
  {32'h3d1d879a, 32'hbcd209b6} /* (21, 1, 23) {real, imag} */,
  {32'hbb368e0e, 32'hbd3db598} /* (21, 1, 22) {real, imag} */,
  {32'h3cb2f558, 32'h3d4228da} /* (21, 1, 21) {real, imag} */,
  {32'hbcf7480f, 32'h3dca7983} /* (21, 1, 20) {real, imag} */,
  {32'h3cbdfc3b, 32'h3c8b346e} /* (21, 1, 19) {real, imag} */,
  {32'hbd9d6379, 32'h3d86f9a4} /* (21, 1, 18) {real, imag} */,
  {32'h3caa645e, 32'hbd2c72fa} /* (21, 1, 17) {real, imag} */,
  {32'h3da78712, 32'h00000000} /* (21, 1, 16) {real, imag} */,
  {32'h3caa645e, 32'h3d2c72fa} /* (21, 1, 15) {real, imag} */,
  {32'hbd9d6379, 32'hbd86f9a4} /* (21, 1, 14) {real, imag} */,
  {32'h3cbdfc3b, 32'hbc8b346e} /* (21, 1, 13) {real, imag} */,
  {32'hbcf7480f, 32'hbdca7983} /* (21, 1, 12) {real, imag} */,
  {32'h3cb2f558, 32'hbd4228da} /* (21, 1, 11) {real, imag} */,
  {32'hbb368e0e, 32'h3d3db598} /* (21, 1, 10) {real, imag} */,
  {32'h3d1d879a, 32'h3cd209b6} /* (21, 1, 9) {real, imag} */,
  {32'hbd8d2ba7, 32'hbd42a8fe} /* (21, 1, 8) {real, imag} */,
  {32'h3dbca11f, 32'hbc686b7c} /* (21, 1, 7) {real, imag} */,
  {32'h3d91a8c3, 32'h3d8aa9d3} /* (21, 1, 6) {real, imag} */,
  {32'h3e80d744, 32'h3d51db61} /* (21, 1, 5) {real, imag} */,
  {32'h3dde13e9, 32'h3e693a30} /* (21, 1, 4) {real, imag} */,
  {32'h3e1a3542, 32'h3e0163f5} /* (21, 1, 3) {real, imag} */,
  {32'h3bc79180, 32'h3f70b41f} /* (21, 1, 2) {real, imag} */,
  {32'hc0631050, 32'hc06ec5da} /* (21, 1, 1) {real, imag} */,
  {32'hc0b1b29b, 32'h00000000} /* (21, 1, 0) {real, imag} */,
  {32'hc06c4589, 32'h4045a4e8} /* (21, 0, 31) {real, imag} */,
  {32'h3e80d046, 32'hbf430249} /* (21, 0, 30) {real, imag} */,
  {32'h3e619e64, 32'h3c9b2a64} /* (21, 0, 29) {real, imag} */,
  {32'hbc8babf0, 32'hbe2716b9} /* (21, 0, 28) {real, imag} */,
  {32'h3da63412, 32'hbce3c34c} /* (21, 0, 27) {real, imag} */,
  {32'hbd745329, 32'hbcdc03bc} /* (21, 0, 26) {real, imag} */,
  {32'hbcaa5fd4, 32'h3daf723a} /* (21, 0, 25) {real, imag} */,
  {32'hbcc182df, 32'h3aee5680} /* (21, 0, 24) {real, imag} */,
  {32'h3d89386d, 32'hbba366ac} /* (21, 0, 23) {real, imag} */,
  {32'h3c7a010b, 32'hbe1d13b6} /* (21, 0, 22) {real, imag} */,
  {32'hbd144a57, 32'h3d722322} /* (21, 0, 21) {real, imag} */,
  {32'h3d3f9fc9, 32'hbd7f0f22} /* (21, 0, 20) {real, imag} */,
  {32'hbc3b46ba, 32'h3cd0075f} /* (21, 0, 19) {real, imag} */,
  {32'h3d16714d, 32'h3bfb7bd0} /* (21, 0, 18) {real, imag} */,
  {32'h3ccc1b98, 32'h3caf4617} /* (21, 0, 17) {real, imag} */,
  {32'hbd80305f, 32'h00000000} /* (21, 0, 16) {real, imag} */,
  {32'h3ccc1b98, 32'hbcaf4617} /* (21, 0, 15) {real, imag} */,
  {32'h3d16714d, 32'hbbfb7bd0} /* (21, 0, 14) {real, imag} */,
  {32'hbc3b46ba, 32'hbcd0075f} /* (21, 0, 13) {real, imag} */,
  {32'h3d3f9fc9, 32'h3d7f0f22} /* (21, 0, 12) {real, imag} */,
  {32'hbd144a57, 32'hbd722322} /* (21, 0, 11) {real, imag} */,
  {32'h3c7a010b, 32'h3e1d13b6} /* (21, 0, 10) {real, imag} */,
  {32'h3d89386d, 32'h3ba366ac} /* (21, 0, 9) {real, imag} */,
  {32'hbcc182df, 32'hbaee5680} /* (21, 0, 8) {real, imag} */,
  {32'hbcaa5fd4, 32'hbdaf723a} /* (21, 0, 7) {real, imag} */,
  {32'hbd745329, 32'h3cdc03bc} /* (21, 0, 6) {real, imag} */,
  {32'h3da63412, 32'h3ce3c34c} /* (21, 0, 5) {real, imag} */,
  {32'hbc8babf0, 32'h3e2716b9} /* (21, 0, 4) {real, imag} */,
  {32'h3e619e64, 32'hbc9b2a64} /* (21, 0, 3) {real, imag} */,
  {32'h3e80d046, 32'h3f430249} /* (21, 0, 2) {real, imag} */,
  {32'hc06c4589, 32'hc045a4e8} /* (21, 0, 1) {real, imag} */,
  {32'hc0aa0cf8, 32'h00000000} /* (21, 0, 0) {real, imag} */,
  {32'hc081f7a3, 32'h400f1b06} /* (20, 31, 31) {real, imag} */,
  {32'h3f49e391, 32'hbf0f5c30} /* (20, 31, 30) {real, imag} */,
  {32'h3d91581d, 32'hbd15fb03} /* (20, 31, 29) {real, imag} */,
  {32'hbd91a406, 32'h3c42bbc0} /* (20, 31, 28) {real, imag} */,
  {32'h3da225ba, 32'h3cbaf6c8} /* (20, 31, 27) {real, imag} */,
  {32'hbc84ed28, 32'h3c98626b} /* (20, 31, 26) {real, imag} */,
  {32'h3bed9738, 32'h3d116b0a} /* (20, 31, 25) {real, imag} */,
  {32'h3c957de6, 32'hbcbb7f6c} /* (20, 31, 24) {real, imag} */,
  {32'hbaa4f400, 32'hbda12106} /* (20, 31, 23) {real, imag} */,
  {32'h3d496a91, 32'h3932ea00} /* (20, 31, 22) {real, imag} */,
  {32'hbc032df8, 32'h3d909272} /* (20, 31, 21) {real, imag} */,
  {32'h3d06063e, 32'h3cb81177} /* (20, 31, 20) {real, imag} */,
  {32'hbc5c13c4, 32'hbcb2fe69} /* (20, 31, 19) {real, imag} */,
  {32'h3ba36522, 32'hbd150e8a} /* (20, 31, 18) {real, imag} */,
  {32'hbc8ffed4, 32'hbad03a00} /* (20, 31, 17) {real, imag} */,
  {32'h39f47040, 32'h00000000} /* (20, 31, 16) {real, imag} */,
  {32'hbc8ffed4, 32'h3ad03a00} /* (20, 31, 15) {real, imag} */,
  {32'h3ba36522, 32'h3d150e8a} /* (20, 31, 14) {real, imag} */,
  {32'hbc5c13c4, 32'h3cb2fe69} /* (20, 31, 13) {real, imag} */,
  {32'h3d06063e, 32'hbcb81177} /* (20, 31, 12) {real, imag} */,
  {32'hbc032df8, 32'hbd909272} /* (20, 31, 11) {real, imag} */,
  {32'h3d496a91, 32'hb932ea00} /* (20, 31, 10) {real, imag} */,
  {32'hbaa4f400, 32'h3da12106} /* (20, 31, 9) {real, imag} */,
  {32'h3c957de6, 32'h3cbb7f6c} /* (20, 31, 8) {real, imag} */,
  {32'h3bed9738, 32'hbd116b0a} /* (20, 31, 7) {real, imag} */,
  {32'hbc84ed28, 32'hbc98626b} /* (20, 31, 6) {real, imag} */,
  {32'h3da225ba, 32'hbcbaf6c8} /* (20, 31, 5) {real, imag} */,
  {32'hbd91a406, 32'hbc42bbc0} /* (20, 31, 4) {real, imag} */,
  {32'h3d91581d, 32'h3d15fb03} /* (20, 31, 3) {real, imag} */,
  {32'h3f49e391, 32'h3f0f5c30} /* (20, 31, 2) {real, imag} */,
  {32'hc081f7a3, 32'hc00f1b06} /* (20, 31, 1) {real, imag} */,
  {32'hc0a31735, 32'h00000000} /* (20, 31, 0) {real, imag} */,
  {32'hc09923b2, 32'h3fefb914} /* (20, 30, 31) {real, imag} */,
  {32'h3fab1562, 32'hbee4ea26} /* (20, 30, 30) {real, imag} */,
  {32'h3b707e90, 32'hbd202925} /* (20, 30, 29) {real, imag} */,
  {32'hbd200f71, 32'h3e060458} /* (20, 30, 28) {real, imag} */,
  {32'h3e326358, 32'h3a21cc70} /* (20, 30, 27) {real, imag} */,
  {32'hbc379acc, 32'hbd15f178} /* (20, 30, 26) {real, imag} */,
  {32'hbb623a80, 32'h3b294fd8} /* (20, 30, 25) {real, imag} */,
  {32'hbd3b8f22, 32'hbc54ed2a} /* (20, 30, 24) {real, imag} */,
  {32'hbd072a2c, 32'h3d98ae31} /* (20, 30, 23) {real, imag} */,
  {32'h3d2d5c4f, 32'hbc314160} /* (20, 30, 22) {real, imag} */,
  {32'h3d4cea78, 32'hbc45b672} /* (20, 30, 21) {real, imag} */,
  {32'h3be24e88, 32'hbd19581a} /* (20, 30, 20) {real, imag} */,
  {32'hbdb5e9c8, 32'hbcdb51d3} /* (20, 30, 19) {real, imag} */,
  {32'h3da87a94, 32'hbd5f1b52} /* (20, 30, 18) {real, imag} */,
  {32'hbd15b250, 32'h3d540760} /* (20, 30, 17) {real, imag} */,
  {32'h3d7bd52e, 32'h00000000} /* (20, 30, 16) {real, imag} */,
  {32'hbd15b250, 32'hbd540760} /* (20, 30, 15) {real, imag} */,
  {32'h3da87a94, 32'h3d5f1b52} /* (20, 30, 14) {real, imag} */,
  {32'hbdb5e9c8, 32'h3cdb51d3} /* (20, 30, 13) {real, imag} */,
  {32'h3be24e88, 32'h3d19581a} /* (20, 30, 12) {real, imag} */,
  {32'h3d4cea78, 32'h3c45b672} /* (20, 30, 11) {real, imag} */,
  {32'h3d2d5c4f, 32'h3c314160} /* (20, 30, 10) {real, imag} */,
  {32'hbd072a2c, 32'hbd98ae31} /* (20, 30, 9) {real, imag} */,
  {32'hbd3b8f22, 32'h3c54ed2a} /* (20, 30, 8) {real, imag} */,
  {32'hbb623a80, 32'hbb294fd8} /* (20, 30, 7) {real, imag} */,
  {32'hbc379acc, 32'h3d15f178} /* (20, 30, 6) {real, imag} */,
  {32'h3e326358, 32'hba21cc70} /* (20, 30, 5) {real, imag} */,
  {32'hbd200f71, 32'hbe060458} /* (20, 30, 4) {real, imag} */,
  {32'h3b707e90, 32'h3d202925} /* (20, 30, 3) {real, imag} */,
  {32'h3fab1562, 32'h3ee4ea26} /* (20, 30, 2) {real, imag} */,
  {32'hc09923b2, 32'hbfefb914} /* (20, 30, 1) {real, imag} */,
  {32'hc0a79342, 32'h00000000} /* (20, 30, 0) {real, imag} */,
  {32'hc09f4b31, 32'h3fd4e3ea} /* (20, 29, 31) {real, imag} */,
  {32'h3fbf427a, 32'hbeaf812b} /* (20, 29, 30) {real, imag} */,
  {32'h3d0e71ed, 32'hbd60ea7a} /* (20, 29, 29) {real, imag} */,
  {32'hbe96abaa, 32'h3dbb02e2} /* (20, 29, 28) {real, imag} */,
  {32'h3dcea7ad, 32'hbd4bd0af} /* (20, 29, 27) {real, imag} */,
  {32'hbca5ec60, 32'hbd2b4360} /* (20, 29, 26) {real, imag} */,
  {32'h3ca4d43b, 32'h3d9b2905} /* (20, 29, 25) {real, imag} */,
  {32'h3d7293f4, 32'h3c20e7d4} /* (20, 29, 24) {real, imag} */,
  {32'hbd2640d5, 32'hbd825a2e} /* (20, 29, 23) {real, imag} */,
  {32'hbd71a449, 32'h3dbe698c} /* (20, 29, 22) {real, imag} */,
  {32'h3d029790, 32'hbdad5b07} /* (20, 29, 21) {real, imag} */,
  {32'h3c40c880, 32'hbd3ca56e} /* (20, 29, 20) {real, imag} */,
  {32'h3b4cfeec, 32'h3cde577c} /* (20, 29, 19) {real, imag} */,
  {32'h3c321158, 32'h3c384f70} /* (20, 29, 18) {real, imag} */,
  {32'h3bd381c0, 32'hbc118934} /* (20, 29, 17) {real, imag} */,
  {32'hbda849e8, 32'h00000000} /* (20, 29, 16) {real, imag} */,
  {32'h3bd381c0, 32'h3c118934} /* (20, 29, 15) {real, imag} */,
  {32'h3c321158, 32'hbc384f70} /* (20, 29, 14) {real, imag} */,
  {32'h3b4cfeec, 32'hbcde577c} /* (20, 29, 13) {real, imag} */,
  {32'h3c40c880, 32'h3d3ca56e} /* (20, 29, 12) {real, imag} */,
  {32'h3d029790, 32'h3dad5b07} /* (20, 29, 11) {real, imag} */,
  {32'hbd71a449, 32'hbdbe698c} /* (20, 29, 10) {real, imag} */,
  {32'hbd2640d5, 32'h3d825a2e} /* (20, 29, 9) {real, imag} */,
  {32'h3d7293f4, 32'hbc20e7d4} /* (20, 29, 8) {real, imag} */,
  {32'h3ca4d43b, 32'hbd9b2905} /* (20, 29, 7) {real, imag} */,
  {32'hbca5ec60, 32'h3d2b4360} /* (20, 29, 6) {real, imag} */,
  {32'h3dcea7ad, 32'h3d4bd0af} /* (20, 29, 5) {real, imag} */,
  {32'hbe96abaa, 32'hbdbb02e2} /* (20, 29, 4) {real, imag} */,
  {32'h3d0e71ed, 32'h3d60ea7a} /* (20, 29, 3) {real, imag} */,
  {32'h3fbf427a, 32'h3eaf812b} /* (20, 29, 2) {real, imag} */,
  {32'hc09f4b31, 32'hbfd4e3ea} /* (20, 29, 1) {real, imag} */,
  {32'hc0a6bc94, 32'h00000000} /* (20, 29, 0) {real, imag} */,
  {32'hc0a3a2ea, 32'h3fb5e290} /* (20, 28, 31) {real, imag} */,
  {32'h3fde483e, 32'hbefcf94b} /* (20, 28, 30) {real, imag} */,
  {32'h3cc7de02, 32'hbd471878} /* (20, 28, 29) {real, imag} */,
  {32'hbeb3607f, 32'h3de1957f} /* (20, 28, 28) {real, imag} */,
  {32'h3d99e8aa, 32'hbd90c1e6} /* (20, 28, 27) {real, imag} */,
  {32'h3dc93618, 32'hbd1d05fb} /* (20, 28, 26) {real, imag} */,
  {32'hbe0699b5, 32'h3d6e2428} /* (20, 28, 25) {real, imag} */,
  {32'hbd45c037, 32'hbddcdb7a} /* (20, 28, 24) {real, imag} */,
  {32'hbcf2690c, 32'hbd3b7d0f} /* (20, 28, 23) {real, imag} */,
  {32'h3c1bf9c2, 32'hbc83dd6a} /* (20, 28, 22) {real, imag} */,
  {32'h3dc2f60d, 32'h3d02298a} /* (20, 28, 21) {real, imag} */,
  {32'hbc0ac2f1, 32'hbd1f0e84} /* (20, 28, 20) {real, imag} */,
  {32'h3d07051b, 32'hbcd70c3c} /* (20, 28, 19) {real, imag} */,
  {32'h3b9b72e8, 32'h3a0d20f0} /* (20, 28, 18) {real, imag} */,
  {32'hbcb3bf93, 32'hbac189e0} /* (20, 28, 17) {real, imag} */,
  {32'hbd87ca1d, 32'h00000000} /* (20, 28, 16) {real, imag} */,
  {32'hbcb3bf93, 32'h3ac189e0} /* (20, 28, 15) {real, imag} */,
  {32'h3b9b72e8, 32'hba0d20f0} /* (20, 28, 14) {real, imag} */,
  {32'h3d07051b, 32'h3cd70c3c} /* (20, 28, 13) {real, imag} */,
  {32'hbc0ac2f1, 32'h3d1f0e84} /* (20, 28, 12) {real, imag} */,
  {32'h3dc2f60d, 32'hbd02298a} /* (20, 28, 11) {real, imag} */,
  {32'h3c1bf9c2, 32'h3c83dd6a} /* (20, 28, 10) {real, imag} */,
  {32'hbcf2690c, 32'h3d3b7d0f} /* (20, 28, 9) {real, imag} */,
  {32'hbd45c037, 32'h3ddcdb7a} /* (20, 28, 8) {real, imag} */,
  {32'hbe0699b5, 32'hbd6e2428} /* (20, 28, 7) {real, imag} */,
  {32'h3dc93618, 32'h3d1d05fb} /* (20, 28, 6) {real, imag} */,
  {32'h3d99e8aa, 32'h3d90c1e6} /* (20, 28, 5) {real, imag} */,
  {32'hbeb3607f, 32'hbde1957f} /* (20, 28, 4) {real, imag} */,
  {32'h3cc7de02, 32'h3d471878} /* (20, 28, 3) {real, imag} */,
  {32'h3fde483e, 32'h3efcf94b} /* (20, 28, 2) {real, imag} */,
  {32'hc0a3a2ea, 32'hbfb5e290} /* (20, 28, 1) {real, imag} */,
  {32'hc0ab9dbe, 32'h00000000} /* (20, 28, 0) {real, imag} */,
  {32'hc0a6a3a9, 32'h3f8ee9a7} /* (20, 27, 31) {real, imag} */,
  {32'h3fe47f0d, 32'hbf034d18} /* (20, 27, 30) {real, imag} */,
  {32'h3d05dc80, 32'h3d4fe343} /* (20, 27, 29) {real, imag} */,
  {32'hbe464c3a, 32'h3ddae1c7} /* (20, 27, 28) {real, imag} */,
  {32'h3e52cc03, 32'hbd62975f} /* (20, 27, 27) {real, imag} */,
  {32'h3dc6ab37, 32'hbd9c27b2} /* (20, 27, 26) {real, imag} */,
  {32'hbdeb9638, 32'hbdd2b0da} /* (20, 27, 25) {real, imag} */,
  {32'hbd127d0c, 32'hbd25296a} /* (20, 27, 24) {real, imag} */,
  {32'h3dc9fc74, 32'h3db3c946} /* (20, 27, 23) {real, imag} */,
  {32'h3dc3fe4c, 32'h3c4caad4} /* (20, 27, 22) {real, imag} */,
  {32'hbc4c27d4, 32'hbcbdadf4} /* (20, 27, 21) {real, imag} */,
  {32'h3b9e9908, 32'h3d69cb3e} /* (20, 27, 20) {real, imag} */,
  {32'h3d2faee0, 32'h3c309b9e} /* (20, 27, 19) {real, imag} */,
  {32'hbccab958, 32'hbd28c4be} /* (20, 27, 18) {real, imag} */,
  {32'hbb11bfe0, 32'hbca8417c} /* (20, 27, 17) {real, imag} */,
  {32'h3c5d43b0, 32'h00000000} /* (20, 27, 16) {real, imag} */,
  {32'hbb11bfe0, 32'h3ca8417c} /* (20, 27, 15) {real, imag} */,
  {32'hbccab958, 32'h3d28c4be} /* (20, 27, 14) {real, imag} */,
  {32'h3d2faee0, 32'hbc309b9e} /* (20, 27, 13) {real, imag} */,
  {32'h3b9e9908, 32'hbd69cb3e} /* (20, 27, 12) {real, imag} */,
  {32'hbc4c27d4, 32'h3cbdadf4} /* (20, 27, 11) {real, imag} */,
  {32'h3dc3fe4c, 32'hbc4caad4} /* (20, 27, 10) {real, imag} */,
  {32'h3dc9fc74, 32'hbdb3c946} /* (20, 27, 9) {real, imag} */,
  {32'hbd127d0c, 32'h3d25296a} /* (20, 27, 8) {real, imag} */,
  {32'hbdeb9638, 32'h3dd2b0da} /* (20, 27, 7) {real, imag} */,
  {32'h3dc6ab37, 32'h3d9c27b2} /* (20, 27, 6) {real, imag} */,
  {32'h3e52cc03, 32'h3d62975f} /* (20, 27, 5) {real, imag} */,
  {32'hbe464c3a, 32'hbddae1c7} /* (20, 27, 4) {real, imag} */,
  {32'h3d05dc80, 32'hbd4fe343} /* (20, 27, 3) {real, imag} */,
  {32'h3fe47f0d, 32'h3f034d18} /* (20, 27, 2) {real, imag} */,
  {32'hc0a6a3a9, 32'hbf8ee9a7} /* (20, 27, 1) {real, imag} */,
  {32'hc0af427e, 32'h00000000} /* (20, 27, 0) {real, imag} */,
  {32'hc0a17475, 32'h3f7077c4} /* (20, 26, 31) {real, imag} */,
  {32'h3fec44b8, 32'hbee82b13} /* (20, 26, 30) {real, imag} */,
  {32'hbd6e5a28, 32'h3d823503} /* (20, 26, 29) {real, imag} */,
  {32'hbe9cbca2, 32'h3d54fd2e} /* (20, 26, 28) {real, imag} */,
  {32'h3e943d7c, 32'hbdea9b62} /* (20, 26, 27) {real, imag} */,
  {32'hbc0abc33, 32'hbe0d7558} /* (20, 26, 26) {real, imag} */,
  {32'hbcfc14f0, 32'hbc00900c} /* (20, 26, 25) {real, imag} */,
  {32'h3c50cb70, 32'hbd46ce72} /* (20, 26, 24) {real, imag} */,
  {32'hbc165e94, 32'h3d882f52} /* (20, 26, 23) {real, imag} */,
  {32'hbdf18fc2, 32'hbd03bc76} /* (20, 26, 22) {real, imag} */,
  {32'h3db3999c, 32'h3cb96b9f} /* (20, 26, 21) {real, imag} */,
  {32'hbc80c544, 32'h3d14d950} /* (20, 26, 20) {real, imag} */,
  {32'h3b608900, 32'hbd2dbd82} /* (20, 26, 19) {real, imag} */,
  {32'hbc547d74, 32'hbd84168a} /* (20, 26, 18) {real, imag} */,
  {32'hbc067543, 32'h3cda5004} /* (20, 26, 17) {real, imag} */,
  {32'hbd83a642, 32'h00000000} /* (20, 26, 16) {real, imag} */,
  {32'hbc067543, 32'hbcda5004} /* (20, 26, 15) {real, imag} */,
  {32'hbc547d74, 32'h3d84168a} /* (20, 26, 14) {real, imag} */,
  {32'h3b608900, 32'h3d2dbd82} /* (20, 26, 13) {real, imag} */,
  {32'hbc80c544, 32'hbd14d950} /* (20, 26, 12) {real, imag} */,
  {32'h3db3999c, 32'hbcb96b9f} /* (20, 26, 11) {real, imag} */,
  {32'hbdf18fc2, 32'h3d03bc76} /* (20, 26, 10) {real, imag} */,
  {32'hbc165e94, 32'hbd882f52} /* (20, 26, 9) {real, imag} */,
  {32'h3c50cb70, 32'h3d46ce72} /* (20, 26, 8) {real, imag} */,
  {32'hbcfc14f0, 32'h3c00900c} /* (20, 26, 7) {real, imag} */,
  {32'hbc0abc33, 32'h3e0d7558} /* (20, 26, 6) {real, imag} */,
  {32'h3e943d7c, 32'h3dea9b62} /* (20, 26, 5) {real, imag} */,
  {32'hbe9cbca2, 32'hbd54fd2e} /* (20, 26, 4) {real, imag} */,
  {32'hbd6e5a28, 32'hbd823503} /* (20, 26, 3) {real, imag} */,
  {32'h3fec44b8, 32'h3ee82b13} /* (20, 26, 2) {real, imag} */,
  {32'hc0a17475, 32'hbf7077c4} /* (20, 26, 1) {real, imag} */,
  {32'hc0a42c09, 32'h00000000} /* (20, 26, 0) {real, imag} */,
  {32'hc09683fd, 32'h3f3514d5} /* (20, 25, 31) {real, imag} */,
  {32'h3fe20683, 32'hbeccb132} /* (20, 25, 30) {real, imag} */,
  {32'h3c3d6dd8, 32'h3e29368e} /* (20, 25, 29) {real, imag} */,
  {32'hbea8fa3c, 32'h3d99f6d5} /* (20, 25, 28) {real, imag} */,
  {32'h3e87eab4, 32'hbe4f7cfd} /* (20, 25, 27) {real, imag} */,
  {32'hbde4a6b2, 32'hbdd36286} /* (20, 25, 26) {real, imag} */,
  {32'h3d2c23a2, 32'h3bf5d3b8} /* (20, 25, 25) {real, imag} */,
  {32'h3db35f24, 32'hbc4c56e0} /* (20, 25, 24) {real, imag} */,
  {32'h3c8a7214, 32'h3c81e39a} /* (20, 25, 23) {real, imag} */,
  {32'hbd97be5b, 32'h3dd33f00} /* (20, 25, 22) {real, imag} */,
  {32'h3de4257e, 32'h3cfc35ff} /* (20, 25, 21) {real, imag} */,
  {32'h3b9367c4, 32'hbd44fb36} /* (20, 25, 20) {real, imag} */,
  {32'hbd3a6dc9, 32'h3c7d6580} /* (20, 25, 19) {real, imag} */,
  {32'h3cc7977b, 32'hbced5ef2} /* (20, 25, 18) {real, imag} */,
  {32'hbd50ce93, 32'h3d7a8924} /* (20, 25, 17) {real, imag} */,
  {32'h3c8febaa, 32'h00000000} /* (20, 25, 16) {real, imag} */,
  {32'hbd50ce93, 32'hbd7a8924} /* (20, 25, 15) {real, imag} */,
  {32'h3cc7977b, 32'h3ced5ef2} /* (20, 25, 14) {real, imag} */,
  {32'hbd3a6dc9, 32'hbc7d6580} /* (20, 25, 13) {real, imag} */,
  {32'h3b9367c4, 32'h3d44fb36} /* (20, 25, 12) {real, imag} */,
  {32'h3de4257e, 32'hbcfc35ff} /* (20, 25, 11) {real, imag} */,
  {32'hbd97be5b, 32'hbdd33f00} /* (20, 25, 10) {real, imag} */,
  {32'h3c8a7214, 32'hbc81e39a} /* (20, 25, 9) {real, imag} */,
  {32'h3db35f24, 32'h3c4c56e0} /* (20, 25, 8) {real, imag} */,
  {32'h3d2c23a2, 32'hbbf5d3b8} /* (20, 25, 7) {real, imag} */,
  {32'hbde4a6b2, 32'h3dd36286} /* (20, 25, 6) {real, imag} */,
  {32'h3e87eab4, 32'h3e4f7cfd} /* (20, 25, 5) {real, imag} */,
  {32'hbea8fa3c, 32'hbd99f6d5} /* (20, 25, 4) {real, imag} */,
  {32'h3c3d6dd8, 32'hbe29368e} /* (20, 25, 3) {real, imag} */,
  {32'h3fe20683, 32'h3eccb132} /* (20, 25, 2) {real, imag} */,
  {32'hc09683fd, 32'hbf3514d5} /* (20, 25, 1) {real, imag} */,
  {32'hc0970893, 32'h00000000} /* (20, 25, 0) {real, imag} */,
  {32'hc083e6e4, 32'h3ec9f4bc} /* (20, 24, 31) {real, imag} */,
  {32'h3fd38d6e, 32'hbee5e0ef} /* (20, 24, 30) {real, imag} */,
  {32'hbd66524e, 32'h3ba399b8} /* (20, 24, 29) {real, imag} */,
  {32'hbe905998, 32'h3c345bca} /* (20, 24, 28) {real, imag} */,
  {32'h3e538bbd, 32'hbe11bb7c} /* (20, 24, 27) {real, imag} */,
  {32'h3d81d84c, 32'hbdc6651a} /* (20, 24, 26) {real, imag} */,
  {32'hbca78d33, 32'h3d52efb8} /* (20, 24, 25) {real, imag} */,
  {32'h3d9d11e3, 32'hbb6c9380} /* (20, 24, 24) {real, imag} */,
  {32'h3d03d01e, 32'h3cc2af9a} /* (20, 24, 23) {real, imag} */,
  {32'hbce32ff8, 32'h3dd42942} /* (20, 24, 22) {real, imag} */,
  {32'hbd62635c, 32'hbd636df3} /* (20, 24, 21) {real, imag} */,
  {32'hbe10be86, 32'hbd895bf9} /* (20, 24, 20) {real, imag} */,
  {32'h3d80979f, 32'hbd8b7a39} /* (20, 24, 19) {real, imag} */,
  {32'hbb3d8bb4, 32'h3d5951fe} /* (20, 24, 18) {real, imag} */,
  {32'hbd885d47, 32'h3d7f3145} /* (20, 24, 17) {real, imag} */,
  {32'hbd13a6ec, 32'h00000000} /* (20, 24, 16) {real, imag} */,
  {32'hbd885d47, 32'hbd7f3145} /* (20, 24, 15) {real, imag} */,
  {32'hbb3d8bb4, 32'hbd5951fe} /* (20, 24, 14) {real, imag} */,
  {32'h3d80979f, 32'h3d8b7a39} /* (20, 24, 13) {real, imag} */,
  {32'hbe10be86, 32'h3d895bf9} /* (20, 24, 12) {real, imag} */,
  {32'hbd62635c, 32'h3d636df3} /* (20, 24, 11) {real, imag} */,
  {32'hbce32ff8, 32'hbdd42942} /* (20, 24, 10) {real, imag} */,
  {32'h3d03d01e, 32'hbcc2af9a} /* (20, 24, 9) {real, imag} */,
  {32'h3d9d11e3, 32'h3b6c9380} /* (20, 24, 8) {real, imag} */,
  {32'hbca78d33, 32'hbd52efb8} /* (20, 24, 7) {real, imag} */,
  {32'h3d81d84c, 32'h3dc6651a} /* (20, 24, 6) {real, imag} */,
  {32'h3e538bbd, 32'h3e11bb7c} /* (20, 24, 5) {real, imag} */,
  {32'hbe905998, 32'hbc345bca} /* (20, 24, 4) {real, imag} */,
  {32'hbd66524e, 32'hbba399b8} /* (20, 24, 3) {real, imag} */,
  {32'h3fd38d6e, 32'h3ee5e0ef} /* (20, 24, 2) {real, imag} */,
  {32'hc083e6e4, 32'hbec9f4bc} /* (20, 24, 1) {real, imag} */,
  {32'hc0879053, 32'h00000000} /* (20, 24, 0) {real, imag} */,
  {32'hc0572b0a, 32'h3e9b6524} /* (20, 23, 31) {real, imag} */,
  {32'h3fb478e9, 32'hbeccb476} /* (20, 23, 30) {real, imag} */,
  {32'hbdbf1738, 32'hbd622f9c} /* (20, 23, 29) {real, imag} */,
  {32'hbe69b93c, 32'hbd02c8be} /* (20, 23, 28) {real, imag} */,
  {32'h3e96b4e4, 32'hbe008958} /* (20, 23, 27) {real, imag} */,
  {32'hbd9bc844, 32'hbdab12b2} /* (20, 23, 26) {real, imag} */,
  {32'hbd10dad0, 32'h3ba0e860} /* (20, 23, 25) {real, imag} */,
  {32'h3cb2443c, 32'hbdd4ad54} /* (20, 23, 24) {real, imag} */,
  {32'hbd9712c1, 32'h3dbe1690} /* (20, 23, 23) {real, imag} */,
  {32'h3defc4d0, 32'hbcc0fccd} /* (20, 23, 22) {real, imag} */,
  {32'hbd2c12a2, 32'hbdd35ef9} /* (20, 23, 21) {real, imag} */,
  {32'h3c81480c, 32'h3c961914} /* (20, 23, 20) {real, imag} */,
  {32'h3c73dfab, 32'hbd6f0d4c} /* (20, 23, 19) {real, imag} */,
  {32'h3d137962, 32'hbd0bcd9f} /* (20, 23, 18) {real, imag} */,
  {32'h3cccbdda, 32'h3d5a08d6} /* (20, 23, 17) {real, imag} */,
  {32'h3ca60664, 32'h00000000} /* (20, 23, 16) {real, imag} */,
  {32'h3cccbdda, 32'hbd5a08d6} /* (20, 23, 15) {real, imag} */,
  {32'h3d137962, 32'h3d0bcd9f} /* (20, 23, 14) {real, imag} */,
  {32'h3c73dfab, 32'h3d6f0d4c} /* (20, 23, 13) {real, imag} */,
  {32'h3c81480c, 32'hbc961914} /* (20, 23, 12) {real, imag} */,
  {32'hbd2c12a2, 32'h3dd35ef9} /* (20, 23, 11) {real, imag} */,
  {32'h3defc4d0, 32'h3cc0fccd} /* (20, 23, 10) {real, imag} */,
  {32'hbd9712c1, 32'hbdbe1690} /* (20, 23, 9) {real, imag} */,
  {32'h3cb2443c, 32'h3dd4ad54} /* (20, 23, 8) {real, imag} */,
  {32'hbd10dad0, 32'hbba0e860} /* (20, 23, 7) {real, imag} */,
  {32'hbd9bc844, 32'h3dab12b2} /* (20, 23, 6) {real, imag} */,
  {32'h3e96b4e4, 32'h3e008958} /* (20, 23, 5) {real, imag} */,
  {32'hbe69b93c, 32'h3d02c8be} /* (20, 23, 4) {real, imag} */,
  {32'hbdbf1738, 32'h3d622f9c} /* (20, 23, 3) {real, imag} */,
  {32'h3fb478e9, 32'h3eccb476} /* (20, 23, 2) {real, imag} */,
  {32'hc0572b0a, 32'hbe9b6524} /* (20, 23, 1) {real, imag} */,
  {32'hc05e9efb, 32'h00000000} /* (20, 23, 0) {real, imag} */,
  {32'hc01dcdbd, 32'h3e3bd170} /* (20, 22, 31) {real, imag} */,
  {32'h3f80ea52, 32'hbe9d36ad} /* (20, 22, 30) {real, imag} */,
  {32'hba3f77c0, 32'h3d3ad6a0} /* (20, 22, 29) {real, imag} */,
  {32'hbe9aebbb, 32'hbd2c4468} /* (20, 22, 28) {real, imag} */,
  {32'h3e92265a, 32'hbe23cb96} /* (20, 22, 27) {real, imag} */,
  {32'hbd3c32c0, 32'h3b35f088} /* (20, 22, 26) {real, imag} */,
  {32'hbc641fec, 32'hbcb4b2a0} /* (20, 22, 25) {real, imag} */,
  {32'hbba02d00, 32'hbdf06dd8} /* (20, 22, 24) {real, imag} */,
  {32'hbd828144, 32'h3d32134b} /* (20, 22, 23) {real, imag} */,
  {32'hbb555f38, 32'hbd0314fd} /* (20, 22, 22) {real, imag} */,
  {32'h3b848fc0, 32'hbd8fadd2} /* (20, 22, 21) {real, imag} */,
  {32'h3d7694d8, 32'hbcfcf21f} /* (20, 22, 20) {real, imag} */,
  {32'h3cff8fde, 32'hbc785a80} /* (20, 22, 19) {real, imag} */,
  {32'h3cde4028, 32'hbb913560} /* (20, 22, 18) {real, imag} */,
  {32'h3d4297ce, 32'hbd38be40} /* (20, 22, 17) {real, imag} */,
  {32'h3d9d4442, 32'h00000000} /* (20, 22, 16) {real, imag} */,
  {32'h3d4297ce, 32'h3d38be40} /* (20, 22, 15) {real, imag} */,
  {32'h3cde4028, 32'h3b913560} /* (20, 22, 14) {real, imag} */,
  {32'h3cff8fde, 32'h3c785a80} /* (20, 22, 13) {real, imag} */,
  {32'h3d7694d8, 32'h3cfcf21f} /* (20, 22, 12) {real, imag} */,
  {32'h3b848fc0, 32'h3d8fadd2} /* (20, 22, 11) {real, imag} */,
  {32'hbb555f38, 32'h3d0314fd} /* (20, 22, 10) {real, imag} */,
  {32'hbd828144, 32'hbd32134b} /* (20, 22, 9) {real, imag} */,
  {32'hbba02d00, 32'h3df06dd8} /* (20, 22, 8) {real, imag} */,
  {32'hbc641fec, 32'h3cb4b2a0} /* (20, 22, 7) {real, imag} */,
  {32'hbd3c32c0, 32'hbb35f088} /* (20, 22, 6) {real, imag} */,
  {32'h3e92265a, 32'h3e23cb96} /* (20, 22, 5) {real, imag} */,
  {32'hbe9aebbb, 32'h3d2c4468} /* (20, 22, 4) {real, imag} */,
  {32'hba3f77c0, 32'hbd3ad6a0} /* (20, 22, 3) {real, imag} */,
  {32'h3f80ea52, 32'h3e9d36ad} /* (20, 22, 2) {real, imag} */,
  {32'hc01dcdbd, 32'hbe3bd170} /* (20, 22, 1) {real, imag} */,
  {32'hc01d4479, 32'h00000000} /* (20, 22, 0) {real, imag} */,
  {32'hbf6624a5, 32'h3d792000} /* (20, 21, 31) {real, imag} */,
  {32'h3ea303a8, 32'hbddf662e} /* (20, 21, 30) {real, imag} */,
  {32'hbd9a3b10, 32'h3e4f760a} /* (20, 21, 29) {real, imag} */,
  {32'hbdab100d, 32'hbd591a4e} /* (20, 21, 28) {real, imag} */,
  {32'h3de6b612, 32'h3c66375c} /* (20, 21, 27) {real, imag} */,
  {32'h3a963878, 32'hbaa17130} /* (20, 21, 26) {real, imag} */,
  {32'h3cad6255, 32'hbd96a914} /* (20, 21, 25) {real, imag} */,
  {32'hbc90001c, 32'hbd2d366c} /* (20, 21, 24) {real, imag} */,
  {32'h3d967dc7, 32'h3caaee82} /* (20, 21, 23) {real, imag} */,
  {32'hbe0cf9d2, 32'hbd76edcb} /* (20, 21, 22) {real, imag} */,
  {32'h3da8563e, 32'hbd882df3} /* (20, 21, 21) {real, imag} */,
  {32'h3e313ba6, 32'h3c50a1c0} /* (20, 21, 20) {real, imag} */,
  {32'hbd4e240e, 32'h3c2c9409} /* (20, 21, 19) {real, imag} */,
  {32'h3d08be72, 32'h3dc30613} /* (20, 21, 18) {real, imag} */,
  {32'hbc953eb3, 32'hbcf865b8} /* (20, 21, 17) {real, imag} */,
  {32'hbde592c7, 32'h00000000} /* (20, 21, 16) {real, imag} */,
  {32'hbc953eb3, 32'h3cf865b8} /* (20, 21, 15) {real, imag} */,
  {32'h3d08be72, 32'hbdc30613} /* (20, 21, 14) {real, imag} */,
  {32'hbd4e240e, 32'hbc2c9409} /* (20, 21, 13) {real, imag} */,
  {32'h3e313ba6, 32'hbc50a1c0} /* (20, 21, 12) {real, imag} */,
  {32'h3da8563e, 32'h3d882df3} /* (20, 21, 11) {real, imag} */,
  {32'hbe0cf9d2, 32'h3d76edcb} /* (20, 21, 10) {real, imag} */,
  {32'h3d967dc7, 32'hbcaaee82} /* (20, 21, 9) {real, imag} */,
  {32'hbc90001c, 32'h3d2d366c} /* (20, 21, 8) {real, imag} */,
  {32'h3cad6255, 32'h3d96a914} /* (20, 21, 7) {real, imag} */,
  {32'h3a963878, 32'h3aa17130} /* (20, 21, 6) {real, imag} */,
  {32'h3de6b612, 32'hbc66375c} /* (20, 21, 5) {real, imag} */,
  {32'hbdab100d, 32'h3d591a4e} /* (20, 21, 4) {real, imag} */,
  {32'hbd9a3b10, 32'hbe4f760a} /* (20, 21, 3) {real, imag} */,
  {32'h3ea303a8, 32'h3ddf662e} /* (20, 21, 2) {real, imag} */,
  {32'hbf6624a5, 32'hbd792000} /* (20, 21, 1) {real, imag} */,
  {32'hbf9957e8, 32'h00000000} /* (20, 21, 0) {real, imag} */,
  {32'h3f979ad2, 32'hbea9ad46} /* (20, 20, 31) {real, imag} */,
  {32'hbef5db26, 32'h3da5b4f0} /* (20, 20, 30) {real, imag} */,
  {32'hbd2932aa, 32'h3d15a9fe} /* (20, 20, 29) {real, imag} */,
  {32'h3aa942c0, 32'hbe5300c4} /* (20, 20, 28) {real, imag} */,
  {32'hbd808ae4, 32'h3da02f62} /* (20, 20, 27) {real, imag} */,
  {32'h3d665e61, 32'hbd09d682} /* (20, 20, 26) {real, imag} */,
  {32'hbc7f94ca, 32'hbdc2a7fd} /* (20, 20, 25) {real, imag} */,
  {32'hbe4cf254, 32'h3de88649} /* (20, 20, 24) {real, imag} */,
  {32'hbda16fa2, 32'hbd2bb0bf} /* (20, 20, 23) {real, imag} */,
  {32'hbd85f384, 32'hbdaf42fc} /* (20, 20, 22) {real, imag} */,
  {32'h3cdb0fad, 32'h3d9a0ada} /* (20, 20, 21) {real, imag} */,
  {32'h3c888282, 32'h3ceaa86c} /* (20, 20, 20) {real, imag} */,
  {32'h3c19f296, 32'h3c99d7d6} /* (20, 20, 19) {real, imag} */,
  {32'h3c85076e, 32'h3c95b1ae} /* (20, 20, 18) {real, imag} */,
  {32'hbca1091d, 32'hbbcb01f4} /* (20, 20, 17) {real, imag} */,
  {32'h3c99fef7, 32'h00000000} /* (20, 20, 16) {real, imag} */,
  {32'hbca1091d, 32'h3bcb01f4} /* (20, 20, 15) {real, imag} */,
  {32'h3c85076e, 32'hbc95b1ae} /* (20, 20, 14) {real, imag} */,
  {32'h3c19f296, 32'hbc99d7d6} /* (20, 20, 13) {real, imag} */,
  {32'h3c888282, 32'hbceaa86c} /* (20, 20, 12) {real, imag} */,
  {32'h3cdb0fad, 32'hbd9a0ada} /* (20, 20, 11) {real, imag} */,
  {32'hbd85f384, 32'h3daf42fc} /* (20, 20, 10) {real, imag} */,
  {32'hbda16fa2, 32'h3d2bb0bf} /* (20, 20, 9) {real, imag} */,
  {32'hbe4cf254, 32'hbde88649} /* (20, 20, 8) {real, imag} */,
  {32'hbc7f94ca, 32'h3dc2a7fd} /* (20, 20, 7) {real, imag} */,
  {32'h3d665e61, 32'h3d09d682} /* (20, 20, 6) {real, imag} */,
  {32'hbd808ae4, 32'hbda02f62} /* (20, 20, 5) {real, imag} */,
  {32'h3aa942c0, 32'h3e5300c4} /* (20, 20, 4) {real, imag} */,
  {32'hbd2932aa, 32'hbd15a9fe} /* (20, 20, 3) {real, imag} */,
  {32'hbef5db26, 32'hbda5b4f0} /* (20, 20, 2) {real, imag} */,
  {32'h3f979ad2, 32'h3ea9ad46} /* (20, 20, 1) {real, imag} */,
  {32'h3e978e10, 32'h00000000} /* (20, 20, 0) {real, imag} */,
  {32'h4029951d, 32'hbf0a6b8e} /* (20, 19, 31) {real, imag} */,
  {32'hbf858203, 32'h3e181488} /* (20, 19, 30) {real, imag} */,
  {32'h3e17ce9b, 32'h3dded765} /* (20, 19, 29) {real, imag} */,
  {32'h3e070d9b, 32'hbd9cc6d9} /* (20, 19, 28) {real, imag} */,
  {32'hbe41a794, 32'h3d816396} /* (20, 19, 27) {real, imag} */,
  {32'hbd689051, 32'h3daa467d} /* (20, 19, 26) {real, imag} */,
  {32'h3ddaa742, 32'h3cb4d26a} /* (20, 19, 25) {real, imag} */,
  {32'h3d056008, 32'h3ddf8f86} /* (20, 19, 24) {real, imag} */,
  {32'hbda5aa88, 32'h3cd7e176} /* (20, 19, 23) {real, imag} */,
  {32'h3d46894d, 32'hbc282950} /* (20, 19, 22) {real, imag} */,
  {32'h3c86d96e, 32'h3d97c782} /* (20, 19, 21) {real, imag} */,
  {32'hbdcaac53, 32'h3d56c6ee} /* (20, 19, 20) {real, imag} */,
  {32'hbd1aa3fe, 32'hbd51ba43} /* (20, 19, 19) {real, imag} */,
  {32'h3c2d22f0, 32'h3cedeec2} /* (20, 19, 18) {real, imag} */,
  {32'hbd08be3d, 32'hbd21f0ee} /* (20, 19, 17) {real, imag} */,
  {32'hbc55914c, 32'h00000000} /* (20, 19, 16) {real, imag} */,
  {32'hbd08be3d, 32'h3d21f0ee} /* (20, 19, 15) {real, imag} */,
  {32'h3c2d22f0, 32'hbcedeec2} /* (20, 19, 14) {real, imag} */,
  {32'hbd1aa3fe, 32'h3d51ba43} /* (20, 19, 13) {real, imag} */,
  {32'hbdcaac53, 32'hbd56c6ee} /* (20, 19, 12) {real, imag} */,
  {32'h3c86d96e, 32'hbd97c782} /* (20, 19, 11) {real, imag} */,
  {32'h3d46894d, 32'h3c282950} /* (20, 19, 10) {real, imag} */,
  {32'hbda5aa88, 32'hbcd7e176} /* (20, 19, 9) {real, imag} */,
  {32'h3d056008, 32'hbddf8f86} /* (20, 19, 8) {real, imag} */,
  {32'h3ddaa742, 32'hbcb4d26a} /* (20, 19, 7) {real, imag} */,
  {32'hbd689051, 32'hbdaa467d} /* (20, 19, 6) {real, imag} */,
  {32'hbe41a794, 32'hbd816396} /* (20, 19, 5) {real, imag} */,
  {32'h3e070d9b, 32'h3d9cc6d9} /* (20, 19, 4) {real, imag} */,
  {32'h3e17ce9b, 32'hbdded765} /* (20, 19, 3) {real, imag} */,
  {32'hbf858203, 32'hbe181488} /* (20, 19, 2) {real, imag} */,
  {32'h4029951d, 32'h3f0a6b8e} /* (20, 19, 1) {real, imag} */,
  {32'h3fa8feb5, 32'h00000000} /* (20, 19, 0) {real, imag} */,
  {32'h40651d40, 32'hbef68438} /* (20, 18, 31) {real, imag} */,
  {32'hbfadab4c, 32'h3e8cf7ea} /* (20, 18, 30) {real, imag} */,
  {32'h3e53a886, 32'h3e1d8a13} /* (20, 18, 29) {real, imag} */,
  {32'h3da7fea6, 32'hbddc6c93} /* (20, 18, 28) {real, imag} */,
  {32'hbdf59b36, 32'h3ddccec5} /* (20, 18, 27) {real, imag} */,
  {32'h3ca061a8, 32'h3ce8b7fe} /* (20, 18, 26) {real, imag} */,
  {32'h3e2d3066, 32'h3da2ca2f} /* (20, 18, 25) {real, imag} */,
  {32'h3d35d6b5, 32'h3e06027f} /* (20, 18, 24) {real, imag} */,
  {32'h3d5b0be7, 32'h3cad76c1} /* (20, 18, 23) {real, imag} */,
  {32'hbd3e0081, 32'h3dc8fda4} /* (20, 18, 22) {real, imag} */,
  {32'h3d848772, 32'h3dcf4a86} /* (20, 18, 21) {real, imag} */,
  {32'h3e1b7e11, 32'hbda97d19} /* (20, 18, 20) {real, imag} */,
  {32'h3d37010c, 32'h3d9b7400} /* (20, 18, 19) {real, imag} */,
  {32'h3c9b1f78, 32'h3da695c7} /* (20, 18, 18) {real, imag} */,
  {32'h3d84f7b2, 32'hbd644420} /* (20, 18, 17) {real, imag} */,
  {32'hbbbf8818, 32'h00000000} /* (20, 18, 16) {real, imag} */,
  {32'h3d84f7b2, 32'h3d644420} /* (20, 18, 15) {real, imag} */,
  {32'h3c9b1f78, 32'hbda695c7} /* (20, 18, 14) {real, imag} */,
  {32'h3d37010c, 32'hbd9b7400} /* (20, 18, 13) {real, imag} */,
  {32'h3e1b7e11, 32'h3da97d19} /* (20, 18, 12) {real, imag} */,
  {32'h3d848772, 32'hbdcf4a86} /* (20, 18, 11) {real, imag} */,
  {32'hbd3e0081, 32'hbdc8fda4} /* (20, 18, 10) {real, imag} */,
  {32'h3d5b0be7, 32'hbcad76c1} /* (20, 18, 9) {real, imag} */,
  {32'h3d35d6b5, 32'hbe06027f} /* (20, 18, 8) {real, imag} */,
  {32'h3e2d3066, 32'hbda2ca2f} /* (20, 18, 7) {real, imag} */,
  {32'h3ca061a8, 32'hbce8b7fe} /* (20, 18, 6) {real, imag} */,
  {32'hbdf59b36, 32'hbddccec5} /* (20, 18, 5) {real, imag} */,
  {32'h3da7fea6, 32'h3ddc6c93} /* (20, 18, 4) {real, imag} */,
  {32'h3e53a886, 32'hbe1d8a13} /* (20, 18, 3) {real, imag} */,
  {32'hbfadab4c, 32'hbe8cf7ea} /* (20, 18, 2) {real, imag} */,
  {32'h40651d40, 32'h3ef68438} /* (20, 18, 1) {real, imag} */,
  {32'h40136f46, 32'h00000000} /* (20, 18, 0) {real, imag} */,
  {32'h40853c97, 32'hbee2edb0} /* (20, 17, 31) {real, imag} */,
  {32'hbfbd7904, 32'h3e96b539} /* (20, 17, 30) {real, imag} */,
  {32'h3c7b6800, 32'h3e348b58} /* (20, 17, 29) {real, imag} */,
  {32'h3df3b150, 32'h3c19faa0} /* (20, 17, 28) {real, imag} */,
  {32'hbd83637a, 32'h3dc5c54d} /* (20, 17, 27) {real, imag} */,
  {32'hbd0d0387, 32'h3d57cb0c} /* (20, 17, 26) {real, imag} */,
  {32'h3db4d180, 32'hbd5abf86} /* (20, 17, 25) {real, imag} */,
  {32'h3c515d50, 32'h3e4bb49a} /* (20, 17, 24) {real, imag} */,
  {32'hbd572ce5, 32'h3cc3d910} /* (20, 17, 23) {real, imag} */,
  {32'hbd8884ae, 32'h3daec4df} /* (20, 17, 22) {real, imag} */,
  {32'hbc9f473c, 32'hbcaa34fc} /* (20, 17, 21) {real, imag} */,
  {32'hbdf32930, 32'h3d0458fa} /* (20, 17, 20) {real, imag} */,
  {32'hbc2b4166, 32'hbd091804} /* (20, 17, 19) {real, imag} */,
  {32'hbdd589d4, 32'h3c944ae6} /* (20, 17, 18) {real, imag} */,
  {32'h3c630888, 32'h3d697dfd} /* (20, 17, 17) {real, imag} */,
  {32'hbc3c6cd6, 32'h00000000} /* (20, 17, 16) {real, imag} */,
  {32'h3c630888, 32'hbd697dfd} /* (20, 17, 15) {real, imag} */,
  {32'hbdd589d4, 32'hbc944ae6} /* (20, 17, 14) {real, imag} */,
  {32'hbc2b4166, 32'h3d091804} /* (20, 17, 13) {real, imag} */,
  {32'hbdf32930, 32'hbd0458fa} /* (20, 17, 12) {real, imag} */,
  {32'hbc9f473c, 32'h3caa34fc} /* (20, 17, 11) {real, imag} */,
  {32'hbd8884ae, 32'hbdaec4df} /* (20, 17, 10) {real, imag} */,
  {32'hbd572ce5, 32'hbcc3d910} /* (20, 17, 9) {real, imag} */,
  {32'h3c515d50, 32'hbe4bb49a} /* (20, 17, 8) {real, imag} */,
  {32'h3db4d180, 32'h3d5abf86} /* (20, 17, 7) {real, imag} */,
  {32'hbd0d0387, 32'hbd57cb0c} /* (20, 17, 6) {real, imag} */,
  {32'hbd83637a, 32'hbdc5c54d} /* (20, 17, 5) {real, imag} */,
  {32'h3df3b150, 32'hbc19faa0} /* (20, 17, 4) {real, imag} */,
  {32'h3c7b6800, 32'hbe348b58} /* (20, 17, 3) {real, imag} */,
  {32'hbfbd7904, 32'hbe96b539} /* (20, 17, 2) {real, imag} */,
  {32'h40853c97, 32'h3ee2edb0} /* (20, 17, 1) {real, imag} */,
  {32'h40376323, 32'h00000000} /* (20, 17, 0) {real, imag} */,
  {32'h408c7d09, 32'hbed91a60} /* (20, 16, 31) {real, imag} */,
  {32'hbfc4cc8f, 32'h3e918204} /* (20, 16, 30) {real, imag} */,
  {32'hbdd577a0, 32'h3d78213f} /* (20, 16, 29) {real, imag} */,
  {32'h3e7ce630, 32'h3bf58c80} /* (20, 16, 28) {real, imag} */,
  {32'hbe333520, 32'h3dd6b5be} /* (20, 16, 27) {real, imag} */,
  {32'hbd7f2f84, 32'hbdb3b473} /* (20, 16, 26) {real, imag} */,
  {32'h3dee110f, 32'hbc03017c} /* (20, 16, 25) {real, imag} */,
  {32'h3bc92e6c, 32'h3d2d16b9} /* (20, 16, 24) {real, imag} */,
  {32'hbc942a8e, 32'h3c09ed88} /* (20, 16, 23) {real, imag} */,
  {32'hbcfe20e9, 32'hbdb634a6} /* (20, 16, 22) {real, imag} */,
  {32'h3c3eae0e, 32'h3cb1f20f} /* (20, 16, 21) {real, imag} */,
  {32'h3c8804ae, 32'h3c1c5570} /* (20, 16, 20) {real, imag} */,
  {32'h3da4f4c1, 32'h3d17759f} /* (20, 16, 19) {real, imag} */,
  {32'hbb5c1ca0, 32'hbc2255b9} /* (20, 16, 18) {real, imag} */,
  {32'h3d21fcb2, 32'hbd1c8789} /* (20, 16, 17) {real, imag} */,
  {32'h3b2b3254, 32'h00000000} /* (20, 16, 16) {real, imag} */,
  {32'h3d21fcb2, 32'h3d1c8789} /* (20, 16, 15) {real, imag} */,
  {32'hbb5c1ca0, 32'h3c2255b9} /* (20, 16, 14) {real, imag} */,
  {32'h3da4f4c1, 32'hbd17759f} /* (20, 16, 13) {real, imag} */,
  {32'h3c8804ae, 32'hbc1c5570} /* (20, 16, 12) {real, imag} */,
  {32'h3c3eae0e, 32'hbcb1f20f} /* (20, 16, 11) {real, imag} */,
  {32'hbcfe20e9, 32'h3db634a6} /* (20, 16, 10) {real, imag} */,
  {32'hbc942a8e, 32'hbc09ed88} /* (20, 16, 9) {real, imag} */,
  {32'h3bc92e6c, 32'hbd2d16b9} /* (20, 16, 8) {real, imag} */,
  {32'h3dee110f, 32'h3c03017c} /* (20, 16, 7) {real, imag} */,
  {32'hbd7f2f84, 32'h3db3b473} /* (20, 16, 6) {real, imag} */,
  {32'hbe333520, 32'hbdd6b5be} /* (20, 16, 5) {real, imag} */,
  {32'h3e7ce630, 32'hbbf58c80} /* (20, 16, 4) {real, imag} */,
  {32'hbdd577a0, 32'hbd78213f} /* (20, 16, 3) {real, imag} */,
  {32'hbfc4cc8f, 32'hbe918204} /* (20, 16, 2) {real, imag} */,
  {32'h408c7d09, 32'h3ed91a60} /* (20, 16, 1) {real, imag} */,
  {32'h404444fc, 32'h00000000} /* (20, 16, 0) {real, imag} */,
  {32'h408e8351, 32'hbece2fc8} /* (20, 15, 31) {real, imag} */,
  {32'hbfbcd816, 32'h3ed1d735} /* (20, 15, 30) {real, imag} */,
  {32'hbdf2803c, 32'h3c9bc054} /* (20, 15, 29) {real, imag} */,
  {32'h3e27e880, 32'hbe2b6ff4} /* (20, 15, 28) {real, imag} */,
  {32'hbea243a4, 32'h3ddcd343} /* (20, 15, 27) {real, imag} */,
  {32'hbdb1d3c8, 32'hbddf68a8} /* (20, 15, 26) {real, imag} */,
  {32'hbd528f45, 32'hbdf60e25} /* (20, 15, 25) {real, imag} */,
  {32'hbe24bf60, 32'h3dc45794} /* (20, 15, 24) {real, imag} */,
  {32'h3d6b5afb, 32'hbd9254f1} /* (20, 15, 23) {real, imag} */,
  {32'hbd5aa450, 32'hbd3293ca} /* (20, 15, 22) {real, imag} */,
  {32'h3d93076a, 32'h3c9febb6} /* (20, 15, 21) {real, imag} */,
  {32'h3d20e8d0, 32'hbdace051} /* (20, 15, 20) {real, imag} */,
  {32'h3c1a2496, 32'hbcbd3ec8} /* (20, 15, 19) {real, imag} */,
  {32'h3d222bd9, 32'h3cbf5ee2} /* (20, 15, 18) {real, imag} */,
  {32'hbdd2cb81, 32'h3d5b949d} /* (20, 15, 17) {real, imag} */,
  {32'h3aa3c5a0, 32'h00000000} /* (20, 15, 16) {real, imag} */,
  {32'hbdd2cb81, 32'hbd5b949d} /* (20, 15, 15) {real, imag} */,
  {32'h3d222bd9, 32'hbcbf5ee2} /* (20, 15, 14) {real, imag} */,
  {32'h3c1a2496, 32'h3cbd3ec8} /* (20, 15, 13) {real, imag} */,
  {32'h3d20e8d0, 32'h3dace051} /* (20, 15, 12) {real, imag} */,
  {32'h3d93076a, 32'hbc9febb6} /* (20, 15, 11) {real, imag} */,
  {32'hbd5aa450, 32'h3d3293ca} /* (20, 15, 10) {real, imag} */,
  {32'h3d6b5afb, 32'h3d9254f1} /* (20, 15, 9) {real, imag} */,
  {32'hbe24bf60, 32'hbdc45794} /* (20, 15, 8) {real, imag} */,
  {32'hbd528f45, 32'h3df60e25} /* (20, 15, 7) {real, imag} */,
  {32'hbdb1d3c8, 32'h3ddf68a8} /* (20, 15, 6) {real, imag} */,
  {32'hbea243a4, 32'hbddcd343} /* (20, 15, 5) {real, imag} */,
  {32'h3e27e880, 32'h3e2b6ff4} /* (20, 15, 4) {real, imag} */,
  {32'hbdf2803c, 32'hbc9bc054} /* (20, 15, 3) {real, imag} */,
  {32'hbfbcd816, 32'hbed1d735} /* (20, 15, 2) {real, imag} */,
  {32'h408e8351, 32'h3ece2fc8} /* (20, 15, 1) {real, imag} */,
  {32'h40411a7f, 32'h00000000} /* (20, 15, 0) {real, imag} */,
  {32'h40792a38, 32'hbea14308} /* (20, 14, 31) {real, imag} */,
  {32'hbfc9684c, 32'h3ea36ec6} /* (20, 14, 30) {real, imag} */,
  {32'hbcf37a40, 32'hbdb825ee} /* (20, 14, 29) {real, imag} */,
  {32'h3e919f18, 32'hbdbb3cbb} /* (20, 14, 28) {real, imag} */,
  {32'hbe61779f, 32'h3dffd84f} /* (20, 14, 27) {real, imag} */,
  {32'hbce3b2e8, 32'h3d9937cc} /* (20, 14, 26) {real, imag} */,
  {32'h3d01bec6, 32'hbd3aa84e} /* (20, 14, 25) {real, imag} */,
  {32'hbd9069c0, 32'h3dbb8717} /* (20, 14, 24) {real, imag} */,
  {32'h3d0a23cd, 32'h3cb8c603} /* (20, 14, 23) {real, imag} */,
  {32'hbd1b9069, 32'hbcea1210} /* (20, 14, 22) {real, imag} */,
  {32'hbd86675e, 32'h3c2675ac} /* (20, 14, 21) {real, imag} */,
  {32'h3d159a85, 32'hbbb878d0} /* (20, 14, 20) {real, imag} */,
  {32'hbe04c135, 32'h3cb061e9} /* (20, 14, 19) {real, imag} */,
  {32'hbd098c61, 32'h3d11e26e} /* (20, 14, 18) {real, imag} */,
  {32'h3cad693a, 32'h3c684c48} /* (20, 14, 17) {real, imag} */,
  {32'hbd426a76, 32'h00000000} /* (20, 14, 16) {real, imag} */,
  {32'h3cad693a, 32'hbc684c48} /* (20, 14, 15) {real, imag} */,
  {32'hbd098c61, 32'hbd11e26e} /* (20, 14, 14) {real, imag} */,
  {32'hbe04c135, 32'hbcb061e9} /* (20, 14, 13) {real, imag} */,
  {32'h3d159a85, 32'h3bb878d0} /* (20, 14, 12) {real, imag} */,
  {32'hbd86675e, 32'hbc2675ac} /* (20, 14, 11) {real, imag} */,
  {32'hbd1b9069, 32'h3cea1210} /* (20, 14, 10) {real, imag} */,
  {32'h3d0a23cd, 32'hbcb8c603} /* (20, 14, 9) {real, imag} */,
  {32'hbd9069c0, 32'hbdbb8717} /* (20, 14, 8) {real, imag} */,
  {32'h3d01bec6, 32'h3d3aa84e} /* (20, 14, 7) {real, imag} */,
  {32'hbce3b2e8, 32'hbd9937cc} /* (20, 14, 6) {real, imag} */,
  {32'hbe61779f, 32'hbdffd84f} /* (20, 14, 5) {real, imag} */,
  {32'h3e919f18, 32'h3dbb3cbb} /* (20, 14, 4) {real, imag} */,
  {32'hbcf37a40, 32'h3db825ee} /* (20, 14, 3) {real, imag} */,
  {32'hbfc9684c, 32'hbea36ec6} /* (20, 14, 2) {real, imag} */,
  {32'h40792a38, 32'h3ea14308} /* (20, 14, 1) {real, imag} */,
  {32'h40334992, 32'h00000000} /* (20, 14, 0) {real, imag} */,
  {32'h404fb1af, 32'hbe3fb158} /* (20, 13, 31) {real, imag} */,
  {32'hbfb3e6c1, 32'h3ea8d8fa} /* (20, 13, 30) {real, imag} */,
  {32'hbccb8412, 32'hbe2cd8a2} /* (20, 13, 29) {real, imag} */,
  {32'h3e80063a, 32'hbcb8d43c} /* (20, 13, 28) {real, imag} */,
  {32'hbe8306dd, 32'h3e400d53} /* (20, 13, 27) {real, imag} */,
  {32'h3d4c3225, 32'h3cf21c6b} /* (20, 13, 26) {real, imag} */,
  {32'h3e00dc35, 32'hbc90dd66} /* (20, 13, 25) {real, imag} */,
  {32'h3bdc05f4, 32'h3cd4e8c8} /* (20, 13, 24) {real, imag} */,
  {32'hbd092fdf, 32'h3df08a3a} /* (20, 13, 23) {real, imag} */,
  {32'hbd9f4419, 32'hbbd9cbd0} /* (20, 13, 22) {real, imag} */,
  {32'h3d3a1c83, 32'h3d9c66ac} /* (20, 13, 21) {real, imag} */,
  {32'h3d43d776, 32'hbcb2de29} /* (20, 13, 20) {real, imag} */,
  {32'hbd2288f8, 32'hbb215050} /* (20, 13, 19) {real, imag} */,
  {32'hbcb3f61e, 32'hbd33c3d3} /* (20, 13, 18) {real, imag} */,
  {32'h3bd7bc88, 32'hbc261ce8} /* (20, 13, 17) {real, imag} */,
  {32'h3cf025c6, 32'h00000000} /* (20, 13, 16) {real, imag} */,
  {32'h3bd7bc88, 32'h3c261ce8} /* (20, 13, 15) {real, imag} */,
  {32'hbcb3f61e, 32'h3d33c3d3} /* (20, 13, 14) {real, imag} */,
  {32'hbd2288f8, 32'h3b215050} /* (20, 13, 13) {real, imag} */,
  {32'h3d43d776, 32'h3cb2de29} /* (20, 13, 12) {real, imag} */,
  {32'h3d3a1c83, 32'hbd9c66ac} /* (20, 13, 11) {real, imag} */,
  {32'hbd9f4419, 32'h3bd9cbd0} /* (20, 13, 10) {real, imag} */,
  {32'hbd092fdf, 32'hbdf08a3a} /* (20, 13, 9) {real, imag} */,
  {32'h3bdc05f4, 32'hbcd4e8c8} /* (20, 13, 8) {real, imag} */,
  {32'h3e00dc35, 32'h3c90dd66} /* (20, 13, 7) {real, imag} */,
  {32'h3d4c3225, 32'hbcf21c6b} /* (20, 13, 6) {real, imag} */,
  {32'hbe8306dd, 32'hbe400d53} /* (20, 13, 5) {real, imag} */,
  {32'h3e80063a, 32'h3cb8d43c} /* (20, 13, 4) {real, imag} */,
  {32'hbccb8412, 32'h3e2cd8a2} /* (20, 13, 3) {real, imag} */,
  {32'hbfb3e6c1, 32'hbea8d8fa} /* (20, 13, 2) {real, imag} */,
  {32'h404fb1af, 32'h3e3fb158} /* (20, 13, 1) {real, imag} */,
  {32'h401b4b16, 32'h00000000} /* (20, 13, 0) {real, imag} */,
  {32'h40134f91, 32'h3e1c064c} /* (20, 12, 31) {real, imag} */,
  {32'hbf8f613c, 32'h3e9a0cce} /* (20, 12, 30) {real, imag} */,
  {32'h3df8eb0f, 32'hbe3c99f2} /* (20, 12, 29) {real, imag} */,
  {32'h3e3183e8, 32'h3d0fc892} /* (20, 12, 28) {real, imag} */,
  {32'hbe9dc1fc, 32'h3dec828e} /* (20, 12, 27) {real, imag} */,
  {32'h3d997804, 32'h3a0039e0} /* (20, 12, 26) {real, imag} */,
  {32'hbd600d12, 32'hbe47baee} /* (20, 12, 25) {real, imag} */,
  {32'hbcb4fd3c, 32'hbd02fb1a} /* (20, 12, 24) {real, imag} */,
  {32'hbb0bcfa0, 32'h3d7d9a35} /* (20, 12, 23) {real, imag} */,
  {32'hbd1cce08, 32'hbbe9b868} /* (20, 12, 22) {real, imag} */,
  {32'h3b005728, 32'h3d91e484} /* (20, 12, 21) {real, imag} */,
  {32'hbd915ab4, 32'h3c552e67} /* (20, 12, 20) {real, imag} */,
  {32'hbb0bf176, 32'hbd719237} /* (20, 12, 19) {real, imag} */,
  {32'h3d15ddaf, 32'h3d87551a} /* (20, 12, 18) {real, imag} */,
  {32'hbc905f8d, 32'hbca84e4f} /* (20, 12, 17) {real, imag} */,
  {32'h3c341622, 32'h00000000} /* (20, 12, 16) {real, imag} */,
  {32'hbc905f8d, 32'h3ca84e4f} /* (20, 12, 15) {real, imag} */,
  {32'h3d15ddaf, 32'hbd87551a} /* (20, 12, 14) {real, imag} */,
  {32'hbb0bf176, 32'h3d719237} /* (20, 12, 13) {real, imag} */,
  {32'hbd915ab4, 32'hbc552e67} /* (20, 12, 12) {real, imag} */,
  {32'h3b005728, 32'hbd91e484} /* (20, 12, 11) {real, imag} */,
  {32'hbd1cce08, 32'h3be9b868} /* (20, 12, 10) {real, imag} */,
  {32'hbb0bcfa0, 32'hbd7d9a35} /* (20, 12, 9) {real, imag} */,
  {32'hbcb4fd3c, 32'h3d02fb1a} /* (20, 12, 8) {real, imag} */,
  {32'hbd600d12, 32'h3e47baee} /* (20, 12, 7) {real, imag} */,
  {32'h3d997804, 32'hba0039e0} /* (20, 12, 6) {real, imag} */,
  {32'hbe9dc1fc, 32'hbdec828e} /* (20, 12, 5) {real, imag} */,
  {32'h3e3183e8, 32'hbd0fc892} /* (20, 12, 4) {real, imag} */,
  {32'h3df8eb0f, 32'h3e3c99f2} /* (20, 12, 3) {real, imag} */,
  {32'hbf8f613c, 32'hbe9a0cce} /* (20, 12, 2) {real, imag} */,
  {32'h40134f91, 32'hbe1c064c} /* (20, 12, 1) {real, imag} */,
  {32'h3fd59810, 32'h00000000} /* (20, 12, 0) {real, imag} */,
  {32'h3f835a4e, 32'h3ecc9598} /* (20, 11, 31) {real, imag} */,
  {32'hbf294aec, 32'hbdb88f8a} /* (20, 11, 30) {real, imag} */,
  {32'h3c9ab0c3, 32'hbda56c40} /* (20, 11, 29) {real, imag} */,
  {32'h3e03e8ea, 32'hbd2c7606} /* (20, 11, 28) {real, imag} */,
  {32'hbe57e4d3, 32'h3e0d2ca5} /* (20, 11, 27) {real, imag} */,
  {32'hbccb92d0, 32'h3d2d02b2} /* (20, 11, 26) {real, imag} */,
  {32'h3d5d7328, 32'h3c02eebc} /* (20, 11, 25) {real, imag} */,
  {32'hbe043dd0, 32'hbda1e5f2} /* (20, 11, 24) {real, imag} */,
  {32'hbde4f9dd, 32'hbd8d1164} /* (20, 11, 23) {real, imag} */,
  {32'h3cd1ff84, 32'h3ca834d6} /* (20, 11, 22) {real, imag} */,
  {32'hbd17f68f, 32'h3cce772d} /* (20, 11, 21) {real, imag} */,
  {32'h3d97f033, 32'h3d2c6a47} /* (20, 11, 20) {real, imag} */,
  {32'hbd3ff89a, 32'h3cf7a73c} /* (20, 11, 19) {real, imag} */,
  {32'hbc12df64, 32'h3a9ebb40} /* (20, 11, 18) {real, imag} */,
  {32'h3d0bf9b4, 32'h3bac057a} /* (20, 11, 17) {real, imag} */,
  {32'hbc190dc8, 32'h00000000} /* (20, 11, 16) {real, imag} */,
  {32'h3d0bf9b4, 32'hbbac057a} /* (20, 11, 15) {real, imag} */,
  {32'hbc12df64, 32'hba9ebb40} /* (20, 11, 14) {real, imag} */,
  {32'hbd3ff89a, 32'hbcf7a73c} /* (20, 11, 13) {real, imag} */,
  {32'h3d97f033, 32'hbd2c6a47} /* (20, 11, 12) {real, imag} */,
  {32'hbd17f68f, 32'hbcce772d} /* (20, 11, 11) {real, imag} */,
  {32'h3cd1ff84, 32'hbca834d6} /* (20, 11, 10) {real, imag} */,
  {32'hbde4f9dd, 32'h3d8d1164} /* (20, 11, 9) {real, imag} */,
  {32'hbe043dd0, 32'h3da1e5f2} /* (20, 11, 8) {real, imag} */,
  {32'h3d5d7328, 32'hbc02eebc} /* (20, 11, 7) {real, imag} */,
  {32'hbccb92d0, 32'hbd2d02b2} /* (20, 11, 6) {real, imag} */,
  {32'hbe57e4d3, 32'hbe0d2ca5} /* (20, 11, 5) {real, imag} */,
  {32'h3e03e8ea, 32'h3d2c7606} /* (20, 11, 4) {real, imag} */,
  {32'h3c9ab0c3, 32'h3da56c40} /* (20, 11, 3) {real, imag} */,
  {32'hbf294aec, 32'h3db88f8a} /* (20, 11, 2) {real, imag} */,
  {32'h3f835a4e, 32'hbecc9598} /* (20, 11, 1) {real, imag} */,
  {32'h3f401980, 32'h00000000} /* (20, 11, 0) {real, imag} */,
  {32'hbf50a6b0, 32'h3f2fe9bc} /* (20, 10, 31) {real, imag} */,
  {32'h3e5d4704, 32'hbe644b56} /* (20, 10, 30) {real, imag} */,
  {32'hbcca43ee, 32'hbdda1272} /* (20, 10, 29) {real, imag} */,
  {32'h3de60bcb, 32'hbd3d6c0c} /* (20, 10, 28) {real, imag} */,
  {32'h3c3c4280, 32'hbd15abc0} /* (20, 10, 27) {real, imag} */,
  {32'h3cff8bcc, 32'hbd54fb56} /* (20, 10, 26) {real, imag} */,
  {32'hbccd4bc0, 32'h3dc0aaf4} /* (20, 10, 25) {real, imag} */,
  {32'h3dd08b1c, 32'hbd257c50} /* (20, 10, 24) {real, imag} */,
  {32'h3dbaee3c, 32'hbb967da8} /* (20, 10, 23) {real, imag} */,
  {32'h3d390a8c, 32'h3da01aaa} /* (20, 10, 22) {real, imag} */,
  {32'hbdd4a402, 32'h3dada9ee} /* (20, 10, 21) {real, imag} */,
  {32'hbb7dcb20, 32'hbd8a53fc} /* (20, 10, 20) {real, imag} */,
  {32'hbc8b1dde, 32'h3d772c26} /* (20, 10, 19) {real, imag} */,
  {32'hbbe0669a, 32'h3d0a6832} /* (20, 10, 18) {real, imag} */,
  {32'hbd45515a, 32'hbbba87c0} /* (20, 10, 17) {real, imag} */,
  {32'hbd84d1a8, 32'h00000000} /* (20, 10, 16) {real, imag} */,
  {32'hbd45515a, 32'h3bba87c0} /* (20, 10, 15) {real, imag} */,
  {32'hbbe0669a, 32'hbd0a6832} /* (20, 10, 14) {real, imag} */,
  {32'hbc8b1dde, 32'hbd772c26} /* (20, 10, 13) {real, imag} */,
  {32'hbb7dcb20, 32'h3d8a53fc} /* (20, 10, 12) {real, imag} */,
  {32'hbdd4a402, 32'hbdada9ee} /* (20, 10, 11) {real, imag} */,
  {32'h3d390a8c, 32'hbda01aaa} /* (20, 10, 10) {real, imag} */,
  {32'h3dbaee3c, 32'h3b967da8} /* (20, 10, 9) {real, imag} */,
  {32'h3dd08b1c, 32'h3d257c50} /* (20, 10, 8) {real, imag} */,
  {32'hbccd4bc0, 32'hbdc0aaf4} /* (20, 10, 7) {real, imag} */,
  {32'h3cff8bcc, 32'h3d54fb56} /* (20, 10, 6) {real, imag} */,
  {32'h3c3c4280, 32'h3d15abc0} /* (20, 10, 5) {real, imag} */,
  {32'h3de60bcb, 32'h3d3d6c0c} /* (20, 10, 4) {real, imag} */,
  {32'hbcca43ee, 32'h3dda1272} /* (20, 10, 3) {real, imag} */,
  {32'h3e5d4704, 32'h3e644b56} /* (20, 10, 2) {real, imag} */,
  {32'hbf50a6b0, 32'hbf2fe9bc} /* (20, 10, 1) {real, imag} */,
  {32'hbf58451b, 32'h00000000} /* (20, 10, 0) {real, imag} */,
  {32'hc00a67a4, 32'h3f86fd42} /* (20, 9, 31) {real, imag} */,
  {32'h3f4f2eae, 32'hbe92eb16} /* (20, 9, 30) {real, imag} */,
  {32'hbd388fb0, 32'h3ccfa560} /* (20, 9, 29) {real, imag} */,
  {32'hbd811694, 32'h3c6d2b08} /* (20, 9, 28) {real, imag} */,
  {32'h3ddbb7a6, 32'hbdc5720e} /* (20, 9, 27) {real, imag} */,
  {32'hbdb3d220, 32'hbd060945} /* (20, 9, 26) {real, imag} */,
  {32'hbd5b022a, 32'h3d8db748} /* (20, 9, 25) {real, imag} */,
  {32'hbc2cc968, 32'hbd9f2ae8} /* (20, 9, 24) {real, imag} */,
  {32'h3d64cf3b, 32'h3d8471c0} /* (20, 9, 23) {real, imag} */,
  {32'h3cb34898, 32'hbb24c848} /* (20, 9, 22) {real, imag} */,
  {32'h3c684ada, 32'hbd3f15e2} /* (20, 9, 21) {real, imag} */,
  {32'hbdae036f, 32'hbc099078} /* (20, 9, 20) {real, imag} */,
  {32'h3c4b21eb, 32'hbcf16c44} /* (20, 9, 19) {real, imag} */,
  {32'h3d14c82c, 32'hbcc334fe} /* (20, 9, 18) {real, imag} */,
  {32'hbd8548b6, 32'hbccd570c} /* (20, 9, 17) {real, imag} */,
  {32'h3ce3b080, 32'h00000000} /* (20, 9, 16) {real, imag} */,
  {32'hbd8548b6, 32'h3ccd570c} /* (20, 9, 15) {real, imag} */,
  {32'h3d14c82c, 32'h3cc334fe} /* (20, 9, 14) {real, imag} */,
  {32'h3c4b21eb, 32'h3cf16c44} /* (20, 9, 13) {real, imag} */,
  {32'hbdae036f, 32'h3c099078} /* (20, 9, 12) {real, imag} */,
  {32'h3c684ada, 32'h3d3f15e2} /* (20, 9, 11) {real, imag} */,
  {32'h3cb34898, 32'h3b24c848} /* (20, 9, 10) {real, imag} */,
  {32'h3d64cf3b, 32'hbd8471c0} /* (20, 9, 9) {real, imag} */,
  {32'hbc2cc968, 32'h3d9f2ae8} /* (20, 9, 8) {real, imag} */,
  {32'hbd5b022a, 32'hbd8db748} /* (20, 9, 7) {real, imag} */,
  {32'hbdb3d220, 32'h3d060945} /* (20, 9, 6) {real, imag} */,
  {32'h3ddbb7a6, 32'h3dc5720e} /* (20, 9, 5) {real, imag} */,
  {32'hbd811694, 32'hbc6d2b08} /* (20, 9, 4) {real, imag} */,
  {32'hbd388fb0, 32'hbccfa560} /* (20, 9, 3) {real, imag} */,
  {32'h3f4f2eae, 32'h3e92eb16} /* (20, 9, 2) {real, imag} */,
  {32'hc00a67a4, 32'hbf86fd42} /* (20, 9, 1) {real, imag} */,
  {32'hc00729cd, 32'h00000000} /* (20, 9, 0) {real, imag} */,
  {32'hc0457701, 32'h3fc9462d} /* (20, 8, 31) {real, imag} */,
  {32'h3f85fa8a, 32'hbef96f7d} /* (20, 8, 30) {real, imag} */,
  {32'hbde0086d, 32'h3d032dfb} /* (20, 8, 29) {real, imag} */,
  {32'hbd0ddfa4, 32'h3c9a4069} /* (20, 8, 28) {real, imag} */,
  {32'h3df34682, 32'hbcaa3f1c} /* (20, 8, 27) {real, imag} */,
  {32'hbde53e34, 32'hbdf07234} /* (20, 8, 26) {real, imag} */,
  {32'h3ca48fc5, 32'h3e5986b6} /* (20, 8, 25) {real, imag} */,
  {32'h3caa812b, 32'hbe3924e4} /* (20, 8, 24) {real, imag} */,
  {32'hbd961d33, 32'hbd4e9ae1} /* (20, 8, 23) {real, imag} */,
  {32'hbd9744d6, 32'h3c99f18a} /* (20, 8, 22) {real, imag} */,
  {32'hbc897519, 32'hbcc10eb2} /* (20, 8, 21) {real, imag} */,
  {32'h3cc3820e, 32'hbcad55e0} /* (20, 8, 20) {real, imag} */,
  {32'h3dd295d3, 32'hbc4a71b8} /* (20, 8, 19) {real, imag} */,
  {32'h3cd1a4de, 32'hbcc39e23} /* (20, 8, 18) {real, imag} */,
  {32'h3cccb20d, 32'h3d69f571} /* (20, 8, 17) {real, imag} */,
  {32'hbcc481e3, 32'h00000000} /* (20, 8, 16) {real, imag} */,
  {32'h3cccb20d, 32'hbd69f571} /* (20, 8, 15) {real, imag} */,
  {32'h3cd1a4de, 32'h3cc39e23} /* (20, 8, 14) {real, imag} */,
  {32'h3dd295d3, 32'h3c4a71b8} /* (20, 8, 13) {real, imag} */,
  {32'h3cc3820e, 32'h3cad55e0} /* (20, 8, 12) {real, imag} */,
  {32'hbc897519, 32'h3cc10eb2} /* (20, 8, 11) {real, imag} */,
  {32'hbd9744d6, 32'hbc99f18a} /* (20, 8, 10) {real, imag} */,
  {32'hbd961d33, 32'h3d4e9ae1} /* (20, 8, 9) {real, imag} */,
  {32'h3caa812b, 32'h3e3924e4} /* (20, 8, 8) {real, imag} */,
  {32'h3ca48fc5, 32'hbe5986b6} /* (20, 8, 7) {real, imag} */,
  {32'hbde53e34, 32'h3df07234} /* (20, 8, 6) {real, imag} */,
  {32'h3df34682, 32'h3caa3f1c} /* (20, 8, 5) {real, imag} */,
  {32'hbd0ddfa4, 32'hbc9a4069} /* (20, 8, 4) {real, imag} */,
  {32'hbde0086d, 32'hbd032dfb} /* (20, 8, 3) {real, imag} */,
  {32'h3f85fa8a, 32'h3ef96f7d} /* (20, 8, 2) {real, imag} */,
  {32'hc0457701, 32'hbfc9462d} /* (20, 8, 1) {real, imag} */,
  {32'hc046e5c6, 32'h00000000} /* (20, 8, 0) {real, imag} */,
  {32'hc06b697f, 32'h3ff8227e} /* (20, 7, 31) {real, imag} */,
  {32'h3f80347d, 32'hbf0eb10b} /* (20, 7, 30) {real, imag} */,
  {32'hbca05e9c, 32'hbe0cdef6} /* (20, 7, 29) {real, imag} */,
  {32'hbd268188, 32'h3d56f456} /* (20, 7, 28) {real, imag} */,
  {32'h3e846a0c, 32'hbcfe4da0} /* (20, 7, 27) {real, imag} */,
  {32'h3cc0f902, 32'hbd8534a6} /* (20, 7, 26) {real, imag} */,
  {32'h3cd7e577, 32'h3d7abad1} /* (20, 7, 25) {real, imag} */,
  {32'h3dbe31a2, 32'hbe2d64b0} /* (20, 7, 24) {real, imag} */,
  {32'hbd821945, 32'h3d2206cf} /* (20, 7, 23) {real, imag} */,
  {32'h3cc9fcdb, 32'hbd1de380} /* (20, 7, 22) {real, imag} */,
  {32'h3c77a620, 32'hbcdb8a27} /* (20, 7, 21) {real, imag} */,
  {32'hbd175042, 32'h3dd26283} /* (20, 7, 20) {real, imag} */,
  {32'h3ca22f7a, 32'hbd603e52} /* (20, 7, 19) {real, imag} */,
  {32'hbc7bb2fe, 32'h3d573d9f} /* (20, 7, 18) {real, imag} */,
  {32'h3c560274, 32'hbdbe3158} /* (20, 7, 17) {real, imag} */,
  {32'h3ac7b2b0, 32'h00000000} /* (20, 7, 16) {real, imag} */,
  {32'h3c560274, 32'h3dbe3158} /* (20, 7, 15) {real, imag} */,
  {32'hbc7bb2fe, 32'hbd573d9f} /* (20, 7, 14) {real, imag} */,
  {32'h3ca22f7a, 32'h3d603e52} /* (20, 7, 13) {real, imag} */,
  {32'hbd175042, 32'hbdd26283} /* (20, 7, 12) {real, imag} */,
  {32'h3c77a620, 32'h3cdb8a27} /* (20, 7, 11) {real, imag} */,
  {32'h3cc9fcdb, 32'h3d1de380} /* (20, 7, 10) {real, imag} */,
  {32'hbd821945, 32'hbd2206cf} /* (20, 7, 9) {real, imag} */,
  {32'h3dbe31a2, 32'h3e2d64b0} /* (20, 7, 8) {real, imag} */,
  {32'h3cd7e577, 32'hbd7abad1} /* (20, 7, 7) {real, imag} */,
  {32'h3cc0f902, 32'h3d8534a6} /* (20, 7, 6) {real, imag} */,
  {32'h3e846a0c, 32'h3cfe4da0} /* (20, 7, 5) {real, imag} */,
  {32'hbd268188, 32'hbd56f456} /* (20, 7, 4) {real, imag} */,
  {32'hbca05e9c, 32'h3e0cdef6} /* (20, 7, 3) {real, imag} */,
  {32'h3f80347d, 32'h3f0eb10b} /* (20, 7, 2) {real, imag} */,
  {32'hc06b697f, 32'hbff8227e} /* (20, 7, 1) {real, imag} */,
  {32'hc0722bee, 32'h00000000} /* (20, 7, 0) {real, imag} */,
  {32'hc0731306, 32'h4019b901} /* (20, 6, 31) {real, imag} */,
  {32'h3f491a31, 32'hbf2fbd16} /* (20, 6, 30) {real, imag} */,
  {32'h3ab953c0, 32'h3d4d60a6} /* (20, 6, 29) {real, imag} */,
  {32'hbd276140, 32'hbd1b0eae} /* (20, 6, 28) {real, imag} */,
  {32'h3e88c814, 32'h3cc9e288} /* (20, 6, 27) {real, imag} */,
  {32'h3c31ed97, 32'hbc5adb68} /* (20, 6, 26) {real, imag} */,
  {32'hbdd196d0, 32'h3d4d0969} /* (20, 6, 25) {real, imag} */,
  {32'h3c010814, 32'hbd3f179e} /* (20, 6, 24) {real, imag} */,
  {32'hbd970194, 32'h3e016077} /* (20, 6, 23) {real, imag} */,
  {32'h3d47c0a1, 32'hbd45e77c} /* (20, 6, 22) {real, imag} */,
  {32'h3d5c3fac, 32'h3ccedda3} /* (20, 6, 21) {real, imag} */,
  {32'hbb22b080, 32'hbd01d7c4} /* (20, 6, 20) {real, imag} */,
  {32'h3c5ef3fe, 32'hbcfbd42c} /* (20, 6, 19) {real, imag} */,
  {32'h3cae49bc, 32'h3da61262} /* (20, 6, 18) {real, imag} */,
  {32'h3c71a82d, 32'h3b946e2e} /* (20, 6, 17) {real, imag} */,
  {32'h3caba05b, 32'h00000000} /* (20, 6, 16) {real, imag} */,
  {32'h3c71a82d, 32'hbb946e2e} /* (20, 6, 15) {real, imag} */,
  {32'h3cae49bc, 32'hbda61262} /* (20, 6, 14) {real, imag} */,
  {32'h3c5ef3fe, 32'h3cfbd42c} /* (20, 6, 13) {real, imag} */,
  {32'hbb22b080, 32'h3d01d7c4} /* (20, 6, 12) {real, imag} */,
  {32'h3d5c3fac, 32'hbccedda3} /* (20, 6, 11) {real, imag} */,
  {32'h3d47c0a1, 32'h3d45e77c} /* (20, 6, 10) {real, imag} */,
  {32'hbd970194, 32'hbe016077} /* (20, 6, 9) {real, imag} */,
  {32'h3c010814, 32'h3d3f179e} /* (20, 6, 8) {real, imag} */,
  {32'hbdd196d0, 32'hbd4d0969} /* (20, 6, 7) {real, imag} */,
  {32'h3c31ed97, 32'h3c5adb68} /* (20, 6, 6) {real, imag} */,
  {32'h3e88c814, 32'hbcc9e288} /* (20, 6, 5) {real, imag} */,
  {32'hbd276140, 32'h3d1b0eae} /* (20, 6, 4) {real, imag} */,
  {32'h3ab953c0, 32'hbd4d60a6} /* (20, 6, 3) {real, imag} */,
  {32'h3f491a31, 32'h3f2fbd16} /* (20, 6, 2) {real, imag} */,
  {32'hc0731306, 32'hc019b901} /* (20, 6, 1) {real, imag} */,
  {32'hc083cbcb, 32'h00000000} /* (20, 6, 0) {real, imag} */,
  {32'hc06bef1d, 32'h4047c3d0} /* (20, 5, 31) {real, imag} */,
  {32'h3e9f980c, 32'hbf534b44} /* (20, 5, 30) {real, imag} */,
  {32'h3d6f42fc, 32'hbdb33d12} /* (20, 5, 29) {real, imag} */,
  {32'h3dcad0ed, 32'hbe38a062} /* (20, 5, 28) {real, imag} */,
  {32'h3e55ca3f, 32'h3d492eb3} /* (20, 5, 27) {real, imag} */,
  {32'h3db3b76b, 32'h3df31c44} /* (20, 5, 26) {real, imag} */,
  {32'hbd13fe08, 32'h3d98adda} /* (20, 5, 25) {real, imag} */,
  {32'hba9e9fa0, 32'hbd43b22a} /* (20, 5, 24) {real, imag} */,
  {32'h3d398567, 32'h3c23132c} /* (20, 5, 23) {real, imag} */,
  {32'hbd8b6b36, 32'hbdced4ca} /* (20, 5, 22) {real, imag} */,
  {32'hbdd50a8a, 32'hbd0aba27} /* (20, 5, 21) {real, imag} */,
  {32'hbcc619a6, 32'hbd34c726} /* (20, 5, 20) {real, imag} */,
  {32'hbd5fa118, 32'h3c03692c} /* (20, 5, 19) {real, imag} */,
  {32'h3dc63796, 32'hbd929b09} /* (20, 5, 18) {real, imag} */,
  {32'h3d8d3a97, 32'h3ce9014a} /* (20, 5, 17) {real, imag} */,
  {32'h3d88c66e, 32'h00000000} /* (20, 5, 16) {real, imag} */,
  {32'h3d8d3a97, 32'hbce9014a} /* (20, 5, 15) {real, imag} */,
  {32'h3dc63796, 32'h3d929b09} /* (20, 5, 14) {real, imag} */,
  {32'hbd5fa118, 32'hbc03692c} /* (20, 5, 13) {real, imag} */,
  {32'hbcc619a6, 32'h3d34c726} /* (20, 5, 12) {real, imag} */,
  {32'hbdd50a8a, 32'h3d0aba27} /* (20, 5, 11) {real, imag} */,
  {32'hbd8b6b36, 32'h3dced4ca} /* (20, 5, 10) {real, imag} */,
  {32'h3d398567, 32'hbc23132c} /* (20, 5, 9) {real, imag} */,
  {32'hba9e9fa0, 32'h3d43b22a} /* (20, 5, 8) {real, imag} */,
  {32'hbd13fe08, 32'hbd98adda} /* (20, 5, 7) {real, imag} */,
  {32'h3db3b76b, 32'hbdf31c44} /* (20, 5, 6) {real, imag} */,
  {32'h3e55ca3f, 32'hbd492eb3} /* (20, 5, 5) {real, imag} */,
  {32'h3dcad0ed, 32'h3e38a062} /* (20, 5, 4) {real, imag} */,
  {32'h3d6f42fc, 32'h3db33d12} /* (20, 5, 3) {real, imag} */,
  {32'h3e9f980c, 32'h3f534b44} /* (20, 5, 2) {real, imag} */,
  {32'hc06bef1d, 32'hc047c3d0} /* (20, 5, 1) {real, imag} */,
  {32'hc09025f4, 32'h00000000} /* (20, 5, 0) {real, imag} */,
  {32'hc05d4e0c, 32'h40702e38} /* (20, 4, 31) {real, imag} */,
  {32'hbe28390c, 32'hbf7a9df2} /* (20, 4, 30) {real, imag} */,
  {32'h3d8dea14, 32'hbe71b47e} /* (20, 4, 29) {real, imag} */,
  {32'h3e3e78fa, 32'hbe672ae0} /* (20, 4, 28) {real, imag} */,
  {32'h3e55dc6d, 32'h3e49b2fb} /* (20, 4, 27) {real, imag} */,
  {32'h3c00f3ac, 32'h3d091ec1} /* (20, 4, 26) {real, imag} */,
  {32'hbd11c25c, 32'hbd7c704c} /* (20, 4, 25) {real, imag} */,
  {32'hbcb27c96, 32'h3c6385f4} /* (20, 4, 24) {real, imag} */,
  {32'h3d429e4c, 32'h3bd65c68} /* (20, 4, 23) {real, imag} */,
  {32'h3c0fc822, 32'h3d667c27} /* (20, 4, 22) {real, imag} */,
  {32'hbd2eba4a, 32'hbd7b80a6} /* (20, 4, 21) {real, imag} */,
  {32'hbb98db7a, 32'h3c68df97} /* (20, 4, 20) {real, imag} */,
  {32'hbd5380c1, 32'h3d8a3ae8} /* (20, 4, 19) {real, imag} */,
  {32'hbc97768e, 32'hbc1e2b4f} /* (20, 4, 18) {real, imag} */,
  {32'hbb065c18, 32'hbdc6ec80} /* (20, 4, 17) {real, imag} */,
  {32'hbce9c3f7, 32'h00000000} /* (20, 4, 16) {real, imag} */,
  {32'hbb065c18, 32'h3dc6ec80} /* (20, 4, 15) {real, imag} */,
  {32'hbc97768e, 32'h3c1e2b4f} /* (20, 4, 14) {real, imag} */,
  {32'hbd5380c1, 32'hbd8a3ae8} /* (20, 4, 13) {real, imag} */,
  {32'hbb98db7a, 32'hbc68df97} /* (20, 4, 12) {real, imag} */,
  {32'hbd2eba4a, 32'h3d7b80a6} /* (20, 4, 11) {real, imag} */,
  {32'h3c0fc822, 32'hbd667c27} /* (20, 4, 10) {real, imag} */,
  {32'h3d429e4c, 32'hbbd65c68} /* (20, 4, 9) {real, imag} */,
  {32'hbcb27c96, 32'hbc6385f4} /* (20, 4, 8) {real, imag} */,
  {32'hbd11c25c, 32'h3d7c704c} /* (20, 4, 7) {real, imag} */,
  {32'h3c00f3ac, 32'hbd091ec1} /* (20, 4, 6) {real, imag} */,
  {32'h3e55dc6d, 32'hbe49b2fb} /* (20, 4, 5) {real, imag} */,
  {32'h3e3e78fa, 32'h3e672ae0} /* (20, 4, 4) {real, imag} */,
  {32'h3d8dea14, 32'h3e71b47e} /* (20, 4, 3) {real, imag} */,
  {32'hbe28390c, 32'h3f7a9df2} /* (20, 4, 2) {real, imag} */,
  {32'hc05d4e0c, 32'hc0702e38} /* (20, 4, 1) {real, imag} */,
  {32'hc0987be6, 32'h00000000} /* (20, 4, 0) {real, imag} */,
  {32'hc050db8a, 32'h407e9913} /* (20, 3, 31) {real, imag} */,
  {32'hbedad868, 32'hbf9a8313} /* (20, 3, 30) {real, imag} */,
  {32'h3c0c7c64, 32'hbe44e81e} /* (20, 3, 29) {real, imag} */,
  {32'h3e1eebfa, 32'hbe8599a8} /* (20, 3, 28) {real, imag} */,
  {32'h3e3e6040, 32'h3e189d2c} /* (20, 3, 27) {real, imag} */,
  {32'h3cb81ca4, 32'h3d04635c} /* (20, 3, 26) {real, imag} */,
  {32'h3d744e7a, 32'hbd77f352} /* (20, 3, 25) {real, imag} */,
  {32'hbd1c3924, 32'hbdfa2f7e} /* (20, 3, 24) {real, imag} */,
  {32'h3d526489, 32'hbc219b44} /* (20, 3, 23) {real, imag} */,
  {32'h3d9f378b, 32'hbddd16d0} /* (20, 3, 22) {real, imag} */,
  {32'h3d4ec8c2, 32'h3dce0f99} /* (20, 3, 21) {real, imag} */,
  {32'hbda24422, 32'h3cf24e59} /* (20, 3, 20) {real, imag} */,
  {32'hbc432283, 32'hbd0dc37c} /* (20, 3, 19) {real, imag} */,
  {32'h3dac780b, 32'hbc940c43} /* (20, 3, 18) {real, imag} */,
  {32'h3d85b589, 32'hbc9f38a2} /* (20, 3, 17) {real, imag} */,
  {32'h3c17d4f8, 32'h00000000} /* (20, 3, 16) {real, imag} */,
  {32'h3d85b589, 32'h3c9f38a2} /* (20, 3, 15) {real, imag} */,
  {32'h3dac780b, 32'h3c940c43} /* (20, 3, 14) {real, imag} */,
  {32'hbc432283, 32'h3d0dc37c} /* (20, 3, 13) {real, imag} */,
  {32'hbda24422, 32'hbcf24e59} /* (20, 3, 12) {real, imag} */,
  {32'h3d4ec8c2, 32'hbdce0f99} /* (20, 3, 11) {real, imag} */,
  {32'h3d9f378b, 32'h3ddd16d0} /* (20, 3, 10) {real, imag} */,
  {32'h3d526489, 32'h3c219b44} /* (20, 3, 9) {real, imag} */,
  {32'hbd1c3924, 32'h3dfa2f7e} /* (20, 3, 8) {real, imag} */,
  {32'h3d744e7a, 32'h3d77f352} /* (20, 3, 7) {real, imag} */,
  {32'h3cb81ca4, 32'hbd04635c} /* (20, 3, 6) {real, imag} */,
  {32'h3e3e6040, 32'hbe189d2c} /* (20, 3, 5) {real, imag} */,
  {32'h3e1eebfa, 32'h3e8599a8} /* (20, 3, 4) {real, imag} */,
  {32'h3c0c7c64, 32'h3e44e81e} /* (20, 3, 3) {real, imag} */,
  {32'hbedad868, 32'h3f9a8313} /* (20, 3, 2) {real, imag} */,
  {32'hc050db8a, 32'hc07e9913} /* (20, 3, 1) {real, imag} */,
  {32'hc0a3e2b8, 32'h00000000} /* (20, 3, 0) {real, imag} */,
  {32'hc053ed5d, 32'h4076213e} /* (20, 2, 31) {real, imag} */,
  {32'hbe77fe48, 32'hbf8785f2} /* (20, 2, 30) {real, imag} */,
  {32'h3d472c89, 32'hbdb6aa2e} /* (20, 2, 29) {real, imag} */,
  {32'h3d858166, 32'hbe8f8087} /* (20, 2, 28) {real, imag} */,
  {32'h3e8d556f, 32'h3ce2ab3c} /* (20, 2, 27) {real, imag} */,
  {32'h3d97aa9c, 32'hbc5ddaf6} /* (20, 2, 26) {real, imag} */,
  {32'h3cbde348, 32'h3d40482c} /* (20, 2, 25) {real, imag} */,
  {32'hbd2ce320, 32'h3d31d62e} /* (20, 2, 24) {real, imag} */,
  {32'h3d46dd62, 32'hbc6e4518} /* (20, 2, 23) {real, imag} */,
  {32'hbb82d158, 32'hbd5c58b4} /* (20, 2, 22) {real, imag} */,
  {32'hba7dd620, 32'hbb89b5d4} /* (20, 2, 21) {real, imag} */,
  {32'hbcc00d12, 32'hbdb87de3} /* (20, 2, 20) {real, imag} */,
  {32'h3d07ced8, 32'hbceb256d} /* (20, 2, 19) {real, imag} */,
  {32'hbd36f220, 32'h3b2127a8} /* (20, 2, 18) {real, imag} */,
  {32'h3ce964ad, 32'hbd05938e} /* (20, 2, 17) {real, imag} */,
  {32'hbc8790d5, 32'h00000000} /* (20, 2, 16) {real, imag} */,
  {32'h3ce964ad, 32'h3d05938e} /* (20, 2, 15) {real, imag} */,
  {32'hbd36f220, 32'hbb2127a8} /* (20, 2, 14) {real, imag} */,
  {32'h3d07ced8, 32'h3ceb256d} /* (20, 2, 13) {real, imag} */,
  {32'hbcc00d12, 32'h3db87de3} /* (20, 2, 12) {real, imag} */,
  {32'hba7dd620, 32'h3b89b5d4} /* (20, 2, 11) {real, imag} */,
  {32'hbb82d158, 32'h3d5c58b4} /* (20, 2, 10) {real, imag} */,
  {32'h3d46dd62, 32'h3c6e4518} /* (20, 2, 9) {real, imag} */,
  {32'hbd2ce320, 32'hbd31d62e} /* (20, 2, 8) {real, imag} */,
  {32'h3cbde348, 32'hbd40482c} /* (20, 2, 7) {real, imag} */,
  {32'h3d97aa9c, 32'h3c5ddaf6} /* (20, 2, 6) {real, imag} */,
  {32'h3e8d556f, 32'hbce2ab3c} /* (20, 2, 5) {real, imag} */,
  {32'h3d858166, 32'h3e8f8087} /* (20, 2, 4) {real, imag} */,
  {32'h3d472c89, 32'h3db6aa2e} /* (20, 2, 3) {real, imag} */,
  {32'hbe77fe48, 32'h3f8785f2} /* (20, 2, 2) {real, imag} */,
  {32'hc053ed5d, 32'hc076213e} /* (20, 2, 1) {real, imag} */,
  {32'hc0aa6a7a, 32'h00000000} /* (20, 2, 0) {real, imag} */,
  {32'hc05d390c, 32'h40625f2e} /* (20, 1, 31) {real, imag} */,
  {32'hbdee8c68, 32'hbf6c5aec} /* (20, 1, 30) {real, imag} */,
  {32'h3e25749a, 32'hbdd83578} /* (20, 1, 29) {real, imag} */,
  {32'h3e28fe0d, 32'hbe8e2907} /* (20, 1, 28) {real, imag} */,
  {32'h3e4acdaf, 32'h3d914d3d} /* (20, 1, 27) {real, imag} */,
  {32'h3def522a, 32'hbd94bb97} /* (20, 1, 26) {real, imag} */,
  {32'hbe067315, 32'h3dad8828} /* (20, 1, 25) {real, imag} */,
  {32'hbdd309d4, 32'h3d5a6b26} /* (20, 1, 24) {real, imag} */,
  {32'hbd9b6558, 32'h3d034e92} /* (20, 1, 23) {real, imag} */,
  {32'h3d2150d3, 32'hbe407668} /* (20, 1, 22) {real, imag} */,
  {32'h3d342b10, 32'hbcf71236} /* (20, 1, 21) {real, imag} */,
  {32'h3cc6e7e9, 32'h3d4f215c} /* (20, 1, 20) {real, imag} */,
  {32'hbc344a80, 32'hbd01f76b} /* (20, 1, 19) {real, imag} */,
  {32'hbc23f567, 32'hbd03b192} /* (20, 1, 18) {real, imag} */,
  {32'hbc64d20c, 32'hbcc3a13c} /* (20, 1, 17) {real, imag} */,
  {32'hbc910a46, 32'h00000000} /* (20, 1, 16) {real, imag} */,
  {32'hbc64d20c, 32'h3cc3a13c} /* (20, 1, 15) {real, imag} */,
  {32'hbc23f567, 32'h3d03b192} /* (20, 1, 14) {real, imag} */,
  {32'hbc344a80, 32'h3d01f76b} /* (20, 1, 13) {real, imag} */,
  {32'h3cc6e7e9, 32'hbd4f215c} /* (20, 1, 12) {real, imag} */,
  {32'h3d342b10, 32'h3cf71236} /* (20, 1, 11) {real, imag} */,
  {32'h3d2150d3, 32'h3e407668} /* (20, 1, 10) {real, imag} */,
  {32'hbd9b6558, 32'hbd034e92} /* (20, 1, 9) {real, imag} */,
  {32'hbdd309d4, 32'hbd5a6b26} /* (20, 1, 8) {real, imag} */,
  {32'hbe067315, 32'hbdad8828} /* (20, 1, 7) {real, imag} */,
  {32'h3def522a, 32'h3d94bb97} /* (20, 1, 6) {real, imag} */,
  {32'h3e4acdaf, 32'hbd914d3d} /* (20, 1, 5) {real, imag} */,
  {32'h3e28fe0d, 32'h3e8e2907} /* (20, 1, 4) {real, imag} */,
  {32'h3e25749a, 32'h3dd83578} /* (20, 1, 3) {real, imag} */,
  {32'hbdee8c68, 32'h3f6c5aec} /* (20, 1, 2) {real, imag} */,
  {32'hc05d390c, 32'hc0625f2e} /* (20, 1, 1) {real, imag} */,
  {32'hc0a4bfdf, 32'h00000000} /* (20, 1, 0) {real, imag} */,
  {32'hc06a6f8a, 32'h403910d2} /* (20, 0, 31) {real, imag} */,
  {32'h3e315638, 32'hbf369ede} /* (20, 0, 30) {real, imag} */,
  {32'h3e0c328b, 32'hbc692694} /* (20, 0, 29) {real, imag} */,
  {32'h3d047b80, 32'hbe18d99e} /* (20, 0, 28) {real, imag} */,
  {32'h3cc53dd0, 32'hbb623b10} /* (20, 0, 27) {real, imag} */,
  {32'hbcfcc9b7, 32'hbd8ef007} /* (20, 0, 26) {real, imag} */,
  {32'hbd9577b1, 32'h3c8a0036} /* (20, 0, 25) {real, imag} */,
  {32'hbcaaf2f5, 32'hbd8e997e} /* (20, 0, 24) {real, imag} */,
  {32'hbd3a59d1, 32'h3d83b693} /* (20, 0, 23) {real, imag} */,
  {32'hbd2b648c, 32'hbda171f0} /* (20, 0, 22) {real, imag} */,
  {32'h3c5d1d58, 32'hbb70d738} /* (20, 0, 21) {real, imag} */,
  {32'hbcacd2ce, 32'hbd34cff2} /* (20, 0, 20) {real, imag} */,
  {32'hbd28b89e, 32'hbca22f96} /* (20, 0, 19) {real, imag} */,
  {32'hbd685a26, 32'hbd192bb5} /* (20, 0, 18) {real, imag} */,
  {32'hbcee4ed3, 32'h3c650b3c} /* (20, 0, 17) {real, imag} */,
  {32'hbc84a64c, 32'h00000000} /* (20, 0, 16) {real, imag} */,
  {32'hbcee4ed3, 32'hbc650b3c} /* (20, 0, 15) {real, imag} */,
  {32'hbd685a26, 32'h3d192bb5} /* (20, 0, 14) {real, imag} */,
  {32'hbd28b89e, 32'h3ca22f96} /* (20, 0, 13) {real, imag} */,
  {32'hbcacd2ce, 32'h3d34cff2} /* (20, 0, 12) {real, imag} */,
  {32'h3c5d1d58, 32'h3b70d738} /* (20, 0, 11) {real, imag} */,
  {32'hbd2b648c, 32'h3da171f0} /* (20, 0, 10) {real, imag} */,
  {32'hbd3a59d1, 32'hbd83b693} /* (20, 0, 9) {real, imag} */,
  {32'hbcaaf2f5, 32'h3d8e997e} /* (20, 0, 8) {real, imag} */,
  {32'hbd9577b1, 32'hbc8a0036} /* (20, 0, 7) {real, imag} */,
  {32'hbcfcc9b7, 32'h3d8ef007} /* (20, 0, 6) {real, imag} */,
  {32'h3cc53dd0, 32'h3b623b10} /* (20, 0, 5) {real, imag} */,
  {32'h3d047b80, 32'h3e18d99e} /* (20, 0, 4) {real, imag} */,
  {32'h3e0c328b, 32'h3c692694} /* (20, 0, 3) {real, imag} */,
  {32'h3e315638, 32'h3f369ede} /* (20, 0, 2) {real, imag} */,
  {32'hc06a6f8a, 32'hc03910d2} /* (20, 0, 1) {real, imag} */,
  {32'hc09efb64, 32'h00000000} /* (20, 0, 0) {real, imag} */,
  {32'hc076fb87, 32'h3ffd39e8} /* (19, 31, 31) {real, imag} */,
  {32'h3f235dba, 32'hbefed87d} /* (19, 31, 30) {real, imag} */,
  {32'h3d3032f2, 32'h3cc0572a} /* (19, 31, 29) {real, imag} */,
  {32'hbd01ffe9, 32'h3aca6b80} /* (19, 31, 28) {real, imag} */,
  {32'h3d9795c1, 32'hbd9b7899} /* (19, 31, 27) {real, imag} */,
  {32'hbd48693c, 32'h3cb15064} /* (19, 31, 26) {real, imag} */,
  {32'hbd280d40, 32'h3c758820} /* (19, 31, 25) {real, imag} */,
  {32'h3d96b18f, 32'hbd32f5a6} /* (19, 31, 24) {real, imag} */,
  {32'h3dddb5b3, 32'h3ceaf9fc} /* (19, 31, 23) {real, imag} */,
  {32'h3c9efee7, 32'hbd9edebf} /* (19, 31, 22) {real, imag} */,
  {32'h3d6851c8, 32'h3c8f2d9c} /* (19, 31, 21) {real, imag} */,
  {32'hbc8dcab0, 32'hbc1ce8da} /* (19, 31, 20) {real, imag} */,
  {32'hbce392f8, 32'hbc9cdabd} /* (19, 31, 19) {real, imag} */,
  {32'h3ba14828, 32'hbc896951} /* (19, 31, 18) {real, imag} */,
  {32'hbc816777, 32'h3bd11074} /* (19, 31, 17) {real, imag} */,
  {32'hbd3b2661, 32'h00000000} /* (19, 31, 16) {real, imag} */,
  {32'hbc816777, 32'hbbd11074} /* (19, 31, 15) {real, imag} */,
  {32'h3ba14828, 32'h3c896951} /* (19, 31, 14) {real, imag} */,
  {32'hbce392f8, 32'h3c9cdabd} /* (19, 31, 13) {real, imag} */,
  {32'hbc8dcab0, 32'h3c1ce8da} /* (19, 31, 12) {real, imag} */,
  {32'h3d6851c8, 32'hbc8f2d9c} /* (19, 31, 11) {real, imag} */,
  {32'h3c9efee7, 32'h3d9edebf} /* (19, 31, 10) {real, imag} */,
  {32'h3dddb5b3, 32'hbceaf9fc} /* (19, 31, 9) {real, imag} */,
  {32'h3d96b18f, 32'h3d32f5a6} /* (19, 31, 8) {real, imag} */,
  {32'hbd280d40, 32'hbc758820} /* (19, 31, 7) {real, imag} */,
  {32'hbd48693c, 32'hbcb15064} /* (19, 31, 6) {real, imag} */,
  {32'h3d9795c1, 32'h3d9b7899} /* (19, 31, 5) {real, imag} */,
  {32'hbd01ffe9, 32'hbaca6b80} /* (19, 31, 4) {real, imag} */,
  {32'h3d3032f2, 32'hbcc0572a} /* (19, 31, 3) {real, imag} */,
  {32'h3f235dba, 32'h3efed87d} /* (19, 31, 2) {real, imag} */,
  {32'hc076fb87, 32'hbffd39e8} /* (19, 31, 1) {real, imag} */,
  {32'hc094785b, 32'h00000000} /* (19, 31, 0) {real, imag} */,
  {32'hc08d91ce, 32'h3fd6ba0c} /* (19, 30, 31) {real, imag} */,
  {32'h3f9936ee, 32'hbef272f4} /* (19, 30, 30) {real, imag} */,
  {32'h3d51c236, 32'hbc0d1b50} /* (19, 30, 29) {real, imag} */,
  {32'hbd46236b, 32'h3d129818} /* (19, 30, 28) {real, imag} */,
  {32'h3d3fc38e, 32'hbdcb0d84} /* (19, 30, 27) {real, imag} */,
  {32'h3d3d58ce, 32'h3b4ad480} /* (19, 30, 26) {real, imag} */,
  {32'h3d0fffa4, 32'h3dff5508} /* (19, 30, 25) {real, imag} */,
  {32'h3d7381e2, 32'h3c3a42d8} /* (19, 30, 24) {real, imag} */,
  {32'h3da6e160, 32'hbdee0cc0} /* (19, 30, 23) {real, imag} */,
  {32'h3bd38d48, 32'hbd5342a8} /* (19, 30, 22) {real, imag} */,
  {32'hbd830a84, 32'hbd83f030} /* (19, 30, 21) {real, imag} */,
  {32'h3cb7d902, 32'h3d1de7ba} /* (19, 30, 20) {real, imag} */,
  {32'h3d2b92cb, 32'h3d3bbcc8} /* (19, 30, 19) {real, imag} */,
  {32'hbbb2534f, 32'hbd6e35e2} /* (19, 30, 18) {real, imag} */,
  {32'hbd6271ee, 32'hbd26eed3} /* (19, 30, 17) {real, imag} */,
  {32'h3d645f63, 32'h00000000} /* (19, 30, 16) {real, imag} */,
  {32'hbd6271ee, 32'h3d26eed3} /* (19, 30, 15) {real, imag} */,
  {32'hbbb2534f, 32'h3d6e35e2} /* (19, 30, 14) {real, imag} */,
  {32'h3d2b92cb, 32'hbd3bbcc8} /* (19, 30, 13) {real, imag} */,
  {32'h3cb7d902, 32'hbd1de7ba} /* (19, 30, 12) {real, imag} */,
  {32'hbd830a84, 32'h3d83f030} /* (19, 30, 11) {real, imag} */,
  {32'h3bd38d48, 32'h3d5342a8} /* (19, 30, 10) {real, imag} */,
  {32'h3da6e160, 32'h3dee0cc0} /* (19, 30, 9) {real, imag} */,
  {32'h3d7381e2, 32'hbc3a42d8} /* (19, 30, 8) {real, imag} */,
  {32'h3d0fffa4, 32'hbdff5508} /* (19, 30, 7) {real, imag} */,
  {32'h3d3d58ce, 32'hbb4ad480} /* (19, 30, 6) {real, imag} */,
  {32'h3d3fc38e, 32'h3dcb0d84} /* (19, 30, 5) {real, imag} */,
  {32'hbd46236b, 32'hbd129818} /* (19, 30, 4) {real, imag} */,
  {32'h3d51c236, 32'h3c0d1b50} /* (19, 30, 3) {real, imag} */,
  {32'h3f9936ee, 32'h3ef272f4} /* (19, 30, 2) {real, imag} */,
  {32'hc08d91ce, 32'hbfd6ba0c} /* (19, 30, 1) {real, imag} */,
  {32'hc09707b5, 32'h00000000} /* (19, 30, 0) {real, imag} */,
  {32'hc0969d16, 32'h3fa75245} /* (19, 29, 31) {real, imag} */,
  {32'h3fb89a72, 32'hbeebdd98} /* (19, 29, 30) {real, imag} */,
  {32'h3c2fd496, 32'hbd96a6ad} /* (19, 29, 29) {real, imag} */,
  {32'hbea47189, 32'h3dc918a1} /* (19, 29, 28) {real, imag} */,
  {32'h3e2182b2, 32'hbc9b1388} /* (19, 29, 27) {real, imag} */,
  {32'h3cca54ee, 32'hbdaba309} /* (19, 29, 26) {real, imag} */,
  {32'hbd8c0232, 32'hbc0b829c} /* (19, 29, 25) {real, imag} */,
  {32'h3aae3990, 32'h3dd1a966} /* (19, 29, 24) {real, imag} */,
  {32'h3cbd2fc0, 32'hbde6f89a} /* (19, 29, 23) {real, imag} */,
  {32'hbc6b0c09, 32'h3d6d1528} /* (19, 29, 22) {real, imag} */,
  {32'h3d310686, 32'hbc01744a} /* (19, 29, 21) {real, imag} */,
  {32'hbd17af6d, 32'h3c3fdb36} /* (19, 29, 20) {real, imag} */,
  {32'h3d34bfdf, 32'h3bfeda38} /* (19, 29, 19) {real, imag} */,
  {32'h3c371b3c, 32'hbda9bcd5} /* (19, 29, 18) {real, imag} */,
  {32'h3abe5ff8, 32'h3b5b9ffe} /* (19, 29, 17) {real, imag} */,
  {32'h3dbb2db0, 32'h00000000} /* (19, 29, 16) {real, imag} */,
  {32'h3abe5ff8, 32'hbb5b9ffe} /* (19, 29, 15) {real, imag} */,
  {32'h3c371b3c, 32'h3da9bcd5} /* (19, 29, 14) {real, imag} */,
  {32'h3d34bfdf, 32'hbbfeda38} /* (19, 29, 13) {real, imag} */,
  {32'hbd17af6d, 32'hbc3fdb36} /* (19, 29, 12) {real, imag} */,
  {32'h3d310686, 32'h3c01744a} /* (19, 29, 11) {real, imag} */,
  {32'hbc6b0c09, 32'hbd6d1528} /* (19, 29, 10) {real, imag} */,
  {32'h3cbd2fc0, 32'h3de6f89a} /* (19, 29, 9) {real, imag} */,
  {32'h3aae3990, 32'hbdd1a966} /* (19, 29, 8) {real, imag} */,
  {32'hbd8c0232, 32'h3c0b829c} /* (19, 29, 7) {real, imag} */,
  {32'h3cca54ee, 32'h3daba309} /* (19, 29, 6) {real, imag} */,
  {32'h3e2182b2, 32'h3c9b1388} /* (19, 29, 5) {real, imag} */,
  {32'hbea47189, 32'hbdc918a1} /* (19, 29, 4) {real, imag} */,
  {32'h3c2fd496, 32'h3d96a6ad} /* (19, 29, 3) {real, imag} */,
  {32'h3fb89a72, 32'h3eebdd98} /* (19, 29, 2) {real, imag} */,
  {32'hc0969d16, 32'hbfa75245} /* (19, 29, 1) {real, imag} */,
  {32'hc095f1d5, 32'h00000000} /* (19, 29, 0) {real, imag} */,
  {32'hc09cd23a, 32'h3f9d2dcf} /* (19, 28, 31) {real, imag} */,
  {32'h3fcf83f8, 32'hbea4066c} /* (19, 28, 30) {real, imag} */,
  {32'h3cebe6e6, 32'hbe33cdba} /* (19, 28, 29) {real, imag} */,
  {32'hbe9608c0, 32'h3d7e7fd6} /* (19, 28, 28) {real, imag} */,
  {32'h3e47af47, 32'hb9994200} /* (19, 28, 27) {real, imag} */,
  {32'h3d988034, 32'hbdf8e296} /* (19, 28, 26) {real, imag} */,
  {32'hbda877dc, 32'hbdb819ea} /* (19, 28, 25) {real, imag} */,
  {32'hbaa09d50, 32'hbd041b71} /* (19, 28, 24) {real, imag} */,
  {32'hbd883e3e, 32'h3abfb7d8} /* (19, 28, 23) {real, imag} */,
  {32'h3d322218, 32'h3dcc7918} /* (19, 28, 22) {real, imag} */,
  {32'h3c006e20, 32'hbd52978a} /* (19, 28, 21) {real, imag} */,
  {32'hbca0a315, 32'hbcf398f6} /* (19, 28, 20) {real, imag} */,
  {32'h3d6fcc85, 32'h3d934809} /* (19, 28, 19) {real, imag} */,
  {32'h3dedca07, 32'hbdfb67d1} /* (19, 28, 18) {real, imag} */,
  {32'hbd9f1e07, 32'hbc88494b} /* (19, 28, 17) {real, imag} */,
  {32'hbcdb10e0, 32'h00000000} /* (19, 28, 16) {real, imag} */,
  {32'hbd9f1e07, 32'h3c88494b} /* (19, 28, 15) {real, imag} */,
  {32'h3dedca07, 32'h3dfb67d1} /* (19, 28, 14) {real, imag} */,
  {32'h3d6fcc85, 32'hbd934809} /* (19, 28, 13) {real, imag} */,
  {32'hbca0a315, 32'h3cf398f6} /* (19, 28, 12) {real, imag} */,
  {32'h3c006e20, 32'h3d52978a} /* (19, 28, 11) {real, imag} */,
  {32'h3d322218, 32'hbdcc7918} /* (19, 28, 10) {real, imag} */,
  {32'hbd883e3e, 32'hbabfb7d8} /* (19, 28, 9) {real, imag} */,
  {32'hbaa09d50, 32'h3d041b71} /* (19, 28, 8) {real, imag} */,
  {32'hbda877dc, 32'h3db819ea} /* (19, 28, 7) {real, imag} */,
  {32'h3d988034, 32'h3df8e296} /* (19, 28, 6) {real, imag} */,
  {32'h3e47af47, 32'h39994200} /* (19, 28, 5) {real, imag} */,
  {32'hbe9608c0, 32'hbd7e7fd6} /* (19, 28, 4) {real, imag} */,
  {32'h3cebe6e6, 32'h3e33cdba} /* (19, 28, 3) {real, imag} */,
  {32'h3fcf83f8, 32'h3ea4066c} /* (19, 28, 2) {real, imag} */,
  {32'hc09cd23a, 32'hbf9d2dcf} /* (19, 28, 1) {real, imag} */,
  {32'hc099e26a, 32'h00000000} /* (19, 28, 0) {real, imag} */,
  {32'hc0991ac2, 32'h3f6c0b70} /* (19, 27, 31) {real, imag} */,
  {32'h3fdebbac, 32'hbecef1f0} /* (19, 27, 30) {real, imag} */,
  {32'hbd0b9763, 32'hbc69ace8} /* (19, 27, 29) {real, imag} */,
  {32'hbe8e6ecb, 32'h3c35ea90} /* (19, 27, 28) {real, imag} */,
  {32'h3ddd4d7a, 32'h3e17a038} /* (19, 27, 27) {real, imag} */,
  {32'h3dc451c0, 32'h3d8495f7} /* (19, 27, 26) {real, imag} */,
  {32'hbc5b6c50, 32'hbcc1caed} /* (19, 27, 25) {real, imag} */,
  {32'h3cbc78ea, 32'hbe128311} /* (19, 27, 24) {real, imag} */,
  {32'h3bfe6eb4, 32'hbc9dcc48} /* (19, 27, 23) {real, imag} */,
  {32'h3c796f34, 32'h3d5fb0ee} /* (19, 27, 22) {real, imag} */,
  {32'hba4ddfc0, 32'hbd891f1a} /* (19, 27, 21) {real, imag} */,
  {32'h3c5de8dd, 32'h3afc3db0} /* (19, 27, 20) {real, imag} */,
  {32'h3d677190, 32'hbd1a2f30} /* (19, 27, 19) {real, imag} */,
  {32'hbd46abce, 32'h3d704386} /* (19, 27, 18) {real, imag} */,
  {32'h3c58d24b, 32'h3cc72c30} /* (19, 27, 17) {real, imag} */,
  {32'h3dac5172, 32'h00000000} /* (19, 27, 16) {real, imag} */,
  {32'h3c58d24b, 32'hbcc72c30} /* (19, 27, 15) {real, imag} */,
  {32'hbd46abce, 32'hbd704386} /* (19, 27, 14) {real, imag} */,
  {32'h3d677190, 32'h3d1a2f30} /* (19, 27, 13) {real, imag} */,
  {32'h3c5de8dd, 32'hbafc3db0} /* (19, 27, 12) {real, imag} */,
  {32'hba4ddfc0, 32'h3d891f1a} /* (19, 27, 11) {real, imag} */,
  {32'h3c796f34, 32'hbd5fb0ee} /* (19, 27, 10) {real, imag} */,
  {32'h3bfe6eb4, 32'h3c9dcc48} /* (19, 27, 9) {real, imag} */,
  {32'h3cbc78ea, 32'h3e128311} /* (19, 27, 8) {real, imag} */,
  {32'hbc5b6c50, 32'h3cc1caed} /* (19, 27, 7) {real, imag} */,
  {32'h3dc451c0, 32'hbd8495f7} /* (19, 27, 6) {real, imag} */,
  {32'h3ddd4d7a, 32'hbe17a038} /* (19, 27, 5) {real, imag} */,
  {32'hbe8e6ecb, 32'hbc35ea90} /* (19, 27, 4) {real, imag} */,
  {32'hbd0b9763, 32'h3c69ace8} /* (19, 27, 3) {real, imag} */,
  {32'h3fdebbac, 32'h3ecef1f0} /* (19, 27, 2) {real, imag} */,
  {32'hc0991ac2, 32'hbf6c0b70} /* (19, 27, 1) {real, imag} */,
  {32'hc09b4138, 32'h00000000} /* (19, 27, 0) {real, imag} */,
  {32'hc0940748, 32'h3f42045b} /* (19, 26, 31) {real, imag} */,
  {32'h3fd7f53e, 32'hbef896e5} /* (19, 26, 30) {real, imag} */,
  {32'hbcc4dea4, 32'h3e06451c} /* (19, 26, 29) {real, imag} */,
  {32'hbea1d98a, 32'hbd08822b} /* (19, 26, 28) {real, imag} */,
  {32'h3e24f27c, 32'hbdb880be} /* (19, 26, 27) {real, imag} */,
  {32'hbcb2ec9e, 32'hbd5e16fe} /* (19, 26, 26) {real, imag} */,
  {32'hbd2167b4, 32'hbce274ca} /* (19, 26, 25) {real, imag} */,
  {32'hbde8023b, 32'hbd36536e} /* (19, 26, 24) {real, imag} */,
  {32'h3b8d5642, 32'hbd8ae54d} /* (19, 26, 23) {real, imag} */,
  {32'h3ce36c5d, 32'h3cefbfc4} /* (19, 26, 22) {real, imag} */,
  {32'h3d8494c5, 32'h3d966074} /* (19, 26, 21) {real, imag} */,
  {32'hbcb87756, 32'hbce215e0} /* (19, 26, 20) {real, imag} */,
  {32'h3d656234, 32'hbd89c95e} /* (19, 26, 19) {real, imag} */,
  {32'hbd8b7a0d, 32'h3aab6010} /* (19, 26, 18) {real, imag} */,
  {32'h3d1b94c2, 32'hbbef8cda} /* (19, 26, 17) {real, imag} */,
  {32'hbcd60978, 32'h00000000} /* (19, 26, 16) {real, imag} */,
  {32'h3d1b94c2, 32'h3bef8cda} /* (19, 26, 15) {real, imag} */,
  {32'hbd8b7a0d, 32'hbaab6010} /* (19, 26, 14) {real, imag} */,
  {32'h3d656234, 32'h3d89c95e} /* (19, 26, 13) {real, imag} */,
  {32'hbcb87756, 32'h3ce215e0} /* (19, 26, 12) {real, imag} */,
  {32'h3d8494c5, 32'hbd966074} /* (19, 26, 11) {real, imag} */,
  {32'h3ce36c5d, 32'hbcefbfc4} /* (19, 26, 10) {real, imag} */,
  {32'h3b8d5642, 32'h3d8ae54d} /* (19, 26, 9) {real, imag} */,
  {32'hbde8023b, 32'h3d36536e} /* (19, 26, 8) {real, imag} */,
  {32'hbd2167b4, 32'h3ce274ca} /* (19, 26, 7) {real, imag} */,
  {32'hbcb2ec9e, 32'h3d5e16fe} /* (19, 26, 6) {real, imag} */,
  {32'h3e24f27c, 32'h3db880be} /* (19, 26, 5) {real, imag} */,
  {32'hbea1d98a, 32'h3d08822b} /* (19, 26, 4) {real, imag} */,
  {32'hbcc4dea4, 32'hbe06451c} /* (19, 26, 3) {real, imag} */,
  {32'h3fd7f53e, 32'h3ef896e5} /* (19, 26, 2) {real, imag} */,
  {32'hc0940748, 32'hbf42045b} /* (19, 26, 1) {real, imag} */,
  {32'hc0969ca8, 32'h00000000} /* (19, 26, 0) {real, imag} */,
  {32'hc08bb26a, 32'h3f2ad46b} /* (19, 25, 31) {real, imag} */,
  {32'h3fcf5bda, 32'hbec1b0a3} /* (19, 25, 30) {real, imag} */,
  {32'hbda61df6, 32'h3ca8de0e} /* (19, 25, 29) {real, imag} */,
  {32'hbecbb264, 32'hbc9e8758} /* (19, 25, 28) {real, imag} */,
  {32'h3e83f70c, 32'hbe881acf} /* (19, 25, 27) {real, imag} */,
  {32'hbdf36280, 32'hbd7b56f0} /* (19, 25, 26) {real, imag} */,
  {32'h3dc5cc90, 32'h3db99f31} /* (19, 25, 25) {real, imag} */,
  {32'h3daf53c4, 32'hbd11d155} /* (19, 25, 24) {real, imag} */,
  {32'hbc639993, 32'hbe31308f} /* (19, 25, 23) {real, imag} */,
  {32'h3db01916, 32'hbbe77b20} /* (19, 25, 22) {real, imag} */,
  {32'h3c641110, 32'hbd3d9292} /* (19, 25, 21) {real, imag} */,
  {32'h3d21107e, 32'hbd550bf8} /* (19, 25, 20) {real, imag} */,
  {32'h3d9501a9, 32'h3d5a5452} /* (19, 25, 19) {real, imag} */,
  {32'hbcffb3e5, 32'hbd0f773a} /* (19, 25, 18) {real, imag} */,
  {32'h3d9102b6, 32'h3d06be8c} /* (19, 25, 17) {real, imag} */,
  {32'hbdb26dd6, 32'h00000000} /* (19, 25, 16) {real, imag} */,
  {32'h3d9102b6, 32'hbd06be8c} /* (19, 25, 15) {real, imag} */,
  {32'hbcffb3e5, 32'h3d0f773a} /* (19, 25, 14) {real, imag} */,
  {32'h3d9501a9, 32'hbd5a5452} /* (19, 25, 13) {real, imag} */,
  {32'h3d21107e, 32'h3d550bf8} /* (19, 25, 12) {real, imag} */,
  {32'h3c641110, 32'h3d3d9292} /* (19, 25, 11) {real, imag} */,
  {32'h3db01916, 32'h3be77b20} /* (19, 25, 10) {real, imag} */,
  {32'hbc639993, 32'h3e31308f} /* (19, 25, 9) {real, imag} */,
  {32'h3daf53c4, 32'h3d11d155} /* (19, 25, 8) {real, imag} */,
  {32'h3dc5cc90, 32'hbdb99f31} /* (19, 25, 7) {real, imag} */,
  {32'hbdf36280, 32'h3d7b56f0} /* (19, 25, 6) {real, imag} */,
  {32'h3e83f70c, 32'h3e881acf} /* (19, 25, 5) {real, imag} */,
  {32'hbecbb264, 32'h3c9e8758} /* (19, 25, 4) {real, imag} */,
  {32'hbda61df6, 32'hbca8de0e} /* (19, 25, 3) {real, imag} */,
  {32'h3fcf5bda, 32'h3ec1b0a3} /* (19, 25, 2) {real, imag} */,
  {32'hc08bb26a, 32'hbf2ad46b} /* (19, 25, 1) {real, imag} */,
  {32'hc0911c77, 32'h00000000} /* (19, 25, 0) {real, imag} */,
  {32'hc0744cd9, 32'h3ebd5e8c} /* (19, 24, 31) {real, imag} */,
  {32'h3fd301f9, 32'hbea1c462} /* (19, 24, 30) {real, imag} */,
  {32'hbe12aa6f, 32'hbd496de2} /* (19, 24, 29) {real, imag} */,
  {32'hbec71592, 32'h3ba99510} /* (19, 24, 28) {real, imag} */,
  {32'h3e883a66, 32'hbe21557e} /* (19, 24, 27) {real, imag} */,
  {32'h3d3d995b, 32'hbdea3105} /* (19, 24, 26) {real, imag} */,
  {32'hbd93a75a, 32'h3dfa6143} /* (19, 24, 25) {real, imag} */,
  {32'hbc032c0c, 32'hbcd05db8} /* (19, 24, 24) {real, imag} */,
  {32'h3dfec978, 32'hbcdf2cd7} /* (19, 24, 23) {real, imag} */,
  {32'hbcdc4018, 32'hbd22f45c} /* (19, 24, 22) {real, imag} */,
  {32'h3d855dda, 32'hbbee1b90} /* (19, 24, 21) {real, imag} */,
  {32'hbc92b9a6, 32'h3d511000} /* (19, 24, 20) {real, imag} */,
  {32'hbcca5400, 32'hbd97263e} /* (19, 24, 19) {real, imag} */,
  {32'hbd27491e, 32'h3b936698} /* (19, 24, 18) {real, imag} */,
  {32'hbcfadc4a, 32'h3dbf8c9d} /* (19, 24, 17) {real, imag} */,
  {32'h3df62dc0, 32'h00000000} /* (19, 24, 16) {real, imag} */,
  {32'hbcfadc4a, 32'hbdbf8c9d} /* (19, 24, 15) {real, imag} */,
  {32'hbd27491e, 32'hbb936698} /* (19, 24, 14) {real, imag} */,
  {32'hbcca5400, 32'h3d97263e} /* (19, 24, 13) {real, imag} */,
  {32'hbc92b9a6, 32'hbd511000} /* (19, 24, 12) {real, imag} */,
  {32'h3d855dda, 32'h3bee1b90} /* (19, 24, 11) {real, imag} */,
  {32'hbcdc4018, 32'h3d22f45c} /* (19, 24, 10) {real, imag} */,
  {32'h3dfec978, 32'h3cdf2cd7} /* (19, 24, 9) {real, imag} */,
  {32'hbc032c0c, 32'h3cd05db8} /* (19, 24, 8) {real, imag} */,
  {32'hbd93a75a, 32'hbdfa6143} /* (19, 24, 7) {real, imag} */,
  {32'h3d3d995b, 32'h3dea3105} /* (19, 24, 6) {real, imag} */,
  {32'h3e883a66, 32'h3e21557e} /* (19, 24, 5) {real, imag} */,
  {32'hbec71592, 32'hbba99510} /* (19, 24, 4) {real, imag} */,
  {32'hbe12aa6f, 32'h3d496de2} /* (19, 24, 3) {real, imag} */,
  {32'h3fd301f9, 32'h3ea1c462} /* (19, 24, 2) {real, imag} */,
  {32'hc0744cd9, 32'hbebd5e8c} /* (19, 24, 1) {real, imag} */,
  {32'hc07c1780, 32'h00000000} /* (19, 24, 0) {real, imag} */,
  {32'hc04b8c67, 32'h3ea63e90} /* (19, 23, 31) {real, imag} */,
  {32'h3fbe36c4, 32'hbeb8c0dd} /* (19, 23, 30) {real, imag} */,
  {32'hbe41a308, 32'hbe3f17ed} /* (19, 23, 29) {real, imag} */,
  {32'hbe81432d, 32'h3e5cd5c3} /* (19, 23, 28) {real, imag} */,
  {32'h3ea6a070, 32'hbd6778f0} /* (19, 23, 27) {real, imag} */,
  {32'hbdc4806d, 32'hbda53ddf} /* (19, 23, 26) {real, imag} */,
  {32'hbd495094, 32'h3beb3ed4} /* (19, 23, 25) {real, imag} */,
  {32'h3d165742, 32'hbdd6738e} /* (19, 23, 24) {real, imag} */,
  {32'h3d93fd33, 32'h3deb9da8} /* (19, 23, 23) {real, imag} */,
  {32'hbc192634, 32'hbd2b4f6c} /* (19, 23, 22) {real, imag} */,
  {32'h3db85053, 32'h3c947ef0} /* (19, 23, 21) {real, imag} */,
  {32'hb9d928a0, 32'h3cfefb9b} /* (19, 23, 20) {real, imag} */,
  {32'hbc568e18, 32'hbcfaf8b2} /* (19, 23, 19) {real, imag} */,
  {32'h3dcda78f, 32'hbd4dad15} /* (19, 23, 18) {real, imag} */,
  {32'hbd680bea, 32'h3c6e1a5e} /* (19, 23, 17) {real, imag} */,
  {32'h3d84a396, 32'h00000000} /* (19, 23, 16) {real, imag} */,
  {32'hbd680bea, 32'hbc6e1a5e} /* (19, 23, 15) {real, imag} */,
  {32'h3dcda78f, 32'h3d4dad15} /* (19, 23, 14) {real, imag} */,
  {32'hbc568e18, 32'h3cfaf8b2} /* (19, 23, 13) {real, imag} */,
  {32'hb9d928a0, 32'hbcfefb9b} /* (19, 23, 12) {real, imag} */,
  {32'h3db85053, 32'hbc947ef0} /* (19, 23, 11) {real, imag} */,
  {32'hbc192634, 32'h3d2b4f6c} /* (19, 23, 10) {real, imag} */,
  {32'h3d93fd33, 32'hbdeb9da8} /* (19, 23, 9) {real, imag} */,
  {32'h3d165742, 32'h3dd6738e} /* (19, 23, 8) {real, imag} */,
  {32'hbd495094, 32'hbbeb3ed4} /* (19, 23, 7) {real, imag} */,
  {32'hbdc4806d, 32'h3da53ddf} /* (19, 23, 6) {real, imag} */,
  {32'h3ea6a070, 32'h3d6778f0} /* (19, 23, 5) {real, imag} */,
  {32'hbe81432d, 32'hbe5cd5c3} /* (19, 23, 4) {real, imag} */,
  {32'hbe41a308, 32'h3e3f17ed} /* (19, 23, 3) {real, imag} */,
  {32'h3fbe36c4, 32'h3eb8c0dd} /* (19, 23, 2) {real, imag} */,
  {32'hc04b8c67, 32'hbea63e90} /* (19, 23, 1) {real, imag} */,
  {32'hc0566e1a, 32'h00000000} /* (19, 23, 0) {real, imag} */,
  {32'hc011d2e7, 32'h3e5b2428} /* (19, 22, 31) {real, imag} */,
  {32'h3f797bab, 32'hbdfe8bfa} /* (19, 22, 30) {real, imag} */,
  {32'hbe39e389, 32'h3d983d6e} /* (19, 22, 29) {real, imag} */,
  {32'hbe2e2d94, 32'hbcfbb686} /* (19, 22, 28) {real, imag} */,
  {32'h3e737156, 32'hbe5d73d9} /* (19, 22, 27) {real, imag} */,
  {32'hbd1a2ee8, 32'hbde29fd8} /* (19, 22, 26) {real, imag} */,
  {32'hbd2123d4, 32'hbc8fcdbe} /* (19, 22, 25) {real, imag} */,
  {32'h3db20b24, 32'hbd813344} /* (19, 22, 24) {real, imag} */,
  {32'hbbbc922c, 32'hbdd7c5ef} /* (19, 22, 23) {real, imag} */,
  {32'h3cc2df0e, 32'hbccc504f} /* (19, 22, 22) {real, imag} */,
  {32'hbd8ab78f, 32'hbe164ae4} /* (19, 22, 21) {real, imag} */,
  {32'h3dc2fb5a, 32'hbca83b09} /* (19, 22, 20) {real, imag} */,
  {32'hbd0ba668, 32'h3d836e55} /* (19, 22, 19) {real, imag} */,
  {32'hbcb42cbc, 32'hbcecf419} /* (19, 22, 18) {real, imag} */,
  {32'hbd4cffb4, 32'h3c8731c0} /* (19, 22, 17) {real, imag} */,
  {32'hbd8cd31a, 32'h00000000} /* (19, 22, 16) {real, imag} */,
  {32'hbd4cffb4, 32'hbc8731c0} /* (19, 22, 15) {real, imag} */,
  {32'hbcb42cbc, 32'h3cecf419} /* (19, 22, 14) {real, imag} */,
  {32'hbd0ba668, 32'hbd836e55} /* (19, 22, 13) {real, imag} */,
  {32'h3dc2fb5a, 32'h3ca83b09} /* (19, 22, 12) {real, imag} */,
  {32'hbd8ab78f, 32'h3e164ae4} /* (19, 22, 11) {real, imag} */,
  {32'h3cc2df0e, 32'h3ccc504f} /* (19, 22, 10) {real, imag} */,
  {32'hbbbc922c, 32'h3dd7c5ef} /* (19, 22, 9) {real, imag} */,
  {32'h3db20b24, 32'h3d813344} /* (19, 22, 8) {real, imag} */,
  {32'hbd2123d4, 32'h3c8fcdbe} /* (19, 22, 7) {real, imag} */,
  {32'hbd1a2ee8, 32'h3de29fd8} /* (19, 22, 6) {real, imag} */,
  {32'h3e737156, 32'h3e5d73d9} /* (19, 22, 5) {real, imag} */,
  {32'hbe2e2d94, 32'h3cfbb686} /* (19, 22, 4) {real, imag} */,
  {32'hbe39e389, 32'hbd983d6e} /* (19, 22, 3) {real, imag} */,
  {32'h3f797bab, 32'h3dfe8bfa} /* (19, 22, 2) {real, imag} */,
  {32'hc011d2e7, 32'hbe5b2428} /* (19, 22, 1) {real, imag} */,
  {32'hc025f4e9, 32'h00000000} /* (19, 22, 0) {real, imag} */,
  {32'hbf3d92b0, 32'h3db9b040} /* (19, 21, 31) {real, imag} */,
  {32'h3ed66136, 32'h3d1250e4} /* (19, 21, 30) {real, imag} */,
  {32'hbdaa6ff6, 32'h3e4a8d5c} /* (19, 21, 29) {real, imag} */,
  {32'hbdddc98d, 32'hbdee9b3b} /* (19, 21, 28) {real, imag} */,
  {32'h3d9e763c, 32'hbd92740b} /* (19, 21, 27) {real, imag} */,
  {32'h3c92396c, 32'h3c6b2a88} /* (19, 21, 26) {real, imag} */,
  {32'h3cd76d46, 32'hbcfd2761} /* (19, 21, 25) {real, imag} */,
  {32'h3d4c8a08, 32'h3c728196} /* (19, 21, 24) {real, imag} */,
  {32'h3d4a3cce, 32'h3cc42464} /* (19, 21, 23) {real, imag} */,
  {32'hbcb9fd7a, 32'hbd1ad586} /* (19, 21, 22) {real, imag} */,
  {32'hbc1450a8, 32'h3cc0f723} /* (19, 21, 21) {real, imag} */,
  {32'h3ce3a296, 32'h3d417c4a} /* (19, 21, 20) {real, imag} */,
  {32'hbc973a12, 32'hbbaf2030} /* (19, 21, 19) {real, imag} */,
  {32'hbc2ca214, 32'hbc0b1740} /* (19, 21, 18) {real, imag} */,
  {32'h3d483e96, 32'h3b1a0438} /* (19, 21, 17) {real, imag} */,
  {32'hbb7c0390, 32'h00000000} /* (19, 21, 16) {real, imag} */,
  {32'h3d483e96, 32'hbb1a0438} /* (19, 21, 15) {real, imag} */,
  {32'hbc2ca214, 32'h3c0b1740} /* (19, 21, 14) {real, imag} */,
  {32'hbc973a12, 32'h3baf2030} /* (19, 21, 13) {real, imag} */,
  {32'h3ce3a296, 32'hbd417c4a} /* (19, 21, 12) {real, imag} */,
  {32'hbc1450a8, 32'hbcc0f723} /* (19, 21, 11) {real, imag} */,
  {32'hbcb9fd7a, 32'h3d1ad586} /* (19, 21, 10) {real, imag} */,
  {32'h3d4a3cce, 32'hbcc42464} /* (19, 21, 9) {real, imag} */,
  {32'h3d4c8a08, 32'hbc728196} /* (19, 21, 8) {real, imag} */,
  {32'h3cd76d46, 32'h3cfd2761} /* (19, 21, 7) {real, imag} */,
  {32'h3c92396c, 32'hbc6b2a88} /* (19, 21, 6) {real, imag} */,
  {32'h3d9e763c, 32'h3d92740b} /* (19, 21, 5) {real, imag} */,
  {32'hbdddc98d, 32'h3dee9b3b} /* (19, 21, 4) {real, imag} */,
  {32'hbdaa6ff6, 32'hbe4a8d5c} /* (19, 21, 3) {real, imag} */,
  {32'h3ed66136, 32'hbd1250e4} /* (19, 21, 2) {real, imag} */,
  {32'hbf3d92b0, 32'hbdb9b040} /* (19, 21, 1) {real, imag} */,
  {32'hbfa06f14, 32'h00000000} /* (19, 21, 0) {real, imag} */,
  {32'h3f8f4b07, 32'hbe729aa0} /* (19, 20, 31) {real, imag} */,
  {32'hbec1062e, 32'h3e3cd662} /* (19, 20, 30) {real, imag} */,
  {32'hbde93d46, 32'h3d1f8c6c} /* (19, 20, 29) {real, imag} */,
  {32'h3e251ba0, 32'hbc892731} /* (19, 20, 28) {real, imag} */,
  {32'hbe16bef8, 32'h3e0b13d5} /* (19, 20, 27) {real, imag} */,
  {32'h3cf76758, 32'h3d481cf9} /* (19, 20, 26) {real, imag} */,
  {32'h3e02774e, 32'h3d43db6a} /* (19, 20, 25) {real, imag} */,
  {32'hbdca3a9d, 32'hbd65e677} /* (19, 20, 24) {real, imag} */,
  {32'hbd5f4bc4, 32'hbdd421bf} /* (19, 20, 23) {real, imag} */,
  {32'hbd53653a, 32'hbcad0c76} /* (19, 20, 22) {real, imag} */,
  {32'hbd1466e4, 32'h3c73b9d0} /* (19, 20, 21) {real, imag} */,
  {32'h3daa04f0, 32'hbcf1d622} /* (19, 20, 20) {real, imag} */,
  {32'h3c5dbf70, 32'h3d76c852} /* (19, 20, 19) {real, imag} */,
  {32'hbb04f1e8, 32'h3da19638} /* (19, 20, 18) {real, imag} */,
  {32'hbd3f4a9d, 32'hbd05a567} /* (19, 20, 17) {real, imag} */,
  {32'h3d816546, 32'h00000000} /* (19, 20, 16) {real, imag} */,
  {32'hbd3f4a9d, 32'h3d05a567} /* (19, 20, 15) {real, imag} */,
  {32'hbb04f1e8, 32'hbda19638} /* (19, 20, 14) {real, imag} */,
  {32'h3c5dbf70, 32'hbd76c852} /* (19, 20, 13) {real, imag} */,
  {32'h3daa04f0, 32'h3cf1d622} /* (19, 20, 12) {real, imag} */,
  {32'hbd1466e4, 32'hbc73b9d0} /* (19, 20, 11) {real, imag} */,
  {32'hbd53653a, 32'h3cad0c76} /* (19, 20, 10) {real, imag} */,
  {32'hbd5f4bc4, 32'h3dd421bf} /* (19, 20, 9) {real, imag} */,
  {32'hbdca3a9d, 32'h3d65e677} /* (19, 20, 8) {real, imag} */,
  {32'h3e02774e, 32'hbd43db6a} /* (19, 20, 7) {real, imag} */,
  {32'h3cf76758, 32'hbd481cf9} /* (19, 20, 6) {real, imag} */,
  {32'hbe16bef8, 32'hbe0b13d5} /* (19, 20, 5) {real, imag} */,
  {32'h3e251ba0, 32'h3c892731} /* (19, 20, 4) {real, imag} */,
  {32'hbde93d46, 32'hbd1f8c6c} /* (19, 20, 3) {real, imag} */,
  {32'hbec1062e, 32'hbe3cd662} /* (19, 20, 2) {real, imag} */,
  {32'h3f8f4b07, 32'h3e729aa0} /* (19, 20, 1) {real, imag} */,
  {32'h3e9412c0, 32'h00000000} /* (19, 20, 0) {real, imag} */,
  {32'h401cfe57, 32'hbec45b00} /* (19, 19, 31) {real, imag} */,
  {32'hbf69ca0c, 32'h3de798ba} /* (19, 19, 30) {real, imag} */,
  {32'hbcd4d7e6, 32'h3e1eeb1c} /* (19, 19, 29) {real, imag} */,
  {32'h3e7be862, 32'hbd604d63} /* (19, 19, 28) {real, imag} */,
  {32'hbe332efa, 32'h3e4bbe60} /* (19, 19, 27) {real, imag} */,
  {32'hbccf52ea, 32'h3df62a7a} /* (19, 19, 26) {real, imag} */,
  {32'h3e02f8ce, 32'hbd6c96f2} /* (19, 19, 25) {real, imag} */,
  {32'h3d60c6a8, 32'h3dabf56c} /* (19, 19, 24) {real, imag} */,
  {32'h3d9da774, 32'hbdc90d06} /* (19, 19, 23) {real, imag} */,
  {32'hbde2a386, 32'h3d33a7f8} /* (19, 19, 22) {real, imag} */,
  {32'hbd52d75a, 32'h3d51c362} /* (19, 19, 21) {real, imag} */,
  {32'h3d09d42e, 32'h3d43e53a} /* (19, 19, 20) {real, imag} */,
  {32'hbd2bf3cc, 32'hbd2138ee} /* (19, 19, 19) {real, imag} */,
  {32'h3b995698, 32'hbc5acac0} /* (19, 19, 18) {real, imag} */,
  {32'h3d649272, 32'h3d417873} /* (19, 19, 17) {real, imag} */,
  {32'h3d696b78, 32'h00000000} /* (19, 19, 16) {real, imag} */,
  {32'h3d649272, 32'hbd417873} /* (19, 19, 15) {real, imag} */,
  {32'h3b995698, 32'h3c5acac0} /* (19, 19, 14) {real, imag} */,
  {32'hbd2bf3cc, 32'h3d2138ee} /* (19, 19, 13) {real, imag} */,
  {32'h3d09d42e, 32'hbd43e53a} /* (19, 19, 12) {real, imag} */,
  {32'hbd52d75a, 32'hbd51c362} /* (19, 19, 11) {real, imag} */,
  {32'hbde2a386, 32'hbd33a7f8} /* (19, 19, 10) {real, imag} */,
  {32'h3d9da774, 32'h3dc90d06} /* (19, 19, 9) {real, imag} */,
  {32'h3d60c6a8, 32'hbdabf56c} /* (19, 19, 8) {real, imag} */,
  {32'h3e02f8ce, 32'h3d6c96f2} /* (19, 19, 7) {real, imag} */,
  {32'hbccf52ea, 32'hbdf62a7a} /* (19, 19, 6) {real, imag} */,
  {32'hbe332efa, 32'hbe4bbe60} /* (19, 19, 5) {real, imag} */,
  {32'h3e7be862, 32'h3d604d63} /* (19, 19, 4) {real, imag} */,
  {32'hbcd4d7e6, 32'hbe1eeb1c} /* (19, 19, 3) {real, imag} */,
  {32'hbf69ca0c, 32'hbde798ba} /* (19, 19, 2) {real, imag} */,
  {32'h401cfe57, 32'h3ec45b00} /* (19, 19, 1) {real, imag} */,
  {32'h3fb1175e, 32'h00000000} /* (19, 19, 0) {real, imag} */,
  {32'h40504838, 32'hbe9bba90} /* (19, 18, 31) {real, imag} */,
  {32'hbfa3ee5e, 32'h3e676b5b} /* (19, 18, 30) {real, imag} */,
  {32'h3dfd5c78, 32'h3e09bfd9} /* (19, 18, 29) {real, imag} */,
  {32'h3e9c2e78, 32'hbd04da62} /* (19, 18, 28) {real, imag} */,
  {32'hbd58d3ba, 32'h3bf8c9f8} /* (19, 18, 27) {real, imag} */,
  {32'hbdaeec81, 32'hbe2af88a} /* (19, 18, 26) {real, imag} */,
  {32'h3d65ff0a, 32'h3cb25188} /* (19, 18, 25) {real, imag} */,
  {32'h3ccefc13, 32'h3e11146f} /* (19, 18, 24) {real, imag} */,
  {32'h3de19d38, 32'hbd953670} /* (19, 18, 23) {real, imag} */,
  {32'h3d0d2e89, 32'h3a10a480} /* (19, 18, 22) {real, imag} */,
  {32'hbde05188, 32'h3e1db0b0} /* (19, 18, 21) {real, imag} */,
  {32'hbcad47a8, 32'h3cec1540} /* (19, 18, 20) {real, imag} */,
  {32'h3d207679, 32'hbd04a3eb} /* (19, 18, 19) {real, imag} */,
  {32'h3da03adc, 32'h3d3040bb} /* (19, 18, 18) {real, imag} */,
  {32'h3d83c3b0, 32'h3c8dc00a} /* (19, 18, 17) {real, imag} */,
  {32'h3b8ca258, 32'h00000000} /* (19, 18, 16) {real, imag} */,
  {32'h3d83c3b0, 32'hbc8dc00a} /* (19, 18, 15) {real, imag} */,
  {32'h3da03adc, 32'hbd3040bb} /* (19, 18, 14) {real, imag} */,
  {32'h3d207679, 32'h3d04a3eb} /* (19, 18, 13) {real, imag} */,
  {32'hbcad47a8, 32'hbcec1540} /* (19, 18, 12) {real, imag} */,
  {32'hbde05188, 32'hbe1db0b0} /* (19, 18, 11) {real, imag} */,
  {32'h3d0d2e89, 32'hba10a480} /* (19, 18, 10) {real, imag} */,
  {32'h3de19d38, 32'h3d953670} /* (19, 18, 9) {real, imag} */,
  {32'h3ccefc13, 32'hbe11146f} /* (19, 18, 8) {real, imag} */,
  {32'h3d65ff0a, 32'hbcb25188} /* (19, 18, 7) {real, imag} */,
  {32'hbdaeec81, 32'h3e2af88a} /* (19, 18, 6) {real, imag} */,
  {32'hbd58d3ba, 32'hbbf8c9f8} /* (19, 18, 5) {real, imag} */,
  {32'h3e9c2e78, 32'h3d04da62} /* (19, 18, 4) {real, imag} */,
  {32'h3dfd5c78, 32'hbe09bfd9} /* (19, 18, 3) {real, imag} */,
  {32'hbfa3ee5e, 32'hbe676b5b} /* (19, 18, 2) {real, imag} */,
  {32'h40504838, 32'h3e9bba90} /* (19, 18, 1) {real, imag} */,
  {32'h4004e4a3, 32'h00000000} /* (19, 18, 0) {real, imag} */,
  {32'h406ca2ae, 32'hbeaffe3f} /* (19, 17, 31) {real, imag} */,
  {32'hbfb7e339, 32'h3e7bf1ba} /* (19, 17, 30) {real, imag} */,
  {32'h3cdf7bba, 32'h3d420f6a} /* (19, 17, 29) {real, imag} */,
  {32'h3e149889, 32'hbdba39ee} /* (19, 17, 28) {real, imag} */,
  {32'hbdb2203b, 32'h3e0f1aa4} /* (19, 17, 27) {real, imag} */,
  {32'hbd658b92, 32'hbb2b7a50} /* (19, 17, 26) {real, imag} */,
  {32'h3df57412, 32'hbd38691c} /* (19, 17, 25) {real, imag} */,
  {32'hbdc57b7d, 32'h3da282a8} /* (19, 17, 24) {real, imag} */,
  {32'h3d7c48ea, 32'h3caeb7c3} /* (19, 17, 23) {real, imag} */,
  {32'h39ad6ec0, 32'h3ddb3b6a} /* (19, 17, 22) {real, imag} */,
  {32'hbd050d64, 32'hbc1a7995} /* (19, 17, 21) {real, imag} */,
  {32'h3c8a6c8e, 32'hbcc327aa} /* (19, 17, 20) {real, imag} */,
  {32'h3dfb4665, 32'hbc58f5b2} /* (19, 17, 19) {real, imag} */,
  {32'hbd5ab622, 32'hbdba4cf1} /* (19, 17, 18) {real, imag} */,
  {32'h3d18e6db, 32'hbdc5c51a} /* (19, 17, 17) {real, imag} */,
  {32'h3db45098, 32'h00000000} /* (19, 17, 16) {real, imag} */,
  {32'h3d18e6db, 32'h3dc5c51a} /* (19, 17, 15) {real, imag} */,
  {32'hbd5ab622, 32'h3dba4cf1} /* (19, 17, 14) {real, imag} */,
  {32'h3dfb4665, 32'h3c58f5b2} /* (19, 17, 13) {real, imag} */,
  {32'h3c8a6c8e, 32'h3cc327aa} /* (19, 17, 12) {real, imag} */,
  {32'hbd050d64, 32'h3c1a7995} /* (19, 17, 11) {real, imag} */,
  {32'h39ad6ec0, 32'hbddb3b6a} /* (19, 17, 10) {real, imag} */,
  {32'h3d7c48ea, 32'hbcaeb7c3} /* (19, 17, 9) {real, imag} */,
  {32'hbdc57b7d, 32'hbda282a8} /* (19, 17, 8) {real, imag} */,
  {32'h3df57412, 32'h3d38691c} /* (19, 17, 7) {real, imag} */,
  {32'hbd658b92, 32'h3b2b7a50} /* (19, 17, 6) {real, imag} */,
  {32'hbdb2203b, 32'hbe0f1aa4} /* (19, 17, 5) {real, imag} */,
  {32'h3e149889, 32'h3dba39ee} /* (19, 17, 4) {real, imag} */,
  {32'h3cdf7bba, 32'hbd420f6a} /* (19, 17, 3) {real, imag} */,
  {32'hbfb7e339, 32'hbe7bf1ba} /* (19, 17, 2) {real, imag} */,
  {32'h406ca2ae, 32'h3eaffe3f} /* (19, 17, 1) {real, imag} */,
  {32'h40276c76, 32'h00000000} /* (19, 17, 0) {real, imag} */,
  {32'h407c2b48, 32'hbec1394c} /* (19, 16, 31) {real, imag} */,
  {32'hbfd00f64, 32'h3e04b824} /* (19, 16, 30) {real, imag} */,
  {32'hbdc29584, 32'hbcb466b5} /* (19, 16, 29) {real, imag} */,
  {32'h3e8875dc, 32'hbd1ac301} /* (19, 16, 28) {real, imag} */,
  {32'hbe458731, 32'h3e14bd42} /* (19, 16, 27) {real, imag} */,
  {32'hbd924f74, 32'h3c92180f} /* (19, 16, 26) {real, imag} */,
  {32'h3d22465f, 32'hbd859075} /* (19, 16, 25) {real, imag} */,
  {32'hbd27b5d9, 32'h3cf75a2b} /* (19, 16, 24) {real, imag} */,
  {32'hbc37cc54, 32'hbdc01b18} /* (19, 16, 23) {real, imag} */,
  {32'h3a99885c, 32'hbdd93e24} /* (19, 16, 22) {real, imag} */,
  {32'hbd982e39, 32'h3dcf2077} /* (19, 16, 21) {real, imag} */,
  {32'hbd25deb6, 32'h3ce91206} /* (19, 16, 20) {real, imag} */,
  {32'hbd278c9d, 32'hbdd05555} /* (19, 16, 19) {real, imag} */,
  {32'h3b821344, 32'h3d59e2c2} /* (19, 16, 18) {real, imag} */,
  {32'hbd7cd8e6, 32'hbd33e872} /* (19, 16, 17) {real, imag} */,
  {32'hbcefffbc, 32'h00000000} /* (19, 16, 16) {real, imag} */,
  {32'hbd7cd8e6, 32'h3d33e872} /* (19, 16, 15) {real, imag} */,
  {32'h3b821344, 32'hbd59e2c2} /* (19, 16, 14) {real, imag} */,
  {32'hbd278c9d, 32'h3dd05555} /* (19, 16, 13) {real, imag} */,
  {32'hbd25deb6, 32'hbce91206} /* (19, 16, 12) {real, imag} */,
  {32'hbd982e39, 32'hbdcf2077} /* (19, 16, 11) {real, imag} */,
  {32'h3a99885c, 32'h3dd93e24} /* (19, 16, 10) {real, imag} */,
  {32'hbc37cc54, 32'h3dc01b18} /* (19, 16, 9) {real, imag} */,
  {32'hbd27b5d9, 32'hbcf75a2b} /* (19, 16, 8) {real, imag} */,
  {32'h3d22465f, 32'h3d859075} /* (19, 16, 7) {real, imag} */,
  {32'hbd924f74, 32'hbc92180f} /* (19, 16, 6) {real, imag} */,
  {32'hbe458731, 32'hbe14bd42} /* (19, 16, 5) {real, imag} */,
  {32'h3e8875dc, 32'h3d1ac301} /* (19, 16, 4) {real, imag} */,
  {32'hbdc29584, 32'h3cb466b5} /* (19, 16, 3) {real, imag} */,
  {32'hbfd00f64, 32'hbe04b824} /* (19, 16, 2) {real, imag} */,
  {32'h407c2b48, 32'h3ec1394c} /* (19, 16, 1) {real, imag} */,
  {32'h402e858c, 32'h00000000} /* (19, 16, 0) {real, imag} */,
  {32'h407b1aee, 32'hbeb54321} /* (19, 15, 31) {real, imag} */,
  {32'hbfe08491, 32'h3e5f4d46} /* (19, 15, 30) {real, imag} */,
  {32'hbd230f1f, 32'hbd486828} /* (19, 15, 29) {real, imag} */,
  {32'h3eb3a454, 32'hbdcf0cd2} /* (19, 15, 28) {real, imag} */,
  {32'hbe55ca22, 32'h3e0c1d30} /* (19, 15, 27) {real, imag} */,
  {32'hbc9b31a4, 32'h3c35210c} /* (19, 15, 26) {real, imag} */,
  {32'hbcde1a66, 32'hbdf2d27a} /* (19, 15, 25) {real, imag} */,
  {32'h3c6b46c8, 32'h3dad4c4a} /* (19, 15, 24) {real, imag} */,
  {32'hbd97631d, 32'hbd02ec9e} /* (19, 15, 23) {real, imag} */,
  {32'h3ab0f370, 32'h3d05e8cb} /* (19, 15, 22) {real, imag} */,
  {32'hbca6c347, 32'h3d24fbc7} /* (19, 15, 21) {real, imag} */,
  {32'hbda1cc52, 32'hbd91febc} /* (19, 15, 20) {real, imag} */,
  {32'h3c227b38, 32'h3ca65ae7} /* (19, 15, 19) {real, imag} */,
  {32'hbc21f1c6, 32'h3dfb285b} /* (19, 15, 18) {real, imag} */,
  {32'hbd2db9b7, 32'h3b65b2c0} /* (19, 15, 17) {real, imag} */,
  {32'h3dbfd88a, 32'h00000000} /* (19, 15, 16) {real, imag} */,
  {32'hbd2db9b7, 32'hbb65b2c0} /* (19, 15, 15) {real, imag} */,
  {32'hbc21f1c6, 32'hbdfb285b} /* (19, 15, 14) {real, imag} */,
  {32'h3c227b38, 32'hbca65ae7} /* (19, 15, 13) {real, imag} */,
  {32'hbda1cc52, 32'h3d91febc} /* (19, 15, 12) {real, imag} */,
  {32'hbca6c347, 32'hbd24fbc7} /* (19, 15, 11) {real, imag} */,
  {32'h3ab0f370, 32'hbd05e8cb} /* (19, 15, 10) {real, imag} */,
  {32'hbd97631d, 32'h3d02ec9e} /* (19, 15, 9) {real, imag} */,
  {32'h3c6b46c8, 32'hbdad4c4a} /* (19, 15, 8) {real, imag} */,
  {32'hbcde1a66, 32'h3df2d27a} /* (19, 15, 7) {real, imag} */,
  {32'hbc9b31a4, 32'hbc35210c} /* (19, 15, 6) {real, imag} */,
  {32'hbe55ca22, 32'hbe0c1d30} /* (19, 15, 5) {real, imag} */,
  {32'h3eb3a454, 32'h3dcf0cd2} /* (19, 15, 4) {real, imag} */,
  {32'hbd230f1f, 32'h3d486828} /* (19, 15, 3) {real, imag} */,
  {32'hbfe08491, 32'hbe5f4d46} /* (19, 15, 2) {real, imag} */,
  {32'h407b1aee, 32'h3eb54321} /* (19, 15, 1) {real, imag} */,
  {32'h403c209e, 32'h00000000} /* (19, 15, 0) {real, imag} */,
  {32'h4065f46a, 32'hbe9335f0} /* (19, 14, 31) {real, imag} */,
  {32'hbfcf520a, 32'h3e79245d} /* (19, 14, 30) {real, imag} */,
  {32'h3d2ab667, 32'hbcb98980} /* (19, 14, 29) {real, imag} */,
  {32'h3e2815f9, 32'hbd95e927} /* (19, 14, 28) {real, imag} */,
  {32'hbe5fb7e6, 32'h3daa9b6c} /* (19, 14, 27) {real, imag} */,
  {32'hbda13975, 32'h3e0ad832} /* (19, 14, 26) {real, imag} */,
  {32'h3d1e9cea, 32'hbdc5e585} /* (19, 14, 25) {real, imag} */,
  {32'hbc3e259e, 32'h3dc06c7f} /* (19, 14, 24) {real, imag} */,
  {32'h3d899b94, 32'hbd317fba} /* (19, 14, 23) {real, imag} */,
  {32'hbd27b1d5, 32'hbd9e6667} /* (19, 14, 22) {real, imag} */,
  {32'hbcd34832, 32'h3d4b4558} /* (19, 14, 21) {real, imag} */,
  {32'hba2622c0, 32'h3c3dfd60} /* (19, 14, 20) {real, imag} */,
  {32'hbd04777f, 32'h3cc7ac78} /* (19, 14, 19) {real, imag} */,
  {32'hbd64c0f8, 32'hbb5daf20} /* (19, 14, 18) {real, imag} */,
  {32'h3c929348, 32'h3d21346d} /* (19, 14, 17) {real, imag} */,
  {32'h3d5c0185, 32'h00000000} /* (19, 14, 16) {real, imag} */,
  {32'h3c929348, 32'hbd21346d} /* (19, 14, 15) {real, imag} */,
  {32'hbd64c0f8, 32'h3b5daf20} /* (19, 14, 14) {real, imag} */,
  {32'hbd04777f, 32'hbcc7ac78} /* (19, 14, 13) {real, imag} */,
  {32'hba2622c0, 32'hbc3dfd60} /* (19, 14, 12) {real, imag} */,
  {32'hbcd34832, 32'hbd4b4558} /* (19, 14, 11) {real, imag} */,
  {32'hbd27b1d5, 32'h3d9e6667} /* (19, 14, 10) {real, imag} */,
  {32'h3d899b94, 32'h3d317fba} /* (19, 14, 9) {real, imag} */,
  {32'hbc3e259e, 32'hbdc06c7f} /* (19, 14, 8) {real, imag} */,
  {32'h3d1e9cea, 32'h3dc5e585} /* (19, 14, 7) {real, imag} */,
  {32'hbda13975, 32'hbe0ad832} /* (19, 14, 6) {real, imag} */,
  {32'hbe5fb7e6, 32'hbdaa9b6c} /* (19, 14, 5) {real, imag} */,
  {32'h3e2815f9, 32'h3d95e927} /* (19, 14, 4) {real, imag} */,
  {32'h3d2ab667, 32'h3cb98980} /* (19, 14, 3) {real, imag} */,
  {32'hbfcf520a, 32'hbe79245d} /* (19, 14, 2) {real, imag} */,
  {32'h4065f46a, 32'h3e9335f0} /* (19, 14, 1) {real, imag} */,
  {32'h402490b1, 32'h00000000} /* (19, 14, 0) {real, imag} */,
  {32'h4041aae5, 32'hbdfdf460} /* (19, 13, 31) {real, imag} */,
  {32'hbfb21a66, 32'h3e45fc9f} /* (19, 13, 30) {real, imag} */,
  {32'h3d82ccb0, 32'hbe77321c} /* (19, 13, 29) {real, imag} */,
  {32'h3e235e2e, 32'hbcd5f32a} /* (19, 13, 28) {real, imag} */,
  {32'hbe6ca15e, 32'h3cba5020} /* (19, 13, 27) {real, imag} */,
  {32'h3d536827, 32'h3da9e68e} /* (19, 13, 26) {real, imag} */,
  {32'hbd3fe7d2, 32'hbcec28d4} /* (19, 13, 25) {real, imag} */,
  {32'hbce68118, 32'h3d0bb74c} /* (19, 13, 24) {real, imag} */,
  {32'h3d9796f0, 32'h3cbaa050} /* (19, 13, 23) {real, imag} */,
  {32'hbdae5e3e, 32'hbe02e785} /* (19, 13, 22) {real, imag} */,
  {32'hbd1fa3cc, 32'h3da55cdb} /* (19, 13, 21) {real, imag} */,
  {32'h3d1fac28, 32'hbcd3286d} /* (19, 13, 20) {real, imag} */,
  {32'hbcd5135c, 32'h3c8e52d1} /* (19, 13, 19) {real, imag} */,
  {32'h3dc4c888, 32'h3e13cb53} /* (19, 13, 18) {real, imag} */,
  {32'h3ce6bd04, 32'hbd2a30c3} /* (19, 13, 17) {real, imag} */,
  {32'h3d856cec, 32'h00000000} /* (19, 13, 16) {real, imag} */,
  {32'h3ce6bd04, 32'h3d2a30c3} /* (19, 13, 15) {real, imag} */,
  {32'h3dc4c888, 32'hbe13cb53} /* (19, 13, 14) {real, imag} */,
  {32'hbcd5135c, 32'hbc8e52d1} /* (19, 13, 13) {real, imag} */,
  {32'h3d1fac28, 32'h3cd3286d} /* (19, 13, 12) {real, imag} */,
  {32'hbd1fa3cc, 32'hbda55cdb} /* (19, 13, 11) {real, imag} */,
  {32'hbdae5e3e, 32'h3e02e785} /* (19, 13, 10) {real, imag} */,
  {32'h3d9796f0, 32'hbcbaa050} /* (19, 13, 9) {real, imag} */,
  {32'hbce68118, 32'hbd0bb74c} /* (19, 13, 8) {real, imag} */,
  {32'hbd3fe7d2, 32'h3cec28d4} /* (19, 13, 7) {real, imag} */,
  {32'h3d536827, 32'hbda9e68e} /* (19, 13, 6) {real, imag} */,
  {32'hbe6ca15e, 32'hbcba5020} /* (19, 13, 5) {real, imag} */,
  {32'h3e235e2e, 32'h3cd5f32a} /* (19, 13, 4) {real, imag} */,
  {32'h3d82ccb0, 32'h3e77321c} /* (19, 13, 3) {real, imag} */,
  {32'hbfb21a66, 32'hbe45fc9f} /* (19, 13, 2) {real, imag} */,
  {32'h4041aae5, 32'h3dfdf460} /* (19, 13, 1) {real, imag} */,
  {32'h4003b053, 32'h00000000} /* (19, 13, 0) {real, imag} */,
  {32'h40082968, 32'h3d70a980} /* (19, 12, 31) {real, imag} */,
  {32'hbf9bb6e6, 32'h3e87dfa8} /* (19, 12, 30) {real, imag} */,
  {32'h3e158b45, 32'hbe4019d1} /* (19, 12, 29) {real, imag} */,
  {32'h3dc32859, 32'hbcbd6071} /* (19, 12, 28) {real, imag} */,
  {32'hbe625364, 32'h3e24f16f} /* (19, 12, 27) {real, imag} */,
  {32'h3dbeafca, 32'h3d1b378f} /* (19, 12, 26) {real, imag} */,
  {32'hbd3f2fca, 32'hbce2357c} /* (19, 12, 25) {real, imag} */,
  {32'hbdef7953, 32'hbcc53582} /* (19, 12, 24) {real, imag} */,
  {32'h3c9b9f58, 32'h3df05f21} /* (19, 12, 23) {real, imag} */,
  {32'hba037e00, 32'hbd44e217} /* (19, 12, 22) {real, imag} */,
  {32'h3cf64c3f, 32'h3d0cafb8} /* (19, 12, 21) {real, imag} */,
  {32'h3d3ead11, 32'hbd7e420d} /* (19, 12, 20) {real, imag} */,
  {32'hbd733ea0, 32'h3db77431} /* (19, 12, 19) {real, imag} */,
  {32'h3d728f94, 32'h3cd02c38} /* (19, 12, 18) {real, imag} */,
  {32'hbd238cb9, 32'hbc5f9f80} /* (19, 12, 17) {real, imag} */,
  {32'hbcb7d42a, 32'h00000000} /* (19, 12, 16) {real, imag} */,
  {32'hbd238cb9, 32'h3c5f9f80} /* (19, 12, 15) {real, imag} */,
  {32'h3d728f94, 32'hbcd02c38} /* (19, 12, 14) {real, imag} */,
  {32'hbd733ea0, 32'hbdb77431} /* (19, 12, 13) {real, imag} */,
  {32'h3d3ead11, 32'h3d7e420d} /* (19, 12, 12) {real, imag} */,
  {32'h3cf64c3f, 32'hbd0cafb8} /* (19, 12, 11) {real, imag} */,
  {32'hba037e00, 32'h3d44e217} /* (19, 12, 10) {real, imag} */,
  {32'h3c9b9f58, 32'hbdf05f21} /* (19, 12, 9) {real, imag} */,
  {32'hbdef7953, 32'h3cc53582} /* (19, 12, 8) {real, imag} */,
  {32'hbd3f2fca, 32'h3ce2357c} /* (19, 12, 7) {real, imag} */,
  {32'h3dbeafca, 32'hbd1b378f} /* (19, 12, 6) {real, imag} */,
  {32'hbe625364, 32'hbe24f16f} /* (19, 12, 5) {real, imag} */,
  {32'h3dc32859, 32'h3cbd6071} /* (19, 12, 4) {real, imag} */,
  {32'h3e158b45, 32'h3e4019d1} /* (19, 12, 3) {real, imag} */,
  {32'hbf9bb6e6, 32'hbe87dfa8} /* (19, 12, 2) {real, imag} */,
  {32'h40082968, 32'hbd70a980} /* (19, 12, 1) {real, imag} */,
  {32'h3fb3c06e, 32'h00000000} /* (19, 12, 0) {real, imag} */,
  {32'h3f736eb0, 32'h3eabbdf8} /* (19, 11, 31) {real, imag} */,
  {32'hbf1b3e2d, 32'h3dc59906} /* (19, 11, 30) {real, imag} */,
  {32'h3e0608c8, 32'hbdb52d08} /* (19, 11, 29) {real, imag} */,
  {32'h3dc2e0a3, 32'hbbf425a0} /* (19, 11, 28) {real, imag} */,
  {32'hbe722a6e, 32'h3ca44704} /* (19, 11, 27) {real, imag} */,
  {32'h3df1e0d9, 32'h3c8d5ac8} /* (19, 11, 26) {real, imag} */,
  {32'hbdec53ae, 32'h3d26eb76} /* (19, 11, 25) {real, imag} */,
  {32'hbd96422f, 32'hbcd29903} /* (19, 11, 24) {real, imag} */,
  {32'h3d39dee0, 32'h3d07dcfa} /* (19, 11, 23) {real, imag} */,
  {32'hbc05b91c, 32'hbda68399} /* (19, 11, 22) {real, imag} */,
  {32'hbd719c58, 32'h3c6573ba} /* (19, 11, 21) {real, imag} */,
  {32'h3d904d70, 32'h3b4bb7c8} /* (19, 11, 20) {real, imag} */,
  {32'hbb5baef4, 32'h3da7b567} /* (19, 11, 19) {real, imag} */,
  {32'h3cdfc734, 32'hbcae8a78} /* (19, 11, 18) {real, imag} */,
  {32'h3b9ed9fc, 32'h3d5185aa} /* (19, 11, 17) {real, imag} */,
  {32'h3dd4dbc8, 32'h00000000} /* (19, 11, 16) {real, imag} */,
  {32'h3b9ed9fc, 32'hbd5185aa} /* (19, 11, 15) {real, imag} */,
  {32'h3cdfc734, 32'h3cae8a78} /* (19, 11, 14) {real, imag} */,
  {32'hbb5baef4, 32'hbda7b567} /* (19, 11, 13) {real, imag} */,
  {32'h3d904d70, 32'hbb4bb7c8} /* (19, 11, 12) {real, imag} */,
  {32'hbd719c58, 32'hbc6573ba} /* (19, 11, 11) {real, imag} */,
  {32'hbc05b91c, 32'h3da68399} /* (19, 11, 10) {real, imag} */,
  {32'h3d39dee0, 32'hbd07dcfa} /* (19, 11, 9) {real, imag} */,
  {32'hbd96422f, 32'h3cd29903} /* (19, 11, 8) {real, imag} */,
  {32'hbdec53ae, 32'hbd26eb76} /* (19, 11, 7) {real, imag} */,
  {32'h3df1e0d9, 32'hbc8d5ac8} /* (19, 11, 6) {real, imag} */,
  {32'hbe722a6e, 32'hbca44704} /* (19, 11, 5) {real, imag} */,
  {32'h3dc2e0a3, 32'h3bf425a0} /* (19, 11, 4) {real, imag} */,
  {32'h3e0608c8, 32'h3db52d08} /* (19, 11, 3) {real, imag} */,
  {32'hbf1b3e2d, 32'hbdc59906} /* (19, 11, 2) {real, imag} */,
  {32'h3f736eb0, 32'hbeabbdf8} /* (19, 11, 1) {real, imag} */,
  {32'h3f088258, 32'h00000000} /* (19, 11, 0) {real, imag} */,
  {32'hbf5cbab1, 32'h3f490ab8} /* (19, 10, 31) {real, imag} */,
  {32'h3eb8218a, 32'hbdaf0352} /* (19, 10, 30) {real, imag} */,
  {32'hba5bcd00, 32'hbd9e78b2} /* (19, 10, 29) {real, imag} */,
  {32'hbd7cccbe, 32'h3b628e30} /* (19, 10, 28) {real, imag} */,
  {32'hbb819bc0, 32'h3ca74d30} /* (19, 10, 27) {real, imag} */,
  {32'h3d9bcd3a, 32'hbd5bd378} /* (19, 10, 26) {real, imag} */,
  {32'hbe056f96, 32'h3dd27b2c} /* (19, 10, 25) {real, imag} */,
  {32'hbc369ffc, 32'hbdc31244} /* (19, 10, 24) {real, imag} */,
  {32'h3d4c59ac, 32'h3e0ef52b} /* (19, 10, 23) {real, imag} */,
  {32'h3d873efc, 32'hbc7a2752} /* (19, 10, 22) {real, imag} */,
  {32'hbcac60b4, 32'h3d606766} /* (19, 10, 21) {real, imag} */,
  {32'hbd1bffe4, 32'hbc25dcac} /* (19, 10, 20) {real, imag} */,
  {32'h3ce0d77e, 32'hbc8a373b} /* (19, 10, 19) {real, imag} */,
  {32'h3cbbd08c, 32'h3d06c71a} /* (19, 10, 18) {real, imag} */,
  {32'hbce5141f, 32'hbd9bf14e} /* (19, 10, 17) {real, imag} */,
  {32'h3d21c48c, 32'h00000000} /* (19, 10, 16) {real, imag} */,
  {32'hbce5141f, 32'h3d9bf14e} /* (19, 10, 15) {real, imag} */,
  {32'h3cbbd08c, 32'hbd06c71a} /* (19, 10, 14) {real, imag} */,
  {32'h3ce0d77e, 32'h3c8a373b} /* (19, 10, 13) {real, imag} */,
  {32'hbd1bffe4, 32'h3c25dcac} /* (19, 10, 12) {real, imag} */,
  {32'hbcac60b4, 32'hbd606766} /* (19, 10, 11) {real, imag} */,
  {32'h3d873efc, 32'h3c7a2752} /* (19, 10, 10) {real, imag} */,
  {32'h3d4c59ac, 32'hbe0ef52b} /* (19, 10, 9) {real, imag} */,
  {32'hbc369ffc, 32'h3dc31244} /* (19, 10, 8) {real, imag} */,
  {32'hbe056f96, 32'hbdd27b2c} /* (19, 10, 7) {real, imag} */,
  {32'h3d9bcd3a, 32'h3d5bd378} /* (19, 10, 6) {real, imag} */,
  {32'hbb819bc0, 32'hbca74d30} /* (19, 10, 5) {real, imag} */,
  {32'hbd7cccbe, 32'hbb628e30} /* (19, 10, 4) {real, imag} */,
  {32'hba5bcd00, 32'h3d9e78b2} /* (19, 10, 3) {real, imag} */,
  {32'h3eb8218a, 32'h3daf0352} /* (19, 10, 2) {real, imag} */,
  {32'hbf5cbab1, 32'hbf490ab8} /* (19, 10, 1) {real, imag} */,
  {32'hbf62157c, 32'h00000000} /* (19, 10, 0) {real, imag} */,
  {32'hc01164b1, 32'h3f840e23} /* (19, 9, 31) {real, imag} */,
  {32'h3f6db53c, 32'hbe56dd12} /* (19, 9, 30) {real, imag} */,
  {32'hbe0b43ca, 32'h3cc786b8} /* (19, 9, 29) {real, imag} */,
  {32'h3ce99f74, 32'hbcd0d088} /* (19, 9, 28) {real, imag} */,
  {32'h3dc3ca6a, 32'h3c89f190} /* (19, 9, 27) {real, imag} */,
  {32'h3cc50728, 32'hbd49743a} /* (19, 9, 26) {real, imag} */,
  {32'hbe3a21e9, 32'h3d0727c0} /* (19, 9, 25) {real, imag} */,
  {32'h3d6a6f40, 32'hbe0f0faf} /* (19, 9, 24) {real, imag} */,
  {32'h3d8002ab, 32'h3da15320} /* (19, 9, 23) {real, imag} */,
  {32'hbe04238a, 32'h3ce7bfb0} /* (19, 9, 22) {real, imag} */,
  {32'h3dd42a09, 32'hbd631a3c} /* (19, 9, 21) {real, imag} */,
  {32'hbb02c2a4, 32'hbd18caea} /* (19, 9, 20) {real, imag} */,
  {32'h3e294946, 32'hbd4f2d3d} /* (19, 9, 19) {real, imag} */,
  {32'hbe010c1f, 32'hbd0717cb} /* (19, 9, 18) {real, imag} */,
  {32'hbd418624, 32'hbc1ecc42} /* (19, 9, 17) {real, imag} */,
  {32'hbd611c59, 32'h00000000} /* (19, 9, 16) {real, imag} */,
  {32'hbd418624, 32'h3c1ecc42} /* (19, 9, 15) {real, imag} */,
  {32'hbe010c1f, 32'h3d0717cb} /* (19, 9, 14) {real, imag} */,
  {32'h3e294946, 32'h3d4f2d3d} /* (19, 9, 13) {real, imag} */,
  {32'hbb02c2a4, 32'h3d18caea} /* (19, 9, 12) {real, imag} */,
  {32'h3dd42a09, 32'h3d631a3c} /* (19, 9, 11) {real, imag} */,
  {32'hbe04238a, 32'hbce7bfb0} /* (19, 9, 10) {real, imag} */,
  {32'h3d8002ab, 32'hbda15320} /* (19, 9, 9) {real, imag} */,
  {32'h3d6a6f40, 32'h3e0f0faf} /* (19, 9, 8) {real, imag} */,
  {32'hbe3a21e9, 32'hbd0727c0} /* (19, 9, 7) {real, imag} */,
  {32'h3cc50728, 32'h3d49743a} /* (19, 9, 6) {real, imag} */,
  {32'h3dc3ca6a, 32'hbc89f190} /* (19, 9, 5) {real, imag} */,
  {32'h3ce99f74, 32'h3cd0d088} /* (19, 9, 4) {real, imag} */,
  {32'hbe0b43ca, 32'hbcc786b8} /* (19, 9, 3) {real, imag} */,
  {32'h3f6db53c, 32'h3e56dd12} /* (19, 9, 2) {real, imag} */,
  {32'hc01164b1, 32'hbf840e23} /* (19, 9, 1) {real, imag} */,
  {32'hbff7d4a4, 32'h00000000} /* (19, 9, 0) {real, imag} */,
  {32'hc03ffaa7, 32'h3fad88fb} /* (19, 8, 31) {real, imag} */,
  {32'h3f76cc3e, 32'hbe912a5c} /* (19, 8, 30) {real, imag} */,
  {32'hbdb411c1, 32'hbb1b04d8} /* (19, 8, 29) {real, imag} */,
  {32'hbdf76aa6, 32'h3d25af66} /* (19, 8, 28) {real, imag} */,
  {32'h3e44ff42, 32'hbd307d97} /* (19, 8, 27) {real, imag} */,
  {32'hbd42e0e9, 32'hbd78e0ee} /* (19, 8, 26) {real, imag} */,
  {32'hbd1f416a, 32'h3c518978} /* (19, 8, 25) {real, imag} */,
  {32'h3dcfe75a, 32'hbd865aea} /* (19, 8, 24) {real, imag} */,
  {32'h3d9bb450, 32'h3d9ed10a} /* (19, 8, 23) {real, imag} */,
  {32'hbe2bb4ff, 32'hbcb3ad39} /* (19, 8, 22) {real, imag} */,
  {32'hbc508450, 32'hbe2fe75e} /* (19, 8, 21) {real, imag} */,
  {32'hbd32c308, 32'hbc1e033a} /* (19, 8, 20) {real, imag} */,
  {32'hbd068084, 32'h3ca38cee} /* (19, 8, 19) {real, imag} */,
  {32'h3c75fb76, 32'hbd833a9a} /* (19, 8, 18) {real, imag} */,
  {32'h3d79782b, 32'h3c83a83c} /* (19, 8, 17) {real, imag} */,
  {32'hbc37dc90, 32'h00000000} /* (19, 8, 16) {real, imag} */,
  {32'h3d79782b, 32'hbc83a83c} /* (19, 8, 15) {real, imag} */,
  {32'h3c75fb76, 32'h3d833a9a} /* (19, 8, 14) {real, imag} */,
  {32'hbd068084, 32'hbca38cee} /* (19, 8, 13) {real, imag} */,
  {32'hbd32c308, 32'h3c1e033a} /* (19, 8, 12) {real, imag} */,
  {32'hbc508450, 32'h3e2fe75e} /* (19, 8, 11) {real, imag} */,
  {32'hbe2bb4ff, 32'h3cb3ad39} /* (19, 8, 10) {real, imag} */,
  {32'h3d9bb450, 32'hbd9ed10a} /* (19, 8, 9) {real, imag} */,
  {32'h3dcfe75a, 32'h3d865aea} /* (19, 8, 8) {real, imag} */,
  {32'hbd1f416a, 32'hbc518978} /* (19, 8, 7) {real, imag} */,
  {32'hbd42e0e9, 32'h3d78e0ee} /* (19, 8, 6) {real, imag} */,
  {32'h3e44ff42, 32'h3d307d97} /* (19, 8, 5) {real, imag} */,
  {32'hbdf76aa6, 32'hbd25af66} /* (19, 8, 4) {real, imag} */,
  {32'hbdb411c1, 32'h3b1b04d8} /* (19, 8, 3) {real, imag} */,
  {32'h3f76cc3e, 32'h3e912a5c} /* (19, 8, 2) {real, imag} */,
  {32'hc03ffaa7, 32'hbfad88fb} /* (19, 8, 1) {real, imag} */,
  {32'hc033073c, 32'h00000000} /* (19, 8, 0) {real, imag} */,
  {32'hc059fd84, 32'h3fe874ee} /* (19, 7, 31) {real, imag} */,
  {32'h3f861c1c, 32'hbf06d418} /* (19, 7, 30) {real, imag} */,
  {32'hbe0a43d3, 32'hbb8c1de8} /* (19, 7, 29) {real, imag} */,
  {32'hbdca1cc0, 32'h3e1b6b27} /* (19, 7, 28) {real, imag} */,
  {32'h3e0929a3, 32'hbd5be488} /* (19, 7, 27) {real, imag} */,
  {32'hbc5fe1a4, 32'h3d2eea88} /* (19, 7, 26) {real, imag} */,
  {32'h3da84f6c, 32'h3d787926} /* (19, 7, 25) {real, imag} */,
  {32'hbc97bc12, 32'hbdf892d6} /* (19, 7, 24) {real, imag} */,
  {32'hbd04f7ce, 32'h3dca3106} /* (19, 7, 23) {real, imag} */,
  {32'h3d8537e4, 32'h3d92a014} /* (19, 7, 22) {real, imag} */,
  {32'h3dea81da, 32'hbe015eec} /* (19, 7, 21) {real, imag} */,
  {32'hbd6b0066, 32'h3dbe7140} /* (19, 7, 20) {real, imag} */,
  {32'hbbb8a970, 32'h3dca7637} /* (19, 7, 19) {real, imag} */,
  {32'h3c588c96, 32'h3c9e8e48} /* (19, 7, 18) {real, imag} */,
  {32'h3d0f3f9a, 32'h3d1a0a8c} /* (19, 7, 17) {real, imag} */,
  {32'hbd3385dc, 32'h00000000} /* (19, 7, 16) {real, imag} */,
  {32'h3d0f3f9a, 32'hbd1a0a8c} /* (19, 7, 15) {real, imag} */,
  {32'h3c588c96, 32'hbc9e8e48} /* (19, 7, 14) {real, imag} */,
  {32'hbbb8a970, 32'hbdca7637} /* (19, 7, 13) {real, imag} */,
  {32'hbd6b0066, 32'hbdbe7140} /* (19, 7, 12) {real, imag} */,
  {32'h3dea81da, 32'h3e015eec} /* (19, 7, 11) {real, imag} */,
  {32'h3d8537e4, 32'hbd92a014} /* (19, 7, 10) {real, imag} */,
  {32'hbd04f7ce, 32'hbdca3106} /* (19, 7, 9) {real, imag} */,
  {32'hbc97bc12, 32'h3df892d6} /* (19, 7, 8) {real, imag} */,
  {32'h3da84f6c, 32'hbd787926} /* (19, 7, 7) {real, imag} */,
  {32'hbc5fe1a4, 32'hbd2eea88} /* (19, 7, 6) {real, imag} */,
  {32'h3e0929a3, 32'h3d5be488} /* (19, 7, 5) {real, imag} */,
  {32'hbdca1cc0, 32'hbe1b6b27} /* (19, 7, 4) {real, imag} */,
  {32'hbe0a43d3, 32'h3b8c1de8} /* (19, 7, 3) {real, imag} */,
  {32'h3f861c1c, 32'h3f06d418} /* (19, 7, 2) {real, imag} */,
  {32'hc059fd84, 32'hbfe874ee} /* (19, 7, 1) {real, imag} */,
  {32'hc060e3ce, 32'h00000000} /* (19, 7, 0) {real, imag} */,
  {32'hc06123f8, 32'h4007f18b} /* (19, 6, 31) {real, imag} */,
  {32'h3f538b6f, 32'hbf38faac} /* (19, 6, 30) {real, imag} */,
  {32'hbd922014, 32'hbd819ca5} /* (19, 6, 29) {real, imag} */,
  {32'hbd281bc0, 32'hb8edc200} /* (19, 6, 28) {real, imag} */,
  {32'h3ddeb268, 32'hbc9e10b0} /* (19, 6, 27) {real, imag} */,
  {32'h3ac7c980, 32'h3c15bf18} /* (19, 6, 26) {real, imag} */,
  {32'h3e18d48a, 32'hbc94ddea} /* (19, 6, 25) {real, imag} */,
  {32'h3cacc0fc, 32'hbe2c5aa2} /* (19, 6, 24) {real, imag} */,
  {32'hbbfe3cfa, 32'hbd26520e} /* (19, 6, 23) {real, imag} */,
  {32'hbd5f4c48, 32'h3dcb4f03} /* (19, 6, 22) {real, imag} */,
  {32'h3c5eddb8, 32'hbce0a6c8} /* (19, 6, 21) {real, imag} */,
  {32'hbd7631e1, 32'h3c1ed667} /* (19, 6, 20) {real, imag} */,
  {32'h3d456a70, 32'hbd4ead7c} /* (19, 6, 19) {real, imag} */,
  {32'h3e0105b0, 32'hbd1793fa} /* (19, 6, 18) {real, imag} */,
  {32'hbd5eda06, 32'hbb9882ba} /* (19, 6, 17) {real, imag} */,
  {32'h3c1efe0f, 32'h00000000} /* (19, 6, 16) {real, imag} */,
  {32'hbd5eda06, 32'h3b9882ba} /* (19, 6, 15) {real, imag} */,
  {32'h3e0105b0, 32'h3d1793fa} /* (19, 6, 14) {real, imag} */,
  {32'h3d456a70, 32'h3d4ead7c} /* (19, 6, 13) {real, imag} */,
  {32'hbd7631e1, 32'hbc1ed667} /* (19, 6, 12) {real, imag} */,
  {32'h3c5eddb8, 32'h3ce0a6c8} /* (19, 6, 11) {real, imag} */,
  {32'hbd5f4c48, 32'hbdcb4f03} /* (19, 6, 10) {real, imag} */,
  {32'hbbfe3cfa, 32'h3d26520e} /* (19, 6, 9) {real, imag} */,
  {32'h3cacc0fc, 32'h3e2c5aa2} /* (19, 6, 8) {real, imag} */,
  {32'h3e18d48a, 32'h3c94ddea} /* (19, 6, 7) {real, imag} */,
  {32'h3ac7c980, 32'hbc15bf18} /* (19, 6, 6) {real, imag} */,
  {32'h3ddeb268, 32'h3c9e10b0} /* (19, 6, 5) {real, imag} */,
  {32'hbd281bc0, 32'h38edc200} /* (19, 6, 4) {real, imag} */,
  {32'hbd922014, 32'h3d819ca5} /* (19, 6, 3) {real, imag} */,
  {32'h3f538b6f, 32'h3f38faac} /* (19, 6, 2) {real, imag} */,
  {32'hc06123f8, 32'hc007f18b} /* (19, 6, 1) {real, imag} */,
  {32'hc07385e8, 32'h00000000} /* (19, 6, 0) {real, imag} */,
  {32'hc058e9f0, 32'h4032516d} /* (19, 5, 31) {real, imag} */,
  {32'h3ddab478, 32'hbf63ad54} /* (19, 5, 30) {real, imag} */,
  {32'h3d89faec, 32'hbe1eb606} /* (19, 5, 29) {real, imag} */,
  {32'h3b68ef80, 32'hbc82aa8c} /* (19, 5, 28) {real, imag} */,
  {32'h3e608bab, 32'h3dfb30b0} /* (19, 5, 27) {real, imag} */,
  {32'h3e4813fa, 32'hbda92f11} /* (19, 5, 26) {real, imag} */,
  {32'hbd79c292, 32'h3ccb7857} /* (19, 5, 25) {real, imag} */,
  {32'h3b3a35b0, 32'hbdb4059c} /* (19, 5, 24) {real, imag} */,
  {32'h3d4189b4, 32'hbcd6f408} /* (19, 5, 23) {real, imag} */,
  {32'h3e0f3ede, 32'hbcbe86ac} /* (19, 5, 22) {real, imag} */,
  {32'h3d8a48a6, 32'hbda67ec4} /* (19, 5, 21) {real, imag} */,
  {32'h3bedb98e, 32'h3d49d398} /* (19, 5, 20) {real, imag} */,
  {32'hbcdd82bc, 32'h3cb4f33a} /* (19, 5, 19) {real, imag} */,
  {32'hbc8870f3, 32'h3dbf1833} /* (19, 5, 18) {real, imag} */,
  {32'hbb5495e4, 32'hbdef6744} /* (19, 5, 17) {real, imag} */,
  {32'h3d57eca9, 32'h00000000} /* (19, 5, 16) {real, imag} */,
  {32'hbb5495e4, 32'h3def6744} /* (19, 5, 15) {real, imag} */,
  {32'hbc8870f3, 32'hbdbf1833} /* (19, 5, 14) {real, imag} */,
  {32'hbcdd82bc, 32'hbcb4f33a} /* (19, 5, 13) {real, imag} */,
  {32'h3bedb98e, 32'hbd49d398} /* (19, 5, 12) {real, imag} */,
  {32'h3d8a48a6, 32'h3da67ec4} /* (19, 5, 11) {real, imag} */,
  {32'h3e0f3ede, 32'h3cbe86ac} /* (19, 5, 10) {real, imag} */,
  {32'h3d4189b4, 32'h3cd6f408} /* (19, 5, 9) {real, imag} */,
  {32'h3b3a35b0, 32'h3db4059c} /* (19, 5, 8) {real, imag} */,
  {32'hbd79c292, 32'hbccb7857} /* (19, 5, 7) {real, imag} */,
  {32'h3e4813fa, 32'h3da92f11} /* (19, 5, 6) {real, imag} */,
  {32'h3e608bab, 32'hbdfb30b0} /* (19, 5, 5) {real, imag} */,
  {32'h3b68ef80, 32'h3c82aa8c} /* (19, 5, 4) {real, imag} */,
  {32'h3d89faec, 32'h3e1eb606} /* (19, 5, 3) {real, imag} */,
  {32'h3ddab478, 32'h3f63ad54} /* (19, 5, 2) {real, imag} */,
  {32'hc058e9f0, 32'hc032516d} /* (19, 5, 1) {real, imag} */,
  {32'hc0813d3e, 32'h00000000} /* (19, 5, 0) {real, imag} */,
  {32'hc043fc7c, 32'h405a2266} /* (19, 4, 31) {real, imag} */,
  {32'hbe9b0a8e, 32'hbf8dce0f} /* (19, 4, 30) {real, imag} */,
  {32'h3dc21060, 32'hbd33aeb8} /* (19, 4, 29) {real, imag} */,
  {32'h3e385d54, 32'hbda32689} /* (19, 4, 28) {real, imag} */,
  {32'h3e73b035, 32'h3e42363d} /* (19, 4, 27) {real, imag} */,
  {32'h3cc6d9b0, 32'hbcfc7962} /* (19, 4, 26) {real, imag} */,
  {32'h3b03c980, 32'h3d877eac} /* (19, 4, 25) {real, imag} */,
  {32'hbd6d48f6, 32'hbcec0cb6} /* (19, 4, 24) {real, imag} */,
  {32'h3d49ba20, 32'h3cc1b78e} /* (19, 4, 23) {real, imag} */,
  {32'h3d8334d1, 32'hbd573a0f} /* (19, 4, 22) {real, imag} */,
  {32'h3d944c40, 32'hbde0f475} /* (19, 4, 21) {real, imag} */,
  {32'h3a781420, 32'h3e122fd4} /* (19, 4, 20) {real, imag} */,
  {32'h3d12d1af, 32'h3c91e5e1} /* (19, 4, 19) {real, imag} */,
  {32'hbcdfe3c4, 32'hbcd3b144} /* (19, 4, 18) {real, imag} */,
  {32'h3d3cdb2a, 32'h3bd19194} /* (19, 4, 17) {real, imag} */,
  {32'h3dfedb80, 32'h00000000} /* (19, 4, 16) {real, imag} */,
  {32'h3d3cdb2a, 32'hbbd19194} /* (19, 4, 15) {real, imag} */,
  {32'hbcdfe3c4, 32'h3cd3b144} /* (19, 4, 14) {real, imag} */,
  {32'h3d12d1af, 32'hbc91e5e1} /* (19, 4, 13) {real, imag} */,
  {32'h3a781420, 32'hbe122fd4} /* (19, 4, 12) {real, imag} */,
  {32'h3d944c40, 32'h3de0f475} /* (19, 4, 11) {real, imag} */,
  {32'h3d8334d1, 32'h3d573a0f} /* (19, 4, 10) {real, imag} */,
  {32'h3d49ba20, 32'hbcc1b78e} /* (19, 4, 9) {real, imag} */,
  {32'hbd6d48f6, 32'h3cec0cb6} /* (19, 4, 8) {real, imag} */,
  {32'h3b03c980, 32'hbd877eac} /* (19, 4, 7) {real, imag} */,
  {32'h3cc6d9b0, 32'h3cfc7962} /* (19, 4, 6) {real, imag} */,
  {32'h3e73b035, 32'hbe42363d} /* (19, 4, 5) {real, imag} */,
  {32'h3e385d54, 32'h3da32689} /* (19, 4, 4) {real, imag} */,
  {32'h3dc21060, 32'h3d33aeb8} /* (19, 4, 3) {real, imag} */,
  {32'hbe9b0a8e, 32'h3f8dce0f} /* (19, 4, 2) {real, imag} */,
  {32'hc043fc7c, 32'hc05a2266} /* (19, 4, 1) {real, imag} */,
  {32'hc08d3c0a, 32'h00000000} /* (19, 4, 0) {real, imag} */,
  {32'hc0379e9f, 32'h406ad55a} /* (19, 3, 31) {real, imag} */,
  {32'hbec5989a, 32'hbfa11b56} /* (19, 3, 30) {real, imag} */,
  {32'h3cdc5e69, 32'hbe4a646e} /* (19, 3, 29) {real, imag} */,
  {32'h3e3c6192, 32'hbe2d91f0} /* (19, 3, 28) {real, imag} */,
  {32'h3e525656, 32'h3e280ae3} /* (19, 3, 27) {real, imag} */,
  {32'hbccdf6b8, 32'h3c8cfec4} /* (19, 3, 26) {real, imag} */,
  {32'hbd88b280, 32'hbd95069a} /* (19, 3, 25) {real, imag} */,
  {32'h3cb42c9f, 32'hb9679000} /* (19, 3, 24) {real, imag} */,
  {32'h3db96370, 32'hbdace434} /* (19, 3, 23) {real, imag} */,
  {32'hbd39189e, 32'hbd49ec9c} /* (19, 3, 22) {real, imag} */,
  {32'h3c8ac41a, 32'h3d2856c0} /* (19, 3, 21) {real, imag} */,
  {32'h3c47ac54, 32'hbcec5895} /* (19, 3, 20) {real, imag} */,
  {32'hbc57a18b, 32'h3da4e87c} /* (19, 3, 19) {real, imag} */,
  {32'h3d8963e2, 32'hbc82dbdc} /* (19, 3, 18) {real, imag} */,
  {32'hbcb086de, 32'hbb2f6d22} /* (19, 3, 17) {real, imag} */,
  {32'hbaaffe80, 32'h00000000} /* (19, 3, 16) {real, imag} */,
  {32'hbcb086de, 32'h3b2f6d22} /* (19, 3, 15) {real, imag} */,
  {32'h3d8963e2, 32'h3c82dbdc} /* (19, 3, 14) {real, imag} */,
  {32'hbc57a18b, 32'hbda4e87c} /* (19, 3, 13) {real, imag} */,
  {32'h3c47ac54, 32'h3cec5895} /* (19, 3, 12) {real, imag} */,
  {32'h3c8ac41a, 32'hbd2856c0} /* (19, 3, 11) {real, imag} */,
  {32'hbd39189e, 32'h3d49ec9c} /* (19, 3, 10) {real, imag} */,
  {32'h3db96370, 32'h3dace434} /* (19, 3, 9) {real, imag} */,
  {32'h3cb42c9f, 32'h39679000} /* (19, 3, 8) {real, imag} */,
  {32'hbd88b280, 32'h3d95069a} /* (19, 3, 7) {real, imag} */,
  {32'hbccdf6b8, 32'hbc8cfec4} /* (19, 3, 6) {real, imag} */,
  {32'h3e525656, 32'hbe280ae3} /* (19, 3, 5) {real, imag} */,
  {32'h3e3c6192, 32'h3e2d91f0} /* (19, 3, 4) {real, imag} */,
  {32'h3cdc5e69, 32'h3e4a646e} /* (19, 3, 3) {real, imag} */,
  {32'hbec5989a, 32'h3fa11b56} /* (19, 3, 2) {real, imag} */,
  {32'hc0379e9f, 32'hc06ad55a} /* (19, 3, 1) {real, imag} */,
  {32'hc08fbc9b, 32'h00000000} /* (19, 3, 0) {real, imag} */,
  {32'hc036a121, 32'h405df71c} /* (19, 2, 31) {real, imag} */,
  {32'hbee9084c, 32'hbf957f2a} /* (19, 2, 30) {real, imag} */,
  {32'h3cf2f560, 32'hbe3e8044} /* (19, 2, 29) {real, imag} */,
  {32'h3d908872, 32'hbe911941} /* (19, 2, 28) {real, imag} */,
  {32'h3e6f5eb8, 32'h3e67f0f8} /* (19, 2, 27) {real, imag} */,
  {32'h3dfb0e83, 32'hbde24b3b} /* (19, 2, 26) {real, imag} */,
  {32'hbd6be798, 32'hbc1356fc} /* (19, 2, 25) {real, imag} */,
  {32'h3e3ba7ae, 32'h3e0f7ae6} /* (19, 2, 24) {real, imag} */,
  {32'h3dabc51c, 32'hbda74150} /* (19, 2, 23) {real, imag} */,
  {32'h3d1bcecb, 32'hbd412ce8} /* (19, 2, 22) {real, imag} */,
  {32'h3d3efff6, 32'h3d08325b} /* (19, 2, 21) {real, imag} */,
  {32'h3d380c9b, 32'hbd32d332} /* (19, 2, 20) {real, imag} */,
  {32'hbd90dd38, 32'hbdde107c} /* (19, 2, 19) {real, imag} */,
  {32'h3c313114, 32'h3c6fe0aa} /* (19, 2, 18) {real, imag} */,
  {32'h3bd187a4, 32'h3cc53a3a} /* (19, 2, 17) {real, imag} */,
  {32'hbc0f347c, 32'h00000000} /* (19, 2, 16) {real, imag} */,
  {32'h3bd187a4, 32'hbcc53a3a} /* (19, 2, 15) {real, imag} */,
  {32'h3c313114, 32'hbc6fe0aa} /* (19, 2, 14) {real, imag} */,
  {32'hbd90dd38, 32'h3dde107c} /* (19, 2, 13) {real, imag} */,
  {32'h3d380c9b, 32'h3d32d332} /* (19, 2, 12) {real, imag} */,
  {32'h3d3efff6, 32'hbd08325b} /* (19, 2, 11) {real, imag} */,
  {32'h3d1bcecb, 32'h3d412ce8} /* (19, 2, 10) {real, imag} */,
  {32'h3dabc51c, 32'h3da74150} /* (19, 2, 9) {real, imag} */,
  {32'h3e3ba7ae, 32'hbe0f7ae6} /* (19, 2, 8) {real, imag} */,
  {32'hbd6be798, 32'h3c1356fc} /* (19, 2, 7) {real, imag} */,
  {32'h3dfb0e83, 32'h3de24b3b} /* (19, 2, 6) {real, imag} */,
  {32'h3e6f5eb8, 32'hbe67f0f8} /* (19, 2, 5) {real, imag} */,
  {32'h3d908872, 32'h3e911941} /* (19, 2, 4) {real, imag} */,
  {32'h3cf2f560, 32'h3e3e8044} /* (19, 2, 3) {real, imag} */,
  {32'hbee9084c, 32'h3f957f2a} /* (19, 2, 2) {real, imag} */,
  {32'hc036a121, 32'hc05df71c} /* (19, 2, 1) {real, imag} */,
  {32'hc096af9f, 32'h00000000} /* (19, 2, 0) {real, imag} */,
  {32'hc0422d01, 32'h404b56be} /* (19, 1, 31) {real, imag} */,
  {32'hbe946f6d, 32'hbf7c0826} /* (19, 1, 30) {real, imag} */,
  {32'h3dd82def, 32'hbdb211c8} /* (19, 1, 29) {real, imag} */,
  {32'h3daf613e, 32'hbe953ef6} /* (19, 1, 28) {real, imag} */,
  {32'h3e54e030, 32'h3dcd7aff} /* (19, 1, 27) {real, imag} */,
  {32'h3e0b5df5, 32'hbe4a3f4c} /* (19, 1, 26) {real, imag} */,
  {32'hbd0482be, 32'h3e151b5a} /* (19, 1, 25) {real, imag} */,
  {32'h3c73ccf8, 32'hbd4a10c6} /* (19, 1, 24) {real, imag} */,
  {32'hbd345bd6, 32'h3d63cd96} /* (19, 1, 23) {real, imag} */,
  {32'hbd8a81f5, 32'hbd67deea} /* (19, 1, 22) {real, imag} */,
  {32'hbdaf594e, 32'h3b989fe4} /* (19, 1, 21) {real, imag} */,
  {32'h3d02541a, 32'hbd424c50} /* (19, 1, 20) {real, imag} */,
  {32'h3d33da3c, 32'hbd1b4c0a} /* (19, 1, 19) {real, imag} */,
  {32'h3d43f24a, 32'hbcdf8965} /* (19, 1, 18) {real, imag} */,
  {32'h3bffb6a9, 32'h3cf27f23} /* (19, 1, 17) {real, imag} */,
  {32'h3d0bc4c1, 32'h00000000} /* (19, 1, 16) {real, imag} */,
  {32'h3bffb6a9, 32'hbcf27f23} /* (19, 1, 15) {real, imag} */,
  {32'h3d43f24a, 32'h3cdf8965} /* (19, 1, 14) {real, imag} */,
  {32'h3d33da3c, 32'h3d1b4c0a} /* (19, 1, 13) {real, imag} */,
  {32'h3d02541a, 32'h3d424c50} /* (19, 1, 12) {real, imag} */,
  {32'hbdaf594e, 32'hbb989fe4} /* (19, 1, 11) {real, imag} */,
  {32'hbd8a81f5, 32'h3d67deea} /* (19, 1, 10) {real, imag} */,
  {32'hbd345bd6, 32'hbd63cd96} /* (19, 1, 9) {real, imag} */,
  {32'h3c73ccf8, 32'h3d4a10c6} /* (19, 1, 8) {real, imag} */,
  {32'hbd0482be, 32'hbe151b5a} /* (19, 1, 7) {real, imag} */,
  {32'h3e0b5df5, 32'h3e4a3f4c} /* (19, 1, 6) {real, imag} */,
  {32'h3e54e030, 32'hbdcd7aff} /* (19, 1, 5) {real, imag} */,
  {32'h3daf613e, 32'h3e953ef6} /* (19, 1, 4) {real, imag} */,
  {32'h3dd82def, 32'h3db211c8} /* (19, 1, 3) {real, imag} */,
  {32'hbe946f6d, 32'h3f7c0826} /* (19, 1, 2) {real, imag} */,
  {32'hc0422d01, 32'hc04b56be} /* (19, 1, 1) {real, imag} */,
  {32'hc097a309, 32'h00000000} /* (19, 1, 0) {real, imag} */,
  {32'hc05214c8, 32'h4027e45c} /* (19, 0, 31) {real, imag} */,
  {32'h3db064c0, 32'hbf3ad0f4} /* (19, 0, 30) {real, imag} */,
  {32'h3d5c66e9, 32'hbd60dc5e} /* (19, 0, 29) {real, imag} */,
  {32'h3cd19244, 32'hbdea71e8} /* (19, 0, 28) {real, imag} */,
  {32'h3d39446c, 32'h3d1397a6} /* (19, 0, 27) {real, imag} */,
  {32'h3ce5a90e, 32'h3c51b11a} /* (19, 0, 26) {real, imag} */,
  {32'hbceebe82, 32'h3d63b6de} /* (19, 0, 25) {real, imag} */,
  {32'hbda81c08, 32'hbd5080b0} /* (19, 0, 24) {real, imag} */,
  {32'hbd074f35, 32'h3c0f6d04} /* (19, 0, 23) {real, imag} */,
  {32'h3c0d469c, 32'h3ba7adc0} /* (19, 0, 22) {real, imag} */,
  {32'h3d132eae, 32'h3cd6ffcc} /* (19, 0, 21) {real, imag} */,
  {32'h3be852e4, 32'hbc073574} /* (19, 0, 20) {real, imag} */,
  {32'h3c8d3a22, 32'h3b1a98e0} /* (19, 0, 19) {real, imag} */,
  {32'h3d1722aa, 32'hbd9b7a99} /* (19, 0, 18) {real, imag} */,
  {32'h3d32dd56, 32'hbcb26d43} /* (19, 0, 17) {real, imag} */,
  {32'h3d60bc9a, 32'h00000000} /* (19, 0, 16) {real, imag} */,
  {32'h3d32dd56, 32'h3cb26d43} /* (19, 0, 15) {real, imag} */,
  {32'h3d1722aa, 32'h3d9b7a99} /* (19, 0, 14) {real, imag} */,
  {32'h3c8d3a22, 32'hbb1a98e0} /* (19, 0, 13) {real, imag} */,
  {32'h3be852e4, 32'h3c073574} /* (19, 0, 12) {real, imag} */,
  {32'h3d132eae, 32'hbcd6ffcc} /* (19, 0, 11) {real, imag} */,
  {32'h3c0d469c, 32'hbba7adc0} /* (19, 0, 10) {real, imag} */,
  {32'hbd074f35, 32'hbc0f6d04} /* (19, 0, 9) {real, imag} */,
  {32'hbda81c08, 32'h3d5080b0} /* (19, 0, 8) {real, imag} */,
  {32'hbceebe82, 32'hbd63b6de} /* (19, 0, 7) {real, imag} */,
  {32'h3ce5a90e, 32'hbc51b11a} /* (19, 0, 6) {real, imag} */,
  {32'h3d39446c, 32'hbd1397a6} /* (19, 0, 5) {real, imag} */,
  {32'h3cd19244, 32'h3dea71e8} /* (19, 0, 4) {real, imag} */,
  {32'h3d5c66e9, 32'h3d60dc5e} /* (19, 0, 3) {real, imag} */,
  {32'h3db064c0, 32'h3f3ad0f4} /* (19, 0, 2) {real, imag} */,
  {32'hc05214c8, 32'hc027e45c} /* (19, 0, 1) {real, imag} */,
  {32'hc0907501, 32'h00000000} /* (19, 0, 0) {real, imag} */,
  {32'hc0485909, 32'h3fcd20fe} /* (18, 31, 31) {real, imag} */,
  {32'h3f1271f9, 32'hbef38109} /* (18, 31, 30) {real, imag} */,
  {32'h3dba7b6b, 32'h3da948ba} /* (18, 31, 29) {real, imag} */,
  {32'hbcc7dad9, 32'hbd2250da} /* (18, 31, 28) {real, imag} */,
  {32'h3d7a7fa2, 32'hbdb5a1ca} /* (18, 31, 27) {real, imag} */,
  {32'h3db42166, 32'h3af498f0} /* (18, 31, 26) {real, imag} */,
  {32'h3d23d509, 32'h3d3a506e} /* (18, 31, 25) {real, imag} */,
  {32'hbd195e25, 32'hbd2f5376} /* (18, 31, 24) {real, imag} */,
  {32'h3d583b66, 32'hbd465e42} /* (18, 31, 23) {real, imag} */,
  {32'hbcd7f8a1, 32'h3d92aaeb} /* (18, 31, 22) {real, imag} */,
  {32'hbc9927f6, 32'h3daaaf50} /* (18, 31, 21) {real, imag} */,
  {32'hbd91b142, 32'hbbdfde88} /* (18, 31, 20) {real, imag} */,
  {32'hbd3cd29a, 32'hbd783bbe} /* (18, 31, 19) {real, imag} */,
  {32'hbbe04298, 32'hbd9245a2} /* (18, 31, 18) {real, imag} */,
  {32'h3d0dbbb2, 32'h3c583d56} /* (18, 31, 17) {real, imag} */,
  {32'h3d1e888c, 32'h00000000} /* (18, 31, 16) {real, imag} */,
  {32'h3d0dbbb2, 32'hbc583d56} /* (18, 31, 15) {real, imag} */,
  {32'hbbe04298, 32'h3d9245a2} /* (18, 31, 14) {real, imag} */,
  {32'hbd3cd29a, 32'h3d783bbe} /* (18, 31, 13) {real, imag} */,
  {32'hbd91b142, 32'h3bdfde88} /* (18, 31, 12) {real, imag} */,
  {32'hbc9927f6, 32'hbdaaaf50} /* (18, 31, 11) {real, imag} */,
  {32'hbcd7f8a1, 32'hbd92aaeb} /* (18, 31, 10) {real, imag} */,
  {32'h3d583b66, 32'h3d465e42} /* (18, 31, 9) {real, imag} */,
  {32'hbd195e25, 32'h3d2f5376} /* (18, 31, 8) {real, imag} */,
  {32'h3d23d509, 32'hbd3a506e} /* (18, 31, 7) {real, imag} */,
  {32'h3db42166, 32'hbaf498f0} /* (18, 31, 6) {real, imag} */,
  {32'h3d7a7fa2, 32'h3db5a1ca} /* (18, 31, 5) {real, imag} */,
  {32'hbcc7dad9, 32'h3d2250da} /* (18, 31, 4) {real, imag} */,
  {32'h3dba7b6b, 32'hbda948ba} /* (18, 31, 3) {real, imag} */,
  {32'h3f1271f9, 32'h3ef38109} /* (18, 31, 2) {real, imag} */,
  {32'hc0485909, 32'hbfcd20fe} /* (18, 31, 1) {real, imag} */,
  {32'hc075da3e, 32'h00000000} /* (18, 31, 0) {real, imag} */,
  {32'hc07420a4, 32'h3fb46214} /* (18, 30, 31) {real, imag} */,
  {32'h3f75fd44, 32'hbec8ebf0} /* (18, 30, 30) {real, imag} */,
  {32'h3dc69b41, 32'h3e5a41e3} /* (18, 30, 29) {real, imag} */,
  {32'hbdc97f33, 32'h3d06de40} /* (18, 30, 28) {real, imag} */,
  {32'h3e51f0e8, 32'hbdca790b} /* (18, 30, 27) {real, imag} */,
  {32'h3d2da416, 32'h3bcfd876} /* (18, 30, 26) {real, imag} */,
  {32'h3d5ff5b2, 32'h3e0f1f64} /* (18, 30, 25) {real, imag} */,
  {32'h3d6782a8, 32'hbdad3ff6} /* (18, 30, 24) {real, imag} */,
  {32'h3d3f9596, 32'hbd85e9d2} /* (18, 30, 23) {real, imag} */,
  {32'hbcbe06a0, 32'h3d908893} /* (18, 30, 22) {real, imag} */,
  {32'hbd71b85d, 32'hbd9ff154} /* (18, 30, 21) {real, imag} */,
  {32'hbd555374, 32'h3c1294d4} /* (18, 30, 20) {real, imag} */,
  {32'h3dfcd8be, 32'h3dc03eb2} /* (18, 30, 19) {real, imag} */,
  {32'h3dbf950a, 32'h3d9d9e82} /* (18, 30, 18) {real, imag} */,
  {32'h3cb9196e, 32'h3c9e6a75} /* (18, 30, 17) {real, imag} */,
  {32'hbd6d8676, 32'h00000000} /* (18, 30, 16) {real, imag} */,
  {32'h3cb9196e, 32'hbc9e6a75} /* (18, 30, 15) {real, imag} */,
  {32'h3dbf950a, 32'hbd9d9e82} /* (18, 30, 14) {real, imag} */,
  {32'h3dfcd8be, 32'hbdc03eb2} /* (18, 30, 13) {real, imag} */,
  {32'hbd555374, 32'hbc1294d4} /* (18, 30, 12) {real, imag} */,
  {32'hbd71b85d, 32'h3d9ff154} /* (18, 30, 11) {real, imag} */,
  {32'hbcbe06a0, 32'hbd908893} /* (18, 30, 10) {real, imag} */,
  {32'h3d3f9596, 32'h3d85e9d2} /* (18, 30, 9) {real, imag} */,
  {32'h3d6782a8, 32'h3dad3ff6} /* (18, 30, 8) {real, imag} */,
  {32'h3d5ff5b2, 32'hbe0f1f64} /* (18, 30, 7) {real, imag} */,
  {32'h3d2da416, 32'hbbcfd876} /* (18, 30, 6) {real, imag} */,
  {32'h3e51f0e8, 32'h3dca790b} /* (18, 30, 5) {real, imag} */,
  {32'hbdc97f33, 32'hbd06de40} /* (18, 30, 4) {real, imag} */,
  {32'h3dc69b41, 32'hbe5a41e3} /* (18, 30, 3) {real, imag} */,
  {32'h3f75fd44, 32'h3ec8ebf0} /* (18, 30, 2) {real, imag} */,
  {32'hc07420a4, 32'hbfb46214} /* (18, 30, 1) {real, imag} */,
  {32'hc07b8391, 32'h00000000} /* (18, 30, 0) {real, imag} */,
  {32'hc081b6ac, 32'h3f8af024} /* (18, 29, 31) {real, imag} */,
  {32'h3f98a024, 32'hbedceb3e} /* (18, 29, 30) {real, imag} */,
  {32'h3ac3b2c0, 32'h3d3c1039} /* (18, 29, 29) {real, imag} */,
  {32'hbe231138, 32'h3df45228} /* (18, 29, 28) {real, imag} */,
  {32'h3dc52f29, 32'h3ce40ab4} /* (18, 29, 27) {real, imag} */,
  {32'h3e279f4c, 32'h3d934cd2} /* (18, 29, 26) {real, imag} */,
  {32'h3c973c95, 32'h3dde25da} /* (18, 29, 25) {real, imag} */,
  {32'h3cdf70df, 32'h3c16e826} /* (18, 29, 24) {real, imag} */,
  {32'hbe075cc7, 32'hbd0a7bd5} /* (18, 29, 23) {real, imag} */,
  {32'h3ce1bf26, 32'hbda8ae9b} /* (18, 29, 22) {real, imag} */,
  {32'hbd527046, 32'hbdc56f68} /* (18, 29, 21) {real, imag} */,
  {32'hbd7ec09d, 32'hbd4fac4a} /* (18, 29, 20) {real, imag} */,
  {32'hbc162eea, 32'hbc92b87f} /* (18, 29, 19) {real, imag} */,
  {32'h3a3d66c8, 32'hbd8754ee} /* (18, 29, 18) {real, imag} */,
  {32'hbbd80fbc, 32'h3cb263a6} /* (18, 29, 17) {real, imag} */,
  {32'h3cb6b657, 32'h00000000} /* (18, 29, 16) {real, imag} */,
  {32'hbbd80fbc, 32'hbcb263a6} /* (18, 29, 15) {real, imag} */,
  {32'h3a3d66c8, 32'h3d8754ee} /* (18, 29, 14) {real, imag} */,
  {32'hbc162eea, 32'h3c92b87f} /* (18, 29, 13) {real, imag} */,
  {32'hbd7ec09d, 32'h3d4fac4a} /* (18, 29, 12) {real, imag} */,
  {32'hbd527046, 32'h3dc56f68} /* (18, 29, 11) {real, imag} */,
  {32'h3ce1bf26, 32'h3da8ae9b} /* (18, 29, 10) {real, imag} */,
  {32'hbe075cc7, 32'h3d0a7bd5} /* (18, 29, 9) {real, imag} */,
  {32'h3cdf70df, 32'hbc16e826} /* (18, 29, 8) {real, imag} */,
  {32'h3c973c95, 32'hbdde25da} /* (18, 29, 7) {real, imag} */,
  {32'h3e279f4c, 32'hbd934cd2} /* (18, 29, 6) {real, imag} */,
  {32'h3dc52f29, 32'hbce40ab4} /* (18, 29, 5) {real, imag} */,
  {32'hbe231138, 32'hbdf45228} /* (18, 29, 4) {real, imag} */,
  {32'h3ac3b2c0, 32'hbd3c1039} /* (18, 29, 3) {real, imag} */,
  {32'h3f98a024, 32'h3edceb3e} /* (18, 29, 2) {real, imag} */,
  {32'hc081b6ac, 32'hbf8af024} /* (18, 29, 1) {real, imag} */,
  {32'hc07e2241, 32'h00000000} /* (18, 29, 0) {real, imag} */,
  {32'hc084f7a1, 32'h3f764337} /* (18, 28, 31) {real, imag} */,
  {32'h3fb80218, 32'hbefb5fc4} /* (18, 28, 30) {real, imag} */,
  {32'h3bfda580, 32'hbd697808} /* (18, 28, 29) {real, imag} */,
  {32'hbe6c614b, 32'h3dd260d8} /* (18, 28, 28) {real, imag} */,
  {32'h3d8b8d82, 32'hbd49c079} /* (18, 28, 27) {real, imag} */,
  {32'h3dfc5082, 32'h3bb95f74} /* (18, 28, 26) {real, imag} */,
  {32'hbd104c32, 32'hbdf2398a} /* (18, 28, 25) {real, imag} */,
  {32'hbbf46cdc, 32'hbdd1a35f} /* (18, 28, 24) {real, imag} */,
  {32'hbc98246c, 32'h3df28c1c} /* (18, 28, 23) {real, imag} */,
  {32'hbdb5f1ca, 32'h3ccea5ea} /* (18, 28, 22) {real, imag} */,
  {32'h3d608428, 32'hbd9c11ee} /* (18, 28, 21) {real, imag} */,
  {32'hbb5cfc94, 32'h3c2bef64} /* (18, 28, 20) {real, imag} */,
  {32'hbd48261e, 32'h3b21f7d0} /* (18, 28, 19) {real, imag} */,
  {32'hbc074b9c, 32'hbd064eb2} /* (18, 28, 18) {real, imag} */,
  {32'hbcd030ff, 32'hbb9b24b0} /* (18, 28, 17) {real, imag} */,
  {32'h3c04fbcc, 32'h00000000} /* (18, 28, 16) {real, imag} */,
  {32'hbcd030ff, 32'h3b9b24b0} /* (18, 28, 15) {real, imag} */,
  {32'hbc074b9c, 32'h3d064eb2} /* (18, 28, 14) {real, imag} */,
  {32'hbd48261e, 32'hbb21f7d0} /* (18, 28, 13) {real, imag} */,
  {32'hbb5cfc94, 32'hbc2bef64} /* (18, 28, 12) {real, imag} */,
  {32'h3d608428, 32'h3d9c11ee} /* (18, 28, 11) {real, imag} */,
  {32'hbdb5f1ca, 32'hbccea5ea} /* (18, 28, 10) {real, imag} */,
  {32'hbc98246c, 32'hbdf28c1c} /* (18, 28, 9) {real, imag} */,
  {32'hbbf46cdc, 32'h3dd1a35f} /* (18, 28, 8) {real, imag} */,
  {32'hbd104c32, 32'h3df2398a} /* (18, 28, 7) {real, imag} */,
  {32'h3dfc5082, 32'hbbb95f74} /* (18, 28, 6) {real, imag} */,
  {32'h3d8b8d82, 32'h3d49c079} /* (18, 28, 5) {real, imag} */,
  {32'hbe6c614b, 32'hbdd260d8} /* (18, 28, 4) {real, imag} */,
  {32'h3bfda580, 32'h3d697808} /* (18, 28, 3) {real, imag} */,
  {32'h3fb80218, 32'h3efb5fc4} /* (18, 28, 2) {real, imag} */,
  {32'hc084f7a1, 32'hbf764337} /* (18, 28, 1) {real, imag} */,
  {32'hc081e0fa, 32'h00000000} /* (18, 28, 0) {real, imag} */,
  {32'hc08429df, 32'h3f28df60} /* (18, 27, 31) {real, imag} */,
  {32'h3fbf1e69, 32'hbf048e8a} /* (18, 27, 30) {real, imag} */,
  {32'h3d1b2b12, 32'hbcb72595} /* (18, 27, 29) {real, imag} */,
  {32'hbe5a7d90, 32'hbd1a921e} /* (18, 27, 28) {real, imag} */,
  {32'h3db7cd00, 32'h3c643ad4} /* (18, 27, 27) {real, imag} */,
  {32'hbd5da1e0, 32'h3dd4785e} /* (18, 27, 26) {real, imag} */,
  {32'h3b8d7cac, 32'hbc865142} /* (18, 27, 25) {real, imag} */,
  {32'hbc976db7, 32'hbddb4484} /* (18, 27, 24) {real, imag} */,
  {32'h3cabea79, 32'hbdc947ce} /* (18, 27, 23) {real, imag} */,
  {32'hbce8078a, 32'h3c876187} /* (18, 27, 22) {real, imag} */,
  {32'h3d6b72eb, 32'hbd9933d4} /* (18, 27, 21) {real, imag} */,
  {32'h3db4beaa, 32'h3d40036c} /* (18, 27, 20) {real, imag} */,
  {32'h3c6d3b8a, 32'hbd1e8303} /* (18, 27, 19) {real, imag} */,
  {32'h3d2c46a4, 32'hbd058394} /* (18, 27, 18) {real, imag} */,
  {32'hbc0ec83e, 32'hbc9c8f2d} /* (18, 27, 17) {real, imag} */,
  {32'h3ca6f2dc, 32'h00000000} /* (18, 27, 16) {real, imag} */,
  {32'hbc0ec83e, 32'h3c9c8f2d} /* (18, 27, 15) {real, imag} */,
  {32'h3d2c46a4, 32'h3d058394} /* (18, 27, 14) {real, imag} */,
  {32'h3c6d3b8a, 32'h3d1e8303} /* (18, 27, 13) {real, imag} */,
  {32'h3db4beaa, 32'hbd40036c} /* (18, 27, 12) {real, imag} */,
  {32'h3d6b72eb, 32'h3d9933d4} /* (18, 27, 11) {real, imag} */,
  {32'hbce8078a, 32'hbc876187} /* (18, 27, 10) {real, imag} */,
  {32'h3cabea79, 32'h3dc947ce} /* (18, 27, 9) {real, imag} */,
  {32'hbc976db7, 32'h3ddb4484} /* (18, 27, 8) {real, imag} */,
  {32'h3b8d7cac, 32'h3c865142} /* (18, 27, 7) {real, imag} */,
  {32'hbd5da1e0, 32'hbdd4785e} /* (18, 27, 6) {real, imag} */,
  {32'h3db7cd00, 32'hbc643ad4} /* (18, 27, 5) {real, imag} */,
  {32'hbe5a7d90, 32'h3d1a921e} /* (18, 27, 4) {real, imag} */,
  {32'h3d1b2b12, 32'h3cb72595} /* (18, 27, 3) {real, imag} */,
  {32'h3fbf1e69, 32'h3f048e8a} /* (18, 27, 2) {real, imag} */,
  {32'hc08429df, 32'hbf28df60} /* (18, 27, 1) {real, imag} */,
  {32'hc081594d, 32'h00000000} /* (18, 27, 0) {real, imag} */,
  {32'hc07dcd48, 32'h3f07282c} /* (18, 26, 31) {real, imag} */,
  {32'h3fb2d5e9, 32'hbf0f3042} /* (18, 26, 30) {real, imag} */,
  {32'hbd233766, 32'hbd0e6d82} /* (18, 26, 29) {real, imag} */,
  {32'hbe898ac8, 32'hbd893597} /* (18, 26, 28) {real, imag} */,
  {32'h3dce28f2, 32'hbcfa29ae} /* (18, 26, 27) {real, imag} */,
  {32'h3cb70e2d, 32'h3d81fe06} /* (18, 26, 26) {real, imag} */,
  {32'h3cd42cec, 32'h3b9a6dc4} /* (18, 26, 25) {real, imag} */,
  {32'h3d451530, 32'hbde32530} /* (18, 26, 24) {real, imag} */,
  {32'hbcf93996, 32'hbd8ad9f6} /* (18, 26, 23) {real, imag} */,
  {32'h3d9fa1de, 32'hbcbfcc56} /* (18, 26, 22) {real, imag} */,
  {32'h3d4226e2, 32'h3c8a424d} /* (18, 26, 21) {real, imag} */,
  {32'h3d7744a3, 32'h3d366ed0} /* (18, 26, 20) {real, imag} */,
  {32'hbdb54612, 32'hbd36315e} /* (18, 26, 19) {real, imag} */,
  {32'h3db08157, 32'hbd332cb6} /* (18, 26, 18) {real, imag} */,
  {32'hbd1e07a1, 32'h3a76d6c0} /* (18, 26, 17) {real, imag} */,
  {32'h3d1d1152, 32'h00000000} /* (18, 26, 16) {real, imag} */,
  {32'hbd1e07a1, 32'hba76d6c0} /* (18, 26, 15) {real, imag} */,
  {32'h3db08157, 32'h3d332cb6} /* (18, 26, 14) {real, imag} */,
  {32'hbdb54612, 32'h3d36315e} /* (18, 26, 13) {real, imag} */,
  {32'h3d7744a3, 32'hbd366ed0} /* (18, 26, 12) {real, imag} */,
  {32'h3d4226e2, 32'hbc8a424d} /* (18, 26, 11) {real, imag} */,
  {32'h3d9fa1de, 32'h3cbfcc56} /* (18, 26, 10) {real, imag} */,
  {32'hbcf93996, 32'h3d8ad9f6} /* (18, 26, 9) {real, imag} */,
  {32'h3d451530, 32'h3de32530} /* (18, 26, 8) {real, imag} */,
  {32'h3cd42cec, 32'hbb9a6dc4} /* (18, 26, 7) {real, imag} */,
  {32'h3cb70e2d, 32'hbd81fe06} /* (18, 26, 6) {real, imag} */,
  {32'h3dce28f2, 32'h3cfa29ae} /* (18, 26, 5) {real, imag} */,
  {32'hbe898ac8, 32'h3d893597} /* (18, 26, 4) {real, imag} */,
  {32'hbd233766, 32'h3d0e6d82} /* (18, 26, 3) {real, imag} */,
  {32'h3fb2d5e9, 32'h3f0f3042} /* (18, 26, 2) {real, imag} */,
  {32'hc07dcd48, 32'hbf07282c} /* (18, 26, 1) {real, imag} */,
  {32'hc0806fe4, 32'h00000000} /* (18, 26, 0) {real, imag} */,
  {32'hc06d031c, 32'h3ed63550} /* (18, 25, 31) {real, imag} */,
  {32'h3fae8b52, 32'hbe815ce8} /* (18, 25, 30) {real, imag} */,
  {32'h3d9e27c2, 32'hbd6d72f1} /* (18, 25, 29) {real, imag} */,
  {32'hbed19550, 32'hbdaa2bb8} /* (18, 25, 28) {real, imag} */,
  {32'h3e718903, 32'hbe858523} /* (18, 25, 27) {real, imag} */,
  {32'hbde5ae0c, 32'hbd681d47} /* (18, 25, 26) {real, imag} */,
  {32'hbce537d8, 32'h3e48df32} /* (18, 25, 25) {real, imag} */,
  {32'h3e15cc26, 32'hbde33ff1} /* (18, 25, 24) {real, imag} */,
  {32'hbd9b6b1f, 32'h3d68c9f6} /* (18, 25, 23) {real, imag} */,
  {32'h3e00da9b, 32'hbe117666} /* (18, 25, 22) {real, imag} */,
  {32'hbd1b14c1, 32'hbdd765b3} /* (18, 25, 21) {real, imag} */,
  {32'hbd5a0de9, 32'h3e394612} /* (18, 25, 20) {real, imag} */,
  {32'h3db36809, 32'hbda15c27} /* (18, 25, 19) {real, imag} */,
  {32'h3c6f905c, 32'h3c86dd74} /* (18, 25, 18) {real, imag} */,
  {32'h3c22831a, 32'h3cabdcb4} /* (18, 25, 17) {real, imag} */,
  {32'h3dc41d80, 32'h00000000} /* (18, 25, 16) {real, imag} */,
  {32'h3c22831a, 32'hbcabdcb4} /* (18, 25, 15) {real, imag} */,
  {32'h3c6f905c, 32'hbc86dd74} /* (18, 25, 14) {real, imag} */,
  {32'h3db36809, 32'h3da15c27} /* (18, 25, 13) {real, imag} */,
  {32'hbd5a0de9, 32'hbe394612} /* (18, 25, 12) {real, imag} */,
  {32'hbd1b14c1, 32'h3dd765b3} /* (18, 25, 11) {real, imag} */,
  {32'h3e00da9b, 32'h3e117666} /* (18, 25, 10) {real, imag} */,
  {32'hbd9b6b1f, 32'hbd68c9f6} /* (18, 25, 9) {real, imag} */,
  {32'h3e15cc26, 32'h3de33ff1} /* (18, 25, 8) {real, imag} */,
  {32'hbce537d8, 32'hbe48df32} /* (18, 25, 7) {real, imag} */,
  {32'hbde5ae0c, 32'h3d681d47} /* (18, 25, 6) {real, imag} */,
  {32'h3e718903, 32'h3e858523} /* (18, 25, 5) {real, imag} */,
  {32'hbed19550, 32'h3daa2bb8} /* (18, 25, 4) {real, imag} */,
  {32'h3d9e27c2, 32'h3d6d72f1} /* (18, 25, 3) {real, imag} */,
  {32'h3fae8b52, 32'h3e815ce8} /* (18, 25, 2) {real, imag} */,
  {32'hc06d031c, 32'hbed63550} /* (18, 25, 1) {real, imag} */,
  {32'hc06b02bc, 32'h00000000} /* (18, 25, 0) {real, imag} */,
  {32'hc04e023e, 32'h3e81a1c8} /* (18, 24, 31) {real, imag} */,
  {32'h3fa2c872, 32'hbe1b0720} /* (18, 24, 30) {real, imag} */,
  {32'hbb4fc8d0, 32'hbdeb1202} /* (18, 24, 29) {real, imag} */,
  {32'hbea4f64b, 32'hbcd247f4} /* (18, 24, 28) {real, imag} */,
  {32'h3e859b66, 32'hbe284f00} /* (18, 24, 27) {real, imag} */,
  {32'hbd8ab50c, 32'hbdb9ecc8} /* (18, 24, 26) {real, imag} */,
  {32'hbbfc6798, 32'h3dd71060} /* (18, 24, 25) {real, imag} */,
  {32'h3dba11eb, 32'hbd1ca4aa} /* (18, 24, 24) {real, imag} */,
  {32'hbdc30f30, 32'hba6d0770} /* (18, 24, 23) {real, imag} */,
  {32'h3c7e0d90, 32'h3d0a6ad2} /* (18, 24, 22) {real, imag} */,
  {32'h3cb456a8, 32'hbddc36fe} /* (18, 24, 21) {real, imag} */,
  {32'h3d9c4b04, 32'h3d81a9c4} /* (18, 24, 20) {real, imag} */,
  {32'h3d4c7434, 32'h3d2d5766} /* (18, 24, 19) {real, imag} */,
  {32'h3ceac914, 32'hbd37ab1b} /* (18, 24, 18) {real, imag} */,
  {32'h3d5983bc, 32'hbc61e479} /* (18, 24, 17) {real, imag} */,
  {32'hbda8d139, 32'h00000000} /* (18, 24, 16) {real, imag} */,
  {32'h3d5983bc, 32'h3c61e479} /* (18, 24, 15) {real, imag} */,
  {32'h3ceac914, 32'h3d37ab1b} /* (18, 24, 14) {real, imag} */,
  {32'h3d4c7434, 32'hbd2d5766} /* (18, 24, 13) {real, imag} */,
  {32'h3d9c4b04, 32'hbd81a9c4} /* (18, 24, 12) {real, imag} */,
  {32'h3cb456a8, 32'h3ddc36fe} /* (18, 24, 11) {real, imag} */,
  {32'h3c7e0d90, 32'hbd0a6ad2} /* (18, 24, 10) {real, imag} */,
  {32'hbdc30f30, 32'h3a6d0770} /* (18, 24, 9) {real, imag} */,
  {32'h3dba11eb, 32'h3d1ca4aa} /* (18, 24, 8) {real, imag} */,
  {32'hbbfc6798, 32'hbdd71060} /* (18, 24, 7) {real, imag} */,
  {32'hbd8ab50c, 32'h3db9ecc8} /* (18, 24, 6) {real, imag} */,
  {32'h3e859b66, 32'h3e284f00} /* (18, 24, 5) {real, imag} */,
  {32'hbea4f64b, 32'h3cd247f4} /* (18, 24, 4) {real, imag} */,
  {32'hbb4fc8d0, 32'h3deb1202} /* (18, 24, 3) {real, imag} */,
  {32'h3fa2c872, 32'h3e1b0720} /* (18, 24, 2) {real, imag} */,
  {32'hc04e023e, 32'hbe81a1c8} /* (18, 24, 1) {real, imag} */,
  {32'hc05568d0, 32'h00000000} /* (18, 24, 0) {real, imag} */,
  {32'hc02c152a, 32'h3e547600} /* (18, 23, 31) {real, imag} */,
  {32'h3f91b6d8, 32'hbe3c5cdc} /* (18, 23, 30) {real, imag} */,
  {32'hbde52a56, 32'hbe007e8b} /* (18, 23, 29) {real, imag} */,
  {32'hbe23a7d6, 32'hbd4b4228} /* (18, 23, 28) {real, imag} */,
  {32'h3e81d14a, 32'hbe112f15} /* (18, 23, 27) {real, imag} */,
  {32'h3db45d4e, 32'hbd850af5} /* (18, 23, 26) {real, imag} */,
  {32'hbd9fd136, 32'hbd160803} /* (18, 23, 25) {real, imag} */,
  {32'h3de8a390, 32'h3be8fe50} /* (18, 23, 24) {real, imag} */,
  {32'hbdda3ec1, 32'h3d0b4763} /* (18, 23, 23) {real, imag} */,
  {32'h3cbc459e, 32'h3d69c690} /* (18, 23, 22) {real, imag} */,
  {32'h3dbf4250, 32'hbd5caf4c} /* (18, 23, 21) {real, imag} */,
  {32'hbcc4dfb6, 32'h3d057f5a} /* (18, 23, 20) {real, imag} */,
  {32'h3c91c4bc, 32'h3d077514} /* (18, 23, 19) {real, imag} */,
  {32'h3ba4bd8c, 32'h3c0cb596} /* (18, 23, 18) {real, imag} */,
  {32'hbcc9700e, 32'hbcf30e84} /* (18, 23, 17) {real, imag} */,
  {32'hbd9f2a8d, 32'h00000000} /* (18, 23, 16) {real, imag} */,
  {32'hbcc9700e, 32'h3cf30e84} /* (18, 23, 15) {real, imag} */,
  {32'h3ba4bd8c, 32'hbc0cb596} /* (18, 23, 14) {real, imag} */,
  {32'h3c91c4bc, 32'hbd077514} /* (18, 23, 13) {real, imag} */,
  {32'hbcc4dfb6, 32'hbd057f5a} /* (18, 23, 12) {real, imag} */,
  {32'h3dbf4250, 32'h3d5caf4c} /* (18, 23, 11) {real, imag} */,
  {32'h3cbc459e, 32'hbd69c690} /* (18, 23, 10) {real, imag} */,
  {32'hbdda3ec1, 32'hbd0b4763} /* (18, 23, 9) {real, imag} */,
  {32'h3de8a390, 32'hbbe8fe50} /* (18, 23, 8) {real, imag} */,
  {32'hbd9fd136, 32'h3d160803} /* (18, 23, 7) {real, imag} */,
  {32'h3db45d4e, 32'h3d850af5} /* (18, 23, 6) {real, imag} */,
  {32'h3e81d14a, 32'h3e112f15} /* (18, 23, 5) {real, imag} */,
  {32'hbe23a7d6, 32'h3d4b4228} /* (18, 23, 4) {real, imag} */,
  {32'hbde52a56, 32'h3e007e8b} /* (18, 23, 3) {real, imag} */,
  {32'h3f91b6d8, 32'h3e3c5cdc} /* (18, 23, 2) {real, imag} */,
  {32'hc02c152a, 32'hbe547600} /* (18, 23, 1) {real, imag} */,
  {32'hc02d7d72, 32'h00000000} /* (18, 23, 0) {real, imag} */,
  {32'hbff92926, 32'h3e2caabe} /* (18, 22, 31) {real, imag} */,
  {32'h3f6643bd, 32'hbcfe2d80} /* (18, 22, 30) {real, imag} */,
  {32'hbe295874, 32'h3d1064bd} /* (18, 22, 29) {real, imag} */,
  {32'hbc396dc8, 32'h3d239474} /* (18, 22, 28) {real, imag} */,
  {32'h3df4131d, 32'hbe43e0b4} /* (18, 22, 27) {real, imag} */,
  {32'hbd0811aa, 32'hbdf6d140} /* (18, 22, 26) {real, imag} */,
  {32'hbe1d7913, 32'hbd436959} /* (18, 22, 25) {real, imag} */,
  {32'h3b9c6c64, 32'h3dae8a30} /* (18, 22, 24) {real, imag} */,
  {32'h3c29f4c0, 32'hbacbca20} /* (18, 22, 23) {real, imag} */,
  {32'h3c8a00cf, 32'hbd37ca14} /* (18, 22, 22) {real, imag} */,
  {32'h3ca15da9, 32'h3c2292b8} /* (18, 22, 21) {real, imag} */,
  {32'hbd07d70b, 32'h3d18f3f6} /* (18, 22, 20) {real, imag} */,
  {32'h3d007c55, 32'hbd9700ce} /* (18, 22, 19) {real, imag} */,
  {32'h3ca0683b, 32'hbc0a7d4a} /* (18, 22, 18) {real, imag} */,
  {32'hbc2653c8, 32'hbd4e98d1} /* (18, 22, 17) {real, imag} */,
  {32'h3d163652, 32'h00000000} /* (18, 22, 16) {real, imag} */,
  {32'hbc2653c8, 32'h3d4e98d1} /* (18, 22, 15) {real, imag} */,
  {32'h3ca0683b, 32'h3c0a7d4a} /* (18, 22, 14) {real, imag} */,
  {32'h3d007c55, 32'h3d9700ce} /* (18, 22, 13) {real, imag} */,
  {32'hbd07d70b, 32'hbd18f3f6} /* (18, 22, 12) {real, imag} */,
  {32'h3ca15da9, 32'hbc2292b8} /* (18, 22, 11) {real, imag} */,
  {32'h3c8a00cf, 32'h3d37ca14} /* (18, 22, 10) {real, imag} */,
  {32'h3c29f4c0, 32'h3acbca20} /* (18, 22, 9) {real, imag} */,
  {32'h3b9c6c64, 32'hbdae8a30} /* (18, 22, 8) {real, imag} */,
  {32'hbe1d7913, 32'h3d436959} /* (18, 22, 7) {real, imag} */,
  {32'hbd0811aa, 32'h3df6d140} /* (18, 22, 6) {real, imag} */,
  {32'h3df4131d, 32'h3e43e0b4} /* (18, 22, 5) {real, imag} */,
  {32'hbc396dc8, 32'hbd239474} /* (18, 22, 4) {real, imag} */,
  {32'hbe295874, 32'hbd1064bd} /* (18, 22, 3) {real, imag} */,
  {32'h3f6643bd, 32'h3cfe2d80} /* (18, 22, 2) {real, imag} */,
  {32'hbff92926, 32'hbe2caabe} /* (18, 22, 1) {real, imag} */,
  {32'hc0034fe4, 32'h00000000} /* (18, 22, 0) {real, imag} */,
  {32'hbf40a4bb, 32'h3e18d112} /* (18, 21, 31) {real, imag} */,
  {32'h3e99ce8e, 32'h3e0634ae} /* (18, 21, 30) {real, imag} */,
  {32'hbdb1785a, 32'h3d1b0220} /* (18, 21, 29) {real, imag} */,
  {32'hbcbca76a, 32'h3d3b7c7a} /* (18, 21, 28) {real, imag} */,
  {32'h3d74c374, 32'hbdebe66e} /* (18, 21, 27) {real, imag} */,
  {32'hbd5cfe1a, 32'h3cbb0956} /* (18, 21, 26) {real, imag} */,
  {32'h3d54aea2, 32'h3d92c276} /* (18, 21, 25) {real, imag} */,
  {32'h3d883785, 32'hbd5f77ac} /* (18, 21, 24) {real, imag} */,
  {32'h3d2076f8, 32'hbd101fcc} /* (18, 21, 23) {real, imag} */,
  {32'h3da9e936, 32'hbd9945f7} /* (18, 21, 22) {real, imag} */,
  {32'h3ca42be0, 32'hbdaa2bfb} /* (18, 21, 21) {real, imag} */,
  {32'h3d4d2e90, 32'h397c4280} /* (18, 21, 20) {real, imag} */,
  {32'h3c1e75a2, 32'h3c610305} /* (18, 21, 19) {real, imag} */,
  {32'hbccbbecc, 32'hbc34f4b0} /* (18, 21, 18) {real, imag} */,
  {32'h3b577d58, 32'h3c939ba8} /* (18, 21, 17) {real, imag} */,
  {32'h3bcd8ca6, 32'h00000000} /* (18, 21, 16) {real, imag} */,
  {32'h3b577d58, 32'hbc939ba8} /* (18, 21, 15) {real, imag} */,
  {32'hbccbbecc, 32'h3c34f4b0} /* (18, 21, 14) {real, imag} */,
  {32'h3c1e75a2, 32'hbc610305} /* (18, 21, 13) {real, imag} */,
  {32'h3d4d2e90, 32'hb97c4280} /* (18, 21, 12) {real, imag} */,
  {32'h3ca42be0, 32'h3daa2bfb} /* (18, 21, 11) {real, imag} */,
  {32'h3da9e936, 32'h3d9945f7} /* (18, 21, 10) {real, imag} */,
  {32'h3d2076f8, 32'h3d101fcc} /* (18, 21, 9) {real, imag} */,
  {32'h3d883785, 32'h3d5f77ac} /* (18, 21, 8) {real, imag} */,
  {32'h3d54aea2, 32'hbd92c276} /* (18, 21, 7) {real, imag} */,
  {32'hbd5cfe1a, 32'hbcbb0956} /* (18, 21, 6) {real, imag} */,
  {32'h3d74c374, 32'h3debe66e} /* (18, 21, 5) {real, imag} */,
  {32'hbcbca76a, 32'hbd3b7c7a} /* (18, 21, 4) {real, imag} */,
  {32'hbdb1785a, 32'hbd1b0220} /* (18, 21, 3) {real, imag} */,
  {32'h3e99ce8e, 32'hbe0634ae} /* (18, 21, 2) {real, imag} */,
  {32'hbf40a4bb, 32'hbe18d112} /* (18, 21, 1) {real, imag} */,
  {32'hbf94b6f6, 32'h00000000} /* (18, 21, 0) {real, imag} */,
  {32'h3f5d2809, 32'hbc98e660} /* (18, 20, 31) {real, imag} */,
  {32'hbebf33f6, 32'h3ea2ba84} /* (18, 20, 30) {real, imag} */,
  {32'hbc644590, 32'h3ca95ab4} /* (18, 20, 29) {real, imag} */,
  {32'h3e6670fd, 32'h3cc4629b} /* (18, 20, 28) {real, imag} */,
  {32'hbdc4ef9c, 32'h3db2d91b} /* (18, 20, 27) {real, imag} */,
  {32'hbe0ec652, 32'h3d76cccf} /* (18, 20, 26) {real, imag} */,
  {32'h3e0f5fa0, 32'hbd9218ce} /* (18, 20, 25) {real, imag} */,
  {32'h3d052613, 32'hbdbf5ed8} /* (18, 20, 24) {real, imag} */,
  {32'hbc7a02d8, 32'h3c63fa6a} /* (18, 20, 23) {real, imag} */,
  {32'h3d0bb436, 32'h3cd2800d} /* (18, 20, 22) {real, imag} */,
  {32'hbd57dbd4, 32'hbcae3fa8} /* (18, 20, 21) {real, imag} */,
  {32'hbd1f98de, 32'hbd3c76c4} /* (18, 20, 20) {real, imag} */,
  {32'h3db9564c, 32'h3b6b0f60} /* (18, 20, 19) {real, imag} */,
  {32'hbc8676a6, 32'h3d398fa9} /* (18, 20, 18) {real, imag} */,
  {32'h3d5a2cb2, 32'hbd32c01d} /* (18, 20, 17) {real, imag} */,
  {32'hbc4b7870, 32'h00000000} /* (18, 20, 16) {real, imag} */,
  {32'h3d5a2cb2, 32'h3d32c01d} /* (18, 20, 15) {real, imag} */,
  {32'hbc8676a6, 32'hbd398fa9} /* (18, 20, 14) {real, imag} */,
  {32'h3db9564c, 32'hbb6b0f60} /* (18, 20, 13) {real, imag} */,
  {32'hbd1f98de, 32'h3d3c76c4} /* (18, 20, 12) {real, imag} */,
  {32'hbd57dbd4, 32'h3cae3fa8} /* (18, 20, 11) {real, imag} */,
  {32'h3d0bb436, 32'hbcd2800d} /* (18, 20, 10) {real, imag} */,
  {32'hbc7a02d8, 32'hbc63fa6a} /* (18, 20, 9) {real, imag} */,
  {32'h3d052613, 32'h3dbf5ed8} /* (18, 20, 8) {real, imag} */,
  {32'h3e0f5fa0, 32'h3d9218ce} /* (18, 20, 7) {real, imag} */,
  {32'hbe0ec652, 32'hbd76cccf} /* (18, 20, 6) {real, imag} */,
  {32'hbdc4ef9c, 32'hbdb2d91b} /* (18, 20, 5) {real, imag} */,
  {32'h3e6670fd, 32'hbcc4629b} /* (18, 20, 4) {real, imag} */,
  {32'hbc644590, 32'hbca95ab4} /* (18, 20, 3) {real, imag} */,
  {32'hbebf33f6, 32'hbea2ba84} /* (18, 20, 2) {real, imag} */,
  {32'h3f5d2809, 32'h3c98e660} /* (18, 20, 1) {real, imag} */,
  {32'h3e1848bc, 32'h00000000} /* (18, 20, 0) {real, imag} */,
  {32'h3ffc919e, 32'hbdf6050c} /* (18, 19, 31) {real, imag} */,
  {32'hbf4dfd48, 32'h3e8b66fa} /* (18, 19, 30) {real, imag} */,
  {32'hbcd09e60, 32'h3d802130} /* (18, 19, 29) {real, imag} */,
  {32'h3ebb2050, 32'hbd877edf} /* (18, 19, 28) {real, imag} */,
  {32'hbe00d0ec, 32'h3e068c87} /* (18, 19, 27) {real, imag} */,
  {32'hbe3a8ea1, 32'h3dcd0b53} /* (18, 19, 26) {real, imag} */,
  {32'h3d3c0cb7, 32'hbce7ae12} /* (18, 19, 25) {real, imag} */,
  {32'hbbee6214, 32'h3d5e2d44} /* (18, 19, 24) {real, imag} */,
  {32'hbc2dc722, 32'h3d8058e3} /* (18, 19, 23) {real, imag} */,
  {32'hbd8dd71e, 32'hbd9d759c} /* (18, 19, 22) {real, imag} */,
  {32'hbde8a810, 32'h3de9cae3} /* (18, 19, 21) {real, imag} */,
  {32'h3c6a88db, 32'hbd01513a} /* (18, 19, 20) {real, imag} */,
  {32'hbd8d975e, 32'hbdaeae05} /* (18, 19, 19) {real, imag} */,
  {32'h3c12a635, 32'h3cea7988} /* (18, 19, 18) {real, imag} */,
  {32'hbb091800, 32'h3cae8af6} /* (18, 19, 17) {real, imag} */,
  {32'h3d5312ea, 32'h00000000} /* (18, 19, 16) {real, imag} */,
  {32'hbb091800, 32'hbcae8af6} /* (18, 19, 15) {real, imag} */,
  {32'h3c12a635, 32'hbcea7988} /* (18, 19, 14) {real, imag} */,
  {32'hbd8d975e, 32'h3daeae05} /* (18, 19, 13) {real, imag} */,
  {32'h3c6a88db, 32'h3d01513a} /* (18, 19, 12) {real, imag} */,
  {32'hbde8a810, 32'hbde9cae3} /* (18, 19, 11) {real, imag} */,
  {32'hbd8dd71e, 32'h3d9d759c} /* (18, 19, 10) {real, imag} */,
  {32'hbc2dc722, 32'hbd8058e3} /* (18, 19, 9) {real, imag} */,
  {32'hbbee6214, 32'hbd5e2d44} /* (18, 19, 8) {real, imag} */,
  {32'h3d3c0cb7, 32'h3ce7ae12} /* (18, 19, 7) {real, imag} */,
  {32'hbe3a8ea1, 32'hbdcd0b53} /* (18, 19, 6) {real, imag} */,
  {32'hbe00d0ec, 32'hbe068c87} /* (18, 19, 5) {real, imag} */,
  {32'h3ebb2050, 32'h3d877edf} /* (18, 19, 4) {real, imag} */,
  {32'hbcd09e60, 32'hbd802130} /* (18, 19, 3) {real, imag} */,
  {32'hbf4dfd48, 32'hbe8b66fa} /* (18, 19, 2) {real, imag} */,
  {32'h3ffc919e, 32'h3df6050c} /* (18, 19, 1) {real, imag} */,
  {32'h3f9a844a, 32'h00000000} /* (18, 19, 0) {real, imag} */,
  {32'h402e6a4d, 32'hbe8f5a98} /* (18, 18, 31) {real, imag} */,
  {32'hbf87dfd6, 32'h3e2dd2f3} /* (18, 18, 30) {real, imag} */,
  {32'h3db50537, 32'hbdcf8424} /* (18, 18, 29) {real, imag} */,
  {32'h3eca0803, 32'hbe0509be} /* (18, 18, 28) {real, imag} */,
  {32'hbe1b5b90, 32'h3ddbfb1a} /* (18, 18, 27) {real, imag} */,
  {32'hbdf47c71, 32'hbd16e156} /* (18, 18, 26) {real, imag} */,
  {32'h3c9a3ea2, 32'hbcf342dc} /* (18, 18, 25) {real, imag} */,
  {32'hbbb2959c, 32'h3d04c33a} /* (18, 18, 24) {real, imag} */,
  {32'hbc836308, 32'h3d8a8e98} /* (18, 18, 23) {real, imag} */,
  {32'hbd7b2d4d, 32'h3cf7aa85} /* (18, 18, 22) {real, imag} */,
  {32'hbd791703, 32'h3d2c0e68} /* (18, 18, 21) {real, imag} */,
  {32'hbce5d630, 32'h3db56018} /* (18, 18, 20) {real, imag} */,
  {32'hbd2cb096, 32'h3cd60f65} /* (18, 18, 19) {real, imag} */,
  {32'h3c5c5cf6, 32'h3c7dcf95} /* (18, 18, 18) {real, imag} */,
  {32'hbb2a7ce0, 32'h3cf4edd8} /* (18, 18, 17) {real, imag} */,
  {32'hbd27c0ff, 32'h00000000} /* (18, 18, 16) {real, imag} */,
  {32'hbb2a7ce0, 32'hbcf4edd8} /* (18, 18, 15) {real, imag} */,
  {32'h3c5c5cf6, 32'hbc7dcf95} /* (18, 18, 14) {real, imag} */,
  {32'hbd2cb096, 32'hbcd60f65} /* (18, 18, 13) {real, imag} */,
  {32'hbce5d630, 32'hbdb56018} /* (18, 18, 12) {real, imag} */,
  {32'hbd791703, 32'hbd2c0e68} /* (18, 18, 11) {real, imag} */,
  {32'hbd7b2d4d, 32'hbcf7aa85} /* (18, 18, 10) {real, imag} */,
  {32'hbc836308, 32'hbd8a8e98} /* (18, 18, 9) {real, imag} */,
  {32'hbbb2959c, 32'hbd04c33a} /* (18, 18, 8) {real, imag} */,
  {32'h3c9a3ea2, 32'h3cf342dc} /* (18, 18, 7) {real, imag} */,
  {32'hbdf47c71, 32'h3d16e156} /* (18, 18, 6) {real, imag} */,
  {32'hbe1b5b90, 32'hbddbfb1a} /* (18, 18, 5) {real, imag} */,
  {32'h3eca0803, 32'h3e0509be} /* (18, 18, 4) {real, imag} */,
  {32'h3db50537, 32'h3dcf8424} /* (18, 18, 3) {real, imag} */,
  {32'hbf87dfd6, 32'hbe2dd2f3} /* (18, 18, 2) {real, imag} */,
  {32'h402e6a4d, 32'h3e8f5a98} /* (18, 18, 1) {real, imag} */,
  {32'h3fe3b4de, 32'h00000000} /* (18, 18, 0) {real, imag} */,
  {32'h4048b463, 32'hbe8bc34d} /* (18, 17, 31) {real, imag} */,
  {32'hbf98d860, 32'h3e2f7f82} /* (18, 17, 30) {real, imag} */,
  {32'h3dae050f, 32'hbddda6ae} /* (18, 17, 29) {real, imag} */,
  {32'h3eaafa66, 32'hbd3a063a} /* (18, 17, 28) {real, imag} */,
  {32'hbe853773, 32'h3e021b1c} /* (18, 17, 27) {real, imag} */,
  {32'hbd5b0054, 32'hbc35642c} /* (18, 17, 26) {real, imag} */,
  {32'h3e0e2973, 32'hbcc0862f} /* (18, 17, 25) {real, imag} */,
  {32'hbdcd9d11, 32'h3bd3b11e} /* (18, 17, 24) {real, imag} */,
  {32'hbcd42e23, 32'hbdbd635a} /* (18, 17, 23) {real, imag} */,
  {32'h3d20905b, 32'hbcc821a0} /* (18, 17, 22) {real, imag} */,
  {32'hbae5a188, 32'h3d37202e} /* (18, 17, 21) {real, imag} */,
  {32'h3ce1054f, 32'hbc337489} /* (18, 17, 20) {real, imag} */,
  {32'hbd0e639e, 32'h3d95bad9} /* (18, 17, 19) {real, imag} */,
  {32'h3da1547d, 32'hbd134890} /* (18, 17, 18) {real, imag} */,
  {32'h3d68300d, 32'hbcdf0b3c} /* (18, 17, 17) {real, imag} */,
  {32'hbbb56fe3, 32'h00000000} /* (18, 17, 16) {real, imag} */,
  {32'h3d68300d, 32'h3cdf0b3c} /* (18, 17, 15) {real, imag} */,
  {32'h3da1547d, 32'h3d134890} /* (18, 17, 14) {real, imag} */,
  {32'hbd0e639e, 32'hbd95bad9} /* (18, 17, 13) {real, imag} */,
  {32'h3ce1054f, 32'h3c337489} /* (18, 17, 12) {real, imag} */,
  {32'hbae5a188, 32'hbd37202e} /* (18, 17, 11) {real, imag} */,
  {32'h3d20905b, 32'h3cc821a0} /* (18, 17, 10) {real, imag} */,
  {32'hbcd42e23, 32'h3dbd635a} /* (18, 17, 9) {real, imag} */,
  {32'hbdcd9d11, 32'hbbd3b11e} /* (18, 17, 8) {real, imag} */,
  {32'h3e0e2973, 32'h3cc0862f} /* (18, 17, 7) {real, imag} */,
  {32'hbd5b0054, 32'h3c35642c} /* (18, 17, 6) {real, imag} */,
  {32'hbe853773, 32'hbe021b1c} /* (18, 17, 5) {real, imag} */,
  {32'h3eaafa66, 32'h3d3a063a} /* (18, 17, 4) {real, imag} */,
  {32'h3dae050f, 32'h3ddda6ae} /* (18, 17, 3) {real, imag} */,
  {32'hbf98d860, 32'hbe2f7f82} /* (18, 17, 2) {real, imag} */,
  {32'h4048b463, 32'h3e8bc34d} /* (18, 17, 1) {real, imag} */,
  {32'h40089bae, 32'h00000000} /* (18, 17, 0) {real, imag} */,
  {32'h405761b8, 32'hbe8511e0} /* (18, 16, 31) {real, imag} */,
  {32'hbfbcb132, 32'h3d6aac00} /* (18, 16, 30) {real, imag} */,
  {32'h3dc402fe, 32'hbd984ce6} /* (18, 16, 29) {real, imag} */,
  {32'h3ea1f033, 32'h3d03b72e} /* (18, 16, 28) {real, imag} */,
  {32'hbea58dd0, 32'h3e0d5af1} /* (18, 16, 27) {real, imag} */,
  {32'hbd7ac634, 32'h3d40802f} /* (18, 16, 26) {real, imag} */,
  {32'h3d6adc82, 32'hbd32a59a} /* (18, 16, 25) {real, imag} */,
  {32'hbddb7e2e, 32'h3dcd7c1c} /* (18, 16, 24) {real, imag} */,
  {32'hbc825a6e, 32'h3d3aa93e} /* (18, 16, 23) {real, imag} */,
  {32'hbd9aadd2, 32'h3dae2cdb} /* (18, 16, 22) {real, imag} */,
  {32'hb9cf9e20, 32'h3d8d3f80} /* (18, 16, 21) {real, imag} */,
  {32'h3e1a4785, 32'hbcdfe39f} /* (18, 16, 20) {real, imag} */,
  {32'hbd7dae2a, 32'h3a3c1c70} /* (18, 16, 19) {real, imag} */,
  {32'hbd267a0f, 32'h3cc07c14} /* (18, 16, 18) {real, imag} */,
  {32'h3c968668, 32'hbcc94128} /* (18, 16, 17) {real, imag} */,
  {32'hbdf19f17, 32'h00000000} /* (18, 16, 16) {real, imag} */,
  {32'h3c968668, 32'h3cc94128} /* (18, 16, 15) {real, imag} */,
  {32'hbd267a0f, 32'hbcc07c14} /* (18, 16, 14) {real, imag} */,
  {32'hbd7dae2a, 32'hba3c1c70} /* (18, 16, 13) {real, imag} */,
  {32'h3e1a4785, 32'h3cdfe39f} /* (18, 16, 12) {real, imag} */,
  {32'hb9cf9e20, 32'hbd8d3f80} /* (18, 16, 11) {real, imag} */,
  {32'hbd9aadd2, 32'hbdae2cdb} /* (18, 16, 10) {real, imag} */,
  {32'hbc825a6e, 32'hbd3aa93e} /* (18, 16, 9) {real, imag} */,
  {32'hbddb7e2e, 32'hbdcd7c1c} /* (18, 16, 8) {real, imag} */,
  {32'h3d6adc82, 32'h3d32a59a} /* (18, 16, 7) {real, imag} */,
  {32'hbd7ac634, 32'hbd40802f} /* (18, 16, 6) {real, imag} */,
  {32'hbea58dd0, 32'hbe0d5af1} /* (18, 16, 5) {real, imag} */,
  {32'h3ea1f033, 32'hbd03b72e} /* (18, 16, 4) {real, imag} */,
  {32'h3dc402fe, 32'h3d984ce6} /* (18, 16, 3) {real, imag} */,
  {32'hbfbcb132, 32'hbd6aac00} /* (18, 16, 2) {real, imag} */,
  {32'h405761b8, 32'h3e8511e0} /* (18, 16, 1) {real, imag} */,
  {32'h401d93aa, 32'h00000000} /* (18, 16, 0) {real, imag} */,
  {32'h40566965, 32'hbe9feacb} /* (18, 15, 31) {real, imag} */,
  {32'hbfbe4800, 32'h3e9c3d48} /* (18, 15, 30) {real, imag} */,
  {32'h3de8710d, 32'hbdd4929e} /* (18, 15, 29) {real, imag} */,
  {32'h3e5294cb, 32'hbc7bdf18} /* (18, 15, 28) {real, imag} */,
  {32'hbe2d9c58, 32'h3e8727c7} /* (18, 15, 27) {real, imag} */,
  {32'h3c707340, 32'hbbf7e130} /* (18, 15, 26) {real, imag} */,
  {32'h3c163130, 32'hbd38cd66} /* (18, 15, 25) {real, imag} */,
  {32'h3d2b99c2, 32'h3d19038c} /* (18, 15, 24) {real, imag} */,
  {32'h3dabe40d, 32'h3d09668c} /* (18, 15, 23) {real, imag} */,
  {32'h3d63f605, 32'h3e0d970c} /* (18, 15, 22) {real, imag} */,
  {32'hbc7531bf, 32'h3e361964} /* (18, 15, 21) {real, imag} */,
  {32'h3ccbf2cf, 32'h3b6b6f74} /* (18, 15, 20) {real, imag} */,
  {32'h3ca27e83, 32'hbc88ad5f} /* (18, 15, 19) {real, imag} */,
  {32'hbd51063e, 32'h3d0c8c62} /* (18, 15, 18) {real, imag} */,
  {32'hbcea7fc6, 32'h3d6ddf2a} /* (18, 15, 17) {real, imag} */,
  {32'h3c0b6784, 32'h00000000} /* (18, 15, 16) {real, imag} */,
  {32'hbcea7fc6, 32'hbd6ddf2a} /* (18, 15, 15) {real, imag} */,
  {32'hbd51063e, 32'hbd0c8c62} /* (18, 15, 14) {real, imag} */,
  {32'h3ca27e83, 32'h3c88ad5f} /* (18, 15, 13) {real, imag} */,
  {32'h3ccbf2cf, 32'hbb6b6f74} /* (18, 15, 12) {real, imag} */,
  {32'hbc7531bf, 32'hbe361964} /* (18, 15, 11) {real, imag} */,
  {32'h3d63f605, 32'hbe0d970c} /* (18, 15, 10) {real, imag} */,
  {32'h3dabe40d, 32'hbd09668c} /* (18, 15, 9) {real, imag} */,
  {32'h3d2b99c2, 32'hbd19038c} /* (18, 15, 8) {real, imag} */,
  {32'h3c163130, 32'h3d38cd66} /* (18, 15, 7) {real, imag} */,
  {32'h3c707340, 32'h3bf7e130} /* (18, 15, 6) {real, imag} */,
  {32'hbe2d9c58, 32'hbe8727c7} /* (18, 15, 5) {real, imag} */,
  {32'h3e5294cb, 32'h3c7bdf18} /* (18, 15, 4) {real, imag} */,
  {32'h3de8710d, 32'h3dd4929e} /* (18, 15, 3) {real, imag} */,
  {32'hbfbe4800, 32'hbe9c3d48} /* (18, 15, 2) {real, imag} */,
  {32'h40566965, 32'h3e9feacb} /* (18, 15, 1) {real, imag} */,
  {32'h4019da1a, 32'h00000000} /* (18, 15, 0) {real, imag} */,
  {32'h4040d2a7, 32'hbe387150} /* (18, 14, 31) {real, imag} */,
  {32'hbfaf9f82, 32'h3eacfa1e} /* (18, 14, 30) {real, imag} */,
  {32'h3e7d7a1a, 32'hbdf7a7fc} /* (18, 14, 29) {real, imag} */,
  {32'h3e55f65a, 32'hbbc27130} /* (18, 14, 28) {real, imag} */,
  {32'hbe7b85e8, 32'h3e77059b} /* (18, 14, 27) {real, imag} */,
  {32'h3dfc1d5f, 32'h3d5748c2} /* (18, 14, 26) {real, imag} */,
  {32'hbd99a45e, 32'hbd99dc36} /* (18, 14, 25) {real, imag} */,
  {32'hbcf88eed, 32'h3ddf7633} /* (18, 14, 24) {real, imag} */,
  {32'hbd554c60, 32'h3d929298} /* (18, 14, 23) {real, imag} */,
  {32'h3d8379b1, 32'hbdaa8153} /* (18, 14, 22) {real, imag} */,
  {32'hbd01040f, 32'h3d146ed4} /* (18, 14, 21) {real, imag} */,
  {32'hbc44ec8d, 32'hbc1386a4} /* (18, 14, 20) {real, imag} */,
  {32'hbb7cf308, 32'hbd8b4bac} /* (18, 14, 19) {real, imag} */,
  {32'hbd8519d7, 32'h3c4287ed} /* (18, 14, 18) {real, imag} */,
  {32'h3d166d2c, 32'hbaae01d8} /* (18, 14, 17) {real, imag} */,
  {32'h3caadbda, 32'h00000000} /* (18, 14, 16) {real, imag} */,
  {32'h3d166d2c, 32'h3aae01d8} /* (18, 14, 15) {real, imag} */,
  {32'hbd8519d7, 32'hbc4287ed} /* (18, 14, 14) {real, imag} */,
  {32'hbb7cf308, 32'h3d8b4bac} /* (18, 14, 13) {real, imag} */,
  {32'hbc44ec8d, 32'h3c1386a4} /* (18, 14, 12) {real, imag} */,
  {32'hbd01040f, 32'hbd146ed4} /* (18, 14, 11) {real, imag} */,
  {32'h3d8379b1, 32'h3daa8153} /* (18, 14, 10) {real, imag} */,
  {32'hbd554c60, 32'hbd929298} /* (18, 14, 9) {real, imag} */,
  {32'hbcf88eed, 32'hbddf7633} /* (18, 14, 8) {real, imag} */,
  {32'hbd99a45e, 32'h3d99dc36} /* (18, 14, 7) {real, imag} */,
  {32'h3dfc1d5f, 32'hbd5748c2} /* (18, 14, 6) {real, imag} */,
  {32'hbe7b85e8, 32'hbe77059b} /* (18, 14, 5) {real, imag} */,
  {32'h3e55f65a, 32'h3bc27130} /* (18, 14, 4) {real, imag} */,
  {32'h3e7d7a1a, 32'h3df7a7fc} /* (18, 14, 3) {real, imag} */,
  {32'hbfaf9f82, 32'hbeacfa1e} /* (18, 14, 2) {real, imag} */,
  {32'h4040d2a7, 32'h3e387150} /* (18, 14, 1) {real, imag} */,
  {32'h400f9b89, 32'h00000000} /* (18, 14, 0) {real, imag} */,
  {32'h40256e97, 32'h3d5ea118} /* (18, 13, 31) {real, imag} */,
  {32'hbf991ee8, 32'h3e76802b} /* (18, 13, 30) {real, imag} */,
  {32'h3e440f78, 32'hbda78f4a} /* (18, 13, 29) {real, imag} */,
  {32'h3db5b066, 32'h3d1a4816} /* (18, 13, 28) {real, imag} */,
  {32'hbe411b8e, 32'h3d8e1cea} /* (18, 13, 27) {real, imag} */,
  {32'h3c5928c0, 32'h3dde7317} /* (18, 13, 26) {real, imag} */,
  {32'hbd29a48b, 32'hbc124d3c} /* (18, 13, 25) {real, imag} */,
  {32'hbd87278f, 32'h3d1224d2} /* (18, 13, 24) {real, imag} */,
  {32'h3d63dfc6, 32'h3d627fcf} /* (18, 13, 23) {real, imag} */,
  {32'hbcf96de0, 32'hbd9215e0} /* (18, 13, 22) {real, imag} */,
  {32'h3b63aac0, 32'h3d4d838a} /* (18, 13, 21) {real, imag} */,
  {32'h3d0c5783, 32'hbd5519fa} /* (18, 13, 20) {real, imag} */,
  {32'h3ca95377, 32'h3dfe9551} /* (18, 13, 19) {real, imag} */,
  {32'hbc597d1b, 32'h3d2937a4} /* (18, 13, 18) {real, imag} */,
  {32'h3c5ac886, 32'h3d6da5cb} /* (18, 13, 17) {real, imag} */,
  {32'hbd730c2e, 32'h00000000} /* (18, 13, 16) {real, imag} */,
  {32'h3c5ac886, 32'hbd6da5cb} /* (18, 13, 15) {real, imag} */,
  {32'hbc597d1b, 32'hbd2937a4} /* (18, 13, 14) {real, imag} */,
  {32'h3ca95377, 32'hbdfe9551} /* (18, 13, 13) {real, imag} */,
  {32'h3d0c5783, 32'h3d5519fa} /* (18, 13, 12) {real, imag} */,
  {32'h3b63aac0, 32'hbd4d838a} /* (18, 13, 11) {real, imag} */,
  {32'hbcf96de0, 32'h3d9215e0} /* (18, 13, 10) {real, imag} */,
  {32'h3d63dfc6, 32'hbd627fcf} /* (18, 13, 9) {real, imag} */,
  {32'hbd87278f, 32'hbd1224d2} /* (18, 13, 8) {real, imag} */,
  {32'hbd29a48b, 32'h3c124d3c} /* (18, 13, 7) {real, imag} */,
  {32'h3c5928c0, 32'hbdde7317} /* (18, 13, 6) {real, imag} */,
  {32'hbe411b8e, 32'hbd8e1cea} /* (18, 13, 5) {real, imag} */,
  {32'h3db5b066, 32'hbd1a4816} /* (18, 13, 4) {real, imag} */,
  {32'h3e440f78, 32'h3da78f4a} /* (18, 13, 3) {real, imag} */,
  {32'hbf991ee8, 32'hbe76802b} /* (18, 13, 2) {real, imag} */,
  {32'h40256e97, 32'hbd5ea118} /* (18, 13, 1) {real, imag} */,
  {32'h3ff5599e, 32'h00000000} /* (18, 13, 0) {real, imag} */,
  {32'h3ff77e12, 32'h3e385a4c} /* (18, 12, 31) {real, imag} */,
  {32'hbf7d76f5, 32'h3e91d79e} /* (18, 12, 30) {real, imag} */,
  {32'h3dc5c33c, 32'hbe1a8b8a} /* (18, 12, 29) {real, imag} */,
  {32'h3da1226a, 32'hbda4750a} /* (18, 12, 28) {real, imag} */,
  {32'hbde2c7ce, 32'h3e05a52a} /* (18, 12, 27) {real, imag} */,
  {32'h3d837200, 32'h3d266d3b} /* (18, 12, 26) {real, imag} */,
  {32'h3d120098, 32'hbdb1256e} /* (18, 12, 25) {real, imag} */,
  {32'hbd103c59, 32'h3be1e4e0} /* (18, 12, 24) {real, imag} */,
  {32'h3d8b5f4d, 32'hbcf3a34b} /* (18, 12, 23) {real, imag} */,
  {32'h3d1ef0c0, 32'h3cff966d} /* (18, 12, 22) {real, imag} */,
  {32'h3d8327f6, 32'h3d898033} /* (18, 12, 21) {real, imag} */,
  {32'hbd211bca, 32'hbccdfedd} /* (18, 12, 20) {real, imag} */,
  {32'h3d8ea538, 32'h3d940567} /* (18, 12, 19) {real, imag} */,
  {32'h3d039707, 32'h3d59efe7} /* (18, 12, 18) {real, imag} */,
  {32'hbd81aa56, 32'h3ca7f0de} /* (18, 12, 17) {real, imag} */,
  {32'hbc63f928, 32'h00000000} /* (18, 12, 16) {real, imag} */,
  {32'hbd81aa56, 32'hbca7f0de} /* (18, 12, 15) {real, imag} */,
  {32'h3d039707, 32'hbd59efe7} /* (18, 12, 14) {real, imag} */,
  {32'h3d8ea538, 32'hbd940567} /* (18, 12, 13) {real, imag} */,
  {32'hbd211bca, 32'h3ccdfedd} /* (18, 12, 12) {real, imag} */,
  {32'h3d8327f6, 32'hbd898033} /* (18, 12, 11) {real, imag} */,
  {32'h3d1ef0c0, 32'hbcff966d} /* (18, 12, 10) {real, imag} */,
  {32'h3d8b5f4d, 32'h3cf3a34b} /* (18, 12, 9) {real, imag} */,
  {32'hbd103c59, 32'hbbe1e4e0} /* (18, 12, 8) {real, imag} */,
  {32'h3d120098, 32'h3db1256e} /* (18, 12, 7) {real, imag} */,
  {32'h3d837200, 32'hbd266d3b} /* (18, 12, 6) {real, imag} */,
  {32'hbde2c7ce, 32'hbe05a52a} /* (18, 12, 5) {real, imag} */,
  {32'h3da1226a, 32'h3da4750a} /* (18, 12, 4) {real, imag} */,
  {32'h3dc5c33c, 32'h3e1a8b8a} /* (18, 12, 3) {real, imag} */,
  {32'hbf7d76f5, 32'hbe91d79e} /* (18, 12, 2) {real, imag} */,
  {32'h3ff77e12, 32'hbe385a4c} /* (18, 12, 1) {real, imag} */,
  {32'h3fac2308, 32'h00000000} /* (18, 12, 0) {real, imag} */,
  {32'h3f6120db, 32'h3ec4f407} /* (18, 11, 31) {real, imag} */,
  {32'hbf135d16, 32'h3e47c4e2} /* (18, 11, 30) {real, imag} */,
  {32'h3e17cfff, 32'hbcd0965f} /* (18, 11, 29) {real, imag} */,
  {32'h3dabfaaa, 32'hbd52e246} /* (18, 11, 28) {real, imag} */,
  {32'hbe0d0edb, 32'h3cb24b18} /* (18, 11, 27) {real, imag} */,
  {32'h3db7ddab, 32'h3dfdce14} /* (18, 11, 26) {real, imag} */,
  {32'hbd7c9a28, 32'h3cdd6262} /* (18, 11, 25) {real, imag} */,
  {32'hbd7e98f6, 32'h3d1a9f24} /* (18, 11, 24) {real, imag} */,
  {32'hbd0b0362, 32'h3d65a01c} /* (18, 11, 23) {real, imag} */,
  {32'h3bc02ee8, 32'hbdc79151} /* (18, 11, 22) {real, imag} */,
  {32'hbde4eb10, 32'h3ddf1691} /* (18, 11, 21) {real, imag} */,
  {32'hbdf02620, 32'hbd63fde0} /* (18, 11, 20) {real, imag} */,
  {32'h3b8026b4, 32'h3c693451} /* (18, 11, 19) {real, imag} */,
  {32'hbcaae252, 32'h3d381d50} /* (18, 11, 18) {real, imag} */,
  {32'h3d3596ee, 32'hbd2e0766} /* (18, 11, 17) {real, imag} */,
  {32'h3cdcd068, 32'h00000000} /* (18, 11, 16) {real, imag} */,
  {32'h3d3596ee, 32'h3d2e0766} /* (18, 11, 15) {real, imag} */,
  {32'hbcaae252, 32'hbd381d50} /* (18, 11, 14) {real, imag} */,
  {32'h3b8026b4, 32'hbc693451} /* (18, 11, 13) {real, imag} */,
  {32'hbdf02620, 32'h3d63fde0} /* (18, 11, 12) {real, imag} */,
  {32'hbde4eb10, 32'hbddf1691} /* (18, 11, 11) {real, imag} */,
  {32'h3bc02ee8, 32'h3dc79151} /* (18, 11, 10) {real, imag} */,
  {32'hbd0b0362, 32'hbd65a01c} /* (18, 11, 9) {real, imag} */,
  {32'hbd7e98f6, 32'hbd1a9f24} /* (18, 11, 8) {real, imag} */,
  {32'hbd7c9a28, 32'hbcdd6262} /* (18, 11, 7) {real, imag} */,
  {32'h3db7ddab, 32'hbdfdce14} /* (18, 11, 6) {real, imag} */,
  {32'hbe0d0edb, 32'hbcb24b18} /* (18, 11, 5) {real, imag} */,
  {32'h3dabfaaa, 32'h3d52e246} /* (18, 11, 4) {real, imag} */,
  {32'h3e17cfff, 32'h3cd0965f} /* (18, 11, 3) {real, imag} */,
  {32'hbf135d16, 32'hbe47c4e2} /* (18, 11, 2) {real, imag} */,
  {32'h3f6120db, 32'hbec4f407} /* (18, 11, 1) {real, imag} */,
  {32'h3f290298, 32'h00000000} /* (18, 11, 0) {real, imag} */,
  {32'hbf46a058, 32'h3f27788e} /* (18, 10, 31) {real, imag} */,
  {32'h3eaa34ba, 32'hbdf113d8} /* (18, 10, 30) {real, imag} */,
  {32'h3d9723d1, 32'h3dcf8aec} /* (18, 10, 29) {real, imag} */,
  {32'hbdcdebe5, 32'hbc23efb0} /* (18, 10, 28) {real, imag} */,
  {32'h3d0b4872, 32'hbbde1470} /* (18, 10, 27) {real, imag} */,
  {32'hbd541c02, 32'h3d7d1c57} /* (18, 10, 26) {real, imag} */,
  {32'hbe1965f3, 32'hbce747ce} /* (18, 10, 25) {real, imag} */,
  {32'hbc864e39, 32'hbbce6aa8} /* (18, 10, 24) {real, imag} */,
  {32'h3b6b8356, 32'hbc358dec} /* (18, 10, 23) {real, imag} */,
  {32'hbd1a2cd8, 32'hbdc18e86} /* (18, 10, 22) {real, imag} */,
  {32'h3ca1576b, 32'hbe0b3cc6} /* (18, 10, 21) {real, imag} */,
  {32'h3d8bcd86, 32'hbc66a75a} /* (18, 10, 20) {real, imag} */,
  {32'hbce60a98, 32'h3cf2d480} /* (18, 10, 19) {real, imag} */,
  {32'hbd05254b, 32'hbd4ec51a} /* (18, 10, 18) {real, imag} */,
  {32'h3d88b779, 32'h3d4eb675} /* (18, 10, 17) {real, imag} */,
  {32'hb9e51380, 32'h00000000} /* (18, 10, 16) {real, imag} */,
  {32'h3d88b779, 32'hbd4eb675} /* (18, 10, 15) {real, imag} */,
  {32'hbd05254b, 32'h3d4ec51a} /* (18, 10, 14) {real, imag} */,
  {32'hbce60a98, 32'hbcf2d480} /* (18, 10, 13) {real, imag} */,
  {32'h3d8bcd86, 32'h3c66a75a} /* (18, 10, 12) {real, imag} */,
  {32'h3ca1576b, 32'h3e0b3cc6} /* (18, 10, 11) {real, imag} */,
  {32'hbd1a2cd8, 32'h3dc18e86} /* (18, 10, 10) {real, imag} */,
  {32'h3b6b8356, 32'h3c358dec} /* (18, 10, 9) {real, imag} */,
  {32'hbc864e39, 32'h3bce6aa8} /* (18, 10, 8) {real, imag} */,
  {32'hbe1965f3, 32'h3ce747ce} /* (18, 10, 7) {real, imag} */,
  {32'hbd541c02, 32'hbd7d1c57} /* (18, 10, 6) {real, imag} */,
  {32'h3d0b4872, 32'h3bde1470} /* (18, 10, 5) {real, imag} */,
  {32'hbdcdebe5, 32'h3c23efb0} /* (18, 10, 4) {real, imag} */,
  {32'h3d9723d1, 32'hbdcf8aec} /* (18, 10, 3) {real, imag} */,
  {32'h3eaa34ba, 32'h3df113d8} /* (18, 10, 2) {real, imag} */,
  {32'hbf46a058, 32'hbf27788e} /* (18, 10, 1) {real, imag} */,
  {32'hbf38ba0c, 32'h00000000} /* (18, 10, 0) {real, imag} */,
  {32'hc0048248, 32'h3f515b04} /* (18, 9, 31) {real, imag} */,
  {32'h3f5b67bd, 32'hbe688f44} /* (18, 9, 30) {real, imag} */,
  {32'hbd31b0bc, 32'h3d19e864} /* (18, 9, 29) {real, imag} */,
  {32'hbd715b12, 32'hbd095474} /* (18, 9, 28) {real, imag} */,
  {32'h3d7bacc4, 32'hbd898f10} /* (18, 9, 27) {real, imag} */,
  {32'h3ca57740, 32'h3dce3b0f} /* (18, 9, 26) {real, imag} */,
  {32'hbdbd818e, 32'hbd47d117} /* (18, 9, 25) {real, imag} */,
  {32'hbdb41698, 32'hbe2063cc} /* (18, 9, 24) {real, imag} */,
  {32'h3cf4591c, 32'hbd8229f8} /* (18, 9, 23) {real, imag} */,
  {32'h3ba22a78, 32'hbd5073f8} /* (18, 9, 22) {real, imag} */,
  {32'h3da0433a, 32'hbde62e66} /* (18, 9, 21) {real, imag} */,
  {32'h3c8d2fde, 32'hbda5c062} /* (18, 9, 20) {real, imag} */,
  {32'hbc8abaf0, 32'h3d7ad498} /* (18, 9, 19) {real, imag} */,
  {32'h3cd4aeb3, 32'hbcde13b5} /* (18, 9, 18) {real, imag} */,
  {32'hbd35f8a1, 32'hbcaa9d9c} /* (18, 9, 17) {real, imag} */,
  {32'hbd753a6a, 32'h00000000} /* (18, 9, 16) {real, imag} */,
  {32'hbd35f8a1, 32'h3caa9d9c} /* (18, 9, 15) {real, imag} */,
  {32'h3cd4aeb3, 32'h3cde13b5} /* (18, 9, 14) {real, imag} */,
  {32'hbc8abaf0, 32'hbd7ad498} /* (18, 9, 13) {real, imag} */,
  {32'h3c8d2fde, 32'h3da5c062} /* (18, 9, 12) {real, imag} */,
  {32'h3da0433a, 32'h3de62e66} /* (18, 9, 11) {real, imag} */,
  {32'h3ba22a78, 32'h3d5073f8} /* (18, 9, 10) {real, imag} */,
  {32'h3cf4591c, 32'h3d8229f8} /* (18, 9, 9) {real, imag} */,
  {32'hbdb41698, 32'h3e2063cc} /* (18, 9, 8) {real, imag} */,
  {32'hbdbd818e, 32'h3d47d117} /* (18, 9, 7) {real, imag} */,
  {32'h3ca57740, 32'hbdce3b0f} /* (18, 9, 6) {real, imag} */,
  {32'h3d7bacc4, 32'h3d898f10} /* (18, 9, 5) {real, imag} */,
  {32'hbd715b12, 32'h3d095474} /* (18, 9, 4) {real, imag} */,
  {32'hbd31b0bc, 32'hbd19e864} /* (18, 9, 3) {real, imag} */,
  {32'h3f5b67bd, 32'h3e688f44} /* (18, 9, 2) {real, imag} */,
  {32'hc0048248, 32'hbf515b04} /* (18, 9, 1) {real, imag} */,
  {32'hbfe0f517, 32'h00000000} /* (18, 9, 0) {real, imag} */,
  {32'hc02d4c32, 32'h3f8c1332} /* (18, 8, 31) {real, imag} */,
  {32'h3f4ed6db, 32'hbe687928} /* (18, 8, 30) {real, imag} */,
  {32'h3cf48742, 32'h3dde3ac2} /* (18, 8, 29) {real, imag} */,
  {32'h3d2992a8, 32'h3c14f858} /* (18, 8, 28) {real, imag} */,
  {32'h3e17cce6, 32'hbdd9a173} /* (18, 8, 27) {real, imag} */,
  {32'h3ce8441a, 32'h3cad4ea2} /* (18, 8, 26) {real, imag} */,
  {32'hbda031d0, 32'h3a6ec3c0} /* (18, 8, 25) {real, imag} */,
  {32'h3ce9c905, 32'hbdc223ff} /* (18, 8, 24) {real, imag} */,
  {32'h3b81dca0, 32'h3c4bc873} /* (18, 8, 23) {real, imag} */,
  {32'hbda537d8, 32'h3ded2487} /* (18, 8, 22) {real, imag} */,
  {32'h3c057bc9, 32'h3d88935a} /* (18, 8, 21) {real, imag} */,
  {32'hbc767bd4, 32'hbbd4f8c8} /* (18, 8, 20) {real, imag} */,
  {32'hbd2a112c, 32'hbbbbc6e0} /* (18, 8, 19) {real, imag} */,
  {32'hbd1d98e0, 32'hbd129e87} /* (18, 8, 18) {real, imag} */,
  {32'hbda621b2, 32'h3bc09366} /* (18, 8, 17) {real, imag} */,
  {32'hbcf5ffd1, 32'h00000000} /* (18, 8, 16) {real, imag} */,
  {32'hbda621b2, 32'hbbc09366} /* (18, 8, 15) {real, imag} */,
  {32'hbd1d98e0, 32'h3d129e87} /* (18, 8, 14) {real, imag} */,
  {32'hbd2a112c, 32'h3bbbc6e0} /* (18, 8, 13) {real, imag} */,
  {32'hbc767bd4, 32'h3bd4f8c8} /* (18, 8, 12) {real, imag} */,
  {32'h3c057bc9, 32'hbd88935a} /* (18, 8, 11) {real, imag} */,
  {32'hbda537d8, 32'hbded2487} /* (18, 8, 10) {real, imag} */,
  {32'h3b81dca0, 32'hbc4bc873} /* (18, 8, 9) {real, imag} */,
  {32'h3ce9c905, 32'h3dc223ff} /* (18, 8, 8) {real, imag} */,
  {32'hbda031d0, 32'hba6ec3c0} /* (18, 8, 7) {real, imag} */,
  {32'h3ce8441a, 32'hbcad4ea2} /* (18, 8, 6) {real, imag} */,
  {32'h3e17cce6, 32'h3dd9a173} /* (18, 8, 5) {real, imag} */,
  {32'h3d2992a8, 32'hbc14f858} /* (18, 8, 4) {real, imag} */,
  {32'h3cf48742, 32'hbdde3ac2} /* (18, 8, 3) {real, imag} */,
  {32'h3f4ed6db, 32'h3e687928} /* (18, 8, 2) {real, imag} */,
  {32'hc02d4c32, 32'hbf8c1332} /* (18, 8, 1) {real, imag} */,
  {32'hc01d1008, 32'h00000000} /* (18, 8, 0) {real, imag} */,
  {32'hc0404dca, 32'h3fb85ac2} /* (18, 7, 31) {real, imag} */,
  {32'h3f7bf831, 32'hbebb8560} /* (18, 7, 30) {real, imag} */,
  {32'hbcd7bd22, 32'h3c5377f4} /* (18, 7, 29) {real, imag} */,
  {32'hbdf96e40, 32'h3da873da} /* (18, 7, 28) {real, imag} */,
  {32'h3cc94628, 32'hbde6903c} /* (18, 7, 27) {real, imag} */,
  {32'hbcf6a238, 32'h3e024004} /* (18, 7, 26) {real, imag} */,
  {32'hbd2548d0, 32'hbcfc75ec} /* (18, 7, 25) {real, imag} */,
  {32'h3d22f349, 32'hbe89482b} /* (18, 7, 24) {real, imag} */,
  {32'h3c8a9529, 32'h3dbdc151} /* (18, 7, 23) {real, imag} */,
  {32'hbcd0a056, 32'h3d070a78} /* (18, 7, 22) {real, imag} */,
  {32'h3d83c6ae, 32'hbd4a9d5a} /* (18, 7, 21) {real, imag} */,
  {32'hbc5fcd0c, 32'hbd6eb741} /* (18, 7, 20) {real, imag} */,
  {32'h3d7fdad7, 32'hbc771958} /* (18, 7, 19) {real, imag} */,
  {32'hbb385620, 32'hbdb83e99} /* (18, 7, 18) {real, imag} */,
  {32'h3cd79c35, 32'h3e048408} /* (18, 7, 17) {real, imag} */,
  {32'h3ce96406, 32'h00000000} /* (18, 7, 16) {real, imag} */,
  {32'h3cd79c35, 32'hbe048408} /* (18, 7, 15) {real, imag} */,
  {32'hbb385620, 32'h3db83e99} /* (18, 7, 14) {real, imag} */,
  {32'h3d7fdad7, 32'h3c771958} /* (18, 7, 13) {real, imag} */,
  {32'hbc5fcd0c, 32'h3d6eb741} /* (18, 7, 12) {real, imag} */,
  {32'h3d83c6ae, 32'h3d4a9d5a} /* (18, 7, 11) {real, imag} */,
  {32'hbcd0a056, 32'hbd070a78} /* (18, 7, 10) {real, imag} */,
  {32'h3c8a9529, 32'hbdbdc151} /* (18, 7, 9) {real, imag} */,
  {32'h3d22f349, 32'h3e89482b} /* (18, 7, 8) {real, imag} */,
  {32'hbd2548d0, 32'h3cfc75ec} /* (18, 7, 7) {real, imag} */,
  {32'hbcf6a238, 32'hbe024004} /* (18, 7, 6) {real, imag} */,
  {32'h3cc94628, 32'h3de6903c} /* (18, 7, 5) {real, imag} */,
  {32'hbdf96e40, 32'hbda873da} /* (18, 7, 4) {real, imag} */,
  {32'hbcd7bd22, 32'hbc5377f4} /* (18, 7, 3) {real, imag} */,
  {32'h3f7bf831, 32'h3ebb8560} /* (18, 7, 2) {real, imag} */,
  {32'hc0404dca, 32'hbfb85ac2} /* (18, 7, 1) {real, imag} */,
  {32'hc03b12ee, 32'h00000000} /* (18, 7, 0) {real, imag} */,
  {32'hc046c8a0, 32'h3feaece2} /* (18, 6, 31) {real, imag} */,
  {32'h3f36498a, 32'hbf33b64e} /* (18, 6, 30) {real, imag} */,
  {32'hbddce935, 32'hbe33bb16} /* (18, 6, 29) {real, imag} */,
  {32'hbd81e822, 32'h3d9ccd1d} /* (18, 6, 28) {real, imag} */,
  {32'h3e3fa193, 32'hbcd274da} /* (18, 6, 27) {real, imag} */,
  {32'h3d94aea1, 32'h3ddefaaa} /* (18, 6, 26) {real, imag} */,
  {32'h3e40601c, 32'h3d04190e} /* (18, 6, 25) {real, imag} */,
  {32'h3dcb0b56, 32'hbe1e402c} /* (18, 6, 24) {real, imag} */,
  {32'hbbbfed22, 32'hbc84956e} /* (18, 6, 23) {real, imag} */,
  {32'h3c27e574, 32'h3c210414} /* (18, 6, 22) {real, imag} */,
  {32'h3cb24219, 32'h3c840349} /* (18, 6, 21) {real, imag} */,
  {32'hbded4122, 32'h3d30e704} /* (18, 6, 20) {real, imag} */,
  {32'h3cc0e910, 32'hbd19b276} /* (18, 6, 19) {real, imag} */,
  {32'hbdc997a9, 32'h3c2a2be6} /* (18, 6, 18) {real, imag} */,
  {32'hbc17b894, 32'h3d16e531} /* (18, 6, 17) {real, imag} */,
  {32'hbb8221f8, 32'h00000000} /* (18, 6, 16) {real, imag} */,
  {32'hbc17b894, 32'hbd16e531} /* (18, 6, 15) {real, imag} */,
  {32'hbdc997a9, 32'hbc2a2be6} /* (18, 6, 14) {real, imag} */,
  {32'h3cc0e910, 32'h3d19b276} /* (18, 6, 13) {real, imag} */,
  {32'hbded4122, 32'hbd30e704} /* (18, 6, 12) {real, imag} */,
  {32'h3cb24219, 32'hbc840349} /* (18, 6, 11) {real, imag} */,
  {32'h3c27e574, 32'hbc210414} /* (18, 6, 10) {real, imag} */,
  {32'hbbbfed22, 32'h3c84956e} /* (18, 6, 9) {real, imag} */,
  {32'h3dcb0b56, 32'h3e1e402c} /* (18, 6, 8) {real, imag} */,
  {32'h3e40601c, 32'hbd04190e} /* (18, 6, 7) {real, imag} */,
  {32'h3d94aea1, 32'hbddefaaa} /* (18, 6, 6) {real, imag} */,
  {32'h3e3fa193, 32'h3cd274da} /* (18, 6, 5) {real, imag} */,
  {32'hbd81e822, 32'hbd9ccd1d} /* (18, 6, 4) {real, imag} */,
  {32'hbddce935, 32'h3e33bb16} /* (18, 6, 3) {real, imag} */,
  {32'h3f36498a, 32'h3f33b64e} /* (18, 6, 2) {real, imag} */,
  {32'hc046c8a0, 32'hbfeaece2} /* (18, 6, 1) {real, imag} */,
  {32'hc04c8518, 32'h00000000} /* (18, 6, 0) {real, imag} */,
  {32'hc02ee7e7, 32'h40173a92} /* (18, 5, 31) {real, imag} */,
  {32'h3e5086e8, 32'hbf595ada} /* (18, 5, 30) {real, imag} */,
  {32'hbb8e2df4, 32'hbd926023} /* (18, 5, 29) {real, imag} */,
  {32'h3d8a676c, 32'hbd40c7e2} /* (18, 5, 28) {real, imag} */,
  {32'h3e1fd6d2, 32'h3d1de413} /* (18, 5, 27) {real, imag} */,
  {32'h3e08d01c, 32'hbd3c0b7c} /* (18, 5, 26) {real, imag} */,
  {32'hbba80044, 32'hbce3cab4} /* (18, 5, 25) {real, imag} */,
  {32'h3d5b15ac, 32'h3cea8f4a} /* (18, 5, 24) {real, imag} */,
  {32'hbd09b546, 32'hbdd49ef2} /* (18, 5, 23) {real, imag} */,
  {32'hbdc2a4e2, 32'h3d80ca76} /* (18, 5, 22) {real, imag} */,
  {32'hbd48a00d, 32'h3dd43f08} /* (18, 5, 21) {real, imag} */,
  {32'h3d6f95a3, 32'hbdbbad7e} /* (18, 5, 20) {real, imag} */,
  {32'h3cb03361, 32'h3cbae7f8} /* (18, 5, 19) {real, imag} */,
  {32'h3abb8490, 32'h3d61cbc4} /* (18, 5, 18) {real, imag} */,
  {32'h3d30e7ec, 32'h3c3fa02e} /* (18, 5, 17) {real, imag} */,
  {32'h3c155fc5, 32'h00000000} /* (18, 5, 16) {real, imag} */,
  {32'h3d30e7ec, 32'hbc3fa02e} /* (18, 5, 15) {real, imag} */,
  {32'h3abb8490, 32'hbd61cbc4} /* (18, 5, 14) {real, imag} */,
  {32'h3cb03361, 32'hbcbae7f8} /* (18, 5, 13) {real, imag} */,
  {32'h3d6f95a3, 32'h3dbbad7e} /* (18, 5, 12) {real, imag} */,
  {32'hbd48a00d, 32'hbdd43f08} /* (18, 5, 11) {real, imag} */,
  {32'hbdc2a4e2, 32'hbd80ca76} /* (18, 5, 10) {real, imag} */,
  {32'hbd09b546, 32'h3dd49ef2} /* (18, 5, 9) {real, imag} */,
  {32'h3d5b15ac, 32'hbcea8f4a} /* (18, 5, 8) {real, imag} */,
  {32'hbba80044, 32'h3ce3cab4} /* (18, 5, 7) {real, imag} */,
  {32'h3e08d01c, 32'h3d3c0b7c} /* (18, 5, 6) {real, imag} */,
  {32'h3e1fd6d2, 32'hbd1de413} /* (18, 5, 5) {real, imag} */,
  {32'h3d8a676c, 32'h3d40c7e2} /* (18, 5, 4) {real, imag} */,
  {32'hbb8e2df4, 32'h3d926023} /* (18, 5, 3) {real, imag} */,
  {32'h3e5086e8, 32'h3f595ada} /* (18, 5, 2) {real, imag} */,
  {32'hc02ee7e7, 32'hc0173a92} /* (18, 5, 1) {real, imag} */,
  {32'hc060977a, 32'h00000000} /* (18, 5, 0) {real, imag} */,
  {32'hc01de71f, 32'h403533e8} /* (18, 4, 31) {real, imag} */,
  {32'hbe560e84, 32'hbf885a4d} /* (18, 4, 30) {real, imag} */,
  {32'h3d6dde58, 32'hbd14c1cc} /* (18, 4, 29) {real, imag} */,
  {32'h3e729189, 32'h3cee158e} /* (18, 4, 28) {real, imag} */,
  {32'h3e4b426d, 32'h3df4ebb6} /* (18, 4, 27) {real, imag} */,
  {32'h3e06917f, 32'h3c27a93e} /* (18, 4, 26) {real, imag} */,
  {32'hbd4b44f0, 32'h3d22ab2c} /* (18, 4, 25) {real, imag} */,
  {32'hbcb14fbd, 32'hbdb0cec7} /* (18, 4, 24) {real, imag} */,
  {32'hbc596700, 32'hbd977a38} /* (18, 4, 23) {real, imag} */,
  {32'hbbc0f968, 32'hbdbaee18} /* (18, 4, 22) {real, imag} */,
  {32'hbc930610, 32'h3c273c84} /* (18, 4, 21) {real, imag} */,
  {32'hbcd4da34, 32'hbca2df66} /* (18, 4, 20) {real, imag} */,
  {32'h3ceef610, 32'h3bbe0080} /* (18, 4, 19) {real, imag} */,
  {32'h3d80f372, 32'hbd9acf57} /* (18, 4, 18) {real, imag} */,
  {32'hbbd976cc, 32'h3d7040b6} /* (18, 4, 17) {real, imag} */,
  {32'h3d6765fb, 32'h00000000} /* (18, 4, 16) {real, imag} */,
  {32'hbbd976cc, 32'hbd7040b6} /* (18, 4, 15) {real, imag} */,
  {32'h3d80f372, 32'h3d9acf57} /* (18, 4, 14) {real, imag} */,
  {32'h3ceef610, 32'hbbbe0080} /* (18, 4, 13) {real, imag} */,
  {32'hbcd4da34, 32'h3ca2df66} /* (18, 4, 12) {real, imag} */,
  {32'hbc930610, 32'hbc273c84} /* (18, 4, 11) {real, imag} */,
  {32'hbbc0f968, 32'h3dbaee18} /* (18, 4, 10) {real, imag} */,
  {32'hbc596700, 32'h3d977a38} /* (18, 4, 9) {real, imag} */,
  {32'hbcb14fbd, 32'h3db0cec7} /* (18, 4, 8) {real, imag} */,
  {32'hbd4b44f0, 32'hbd22ab2c} /* (18, 4, 7) {real, imag} */,
  {32'h3e06917f, 32'hbc27a93e} /* (18, 4, 6) {real, imag} */,
  {32'h3e4b426d, 32'hbdf4ebb6} /* (18, 4, 5) {real, imag} */,
  {32'h3e729189, 32'hbcee158e} /* (18, 4, 4) {real, imag} */,
  {32'h3d6dde58, 32'h3d14c1cc} /* (18, 4, 3) {real, imag} */,
  {32'hbe560e84, 32'h3f885a4d} /* (18, 4, 2) {real, imag} */,
  {32'hc01de71f, 32'hc03533e8} /* (18, 4, 1) {real, imag} */,
  {32'hc067928d, 32'h00000000} /* (18, 4, 0) {real, imag} */,
  {32'hc017395a, 32'h403c9420} /* (18, 3, 31) {real, imag} */,
  {32'hbeb1b311, 32'hbf941cf2} /* (18, 3, 30) {real, imag} */,
  {32'h3cc9949c, 32'hbd2f5a0b} /* (18, 3, 29) {real, imag} */,
  {32'h3d852b4b, 32'hbe08bd40} /* (18, 3, 28) {real, imag} */,
  {32'h3e81621d, 32'h3de9697b} /* (18, 3, 27) {real, imag} */,
  {32'h3c92e878, 32'hbd3198bc} /* (18, 3, 26) {real, imag} */,
  {32'hbc42c1b0, 32'h3dc0416e} /* (18, 3, 25) {real, imag} */,
  {32'h3d74532c, 32'hbd143dc6} /* (18, 3, 24) {real, imag} */,
  {32'hbd106a19, 32'hbd785d41} /* (18, 3, 23) {real, imag} */,
  {32'hbcb67196, 32'hbd968b61} /* (18, 3, 22) {real, imag} */,
  {32'h3e039d34, 32'h3b3748b0} /* (18, 3, 21) {real, imag} */,
  {32'h3bf60b58, 32'hbceedd63} /* (18, 3, 20) {real, imag} */,
  {32'hbc1c461a, 32'hbcaf324f} /* (18, 3, 19) {real, imag} */,
  {32'h3bfcbc9b, 32'h3ca720ca} /* (18, 3, 18) {real, imag} */,
  {32'h3a246940, 32'h3c72a49b} /* (18, 3, 17) {real, imag} */,
  {32'h3d38b576, 32'h00000000} /* (18, 3, 16) {real, imag} */,
  {32'h3a246940, 32'hbc72a49b} /* (18, 3, 15) {real, imag} */,
  {32'h3bfcbc9b, 32'hbca720ca} /* (18, 3, 14) {real, imag} */,
  {32'hbc1c461a, 32'h3caf324f} /* (18, 3, 13) {real, imag} */,
  {32'h3bf60b58, 32'h3ceedd63} /* (18, 3, 12) {real, imag} */,
  {32'h3e039d34, 32'hbb3748b0} /* (18, 3, 11) {real, imag} */,
  {32'hbcb67196, 32'h3d968b61} /* (18, 3, 10) {real, imag} */,
  {32'hbd106a19, 32'h3d785d41} /* (18, 3, 9) {real, imag} */,
  {32'h3d74532c, 32'h3d143dc6} /* (18, 3, 8) {real, imag} */,
  {32'hbc42c1b0, 32'hbdc0416e} /* (18, 3, 7) {real, imag} */,
  {32'h3c92e878, 32'h3d3198bc} /* (18, 3, 6) {real, imag} */,
  {32'h3e81621d, 32'hbde9697b} /* (18, 3, 5) {real, imag} */,
  {32'h3d852b4b, 32'h3e08bd40} /* (18, 3, 4) {real, imag} */,
  {32'h3cc9949c, 32'h3d2f5a0b} /* (18, 3, 3) {real, imag} */,
  {32'hbeb1b311, 32'h3f941cf2} /* (18, 3, 2) {real, imag} */,
  {32'hc017395a, 32'hc03c9420} /* (18, 3, 1) {real, imag} */,
  {32'hc0655107, 32'h00000000} /* (18, 3, 0) {real, imag} */,
  {32'hc0133630, 32'h40398ede} /* (18, 2, 31) {real, imag} */,
  {32'hbed4f5b7, 32'hbf8a9220} /* (18, 2, 30) {real, imag} */,
  {32'h3df86db3, 32'hbcc31cd8} /* (18, 2, 29) {real, imag} */,
  {32'h3dd3bbc3, 32'hbe83f6ee} /* (18, 2, 28) {real, imag} */,
  {32'h3e2253d8, 32'h3e2a7d92} /* (18, 2, 27) {real, imag} */,
  {32'hbb0304a0, 32'hbcf2264a} /* (18, 2, 26) {real, imag} */,
  {32'hbd6aa5da, 32'h3c3121d8} /* (18, 2, 25) {real, imag} */,
  {32'h3d5ee9fe, 32'h3a2e1b40} /* (18, 2, 24) {real, imag} */,
  {32'h3dc1df95, 32'hbdc5561e} /* (18, 2, 23) {real, imag} */,
  {32'h3d67415c, 32'hbcf9a1b3} /* (18, 2, 22) {real, imag} */,
  {32'h3dd13a3c, 32'h3bfc1d00} /* (18, 2, 21) {real, imag} */,
  {32'hbc1a2532, 32'hbd9b39b0} /* (18, 2, 20) {real, imag} */,
  {32'h3d7eda64, 32'h3cce66be} /* (18, 2, 19) {real, imag} */,
  {32'hbdfed610, 32'hbd2ce3ad} /* (18, 2, 18) {real, imag} */,
  {32'h3d4cd323, 32'hbc614196} /* (18, 2, 17) {real, imag} */,
  {32'h3cb8a754, 32'h00000000} /* (18, 2, 16) {real, imag} */,
  {32'h3d4cd323, 32'h3c614196} /* (18, 2, 15) {real, imag} */,
  {32'hbdfed610, 32'h3d2ce3ad} /* (18, 2, 14) {real, imag} */,
  {32'h3d7eda64, 32'hbcce66be} /* (18, 2, 13) {real, imag} */,
  {32'hbc1a2532, 32'h3d9b39b0} /* (18, 2, 12) {real, imag} */,
  {32'h3dd13a3c, 32'hbbfc1d00} /* (18, 2, 11) {real, imag} */,
  {32'h3d67415c, 32'h3cf9a1b3} /* (18, 2, 10) {real, imag} */,
  {32'h3dc1df95, 32'h3dc5561e} /* (18, 2, 9) {real, imag} */,
  {32'h3d5ee9fe, 32'hba2e1b40} /* (18, 2, 8) {real, imag} */,
  {32'hbd6aa5da, 32'hbc3121d8} /* (18, 2, 7) {real, imag} */,
  {32'hbb0304a0, 32'h3cf2264a} /* (18, 2, 6) {real, imag} */,
  {32'h3e2253d8, 32'hbe2a7d92} /* (18, 2, 5) {real, imag} */,
  {32'h3dd3bbc3, 32'h3e83f6ee} /* (18, 2, 4) {real, imag} */,
  {32'h3df86db3, 32'h3cc31cd8} /* (18, 2, 3) {real, imag} */,
  {32'hbed4f5b7, 32'h3f8a9220} /* (18, 2, 2) {real, imag} */,
  {32'hc0133630, 32'hc0398ede} /* (18, 2, 1) {real, imag} */,
  {32'hc0727bbf, 32'h00000000} /* (18, 2, 0) {real, imag} */,
  {32'hc01bec4f, 32'h402afb01} /* (18, 1, 31) {real, imag} */,
  {32'hbe96a812, 32'hbf7df188} /* (18, 1, 30) {real, imag} */,
  {32'h3e081d22, 32'h3daffa3a} /* (18, 1, 29) {real, imag} */,
  {32'h3cb27aa9, 32'hbe91f218} /* (18, 1, 28) {real, imag} */,
  {32'h3e1e144a, 32'h3e0d1c63} /* (18, 1, 27) {real, imag} */,
  {32'h3e192cc0, 32'hbd806d78} /* (18, 1, 26) {real, imag} */,
  {32'h3cc137f6, 32'hbc158276} /* (18, 1, 25) {real, imag} */,
  {32'h3dd2e7b4, 32'hbcae8fe4} /* (18, 1, 24) {real, imag} */,
  {32'h3cd8c1ad, 32'h3c8737a7} /* (18, 1, 23) {real, imag} */,
  {32'h3c82358f, 32'h3cf48784} /* (18, 1, 22) {real, imag} */,
  {32'h3c6ca704, 32'hbba2a7b8} /* (18, 1, 21) {real, imag} */,
  {32'h3c2ad9b2, 32'h3cf2a36a} /* (18, 1, 20) {real, imag} */,
  {32'hbcd81014, 32'h3d4437d8} /* (18, 1, 19) {real, imag} */,
  {32'hbd0236b5, 32'h3b55d190} /* (18, 1, 18) {real, imag} */,
  {32'h3cd364e1, 32'h3ce5a60d} /* (18, 1, 17) {real, imag} */,
  {32'h3bf0ad5c, 32'h00000000} /* (18, 1, 16) {real, imag} */,
  {32'h3cd364e1, 32'hbce5a60d} /* (18, 1, 15) {real, imag} */,
  {32'hbd0236b5, 32'hbb55d190} /* (18, 1, 14) {real, imag} */,
  {32'hbcd81014, 32'hbd4437d8} /* (18, 1, 13) {real, imag} */,
  {32'h3c2ad9b2, 32'hbcf2a36a} /* (18, 1, 12) {real, imag} */,
  {32'h3c6ca704, 32'h3ba2a7b8} /* (18, 1, 11) {real, imag} */,
  {32'h3c82358f, 32'hbcf48784} /* (18, 1, 10) {real, imag} */,
  {32'h3cd8c1ad, 32'hbc8737a7} /* (18, 1, 9) {real, imag} */,
  {32'h3dd2e7b4, 32'h3cae8fe4} /* (18, 1, 8) {real, imag} */,
  {32'h3cc137f6, 32'h3c158276} /* (18, 1, 7) {real, imag} */,
  {32'h3e192cc0, 32'h3d806d78} /* (18, 1, 6) {real, imag} */,
  {32'h3e1e144a, 32'hbe0d1c63} /* (18, 1, 5) {real, imag} */,
  {32'h3cb27aa9, 32'h3e91f218} /* (18, 1, 4) {real, imag} */,
  {32'h3e081d22, 32'hbdaffa3a} /* (18, 1, 3) {real, imag} */,
  {32'hbe96a812, 32'h3f7df188} /* (18, 1, 2) {real, imag} */,
  {32'hc01bec4f, 32'hc02afb01} /* (18, 1, 1) {real, imag} */,
  {32'hc0794a06, 32'h00000000} /* (18, 1, 0) {real, imag} */,
  {32'hc02a71c4, 32'h400b0ae4} /* (18, 0, 31) {real, imag} */,
  {32'h3ca56ae0, 32'hbf34e6a2} /* (18, 0, 30) {real, imag} */,
  {32'h3c3bdd10, 32'h3d676d34} /* (18, 0, 29) {real, imag} */,
  {32'hbbdd8840, 32'hbe18d88c} /* (18, 0, 28) {real, imag} */,
  {32'h3dac61fa, 32'hbc76d090} /* (18, 0, 27) {real, imag} */,
  {32'hbabc1230, 32'hbd1d74e1} /* (18, 0, 26) {real, imag} */,
  {32'h3c931ddb, 32'h3cc4f868} /* (18, 0, 25) {real, imag} */,
  {32'h3d6fdc78, 32'hbdb14b32} /* (18, 0, 24) {real, imag} */,
  {32'hbb74823c, 32'h3d792196} /* (18, 0, 23) {real, imag} */,
  {32'h3c88c5a7, 32'hbd466b32} /* (18, 0, 22) {real, imag} */,
  {32'hbc91cf74, 32'hbd08caff} /* (18, 0, 21) {real, imag} */,
  {32'h3d7fb774, 32'hbcd1acbd} /* (18, 0, 20) {real, imag} */,
  {32'h3d8e445b, 32'h3c91eb1c} /* (18, 0, 19) {real, imag} */,
  {32'h3d189fe5, 32'h3cee0e38} /* (18, 0, 18) {real, imag} */,
  {32'h3c847792, 32'hbbc50b92} /* (18, 0, 17) {real, imag} */,
  {32'hbca83c14, 32'h00000000} /* (18, 0, 16) {real, imag} */,
  {32'h3c847792, 32'h3bc50b92} /* (18, 0, 15) {real, imag} */,
  {32'h3d189fe5, 32'hbcee0e38} /* (18, 0, 14) {real, imag} */,
  {32'h3d8e445b, 32'hbc91eb1c} /* (18, 0, 13) {real, imag} */,
  {32'h3d7fb774, 32'h3cd1acbd} /* (18, 0, 12) {real, imag} */,
  {32'hbc91cf74, 32'h3d08caff} /* (18, 0, 11) {real, imag} */,
  {32'h3c88c5a7, 32'h3d466b32} /* (18, 0, 10) {real, imag} */,
  {32'hbb74823c, 32'hbd792196} /* (18, 0, 9) {real, imag} */,
  {32'h3d6fdc78, 32'h3db14b32} /* (18, 0, 8) {real, imag} */,
  {32'h3c931ddb, 32'hbcc4f868} /* (18, 0, 7) {real, imag} */,
  {32'hbabc1230, 32'h3d1d74e1} /* (18, 0, 6) {real, imag} */,
  {32'h3dac61fa, 32'h3c76d090} /* (18, 0, 5) {real, imag} */,
  {32'hbbdd8840, 32'h3e18d88c} /* (18, 0, 4) {real, imag} */,
  {32'h3c3bdd10, 32'hbd676d34} /* (18, 0, 3) {real, imag} */,
  {32'h3ca56ae0, 32'h3f34e6a2} /* (18, 0, 2) {real, imag} */,
  {32'hc02a71c4, 32'hc00b0ae4} /* (18, 0, 1) {real, imag} */,
  {32'hc067dd84, 32'h00000000} /* (18, 0, 0) {real, imag} */,
  {32'hc007eb98, 32'h3f8ad737} /* (17, 31, 31) {real, imag} */,
  {32'h3ee92877, 32'hbef23056} /* (17, 31, 30) {real, imag} */,
  {32'h3d46adae, 32'h3d1737b6} /* (17, 31, 29) {real, imag} */,
  {32'hbd041f2a, 32'h3c8e6fd0} /* (17, 31, 28) {real, imag} */,
  {32'h3d78ecf2, 32'hbd385544} /* (17, 31, 27) {real, imag} */,
  {32'h3d5eb6eb, 32'h3b734710} /* (17, 31, 26) {real, imag} */,
  {32'h3c880512, 32'h3bd38388} /* (17, 31, 25) {real, imag} */,
  {32'hbcf85a89, 32'hbd511308} /* (17, 31, 24) {real, imag} */,
  {32'hbaa77fd0, 32'h3c8912d2} /* (17, 31, 23) {real, imag} */,
  {32'h3c3108f0, 32'h3ce23736} /* (17, 31, 22) {real, imag} */,
  {32'h3d827b4c, 32'hbd6b62df} /* (17, 31, 21) {real, imag} */,
  {32'hbc0e136c, 32'h3b927b60} /* (17, 31, 20) {real, imag} */,
  {32'h3cf8a8a5, 32'h3c6c3ff7} /* (17, 31, 19) {real, imag} */,
  {32'hbd957e63, 32'hbbb5ba78} /* (17, 31, 18) {real, imag} */,
  {32'h3d34a4f0, 32'hbc5a37e2} /* (17, 31, 17) {real, imag} */,
  {32'hbb8674ac, 32'h00000000} /* (17, 31, 16) {real, imag} */,
  {32'h3d34a4f0, 32'h3c5a37e2} /* (17, 31, 15) {real, imag} */,
  {32'hbd957e63, 32'h3bb5ba78} /* (17, 31, 14) {real, imag} */,
  {32'h3cf8a8a5, 32'hbc6c3ff7} /* (17, 31, 13) {real, imag} */,
  {32'hbc0e136c, 32'hbb927b60} /* (17, 31, 12) {real, imag} */,
  {32'h3d827b4c, 32'h3d6b62df} /* (17, 31, 11) {real, imag} */,
  {32'h3c3108f0, 32'hbce23736} /* (17, 31, 10) {real, imag} */,
  {32'hbaa77fd0, 32'hbc8912d2} /* (17, 31, 9) {real, imag} */,
  {32'hbcf85a89, 32'h3d511308} /* (17, 31, 8) {real, imag} */,
  {32'h3c880512, 32'hbbd38388} /* (17, 31, 7) {real, imag} */,
  {32'h3d5eb6eb, 32'hbb734710} /* (17, 31, 6) {real, imag} */,
  {32'h3d78ecf2, 32'h3d385544} /* (17, 31, 5) {real, imag} */,
  {32'hbd041f2a, 32'hbc8e6fd0} /* (17, 31, 4) {real, imag} */,
  {32'h3d46adae, 32'hbd1737b6} /* (17, 31, 3) {real, imag} */,
  {32'h3ee92877, 32'h3ef23056} /* (17, 31, 2) {real, imag} */,
  {32'hc007eb98, 32'hbf8ad737} /* (17, 31, 1) {real, imag} */,
  {32'hc02253aa, 32'h00000000} /* (17, 31, 0) {real, imag} */,
  {32'hc02d42b2, 32'h3f41df68} /* (17, 30, 31) {real, imag} */,
  {32'h3f4b3d3f, 32'hbed27684} /* (17, 30, 30) {real, imag} */,
  {32'h3cbfac50, 32'h3d9cb4a4} /* (17, 30, 29) {real, imag} */,
  {32'hbdd09e50, 32'h3ddc7b26} /* (17, 30, 28) {real, imag} */,
  {32'h3e81cff2, 32'hbd25bc6c} /* (17, 30, 27) {real, imag} */,
  {32'h3d86666c, 32'hbda58990} /* (17, 30, 26) {real, imag} */,
  {32'h3d2b689c, 32'hbc968a88} /* (17, 30, 25) {real, imag} */,
  {32'h3d9ef7b0, 32'hbe065407} /* (17, 30, 24) {real, imag} */,
  {32'hbd83e182, 32'h3d99d4ac} /* (17, 30, 23) {real, imag} */,
  {32'h3d2673df, 32'h3d25b215} /* (17, 30, 22) {real, imag} */,
  {32'h3d2baea4, 32'hbcb4f328} /* (17, 30, 21) {real, imag} */,
  {32'hbc336ddc, 32'h3d5c08f4} /* (17, 30, 20) {real, imag} */,
  {32'h3c534bec, 32'h3cf65f81} /* (17, 30, 19) {real, imag} */,
  {32'hbcdb8596, 32'hbba7d0cc} /* (17, 30, 18) {real, imag} */,
  {32'hbc4cfe44, 32'h3d08682c} /* (17, 30, 17) {real, imag} */,
  {32'hbc3fc278, 32'h00000000} /* (17, 30, 16) {real, imag} */,
  {32'hbc4cfe44, 32'hbd08682c} /* (17, 30, 15) {real, imag} */,
  {32'hbcdb8596, 32'h3ba7d0cc} /* (17, 30, 14) {real, imag} */,
  {32'h3c534bec, 32'hbcf65f81} /* (17, 30, 13) {real, imag} */,
  {32'hbc336ddc, 32'hbd5c08f4} /* (17, 30, 12) {real, imag} */,
  {32'h3d2baea4, 32'h3cb4f328} /* (17, 30, 11) {real, imag} */,
  {32'h3d2673df, 32'hbd25b215} /* (17, 30, 10) {real, imag} */,
  {32'hbd83e182, 32'hbd99d4ac} /* (17, 30, 9) {real, imag} */,
  {32'h3d9ef7b0, 32'h3e065407} /* (17, 30, 8) {real, imag} */,
  {32'h3d2b689c, 32'h3c968a88} /* (17, 30, 7) {real, imag} */,
  {32'h3d86666c, 32'h3da58990} /* (17, 30, 6) {real, imag} */,
  {32'h3e81cff2, 32'h3d25bc6c} /* (17, 30, 5) {real, imag} */,
  {32'hbdd09e50, 32'hbddc7b26} /* (17, 30, 4) {real, imag} */,
  {32'h3cbfac50, 32'hbd9cb4a4} /* (17, 30, 3) {real, imag} */,
  {32'h3f4b3d3f, 32'h3ed27684} /* (17, 30, 2) {real, imag} */,
  {32'hc02d42b2, 32'hbf41df68} /* (17, 30, 1) {real, imag} */,
  {32'hc02e1a99, 32'h00000000} /* (17, 30, 0) {real, imag} */,
  {32'hc0442b02, 32'h3f27b7e8} /* (17, 29, 31) {real, imag} */,
  {32'h3f833d6f, 32'hbead2b6b} /* (17, 29, 30) {real, imag} */,
  {32'hbda52ede, 32'h3dc850a8} /* (17, 29, 29) {real, imag} */,
  {32'hbe3ce1c0, 32'h3de30058} /* (17, 29, 28) {real, imag} */,
  {32'h3e4f0498, 32'hbd1492f0} /* (17, 29, 27) {real, imag} */,
  {32'h3dfcf2ca, 32'hbbd47620} /* (17, 29, 26) {real, imag} */,
  {32'hbd60a7f7, 32'h3abc9980} /* (17, 29, 25) {real, imag} */,
  {32'h3d328b52, 32'hbcacb088} /* (17, 29, 24) {real, imag} */,
  {32'hbde5019e, 32'hbdacf9b8} /* (17, 29, 23) {real, imag} */,
  {32'h3dbbea76, 32'h3d066546} /* (17, 29, 22) {real, imag} */,
  {32'hbc9fc100, 32'hbbc91cf0} /* (17, 29, 21) {real, imag} */,
  {32'hbdcd4bdc, 32'h3a95cb98} /* (17, 29, 20) {real, imag} */,
  {32'h3c06b8a9, 32'h3d0bdc08} /* (17, 29, 19) {real, imag} */,
  {32'hbc0e3b44, 32'hbcc0fd4a} /* (17, 29, 18) {real, imag} */,
  {32'hbcb8262d, 32'h3ca6156a} /* (17, 29, 17) {real, imag} */,
  {32'hbdde41b4, 32'h00000000} /* (17, 29, 16) {real, imag} */,
  {32'hbcb8262d, 32'hbca6156a} /* (17, 29, 15) {real, imag} */,
  {32'hbc0e3b44, 32'h3cc0fd4a} /* (17, 29, 14) {real, imag} */,
  {32'h3c06b8a9, 32'hbd0bdc08} /* (17, 29, 13) {real, imag} */,
  {32'hbdcd4bdc, 32'hba95cb98} /* (17, 29, 12) {real, imag} */,
  {32'hbc9fc100, 32'h3bc91cf0} /* (17, 29, 11) {real, imag} */,
  {32'h3dbbea76, 32'hbd066546} /* (17, 29, 10) {real, imag} */,
  {32'hbde5019e, 32'h3dacf9b8} /* (17, 29, 9) {real, imag} */,
  {32'h3d328b52, 32'h3cacb088} /* (17, 29, 8) {real, imag} */,
  {32'hbd60a7f7, 32'hbabc9980} /* (17, 29, 7) {real, imag} */,
  {32'h3dfcf2ca, 32'h3bd47620} /* (17, 29, 6) {real, imag} */,
  {32'h3e4f0498, 32'h3d1492f0} /* (17, 29, 5) {real, imag} */,
  {32'hbe3ce1c0, 32'hbde30058} /* (17, 29, 4) {real, imag} */,
  {32'hbda52ede, 32'hbdc850a8} /* (17, 29, 3) {real, imag} */,
  {32'h3f833d6f, 32'h3ead2b6b} /* (17, 29, 2) {real, imag} */,
  {32'hc0442b02, 32'hbf27b7e8} /* (17, 29, 1) {real, imag} */,
  {32'hc03331de, 32'h00000000} /* (17, 29, 0) {real, imag} */,
  {32'hc049b455, 32'h3f13a116} /* (17, 28, 31) {real, imag} */,
  {32'h3f82c906, 32'hbecf5d1a} /* (17, 28, 30) {real, imag} */,
  {32'hbc60cd28, 32'hbca8bce7} /* (17, 28, 29) {real, imag} */,
  {32'hbe261405, 32'h3d6b8e36} /* (17, 28, 28) {real, imag} */,
  {32'h3e0b90b6, 32'hbd5211ec} /* (17, 28, 27) {real, imag} */,
  {32'h3e0ab31d, 32'h3c13387a} /* (17, 28, 26) {real, imag} */,
  {32'hbbfe3508, 32'hbd15e397} /* (17, 28, 25) {real, imag} */,
  {32'h3cbbcf82, 32'hbcc6b734} /* (17, 28, 24) {real, imag} */,
  {32'h3d820c4a, 32'h3cfb97e1} /* (17, 28, 23) {real, imag} */,
  {32'h3c85858f, 32'h3c048348} /* (17, 28, 22) {real, imag} */,
  {32'h3d592726, 32'hbd903352} /* (17, 28, 21) {real, imag} */,
  {32'h3d029686, 32'hbd102d8a} /* (17, 28, 20) {real, imag} */,
  {32'hbcea213c, 32'hbb07ff30} /* (17, 28, 19) {real, imag} */,
  {32'hbd289712, 32'h3d1e3766} /* (17, 28, 18) {real, imag} */,
  {32'h3cbfa640, 32'h3c4cb87a} /* (17, 28, 17) {real, imag} */,
  {32'hbcaa09f0, 32'h00000000} /* (17, 28, 16) {real, imag} */,
  {32'h3cbfa640, 32'hbc4cb87a} /* (17, 28, 15) {real, imag} */,
  {32'hbd289712, 32'hbd1e3766} /* (17, 28, 14) {real, imag} */,
  {32'hbcea213c, 32'h3b07ff30} /* (17, 28, 13) {real, imag} */,
  {32'h3d029686, 32'h3d102d8a} /* (17, 28, 12) {real, imag} */,
  {32'h3d592726, 32'h3d903352} /* (17, 28, 11) {real, imag} */,
  {32'h3c85858f, 32'hbc048348} /* (17, 28, 10) {real, imag} */,
  {32'h3d820c4a, 32'hbcfb97e1} /* (17, 28, 9) {real, imag} */,
  {32'h3cbbcf82, 32'h3cc6b734} /* (17, 28, 8) {real, imag} */,
  {32'hbbfe3508, 32'h3d15e397} /* (17, 28, 7) {real, imag} */,
  {32'h3e0ab31d, 32'hbc13387a} /* (17, 28, 6) {real, imag} */,
  {32'h3e0b90b6, 32'h3d5211ec} /* (17, 28, 5) {real, imag} */,
  {32'hbe261405, 32'hbd6b8e36} /* (17, 28, 4) {real, imag} */,
  {32'hbc60cd28, 32'h3ca8bce7} /* (17, 28, 3) {real, imag} */,
  {32'h3f82c906, 32'h3ecf5d1a} /* (17, 28, 2) {real, imag} */,
  {32'hc049b455, 32'hbf13a116} /* (17, 28, 1) {real, imag} */,
  {32'hc032fd44, 32'h00000000} /* (17, 28, 0) {real, imag} */,
  {32'hc0485a97, 32'h3eca91b0} /* (17, 27, 31) {real, imag} */,
  {32'h3f8e1bec, 32'hbefb8640} /* (17, 27, 30) {real, imag} */,
  {32'hbd9c4d4c, 32'hbd982448} /* (17, 27, 29) {real, imag} */,
  {32'hbe6f6663, 32'h3e55609b} /* (17, 27, 28) {real, imag} */,
  {32'h3e269661, 32'hbd818300} /* (17, 27, 27) {real, imag} */,
  {32'h3da0b19d, 32'h3d95784d} /* (17, 27, 26) {real, imag} */,
  {32'hbb802130, 32'hbb839060} /* (17, 27, 25) {real, imag} */,
  {32'h3de4de15, 32'hbc6a37b8} /* (17, 27, 24) {real, imag} */,
  {32'h3de6efa0, 32'hbd1190d9} /* (17, 27, 23) {real, imag} */,
  {32'h3b878b90, 32'hbcb9ae24} /* (17, 27, 22) {real, imag} */,
  {32'h3daed4e4, 32'hbda5d49f} /* (17, 27, 21) {real, imag} */,
  {32'h3da93fc8, 32'h3d412a66} /* (17, 27, 20) {real, imag} */,
  {32'h3d0d7c0d, 32'h3d3e3b83} /* (17, 27, 19) {real, imag} */,
  {32'hbd0e2494, 32'hbd5cc7f8} /* (17, 27, 18) {real, imag} */,
  {32'h3cb86bc4, 32'h3da2d629} /* (17, 27, 17) {real, imag} */,
  {32'h3c79036c, 32'h00000000} /* (17, 27, 16) {real, imag} */,
  {32'h3cb86bc4, 32'hbda2d629} /* (17, 27, 15) {real, imag} */,
  {32'hbd0e2494, 32'h3d5cc7f8} /* (17, 27, 14) {real, imag} */,
  {32'h3d0d7c0d, 32'hbd3e3b83} /* (17, 27, 13) {real, imag} */,
  {32'h3da93fc8, 32'hbd412a66} /* (17, 27, 12) {real, imag} */,
  {32'h3daed4e4, 32'h3da5d49f} /* (17, 27, 11) {real, imag} */,
  {32'h3b878b90, 32'h3cb9ae24} /* (17, 27, 10) {real, imag} */,
  {32'h3de6efa0, 32'h3d1190d9} /* (17, 27, 9) {real, imag} */,
  {32'h3de4de15, 32'h3c6a37b8} /* (17, 27, 8) {real, imag} */,
  {32'hbb802130, 32'h3b839060} /* (17, 27, 7) {real, imag} */,
  {32'h3da0b19d, 32'hbd95784d} /* (17, 27, 6) {real, imag} */,
  {32'h3e269661, 32'h3d818300} /* (17, 27, 5) {real, imag} */,
  {32'hbe6f6663, 32'hbe55609b} /* (17, 27, 4) {real, imag} */,
  {32'hbd9c4d4c, 32'h3d982448} /* (17, 27, 3) {real, imag} */,
  {32'h3f8e1bec, 32'h3efb8640} /* (17, 27, 2) {real, imag} */,
  {32'hc0485a97, 32'hbeca91b0} /* (17, 27, 1) {real, imag} */,
  {32'hc039a72c, 32'h00000000} /* (17, 27, 0) {real, imag} */,
  {32'hc036c6ed, 32'h3e5e930c} /* (17, 26, 31) {real, imag} */,
  {32'h3f863e36, 32'hbed983a2} /* (17, 26, 30) {real, imag} */,
  {32'hbcff52aa, 32'h3c1b2fae} /* (17, 26, 29) {real, imag} */,
  {32'hbe8aa62a, 32'hbd899e88} /* (17, 26, 28) {real, imag} */,
  {32'h3e1b4574, 32'hbd105f0a} /* (17, 26, 27) {real, imag} */,
  {32'hbc47eee8, 32'h3caa3c5a} /* (17, 26, 26) {real, imag} */,
  {32'hbce3ddc3, 32'h3d847b48} /* (17, 26, 25) {real, imag} */,
  {32'h3da5a7d9, 32'hbd0ae5b0} /* (17, 26, 24) {real, imag} */,
  {32'h3b1f6284, 32'hbdb7098c} /* (17, 26, 23) {real, imag} */,
  {32'hbc8d836e, 32'h3c710160} /* (17, 26, 22) {real, imag} */,
  {32'hbaaa6b40, 32'hbd4d9663} /* (17, 26, 21) {real, imag} */,
  {32'h3cca36b1, 32'h3d9bde85} /* (17, 26, 20) {real, imag} */,
  {32'hbd6983a5, 32'hbd69db0c} /* (17, 26, 19) {real, imag} */,
  {32'h3d078993, 32'hbd3a5a38} /* (17, 26, 18) {real, imag} */,
  {32'hbbce3840, 32'h3d0f6928} /* (17, 26, 17) {real, imag} */,
  {32'hbda2ad36, 32'h00000000} /* (17, 26, 16) {real, imag} */,
  {32'hbbce3840, 32'hbd0f6928} /* (17, 26, 15) {real, imag} */,
  {32'h3d078993, 32'h3d3a5a38} /* (17, 26, 14) {real, imag} */,
  {32'hbd6983a5, 32'h3d69db0c} /* (17, 26, 13) {real, imag} */,
  {32'h3cca36b1, 32'hbd9bde85} /* (17, 26, 12) {real, imag} */,
  {32'hbaaa6b40, 32'h3d4d9663} /* (17, 26, 11) {real, imag} */,
  {32'hbc8d836e, 32'hbc710160} /* (17, 26, 10) {real, imag} */,
  {32'h3b1f6284, 32'h3db7098c} /* (17, 26, 9) {real, imag} */,
  {32'h3da5a7d9, 32'h3d0ae5b0} /* (17, 26, 8) {real, imag} */,
  {32'hbce3ddc3, 32'hbd847b48} /* (17, 26, 7) {real, imag} */,
  {32'hbc47eee8, 32'hbcaa3c5a} /* (17, 26, 6) {real, imag} */,
  {32'h3e1b4574, 32'h3d105f0a} /* (17, 26, 5) {real, imag} */,
  {32'hbe8aa62a, 32'h3d899e88} /* (17, 26, 4) {real, imag} */,
  {32'hbcff52aa, 32'hbc1b2fae} /* (17, 26, 3) {real, imag} */,
  {32'h3f863e36, 32'h3ed983a2} /* (17, 26, 2) {real, imag} */,
  {32'hc036c6ed, 32'hbe5e930c} /* (17, 26, 1) {real, imag} */,
  {32'hc0341ed8, 32'h00000000} /* (17, 26, 0) {real, imag} */,
  {32'hc02d0265, 32'h3e3a0450} /* (17, 25, 31) {real, imag} */,
  {32'h3f62a15b, 32'hbe913080} /* (17, 25, 30) {real, imag} */,
  {32'hbc6a0a64, 32'hbd0c734c} /* (17, 25, 29) {real, imag} */,
  {32'hbe95efc8, 32'hbd95e1ae} /* (17, 25, 28) {real, imag} */,
  {32'h3e4d33a7, 32'hbda05907} /* (17, 25, 27) {real, imag} */,
  {32'h3d8d40c4, 32'hbd246e98} /* (17, 25, 26) {real, imag} */,
  {32'hbdcfbaa6, 32'h3c95d318} /* (17, 25, 25) {real, imag} */,
  {32'h3e4c7dc4, 32'hbe191f6e} /* (17, 25, 24) {real, imag} */,
  {32'h3c8cdea0, 32'h3d2d4989} /* (17, 25, 23) {real, imag} */,
  {32'hbc8c7c4a, 32'hbcc7bf23} /* (17, 25, 22) {real, imag} */,
  {32'h3c1e14b5, 32'hbd72fd40} /* (17, 25, 21) {real, imag} */,
  {32'h3bd690fe, 32'hbc91aeea} /* (17, 25, 20) {real, imag} */,
  {32'hbd6c3a14, 32'hbd06a02a} /* (17, 25, 19) {real, imag} */,
  {32'h3cd23462, 32'hbd8ce112} /* (17, 25, 18) {real, imag} */,
  {32'h3ba34df1, 32'h3b745620} /* (17, 25, 17) {real, imag} */,
  {32'hbcac9c20, 32'h00000000} /* (17, 25, 16) {real, imag} */,
  {32'h3ba34df1, 32'hbb745620} /* (17, 25, 15) {real, imag} */,
  {32'h3cd23462, 32'h3d8ce112} /* (17, 25, 14) {real, imag} */,
  {32'hbd6c3a14, 32'h3d06a02a} /* (17, 25, 13) {real, imag} */,
  {32'h3bd690fe, 32'h3c91aeea} /* (17, 25, 12) {real, imag} */,
  {32'h3c1e14b5, 32'h3d72fd40} /* (17, 25, 11) {real, imag} */,
  {32'hbc8c7c4a, 32'h3cc7bf23} /* (17, 25, 10) {real, imag} */,
  {32'h3c8cdea0, 32'hbd2d4989} /* (17, 25, 9) {real, imag} */,
  {32'h3e4c7dc4, 32'h3e191f6e} /* (17, 25, 8) {real, imag} */,
  {32'hbdcfbaa6, 32'hbc95d318} /* (17, 25, 7) {real, imag} */,
  {32'h3d8d40c4, 32'h3d246e98} /* (17, 25, 6) {real, imag} */,
  {32'h3e4d33a7, 32'h3da05907} /* (17, 25, 5) {real, imag} */,
  {32'hbe95efc8, 32'h3d95e1ae} /* (17, 25, 4) {real, imag} */,
  {32'hbc6a0a64, 32'h3d0c734c} /* (17, 25, 3) {real, imag} */,
  {32'h3f62a15b, 32'h3e913080} /* (17, 25, 2) {real, imag} */,
  {32'hc02d0265, 32'hbe3a0450} /* (17, 25, 1) {real, imag} */,
  {32'hc0267050, 32'h00000000} /* (17, 25, 0) {real, imag} */,
  {32'hc01bd1a1, 32'h3e13a3aa} /* (17, 24, 31) {real, imag} */,
  {32'h3f6eebca, 32'hbdd06dc8} /* (17, 24, 30) {real, imag} */,
  {32'hbd573c2b, 32'hbd8c6d8b} /* (17, 24, 29) {real, imag} */,
  {32'hbea41372, 32'hbd855d47} /* (17, 24, 28) {real, imag} */,
  {32'h3e8d1d00, 32'hbe4e9952} /* (17, 24, 27) {real, imag} */,
  {32'hbd7b5dfc, 32'hbd80e818} /* (17, 24, 26) {real, imag} */,
  {32'hbd756b66, 32'h3cfc43df} /* (17, 24, 25) {real, imag} */,
  {32'h3e8ba308, 32'h3ad34960} /* (17, 24, 24) {real, imag} */,
  {32'hbd8b614b, 32'hbd514fa8} /* (17, 24, 23) {real, imag} */,
  {32'hba6a5580, 32'h3d3e24ce} /* (17, 24, 22) {real, imag} */,
  {32'h3d64146a, 32'hbdf0b728} /* (17, 24, 21) {real, imag} */,
  {32'hbd6061e2, 32'hbbdd2930} /* (17, 24, 20) {real, imag} */,
  {32'h3d650844, 32'hbd0598de} /* (17, 24, 19) {real, imag} */,
  {32'h3b884fe7, 32'hbdea6ea4} /* (17, 24, 18) {real, imag} */,
  {32'h3d255e6a, 32'hbb92a828} /* (17, 24, 17) {real, imag} */,
  {32'hbdeb9f86, 32'h00000000} /* (17, 24, 16) {real, imag} */,
  {32'h3d255e6a, 32'h3b92a828} /* (17, 24, 15) {real, imag} */,
  {32'h3b884fe7, 32'h3dea6ea4} /* (17, 24, 14) {real, imag} */,
  {32'h3d650844, 32'h3d0598de} /* (17, 24, 13) {real, imag} */,
  {32'hbd6061e2, 32'h3bdd2930} /* (17, 24, 12) {real, imag} */,
  {32'h3d64146a, 32'h3df0b728} /* (17, 24, 11) {real, imag} */,
  {32'hba6a5580, 32'hbd3e24ce} /* (17, 24, 10) {real, imag} */,
  {32'hbd8b614b, 32'h3d514fa8} /* (17, 24, 9) {real, imag} */,
  {32'h3e8ba308, 32'hbad34960} /* (17, 24, 8) {real, imag} */,
  {32'hbd756b66, 32'hbcfc43df} /* (17, 24, 7) {real, imag} */,
  {32'hbd7b5dfc, 32'h3d80e818} /* (17, 24, 6) {real, imag} */,
  {32'h3e8d1d00, 32'h3e4e9952} /* (17, 24, 5) {real, imag} */,
  {32'hbea41372, 32'h3d855d47} /* (17, 24, 4) {real, imag} */,
  {32'hbd573c2b, 32'h3d8c6d8b} /* (17, 24, 3) {real, imag} */,
  {32'h3f6eebca, 32'h3dd06dc8} /* (17, 24, 2) {real, imag} */,
  {32'hc01bd1a1, 32'hbe13a3aa} /* (17, 24, 1) {real, imag} */,
  {32'hc02119f2, 32'h00000000} /* (17, 24, 0) {real, imag} */,
  {32'hc002a5b2, 32'h3dcd63fc} /* (17, 23, 31) {real, imag} */,
  {32'h3f5cbc47, 32'hbd9026d3} /* (17, 23, 30) {real, imag} */,
  {32'h3d973eb6, 32'h3c6192c4} /* (17, 23, 29) {real, imag} */,
  {32'hbe0a1cac, 32'hbdb4e9f6} /* (17, 23, 28) {real, imag} */,
  {32'h3e628513, 32'hbe153120} /* (17, 23, 27) {real, imag} */,
  {32'hbcfc3828, 32'hbdcbc754} /* (17, 23, 26) {real, imag} */,
  {32'hbcd80864, 32'hba850780} /* (17, 23, 25) {real, imag} */,
  {32'h3d8d461b, 32'hbd075e82} /* (17, 23, 24) {real, imag} */,
  {32'hbc870360, 32'hbd6228f4} /* (17, 23, 23) {real, imag} */,
  {32'hbccd920a, 32'h3d87722a} /* (17, 23, 22) {real, imag} */,
  {32'hbccaf3ba, 32'h3ddb51f4} /* (17, 23, 21) {real, imag} */,
  {32'h3c96cea6, 32'hbc87cb7c} /* (17, 23, 20) {real, imag} */,
  {32'h3cd1b28b, 32'h3bfde608} /* (17, 23, 19) {real, imag} */,
  {32'hbd4a69f8, 32'hbc903dc0} /* (17, 23, 18) {real, imag} */,
  {32'h3d02a77c, 32'h3d31ea48} /* (17, 23, 17) {real, imag} */,
  {32'h3cbd31db, 32'h00000000} /* (17, 23, 16) {real, imag} */,
  {32'h3d02a77c, 32'hbd31ea48} /* (17, 23, 15) {real, imag} */,
  {32'hbd4a69f8, 32'h3c903dc0} /* (17, 23, 14) {real, imag} */,
  {32'h3cd1b28b, 32'hbbfde608} /* (17, 23, 13) {real, imag} */,
  {32'h3c96cea6, 32'h3c87cb7c} /* (17, 23, 12) {real, imag} */,
  {32'hbccaf3ba, 32'hbddb51f4} /* (17, 23, 11) {real, imag} */,
  {32'hbccd920a, 32'hbd87722a} /* (17, 23, 10) {real, imag} */,
  {32'hbc870360, 32'h3d6228f4} /* (17, 23, 9) {real, imag} */,
  {32'h3d8d461b, 32'h3d075e82} /* (17, 23, 8) {real, imag} */,
  {32'hbcd80864, 32'h3a850780} /* (17, 23, 7) {real, imag} */,
  {32'hbcfc3828, 32'h3dcbc754} /* (17, 23, 6) {real, imag} */,
  {32'h3e628513, 32'h3e153120} /* (17, 23, 5) {real, imag} */,
  {32'hbe0a1cac, 32'h3db4e9f6} /* (17, 23, 4) {real, imag} */,
  {32'h3d973eb6, 32'hbc6192c4} /* (17, 23, 3) {real, imag} */,
  {32'h3f5cbc47, 32'h3d9026d3} /* (17, 23, 2) {real, imag} */,
  {32'hc002a5b2, 32'hbdcd63fc} /* (17, 23, 1) {real, imag} */,
  {32'hc006929d, 32'h00000000} /* (17, 23, 0) {real, imag} */,
  {32'hbfb6a6f2, 32'h3dfd9fc8} /* (17, 22, 31) {real, imag} */,
  {32'h3f222d97, 32'hbdfdff52} /* (17, 22, 30) {real, imag} */,
  {32'hbd8e5dd4, 32'hbb882e98} /* (17, 22, 29) {real, imag} */,
  {32'hbde48000, 32'h3cdf477c} /* (17, 22, 28) {real, imag} */,
  {32'h3ddd4116, 32'hbdf7cc4b} /* (17, 22, 27) {real, imag} */,
  {32'hbcf715fc, 32'h3c645de8} /* (17, 22, 26) {real, imag} */,
  {32'hbd71f071, 32'h3d268e6e} /* (17, 22, 25) {real, imag} */,
  {32'h3ccf14f0, 32'hbd866dc1} /* (17, 22, 24) {real, imag} */,
  {32'h3d2e37a6, 32'hbc641454} /* (17, 22, 23) {real, imag} */,
  {32'hbcdcb172, 32'h3d717a8e} /* (17, 22, 22) {real, imag} */,
  {32'h3e046cb2, 32'hba1570c0} /* (17, 22, 21) {real, imag} */,
  {32'h3c7672b0, 32'h3d04422c} /* (17, 22, 20) {real, imag} */,
  {32'h3b3e0d70, 32'hbb3a41b0} /* (17, 22, 19) {real, imag} */,
  {32'hbc6aec98, 32'hbd05fb66} /* (17, 22, 18) {real, imag} */,
  {32'hbbe8c940, 32'h3d2f164b} /* (17, 22, 17) {real, imag} */,
  {32'hbd6bf93b, 32'h00000000} /* (17, 22, 16) {real, imag} */,
  {32'hbbe8c940, 32'hbd2f164b} /* (17, 22, 15) {real, imag} */,
  {32'hbc6aec98, 32'h3d05fb66} /* (17, 22, 14) {real, imag} */,
  {32'h3b3e0d70, 32'h3b3a41b0} /* (17, 22, 13) {real, imag} */,
  {32'h3c7672b0, 32'hbd04422c} /* (17, 22, 12) {real, imag} */,
  {32'h3e046cb2, 32'h3a1570c0} /* (17, 22, 11) {real, imag} */,
  {32'hbcdcb172, 32'hbd717a8e} /* (17, 22, 10) {real, imag} */,
  {32'h3d2e37a6, 32'h3c641454} /* (17, 22, 9) {real, imag} */,
  {32'h3ccf14f0, 32'h3d866dc1} /* (17, 22, 8) {real, imag} */,
  {32'hbd71f071, 32'hbd268e6e} /* (17, 22, 7) {real, imag} */,
  {32'hbcf715fc, 32'hbc645de8} /* (17, 22, 6) {real, imag} */,
  {32'h3ddd4116, 32'h3df7cc4b} /* (17, 22, 5) {real, imag} */,
  {32'hbde48000, 32'hbcdf477c} /* (17, 22, 4) {real, imag} */,
  {32'hbd8e5dd4, 32'h3b882e98} /* (17, 22, 3) {real, imag} */,
  {32'h3f222d97, 32'h3dfdff52} /* (17, 22, 2) {real, imag} */,
  {32'hbfb6a6f2, 32'hbdfd9fc8} /* (17, 22, 1) {real, imag} */,
  {32'hbfc53cf2, 32'h00000000} /* (17, 22, 0) {real, imag} */,
  {32'hbf13be73, 32'h3e423bf8} /* (17, 21, 31) {real, imag} */,
  {32'h3e7ee008, 32'h3e20e656} /* (17, 21, 30) {real, imag} */,
  {32'hbd11387c, 32'h3d037dd8} /* (17, 21, 29) {real, imag} */,
  {32'hbcb9e563, 32'hbc256bd8} /* (17, 21, 28) {real, imag} */,
  {32'h3daa7e9f, 32'hbd9738f3} /* (17, 21, 27) {real, imag} */,
  {32'hbcb9ae31, 32'hbd2b94da} /* (17, 21, 26) {real, imag} */,
  {32'h3b4213c0, 32'h3de3b12f} /* (17, 21, 25) {real, imag} */,
  {32'h3d2bab7d, 32'hbc1c9d20} /* (17, 21, 24) {real, imag} */,
  {32'h3d1f4e9c, 32'h3b16109a} /* (17, 21, 23) {real, imag} */,
  {32'hbc36d078, 32'hbd863d3a} /* (17, 21, 22) {real, imag} */,
  {32'hbc93b302, 32'hbdfc4d5a} /* (17, 21, 21) {real, imag} */,
  {32'hbd200c06, 32'hbd06c857} /* (17, 21, 20) {real, imag} */,
  {32'h3cdce098, 32'h3b30901e} /* (17, 21, 19) {real, imag} */,
  {32'hbafaeb00, 32'hbab715e0} /* (17, 21, 18) {real, imag} */,
  {32'hbc336ecb, 32'h3c979fd5} /* (17, 21, 17) {real, imag} */,
  {32'hbd6c9c49, 32'h00000000} /* (17, 21, 16) {real, imag} */,
  {32'hbc336ecb, 32'hbc979fd5} /* (17, 21, 15) {real, imag} */,
  {32'hbafaeb00, 32'h3ab715e0} /* (17, 21, 14) {real, imag} */,
  {32'h3cdce098, 32'hbb30901e} /* (17, 21, 13) {real, imag} */,
  {32'hbd200c06, 32'h3d06c857} /* (17, 21, 12) {real, imag} */,
  {32'hbc93b302, 32'h3dfc4d5a} /* (17, 21, 11) {real, imag} */,
  {32'hbc36d078, 32'h3d863d3a} /* (17, 21, 10) {real, imag} */,
  {32'h3d1f4e9c, 32'hbb16109a} /* (17, 21, 9) {real, imag} */,
  {32'h3d2bab7d, 32'h3c1c9d20} /* (17, 21, 8) {real, imag} */,
  {32'h3b4213c0, 32'hbde3b12f} /* (17, 21, 7) {real, imag} */,
  {32'hbcb9ae31, 32'h3d2b94da} /* (17, 21, 6) {real, imag} */,
  {32'h3daa7e9f, 32'h3d9738f3} /* (17, 21, 5) {real, imag} */,
  {32'hbcb9e563, 32'h3c256bd8} /* (17, 21, 4) {real, imag} */,
  {32'hbd11387c, 32'hbd037dd8} /* (17, 21, 3) {real, imag} */,
  {32'h3e7ee008, 32'hbe20e656} /* (17, 21, 2) {real, imag} */,
  {32'hbf13be73, 32'hbe423bf8} /* (17, 21, 1) {real, imag} */,
  {32'hbf493ea5, 32'h00000000} /* (17, 21, 0) {real, imag} */,
  {32'h3f082723, 32'h3d9a8d24} /* (17, 20, 31) {real, imag} */,
  {32'hbe8e11b5, 32'h3e951656} /* (17, 20, 30) {real, imag} */,
  {32'h3d0eaeb0, 32'hbde2e051} /* (17, 20, 29) {real, imag} */,
  {32'h3e3d9a18, 32'hbd599f0c} /* (17, 20, 28) {real, imag} */,
  {32'hbd3a6faa, 32'hbd6a2e6c} /* (17, 20, 27) {real, imag} */,
  {32'h3ca3cabc, 32'hbd494b87} /* (17, 20, 26) {real, imag} */,
  {32'h3d68d301, 32'h3d2271d4} /* (17, 20, 25) {real, imag} */,
  {32'hbdc63bb6, 32'h3cd6de60} /* (17, 20, 24) {real, imag} */,
  {32'hbd25a188, 32'hbb89c304} /* (17, 20, 23) {real, imag} */,
  {32'hbd4364d0, 32'hbde8d26c} /* (17, 20, 22) {real, imag} */,
  {32'hbd8dcdb0, 32'h3dc288a1} /* (17, 20, 21) {real, imag} */,
  {32'h3c628222, 32'h3d759382} /* (17, 20, 20) {real, imag} */,
  {32'hbbd5c062, 32'h3c099d14} /* (17, 20, 19) {real, imag} */,
  {32'hbd631dac, 32'h3da12ffb} /* (17, 20, 18) {real, imag} */,
  {32'h3d88eff9, 32'h3cf2a65b} /* (17, 20, 17) {real, imag} */,
  {32'hbbc571a1, 32'h00000000} /* (17, 20, 16) {real, imag} */,
  {32'h3d88eff9, 32'hbcf2a65b} /* (17, 20, 15) {real, imag} */,
  {32'hbd631dac, 32'hbda12ffb} /* (17, 20, 14) {real, imag} */,
  {32'hbbd5c062, 32'hbc099d14} /* (17, 20, 13) {real, imag} */,
  {32'h3c628222, 32'hbd759382} /* (17, 20, 12) {real, imag} */,
  {32'hbd8dcdb0, 32'hbdc288a1} /* (17, 20, 11) {real, imag} */,
  {32'hbd4364d0, 32'h3de8d26c} /* (17, 20, 10) {real, imag} */,
  {32'hbd25a188, 32'h3b89c304} /* (17, 20, 9) {real, imag} */,
  {32'hbdc63bb6, 32'hbcd6de60} /* (17, 20, 8) {real, imag} */,
  {32'h3d68d301, 32'hbd2271d4} /* (17, 20, 7) {real, imag} */,
  {32'h3ca3cabc, 32'h3d494b87} /* (17, 20, 6) {real, imag} */,
  {32'hbd3a6faa, 32'h3d6a2e6c} /* (17, 20, 5) {real, imag} */,
  {32'h3e3d9a18, 32'h3d599f0c} /* (17, 20, 4) {real, imag} */,
  {32'h3d0eaeb0, 32'h3de2e051} /* (17, 20, 3) {real, imag} */,
  {32'hbe8e11b5, 32'hbe951656} /* (17, 20, 2) {real, imag} */,
  {32'h3f082723, 32'hbd9a8d24} /* (17, 20, 1) {real, imag} */,
  {32'h3e4a9a04, 32'h00000000} /* (17, 20, 0) {real, imag} */,
  {32'h3fb0507e, 32'hbe2b9e52} /* (17, 19, 31) {real, imag} */,
  {32'hbf12c24a, 32'h3e9bbd16} /* (17, 19, 30) {real, imag} */,
  {32'h3e01c857, 32'h3dcdbe76} /* (17, 19, 29) {real, imag} */,
  {32'h3e5c6bb2, 32'hbce21baa} /* (17, 19, 28) {real, imag} */,
  {32'hbdd59792, 32'h3ce512c4} /* (17, 19, 27) {real, imag} */,
  {32'hbdb7d8c2, 32'h3d1eeff4} /* (17, 19, 26) {real, imag} */,
  {32'h3d5d7a48, 32'hbd7feb64} /* (17, 19, 25) {real, imag} */,
  {32'h3d321950, 32'h3dfb6416} /* (17, 19, 24) {real, imag} */,
  {32'hbd40598a, 32'h3d0af076} /* (17, 19, 23) {real, imag} */,
  {32'h3be661d8, 32'h3dada6cf} /* (17, 19, 22) {real, imag} */,
  {32'h3cc70dec, 32'h3c6b2bdc} /* (17, 19, 21) {real, imag} */,
  {32'h3d2a9ffc, 32'h3b0bdda0} /* (17, 19, 20) {real, imag} */,
  {32'h3d055047, 32'h3d27926a} /* (17, 19, 19) {real, imag} */,
  {32'h3d10bb41, 32'hbc98994c} /* (17, 19, 18) {real, imag} */,
  {32'h3bc992c0, 32'hbd509132} /* (17, 19, 17) {real, imag} */,
  {32'hbd492a1c, 32'h00000000} /* (17, 19, 16) {real, imag} */,
  {32'h3bc992c0, 32'h3d509132} /* (17, 19, 15) {real, imag} */,
  {32'h3d10bb41, 32'h3c98994c} /* (17, 19, 14) {real, imag} */,
  {32'h3d055047, 32'hbd27926a} /* (17, 19, 13) {real, imag} */,
  {32'h3d2a9ffc, 32'hbb0bdda0} /* (17, 19, 12) {real, imag} */,
  {32'h3cc70dec, 32'hbc6b2bdc} /* (17, 19, 11) {real, imag} */,
  {32'h3be661d8, 32'hbdada6cf} /* (17, 19, 10) {real, imag} */,
  {32'hbd40598a, 32'hbd0af076} /* (17, 19, 9) {real, imag} */,
  {32'h3d321950, 32'hbdfb6416} /* (17, 19, 8) {real, imag} */,
  {32'h3d5d7a48, 32'h3d7feb64} /* (17, 19, 7) {real, imag} */,
  {32'hbdb7d8c2, 32'hbd1eeff4} /* (17, 19, 6) {real, imag} */,
  {32'hbdd59792, 32'hbce512c4} /* (17, 19, 5) {real, imag} */,
  {32'h3e5c6bb2, 32'h3ce21baa} /* (17, 19, 4) {real, imag} */,
  {32'h3e01c857, 32'hbdcdbe76} /* (17, 19, 3) {real, imag} */,
  {32'hbf12c24a, 32'hbe9bbd16} /* (17, 19, 2) {real, imag} */,
  {32'h3fb0507e, 32'h3e2b9e52} /* (17, 19, 1) {real, imag} */,
  {32'h3f558985, 32'h00000000} /* (17, 19, 0) {real, imag} */,
  {32'h3ff6ea8b, 32'hbd985a5c} /* (17, 18, 31) {real, imag} */,
  {32'hbf46fae7, 32'h3e103e86} /* (17, 18, 30) {real, imag} */,
  {32'h3e1b9db6, 32'h3d607688} /* (17, 18, 29) {real, imag} */,
  {32'h3e83997b, 32'hbc25c120} /* (17, 18, 28) {real, imag} */,
  {32'hbe882440, 32'h3e373e44} /* (17, 18, 27) {real, imag} */,
  {32'hbe0a09ab, 32'h3d449394} /* (17, 18, 26) {real, imag} */,
  {32'h3db1a52d, 32'hbcbfffe9} /* (17, 18, 25) {real, imag} */,
  {32'h3cbd5a7e, 32'h3e414130} /* (17, 18, 24) {real, imag} */,
  {32'hbd939512, 32'hbcdb2648} /* (17, 18, 23) {real, imag} */,
  {32'h3d4d27f3, 32'hbd5248e4} /* (17, 18, 22) {real, imag} */,
  {32'h3d80a3b7, 32'h3d885f24} /* (17, 18, 21) {real, imag} */,
  {32'hbda9799e, 32'hbcd71ed3} /* (17, 18, 20) {real, imag} */,
  {32'h3c59e09f, 32'hbd1fe472} /* (17, 18, 19) {real, imag} */,
  {32'h3d23c847, 32'hbd3403ce} /* (17, 18, 18) {real, imag} */,
  {32'hbd76f822, 32'hbdb037a3} /* (17, 18, 17) {real, imag} */,
  {32'h3d8409b7, 32'h00000000} /* (17, 18, 16) {real, imag} */,
  {32'hbd76f822, 32'h3db037a3} /* (17, 18, 15) {real, imag} */,
  {32'h3d23c847, 32'h3d3403ce} /* (17, 18, 14) {real, imag} */,
  {32'h3c59e09f, 32'h3d1fe472} /* (17, 18, 13) {real, imag} */,
  {32'hbda9799e, 32'h3cd71ed3} /* (17, 18, 12) {real, imag} */,
  {32'h3d80a3b7, 32'hbd885f24} /* (17, 18, 11) {real, imag} */,
  {32'h3d4d27f3, 32'h3d5248e4} /* (17, 18, 10) {real, imag} */,
  {32'hbd939512, 32'h3cdb2648} /* (17, 18, 9) {real, imag} */,
  {32'h3cbd5a7e, 32'hbe414130} /* (17, 18, 8) {real, imag} */,
  {32'h3db1a52d, 32'h3cbfffe9} /* (17, 18, 7) {real, imag} */,
  {32'hbe0a09ab, 32'hbd449394} /* (17, 18, 6) {real, imag} */,
  {32'hbe882440, 32'hbe373e44} /* (17, 18, 5) {real, imag} */,
  {32'h3e83997b, 32'h3c25c120} /* (17, 18, 4) {real, imag} */,
  {32'h3e1b9db6, 32'hbd607688} /* (17, 18, 3) {real, imag} */,
  {32'hbf46fae7, 32'hbe103e86} /* (17, 18, 2) {real, imag} */,
  {32'h3ff6ea8b, 32'h3d985a5c} /* (17, 18, 1) {real, imag} */,
  {32'h3fb89718, 32'h00000000} /* (17, 18, 0) {real, imag} */,
  {32'h4009c7bf, 32'hbd6f1a88} /* (17, 17, 31) {real, imag} */,
  {32'hbf881b14, 32'h3d855c48} /* (17, 17, 30) {real, imag} */,
  {32'h3e70843e, 32'hbd788e00} /* (17, 17, 29) {real, imag} */,
  {32'h3e865f67, 32'hbca2b3c4} /* (17, 17, 28) {real, imag} */,
  {32'hbe980553, 32'h3e010dd2} /* (17, 17, 27) {real, imag} */,
  {32'hbe0721ff, 32'hbda53c66} /* (17, 17, 26) {real, imag} */,
  {32'h3dc7fa53, 32'h3cb87623} /* (17, 17, 25) {real, imag} */,
  {32'hbd3d3c50, 32'h3d4bfcc6} /* (17, 17, 24) {real, imag} */,
  {32'hbbbdda28, 32'h3bcb19a4} /* (17, 17, 23) {real, imag} */,
  {32'hbcdbc2b4, 32'h3d841422} /* (17, 17, 22) {real, imag} */,
  {32'hbd3a1e73, 32'h3cd9ab04} /* (17, 17, 21) {real, imag} */,
  {32'hbb97ae94, 32'hbe009b53} /* (17, 17, 20) {real, imag} */,
  {32'h3dd7c057, 32'h3d085f2d} /* (17, 17, 19) {real, imag} */,
  {32'hbd32dad2, 32'h3d9d594d} /* (17, 17, 18) {real, imag} */,
  {32'h3c312ccc, 32'hbae42720} /* (17, 17, 17) {real, imag} */,
  {32'h3d698b5a, 32'h00000000} /* (17, 17, 16) {real, imag} */,
  {32'h3c312ccc, 32'h3ae42720} /* (17, 17, 15) {real, imag} */,
  {32'hbd32dad2, 32'hbd9d594d} /* (17, 17, 14) {real, imag} */,
  {32'h3dd7c057, 32'hbd085f2d} /* (17, 17, 13) {real, imag} */,
  {32'hbb97ae94, 32'h3e009b53} /* (17, 17, 12) {real, imag} */,
  {32'hbd3a1e73, 32'hbcd9ab04} /* (17, 17, 11) {real, imag} */,
  {32'hbcdbc2b4, 32'hbd841422} /* (17, 17, 10) {real, imag} */,
  {32'hbbbdda28, 32'hbbcb19a4} /* (17, 17, 9) {real, imag} */,
  {32'hbd3d3c50, 32'hbd4bfcc6} /* (17, 17, 8) {real, imag} */,
  {32'h3dc7fa53, 32'hbcb87623} /* (17, 17, 7) {real, imag} */,
  {32'hbe0721ff, 32'h3da53c66} /* (17, 17, 6) {real, imag} */,
  {32'hbe980553, 32'hbe010dd2} /* (17, 17, 5) {real, imag} */,
  {32'h3e865f67, 32'h3ca2b3c4} /* (17, 17, 4) {real, imag} */,
  {32'h3e70843e, 32'h3d788e00} /* (17, 17, 3) {real, imag} */,
  {32'hbf881b14, 32'hbd855c48} /* (17, 17, 2) {real, imag} */,
  {32'h4009c7bf, 32'h3d6f1a88} /* (17, 17, 1) {real, imag} */,
  {32'h3fe193d6, 32'h00000000} /* (17, 17, 0) {real, imag} */,
  {32'h4014a63e, 32'hbe23f8b0} /* (17, 16, 31) {real, imag} */,
  {32'hbf9100b0, 32'h3e1814f8} /* (17, 16, 30) {real, imag} */,
  {32'h3e200772, 32'hbe1f8f7a} /* (17, 16, 29) {real, imag} */,
  {32'h3e96f416, 32'h3c3cea8c} /* (17, 16, 28) {real, imag} */,
  {32'hbe9b584b, 32'h3e32e98c} /* (17, 16, 27) {real, imag} */,
  {32'h3cf7555b, 32'hbd92685e} /* (17, 16, 26) {real, imag} */,
  {32'h3d5e3a04, 32'h3d324f18} /* (17, 16, 25) {real, imag} */,
  {32'hbcfdb244, 32'h3d6ebd45} /* (17, 16, 24) {real, imag} */,
  {32'h3d7460bf, 32'h3b822da8} /* (17, 16, 23) {real, imag} */,
  {32'hbd4fd83a, 32'h3d87f6fd} /* (17, 16, 22) {real, imag} */,
  {32'h3db065b6, 32'hbc74366b} /* (17, 16, 21) {real, imag} */,
  {32'hbd453334, 32'h3d0c7298} /* (17, 16, 20) {real, imag} */,
  {32'hbc844f79, 32'hbbc5c296} /* (17, 16, 19) {real, imag} */,
  {32'h3dba90ed, 32'h3c807334} /* (17, 16, 18) {real, imag} */,
  {32'hbdd37982, 32'h3d110d62} /* (17, 16, 17) {real, imag} */,
  {32'h3d59a181, 32'h00000000} /* (17, 16, 16) {real, imag} */,
  {32'hbdd37982, 32'hbd110d62} /* (17, 16, 15) {real, imag} */,
  {32'h3dba90ed, 32'hbc807334} /* (17, 16, 14) {real, imag} */,
  {32'hbc844f79, 32'h3bc5c296} /* (17, 16, 13) {real, imag} */,
  {32'hbd453334, 32'hbd0c7298} /* (17, 16, 12) {real, imag} */,
  {32'h3db065b6, 32'h3c74366b} /* (17, 16, 11) {real, imag} */,
  {32'hbd4fd83a, 32'hbd87f6fd} /* (17, 16, 10) {real, imag} */,
  {32'h3d7460bf, 32'hbb822da8} /* (17, 16, 9) {real, imag} */,
  {32'hbcfdb244, 32'hbd6ebd45} /* (17, 16, 8) {real, imag} */,
  {32'h3d5e3a04, 32'hbd324f18} /* (17, 16, 7) {real, imag} */,
  {32'h3cf7555b, 32'h3d92685e} /* (17, 16, 6) {real, imag} */,
  {32'hbe9b584b, 32'hbe32e98c} /* (17, 16, 5) {real, imag} */,
  {32'h3e96f416, 32'hbc3cea8c} /* (17, 16, 4) {real, imag} */,
  {32'h3e200772, 32'h3e1f8f7a} /* (17, 16, 3) {real, imag} */,
  {32'hbf9100b0, 32'hbe1814f8} /* (17, 16, 2) {real, imag} */,
  {32'h4014a63e, 32'h3e23f8b0} /* (17, 16, 1) {real, imag} */,
  {32'h3fcb3a74, 32'h00000000} /* (17, 16, 0) {real, imag} */,
  {32'h400ea75f, 32'hbc87e170} /* (17, 15, 31) {real, imag} */,
  {32'hbf86ffc0, 32'h3e62f834} /* (17, 15, 30) {real, imag} */,
  {32'h3df88c69, 32'hbdd297d8} /* (17, 15, 29) {real, imag} */,
  {32'h3e48271a, 32'h3d749e92} /* (17, 15, 28) {real, imag} */,
  {32'hbea66c2f, 32'h3e851564} /* (17, 15, 27) {real, imag} */,
  {32'hbd35874c, 32'hbe5e4ed9} /* (17, 15, 26) {real, imag} */,
  {32'h3dcb0b65, 32'hbbcefb9c} /* (17, 15, 25) {real, imag} */,
  {32'hbe1d26be, 32'h3dad16cb} /* (17, 15, 24) {real, imag} */,
  {32'hbda3a69a, 32'hbd1b1902} /* (17, 15, 23) {real, imag} */,
  {32'h3d92d136, 32'hbb1fbb30} /* (17, 15, 22) {real, imag} */,
  {32'h3cb3ed22, 32'h3dcc079f} /* (17, 15, 21) {real, imag} */,
  {32'h3d87f0d5, 32'hbd0e0343} /* (17, 15, 20) {real, imag} */,
  {32'h3c3d7f78, 32'hbd14405f} /* (17, 15, 19) {real, imag} */,
  {32'h3c8e7a8b, 32'h3cbe4121} /* (17, 15, 18) {real, imag} */,
  {32'hbb2eca72, 32'hbdb31a04} /* (17, 15, 17) {real, imag} */,
  {32'h3ce6000b, 32'h00000000} /* (17, 15, 16) {real, imag} */,
  {32'hbb2eca72, 32'h3db31a04} /* (17, 15, 15) {real, imag} */,
  {32'h3c8e7a8b, 32'hbcbe4121} /* (17, 15, 14) {real, imag} */,
  {32'h3c3d7f78, 32'h3d14405f} /* (17, 15, 13) {real, imag} */,
  {32'h3d87f0d5, 32'h3d0e0343} /* (17, 15, 12) {real, imag} */,
  {32'h3cb3ed22, 32'hbdcc079f} /* (17, 15, 11) {real, imag} */,
  {32'h3d92d136, 32'h3b1fbb30} /* (17, 15, 10) {real, imag} */,
  {32'hbda3a69a, 32'h3d1b1902} /* (17, 15, 9) {real, imag} */,
  {32'hbe1d26be, 32'hbdad16cb} /* (17, 15, 8) {real, imag} */,
  {32'h3dcb0b65, 32'h3bcefb9c} /* (17, 15, 7) {real, imag} */,
  {32'hbd35874c, 32'h3e5e4ed9} /* (17, 15, 6) {real, imag} */,
  {32'hbea66c2f, 32'hbe851564} /* (17, 15, 5) {real, imag} */,
  {32'h3e48271a, 32'hbd749e92} /* (17, 15, 4) {real, imag} */,
  {32'h3df88c69, 32'h3dd297d8} /* (17, 15, 3) {real, imag} */,
  {32'hbf86ffc0, 32'hbe62f834} /* (17, 15, 2) {real, imag} */,
  {32'h400ea75f, 32'h3c87e170} /* (17, 15, 1) {real, imag} */,
  {32'h3fdc9a3e, 32'h00000000} /* (17, 15, 0) {real, imag} */,
  {32'h40060e09, 32'h3c675e60} /* (17, 14, 31) {real, imag} */,
  {32'hbf6b83c1, 32'h3e0ace8a} /* (17, 14, 30) {real, imag} */,
  {32'h3e0e95c6, 32'hbd0ac680} /* (17, 14, 29) {real, imag} */,
  {32'h3dd08e54, 32'h3d7feb28} /* (17, 14, 28) {real, imag} */,
  {32'hbed188da, 32'h3e6180f6} /* (17, 14, 27) {real, imag} */,
  {32'h3d8b9022, 32'h3d8ee846} /* (17, 14, 26) {real, imag} */,
  {32'hbda3a4bf, 32'hbd03e594} /* (17, 14, 25) {real, imag} */,
  {32'hbd453995, 32'h3dd3e9e1} /* (17, 14, 24) {real, imag} */,
  {32'h3d944fde, 32'hbd3e8674} /* (17, 14, 23) {real, imag} */,
  {32'h3d42bd95, 32'h3d76de14} /* (17, 14, 22) {real, imag} */,
  {32'h3c9ac0ab, 32'h3d2d0158} /* (17, 14, 21) {real, imag} */,
  {32'hbd657df4, 32'hbd1fc802} /* (17, 14, 20) {real, imag} */,
  {32'h3cc3be10, 32'h3bdd90a8} /* (17, 14, 19) {real, imag} */,
  {32'hbd17c259, 32'hbe0aafae} /* (17, 14, 18) {real, imag} */,
  {32'h3c3102e8, 32'h3c9367fc} /* (17, 14, 17) {real, imag} */,
  {32'hbd4cfe06, 32'h00000000} /* (17, 14, 16) {real, imag} */,
  {32'h3c3102e8, 32'hbc9367fc} /* (17, 14, 15) {real, imag} */,
  {32'hbd17c259, 32'h3e0aafae} /* (17, 14, 14) {real, imag} */,
  {32'h3cc3be10, 32'hbbdd90a8} /* (17, 14, 13) {real, imag} */,
  {32'hbd657df4, 32'h3d1fc802} /* (17, 14, 12) {real, imag} */,
  {32'h3c9ac0ab, 32'hbd2d0158} /* (17, 14, 11) {real, imag} */,
  {32'h3d42bd95, 32'hbd76de14} /* (17, 14, 10) {real, imag} */,
  {32'h3d944fde, 32'h3d3e8674} /* (17, 14, 9) {real, imag} */,
  {32'hbd453995, 32'hbdd3e9e1} /* (17, 14, 8) {real, imag} */,
  {32'hbda3a4bf, 32'h3d03e594} /* (17, 14, 7) {real, imag} */,
  {32'h3d8b9022, 32'hbd8ee846} /* (17, 14, 6) {real, imag} */,
  {32'hbed188da, 32'hbe6180f6} /* (17, 14, 5) {real, imag} */,
  {32'h3dd08e54, 32'hbd7feb28} /* (17, 14, 4) {real, imag} */,
  {32'h3e0e95c6, 32'h3d0ac680} /* (17, 14, 3) {real, imag} */,
  {32'hbf6b83c1, 32'hbe0ace8a} /* (17, 14, 2) {real, imag} */,
  {32'h40060e09, 32'hbc675e60} /* (17, 14, 1) {real, imag} */,
  {32'h3fcd56ea, 32'h00000000} /* (17, 14, 0) {real, imag} */,
  {32'h3fdc9050, 32'h3e2805d2} /* (17, 13, 31) {real, imag} */,
  {32'hbf6a938e, 32'h3e3a1395} /* (17, 13, 30) {real, imag} */,
  {32'h3e66a8e5, 32'hbdf555e6} /* (17, 13, 29) {real, imag} */,
  {32'h3d263f90, 32'h3d79aed7} /* (17, 13, 28) {real, imag} */,
  {32'hbe6e105b, 32'h3e559fac} /* (17, 13, 27) {real, imag} */,
  {32'hbbf177d8, 32'hbb339758} /* (17, 13, 26) {real, imag} */,
  {32'hbdbe5054, 32'hbd514b58} /* (17, 13, 25) {real, imag} */,
  {32'h3d7a6e74, 32'h3dbb07aa} /* (17, 13, 24) {real, imag} */,
  {32'h3d4a9b1c, 32'h3cdfc264} /* (17, 13, 23) {real, imag} */,
  {32'h3d1eeae3, 32'hbcf69f17} /* (17, 13, 22) {real, imag} */,
  {32'hbaf56b40, 32'hbd5a279b} /* (17, 13, 21) {real, imag} */,
  {32'hbd0a5788, 32'hbd2aad40} /* (17, 13, 20) {real, imag} */,
  {32'h3d3c3cff, 32'h3c0fc7f2} /* (17, 13, 19) {real, imag} */,
  {32'hbc2f3864, 32'hbd2bc2b6} /* (17, 13, 18) {real, imag} */,
  {32'h3c2fd1dc, 32'hbb9302b0} /* (17, 13, 17) {real, imag} */,
  {32'h3df5c082, 32'h00000000} /* (17, 13, 16) {real, imag} */,
  {32'h3c2fd1dc, 32'h3b9302b0} /* (17, 13, 15) {real, imag} */,
  {32'hbc2f3864, 32'h3d2bc2b6} /* (17, 13, 14) {real, imag} */,
  {32'h3d3c3cff, 32'hbc0fc7f2} /* (17, 13, 13) {real, imag} */,
  {32'hbd0a5788, 32'h3d2aad40} /* (17, 13, 12) {real, imag} */,
  {32'hbaf56b40, 32'h3d5a279b} /* (17, 13, 11) {real, imag} */,
  {32'h3d1eeae3, 32'h3cf69f17} /* (17, 13, 10) {real, imag} */,
  {32'h3d4a9b1c, 32'hbcdfc264} /* (17, 13, 9) {real, imag} */,
  {32'h3d7a6e74, 32'hbdbb07aa} /* (17, 13, 8) {real, imag} */,
  {32'hbdbe5054, 32'h3d514b58} /* (17, 13, 7) {real, imag} */,
  {32'hbbf177d8, 32'h3b339758} /* (17, 13, 6) {real, imag} */,
  {32'hbe6e105b, 32'hbe559fac} /* (17, 13, 5) {real, imag} */,
  {32'h3d263f90, 32'hbd79aed7} /* (17, 13, 4) {real, imag} */,
  {32'h3e66a8e5, 32'h3df555e6} /* (17, 13, 3) {real, imag} */,
  {32'hbf6a938e, 32'hbe3a1395} /* (17, 13, 2) {real, imag} */,
  {32'h3fdc9050, 32'hbe2805d2} /* (17, 13, 1) {real, imag} */,
  {32'h3fcdb3b6, 32'h00000000} /* (17, 13, 0) {real, imag} */,
  {32'h3fb52806, 32'h3e268d5e} /* (17, 12, 31) {real, imag} */,
  {32'hbf4b3daa, 32'h3e325f06} /* (17, 12, 30) {real, imag} */,
  {32'h3e78ed10, 32'h3cb090cc} /* (17, 12, 29) {real, imag} */,
  {32'h3e00ff42, 32'h3c4da128} /* (17, 12, 28) {real, imag} */,
  {32'hbe2b0bfa, 32'h3ceb0897} /* (17, 12, 27) {real, imag} */,
  {32'hbdc3ff6b, 32'h3d4a60ed} /* (17, 12, 26) {real, imag} */,
  {32'hbd587063, 32'hbe26cead} /* (17, 12, 25) {real, imag} */,
  {32'hbe03dffc, 32'h3e0317d0} /* (17, 12, 24) {real, imag} */,
  {32'h3daaef27, 32'hbd30bca4} /* (17, 12, 23) {real, imag} */,
  {32'h3c78434a, 32'hbd049a34} /* (17, 12, 22) {real, imag} */,
  {32'hbd28556e, 32'h3a4f6f80} /* (17, 12, 21) {real, imag} */,
  {32'hbba63054, 32'h3b9bb10c} /* (17, 12, 20) {real, imag} */,
  {32'h3d00c4ac, 32'h3ca86432} /* (17, 12, 19) {real, imag} */,
  {32'hbd812509, 32'hbcf98d34} /* (17, 12, 18) {real, imag} */,
  {32'hbd546872, 32'h3d7a6946} /* (17, 12, 17) {real, imag} */,
  {32'h3c06ebbe, 32'h00000000} /* (17, 12, 16) {real, imag} */,
  {32'hbd546872, 32'hbd7a6946} /* (17, 12, 15) {real, imag} */,
  {32'hbd812509, 32'h3cf98d34} /* (17, 12, 14) {real, imag} */,
  {32'h3d00c4ac, 32'hbca86432} /* (17, 12, 13) {real, imag} */,
  {32'hbba63054, 32'hbb9bb10c} /* (17, 12, 12) {real, imag} */,
  {32'hbd28556e, 32'hba4f6f80} /* (17, 12, 11) {real, imag} */,
  {32'h3c78434a, 32'h3d049a34} /* (17, 12, 10) {real, imag} */,
  {32'h3daaef27, 32'h3d30bca4} /* (17, 12, 9) {real, imag} */,
  {32'hbe03dffc, 32'hbe0317d0} /* (17, 12, 8) {real, imag} */,
  {32'hbd587063, 32'h3e26cead} /* (17, 12, 7) {real, imag} */,
  {32'hbdc3ff6b, 32'hbd4a60ed} /* (17, 12, 6) {real, imag} */,
  {32'hbe2b0bfa, 32'hbceb0897} /* (17, 12, 5) {real, imag} */,
  {32'h3e00ff42, 32'hbc4da128} /* (17, 12, 4) {real, imag} */,
  {32'h3e78ed10, 32'hbcb090cc} /* (17, 12, 3) {real, imag} */,
  {32'hbf4b3daa, 32'hbe325f06} /* (17, 12, 2) {real, imag} */,
  {32'h3fb52806, 32'hbe268d5e} /* (17, 12, 1) {real, imag} */,
  {32'h3fb1be64, 32'h00000000} /* (17, 12, 0) {real, imag} */,
  {32'h3f45eac7, 32'h3ea46d74} /* (17, 11, 31) {real, imag} */,
  {32'hbee30656, 32'h3e4a42c8} /* (17, 11, 30) {real, imag} */,
  {32'h3e31d2ff, 32'h3c97c451} /* (17, 11, 29) {real, imag} */,
  {32'h3d12e20e, 32'hbda29a8e} /* (17, 11, 28) {real, imag} */,
  {32'hbd930801, 32'h3de7cc2b} /* (17, 11, 27) {real, imag} */,
  {32'hbd3e3e2c, 32'hbc87db8a} /* (17, 11, 26) {real, imag} */,
  {32'h3d644ed3, 32'h3c0e8db0} /* (17, 11, 25) {real, imag} */,
  {32'hbd9f4054, 32'h3e8d8e11} /* (17, 11, 24) {real, imag} */,
  {32'h3d478408, 32'h3c7223ec} /* (17, 11, 23) {real, imag} */,
  {32'hbd998ab6, 32'h3d8a5b3e} /* (17, 11, 22) {real, imag} */,
  {32'h3d64037b, 32'hbd86188a} /* (17, 11, 21) {real, imag} */,
  {32'hbc7f7578, 32'h3c7012d9} /* (17, 11, 20) {real, imag} */,
  {32'h3bf6ce30, 32'h3c4ceae8} /* (17, 11, 19) {real, imag} */,
  {32'h3d8f4514, 32'h3d5267b4} /* (17, 11, 18) {real, imag} */,
  {32'hbce3cf1c, 32'hbcc265fd} /* (17, 11, 17) {real, imag} */,
  {32'hbe2d088b, 32'h00000000} /* (17, 11, 16) {real, imag} */,
  {32'hbce3cf1c, 32'h3cc265fd} /* (17, 11, 15) {real, imag} */,
  {32'h3d8f4514, 32'hbd5267b4} /* (17, 11, 14) {real, imag} */,
  {32'h3bf6ce30, 32'hbc4ceae8} /* (17, 11, 13) {real, imag} */,
  {32'hbc7f7578, 32'hbc7012d9} /* (17, 11, 12) {real, imag} */,
  {32'h3d64037b, 32'h3d86188a} /* (17, 11, 11) {real, imag} */,
  {32'hbd998ab6, 32'hbd8a5b3e} /* (17, 11, 10) {real, imag} */,
  {32'h3d478408, 32'hbc7223ec} /* (17, 11, 9) {real, imag} */,
  {32'hbd9f4054, 32'hbe8d8e11} /* (17, 11, 8) {real, imag} */,
  {32'h3d644ed3, 32'hbc0e8db0} /* (17, 11, 7) {real, imag} */,
  {32'hbd3e3e2c, 32'h3c87db8a} /* (17, 11, 6) {real, imag} */,
  {32'hbd930801, 32'hbde7cc2b} /* (17, 11, 5) {real, imag} */,
  {32'h3d12e20e, 32'h3da29a8e} /* (17, 11, 4) {real, imag} */,
  {32'h3e31d2ff, 32'hbc97c451} /* (17, 11, 3) {real, imag} */,
  {32'hbee30656, 32'hbe4a42c8} /* (17, 11, 2) {real, imag} */,
  {32'h3f45eac7, 32'hbea46d74} /* (17, 11, 1) {real, imag} */,
  {32'h3f498ff5, 32'h00000000} /* (17, 11, 0) {real, imag} */,
  {32'hbf2abf33, 32'h3f04f355} /* (17, 10, 31) {real, imag} */,
  {32'h3da17488, 32'hbd281cdd} /* (17, 10, 30) {real, imag} */,
  {32'h3da5acdc, 32'h3df3c40e} /* (17, 10, 29) {real, imag} */,
  {32'hbdc86064, 32'hbdac9e55} /* (17, 10, 28) {real, imag} */,
  {32'h3d0b9c1c, 32'hbb8e2390} /* (17, 10, 27) {real, imag} */,
  {32'h3d576b46, 32'hbb95d880} /* (17, 10, 26) {real, imag} */,
  {32'h3d097e23, 32'h3b925464} /* (17, 10, 25) {real, imag} */,
  {32'h3e1b5986, 32'hbd1784ba} /* (17, 10, 24) {real, imag} */,
  {32'hbd2d593c, 32'hbc32da34} /* (17, 10, 23) {real, imag} */,
  {32'hbca043d6, 32'h3c4bed90} /* (17, 10, 22) {real, imag} */,
  {32'hbbc6cad0, 32'h3d52033b} /* (17, 10, 21) {real, imag} */,
  {32'hbdb09d6e, 32'h3d2cc130} /* (17, 10, 20) {real, imag} */,
  {32'h3d214e05, 32'h3dd6a1b4} /* (17, 10, 19) {real, imag} */,
  {32'hbd8a42d9, 32'h3d2897be} /* (17, 10, 18) {real, imag} */,
  {32'hbd05b654, 32'h3cfbaba2} /* (17, 10, 17) {real, imag} */,
  {32'hbcf125fa, 32'h00000000} /* (17, 10, 16) {real, imag} */,
  {32'hbd05b654, 32'hbcfbaba2} /* (17, 10, 15) {real, imag} */,
  {32'hbd8a42d9, 32'hbd2897be} /* (17, 10, 14) {real, imag} */,
  {32'h3d214e05, 32'hbdd6a1b4} /* (17, 10, 13) {real, imag} */,
  {32'hbdb09d6e, 32'hbd2cc130} /* (17, 10, 12) {real, imag} */,
  {32'hbbc6cad0, 32'hbd52033b} /* (17, 10, 11) {real, imag} */,
  {32'hbca043d6, 32'hbc4bed90} /* (17, 10, 10) {real, imag} */,
  {32'hbd2d593c, 32'h3c32da34} /* (17, 10, 9) {real, imag} */,
  {32'h3e1b5986, 32'h3d1784ba} /* (17, 10, 8) {real, imag} */,
  {32'h3d097e23, 32'hbb925464} /* (17, 10, 7) {real, imag} */,
  {32'h3d576b46, 32'h3b95d880} /* (17, 10, 6) {real, imag} */,
  {32'h3d0b9c1c, 32'h3b8e2390} /* (17, 10, 5) {real, imag} */,
  {32'hbdc86064, 32'h3dac9e55} /* (17, 10, 4) {real, imag} */,
  {32'h3da5acdc, 32'hbdf3c40e} /* (17, 10, 3) {real, imag} */,
  {32'h3da17488, 32'h3d281cdd} /* (17, 10, 2) {real, imag} */,
  {32'hbf2abf33, 32'hbf04f355} /* (17, 10, 1) {real, imag} */,
  {32'hbe876446, 32'h00000000} /* (17, 10, 0) {real, imag} */,
  {32'hbfc1ac54, 32'h3f146a28} /* (17, 9, 31) {real, imag} */,
  {32'h3f09e449, 32'hbe1f7fa8} /* (17, 9, 30) {real, imag} */,
  {32'hbde425ac, 32'h3dea709e} /* (17, 9, 29) {real, imag} */,
  {32'h3c13f150, 32'h3c9fb9aa} /* (17, 9, 28) {real, imag} */,
  {32'h3cba7e68, 32'h3c107768} /* (17, 9, 27) {real, imag} */,
  {32'hbdf58972, 32'hbc948a80} /* (17, 9, 26) {real, imag} */,
  {32'hbcc0cda2, 32'h3dbb240c} /* (17, 9, 25) {real, imag} */,
  {32'h3d798ac2, 32'hbda1af17} /* (17, 9, 24) {real, imag} */,
  {32'hbbf8f8b0, 32'hbd0eac36} /* (17, 9, 23) {real, imag} */,
  {32'h3d573d8b, 32'h3caebb65} /* (17, 9, 22) {real, imag} */,
  {32'h3da1a650, 32'hbdcb45c0} /* (17, 9, 21) {real, imag} */,
  {32'hbd7e28b9, 32'h3b22a71c} /* (17, 9, 20) {real, imag} */,
  {32'hbc2da776, 32'h3d4c529a} /* (17, 9, 19) {real, imag} */,
  {32'hb9ac4540, 32'hbd997b07} /* (17, 9, 18) {real, imag} */,
  {32'h3c1d10d2, 32'hbd954d4c} /* (17, 9, 17) {real, imag} */,
  {32'h3bf6110c, 32'h00000000} /* (17, 9, 16) {real, imag} */,
  {32'h3c1d10d2, 32'h3d954d4c} /* (17, 9, 15) {real, imag} */,
  {32'hb9ac4540, 32'h3d997b07} /* (17, 9, 14) {real, imag} */,
  {32'hbc2da776, 32'hbd4c529a} /* (17, 9, 13) {real, imag} */,
  {32'hbd7e28b9, 32'hbb22a71c} /* (17, 9, 12) {real, imag} */,
  {32'h3da1a650, 32'h3dcb45c0} /* (17, 9, 11) {real, imag} */,
  {32'h3d573d8b, 32'hbcaebb65} /* (17, 9, 10) {real, imag} */,
  {32'hbbf8f8b0, 32'h3d0eac36} /* (17, 9, 9) {real, imag} */,
  {32'h3d798ac2, 32'h3da1af17} /* (17, 9, 8) {real, imag} */,
  {32'hbcc0cda2, 32'hbdbb240c} /* (17, 9, 7) {real, imag} */,
  {32'hbdf58972, 32'h3c948a80} /* (17, 9, 6) {real, imag} */,
  {32'h3cba7e68, 32'hbc107768} /* (17, 9, 5) {real, imag} */,
  {32'h3c13f150, 32'hbc9fb9aa} /* (17, 9, 4) {real, imag} */,
  {32'hbde425ac, 32'hbdea709e} /* (17, 9, 3) {real, imag} */,
  {32'h3f09e449, 32'h3e1f7fa8} /* (17, 9, 2) {real, imag} */,
  {32'hbfc1ac54, 32'hbf146a28} /* (17, 9, 1) {real, imag} */,
  {32'hbf716984, 32'h00000000} /* (17, 9, 0) {real, imag} */,
  {32'hc001ec33, 32'h3f39d1de} /* (17, 8, 31) {real, imag} */,
  {32'h3f2a9b16, 32'hbe89b6ce} /* (17, 8, 30) {real, imag} */,
  {32'hbddac762, 32'h3db32741} /* (17, 8, 29) {real, imag} */,
  {32'h3d1e9cf0, 32'hbdaa3fdd} /* (17, 8, 28) {real, imag} */,
  {32'h3d55e068, 32'h3c30e9b8} /* (17, 8, 27) {real, imag} */,
  {32'hbd07fd9c, 32'h3de208fc} /* (17, 8, 26) {real, imag} */,
  {32'hbe23766c, 32'h3d7d7860} /* (17, 8, 25) {real, imag} */,
  {32'h3d9d3498, 32'hbd466197} /* (17, 8, 24) {real, imag} */,
  {32'hbcace50d, 32'hbd0887bc} /* (17, 8, 23) {real, imag} */,
  {32'h3e220ca4, 32'hbd9c2a35} /* (17, 8, 22) {real, imag} */,
  {32'h3d034afa, 32'h3db1bf94} /* (17, 8, 21) {real, imag} */,
  {32'h3d8fb01b, 32'h3c15e1c8} /* (17, 8, 20) {real, imag} */,
  {32'hbce4111c, 32'hbd194b44} /* (17, 8, 19) {real, imag} */,
  {32'h3c87a5f4, 32'h3c7d0070} /* (17, 8, 18) {real, imag} */,
  {32'hbdba7651, 32'hbcaff336} /* (17, 8, 17) {real, imag} */,
  {32'h3d5d4780, 32'h00000000} /* (17, 8, 16) {real, imag} */,
  {32'hbdba7651, 32'h3caff336} /* (17, 8, 15) {real, imag} */,
  {32'h3c87a5f4, 32'hbc7d0070} /* (17, 8, 14) {real, imag} */,
  {32'hbce4111c, 32'h3d194b44} /* (17, 8, 13) {real, imag} */,
  {32'h3d8fb01b, 32'hbc15e1c8} /* (17, 8, 12) {real, imag} */,
  {32'h3d034afa, 32'hbdb1bf94} /* (17, 8, 11) {real, imag} */,
  {32'h3e220ca4, 32'h3d9c2a35} /* (17, 8, 10) {real, imag} */,
  {32'hbcace50d, 32'h3d0887bc} /* (17, 8, 9) {real, imag} */,
  {32'h3d9d3498, 32'h3d466197} /* (17, 8, 8) {real, imag} */,
  {32'hbe23766c, 32'hbd7d7860} /* (17, 8, 7) {real, imag} */,
  {32'hbd07fd9c, 32'hbde208fc} /* (17, 8, 6) {real, imag} */,
  {32'h3d55e068, 32'hbc30e9b8} /* (17, 8, 5) {real, imag} */,
  {32'h3d1e9cf0, 32'h3daa3fdd} /* (17, 8, 4) {real, imag} */,
  {32'hbddac762, 32'hbdb32741} /* (17, 8, 3) {real, imag} */,
  {32'h3f2a9b16, 32'h3e89b6ce} /* (17, 8, 2) {real, imag} */,
  {32'hc001ec33, 32'hbf39d1de} /* (17, 8, 1) {real, imag} */,
  {32'hbfc992a0, 32'h00000000} /* (17, 8, 0) {real, imag} */,
  {32'hc011af73, 32'h3f7b6594} /* (17, 7, 31) {real, imag} */,
  {32'h3f265415, 32'hbec11770} /* (17, 7, 30) {real, imag} */,
  {32'hbd75c959, 32'h3d6fe26a} /* (17, 7, 29) {real, imag} */,
  {32'hbdd68f79, 32'h3dfcdeb2} /* (17, 7, 28) {real, imag} */,
  {32'h3e624e79, 32'hbdbf5c15} /* (17, 7, 27) {real, imag} */,
  {32'h3caa2fea, 32'h3e332cde} /* (17, 7, 26) {real, imag} */,
  {32'hbd37d7bc, 32'hbb327200} /* (17, 7, 25) {real, imag} */,
  {32'h3de30000, 32'hbc9faf70} /* (17, 7, 24) {real, imag} */,
  {32'h3e1cf546, 32'h3ccacbda} /* (17, 7, 23) {real, imag} */,
  {32'hbd3ec6d5, 32'hbd87f47a} /* (17, 7, 22) {real, imag} */,
  {32'hbcaa9380, 32'h3d2f33a2} /* (17, 7, 21) {real, imag} */,
  {32'h3cb7fb5a, 32'h3cd39ca2} /* (17, 7, 20) {real, imag} */,
  {32'h3d05a654, 32'hbd877c39} /* (17, 7, 19) {real, imag} */,
  {32'h3d478d77, 32'hbb903d30} /* (17, 7, 18) {real, imag} */,
  {32'hbbed25e9, 32'h3da575e5} /* (17, 7, 17) {real, imag} */,
  {32'h3dc1c11c, 32'h00000000} /* (17, 7, 16) {real, imag} */,
  {32'hbbed25e9, 32'hbda575e5} /* (17, 7, 15) {real, imag} */,
  {32'h3d478d77, 32'h3b903d30} /* (17, 7, 14) {real, imag} */,
  {32'h3d05a654, 32'h3d877c39} /* (17, 7, 13) {real, imag} */,
  {32'h3cb7fb5a, 32'hbcd39ca2} /* (17, 7, 12) {real, imag} */,
  {32'hbcaa9380, 32'hbd2f33a2} /* (17, 7, 11) {real, imag} */,
  {32'hbd3ec6d5, 32'h3d87f47a} /* (17, 7, 10) {real, imag} */,
  {32'h3e1cf546, 32'hbccacbda} /* (17, 7, 9) {real, imag} */,
  {32'h3de30000, 32'h3c9faf70} /* (17, 7, 8) {real, imag} */,
  {32'hbd37d7bc, 32'h3b327200} /* (17, 7, 7) {real, imag} */,
  {32'h3caa2fea, 32'hbe332cde} /* (17, 7, 6) {real, imag} */,
  {32'h3e624e79, 32'h3dbf5c15} /* (17, 7, 5) {real, imag} */,
  {32'hbdd68f79, 32'hbdfcdeb2} /* (17, 7, 4) {real, imag} */,
  {32'hbd75c959, 32'hbd6fe26a} /* (17, 7, 3) {real, imag} */,
  {32'h3f265415, 32'h3ec11770} /* (17, 7, 2) {real, imag} */,
  {32'hc011af73, 32'hbf7b6594} /* (17, 7, 1) {real, imag} */,
  {32'hc00588ca, 32'h00000000} /* (17, 7, 0) {real, imag} */,
  {32'hc01250b1, 32'h3f9bcfa8} /* (17, 6, 31) {real, imag} */,
  {32'h3f1716c9, 32'hbed22a1e} /* (17, 6, 30) {real, imag} */,
  {32'hbdc2013a, 32'h3c9308cb} /* (17, 6, 29) {real, imag} */,
  {32'hbdb0bf4a, 32'h3d405354} /* (17, 6, 28) {real, imag} */,
  {32'h3e7bbe72, 32'h3c0f35c2} /* (17, 6, 27) {real, imag} */,
  {32'h3e07894c, 32'h3dcf6074} /* (17, 6, 26) {real, imag} */,
  {32'h3b513f98, 32'h3c8668f3} /* (17, 6, 25) {real, imag} */,
  {32'h3d397fde, 32'hbe2ccfe1} /* (17, 6, 24) {real, imag} */,
  {32'hbcaf5e02, 32'h3d227b78} /* (17, 6, 23) {real, imag} */,
  {32'h3bd9e1e2, 32'h3d65288e} /* (17, 6, 22) {real, imag} */,
  {32'hbca05fda, 32'hbe1d1f4d} /* (17, 6, 21) {real, imag} */,
  {32'hbbe0d79c, 32'hbd66b78a} /* (17, 6, 20) {real, imag} */,
  {32'h3dcea7da, 32'h3d4c9b5c} /* (17, 6, 19) {real, imag} */,
  {32'hb9cdd580, 32'h3bbd7b3c} /* (17, 6, 18) {real, imag} */,
  {32'hbd2d5138, 32'h3930eb80} /* (17, 6, 17) {real, imag} */,
  {32'h3c65e090, 32'h00000000} /* (17, 6, 16) {real, imag} */,
  {32'hbd2d5138, 32'hb930eb80} /* (17, 6, 15) {real, imag} */,
  {32'hb9cdd580, 32'hbbbd7b3c} /* (17, 6, 14) {real, imag} */,
  {32'h3dcea7da, 32'hbd4c9b5c} /* (17, 6, 13) {real, imag} */,
  {32'hbbe0d79c, 32'h3d66b78a} /* (17, 6, 12) {real, imag} */,
  {32'hbca05fda, 32'h3e1d1f4d} /* (17, 6, 11) {real, imag} */,
  {32'h3bd9e1e2, 32'hbd65288e} /* (17, 6, 10) {real, imag} */,
  {32'hbcaf5e02, 32'hbd227b78} /* (17, 6, 9) {real, imag} */,
  {32'h3d397fde, 32'h3e2ccfe1} /* (17, 6, 8) {real, imag} */,
  {32'h3b513f98, 32'hbc8668f3} /* (17, 6, 7) {real, imag} */,
  {32'h3e07894c, 32'hbdcf6074} /* (17, 6, 6) {real, imag} */,
  {32'h3e7bbe72, 32'hbc0f35c2} /* (17, 6, 5) {real, imag} */,
  {32'hbdb0bf4a, 32'hbd405354} /* (17, 6, 4) {real, imag} */,
  {32'hbdc2013a, 32'hbc9308cb} /* (17, 6, 3) {real, imag} */,
  {32'h3f1716c9, 32'h3ed22a1e} /* (17, 6, 2) {real, imag} */,
  {32'hc01250b1, 32'hbf9bcfa8} /* (17, 6, 1) {real, imag} */,
  {32'hc0139320, 32'h00000000} /* (17, 6, 0) {real, imag} */,
  {32'hbffb552a, 32'h3fd553d6} /* (17, 5, 31) {real, imag} */,
  {32'h3de1bf04, 32'hbf201d84} /* (17, 5, 30) {real, imag} */,
  {32'hbd2352c8, 32'h3d2e8af0} /* (17, 5, 29) {real, imag} */,
  {32'h3e28a59d, 32'hbc3b53b0} /* (17, 5, 28) {real, imag} */,
  {32'h3de9cc16, 32'h3d2b1b84} /* (17, 5, 27) {real, imag} */,
  {32'h3d9d635b, 32'h3dce357b} /* (17, 5, 26) {real, imag} */,
  {32'h3d3b2a19, 32'hbd4703ea} /* (17, 5, 25) {real, imag} */,
  {32'hbda65265, 32'hbded30c9} /* (17, 5, 24) {real, imag} */,
  {32'hbc1d1530, 32'hbc36c06c} /* (17, 5, 23) {real, imag} */,
  {32'hbbf35020, 32'h3db72697} /* (17, 5, 22) {real, imag} */,
  {32'h3d881374, 32'hbd5b4cfa} /* (17, 5, 21) {real, imag} */,
  {32'h3b822628, 32'h3c1f79ea} /* (17, 5, 20) {real, imag} */,
  {32'hbd25c5e9, 32'h3d8ae2d6} /* (17, 5, 19) {real, imag} */,
  {32'hbd152024, 32'h3d20ec48} /* (17, 5, 18) {real, imag} */,
  {32'h3c56a7dd, 32'h3d4a653a} /* (17, 5, 17) {real, imag} */,
  {32'hbd12c157, 32'h00000000} /* (17, 5, 16) {real, imag} */,
  {32'h3c56a7dd, 32'hbd4a653a} /* (17, 5, 15) {real, imag} */,
  {32'hbd152024, 32'hbd20ec48} /* (17, 5, 14) {real, imag} */,
  {32'hbd25c5e9, 32'hbd8ae2d6} /* (17, 5, 13) {real, imag} */,
  {32'h3b822628, 32'hbc1f79ea} /* (17, 5, 12) {real, imag} */,
  {32'h3d881374, 32'h3d5b4cfa} /* (17, 5, 11) {real, imag} */,
  {32'hbbf35020, 32'hbdb72697} /* (17, 5, 10) {real, imag} */,
  {32'hbc1d1530, 32'h3c36c06c} /* (17, 5, 9) {real, imag} */,
  {32'hbda65265, 32'h3ded30c9} /* (17, 5, 8) {real, imag} */,
  {32'h3d3b2a19, 32'h3d4703ea} /* (17, 5, 7) {real, imag} */,
  {32'h3d9d635b, 32'hbdce357b} /* (17, 5, 6) {real, imag} */,
  {32'h3de9cc16, 32'hbd2b1b84} /* (17, 5, 5) {real, imag} */,
  {32'h3e28a59d, 32'h3c3b53b0} /* (17, 5, 4) {real, imag} */,
  {32'hbd2352c8, 32'hbd2e8af0} /* (17, 5, 3) {real, imag} */,
  {32'h3de1bf04, 32'h3f201d84} /* (17, 5, 2) {real, imag} */,
  {32'hbffb552a, 32'hbfd553d6} /* (17, 5, 1) {real, imag} */,
  {32'hc01cb4bc, 32'h00000000} /* (17, 5, 0) {real, imag} */,
  {32'hbfdab882, 32'h3ffff7d5} /* (17, 4, 31) {real, imag} */,
  {32'hbe936a08, 32'hbf3dcaf5} /* (17, 4, 30) {real, imag} */,
  {32'h3d1f6f0e, 32'h3c3f044a} /* (17, 4, 29) {real, imag} */,
  {32'h3e8675be, 32'hbd7659f0} /* (17, 4, 28) {real, imag} */,
  {32'h3e57a466, 32'h3e50191b} /* (17, 4, 27) {real, imag} */,
  {32'hbdc347c8, 32'h3c7b7e1a} /* (17, 4, 26) {real, imag} */,
  {32'h3d17e6b3, 32'h3d064b8b} /* (17, 4, 25) {real, imag} */,
  {32'hbda9fc7e, 32'hbdbf31ef} /* (17, 4, 24) {real, imag} */,
  {32'h3d4b83fb, 32'h3ae2fbb0} /* (17, 4, 23) {real, imag} */,
  {32'hbd4a0ff2, 32'hbda953e1} /* (17, 4, 22) {real, imag} */,
  {32'hbafaabf0, 32'hbd380f8f} /* (17, 4, 21) {real, imag} */,
  {32'h3de8a025, 32'hbca96e1a} /* (17, 4, 20) {real, imag} */,
  {32'hbce62fe8, 32'h3d0fac7a} /* (17, 4, 19) {real, imag} */,
  {32'h3c4df0e0, 32'hbb8681f0} /* (17, 4, 18) {real, imag} */,
  {32'hbd886e92, 32'h3d7a7ad2} /* (17, 4, 17) {real, imag} */,
  {32'h3d49ba34, 32'h00000000} /* (17, 4, 16) {real, imag} */,
  {32'hbd886e92, 32'hbd7a7ad2} /* (17, 4, 15) {real, imag} */,
  {32'h3c4df0e0, 32'h3b8681f0} /* (17, 4, 14) {real, imag} */,
  {32'hbce62fe8, 32'hbd0fac7a} /* (17, 4, 13) {real, imag} */,
  {32'h3de8a025, 32'h3ca96e1a} /* (17, 4, 12) {real, imag} */,
  {32'hbafaabf0, 32'h3d380f8f} /* (17, 4, 11) {real, imag} */,
  {32'hbd4a0ff2, 32'h3da953e1} /* (17, 4, 10) {real, imag} */,
  {32'h3d4b83fb, 32'hbae2fbb0} /* (17, 4, 9) {real, imag} */,
  {32'hbda9fc7e, 32'h3dbf31ef} /* (17, 4, 8) {real, imag} */,
  {32'h3d17e6b3, 32'hbd064b8b} /* (17, 4, 7) {real, imag} */,
  {32'hbdc347c8, 32'hbc7b7e1a} /* (17, 4, 6) {real, imag} */,
  {32'h3e57a466, 32'hbe50191b} /* (17, 4, 5) {real, imag} */,
  {32'h3e8675be, 32'h3d7659f0} /* (17, 4, 4) {real, imag} */,
  {32'h3d1f6f0e, 32'hbc3f044a} /* (17, 4, 3) {real, imag} */,
  {32'hbe936a08, 32'h3f3dcaf5} /* (17, 4, 2) {real, imag} */,
  {32'hbfdab882, 32'hbffff7d5} /* (17, 4, 1) {real, imag} */,
  {32'hc0158ece, 32'h00000000} /* (17, 4, 0) {real, imag} */,
  {32'hbfe0f38d, 32'h4011965f} /* (17, 3, 31) {real, imag} */,
  {32'hbead3484, 32'hbf718cae} /* (17, 3, 30) {real, imag} */,
  {32'h3e512bb7, 32'h3e3a35be} /* (17, 3, 29) {real, imag} */,
  {32'h3e4ce992, 32'hbe1374fc} /* (17, 3, 28) {real, imag} */,
  {32'h3e187c8c, 32'h3e988bda} /* (17, 3, 27) {real, imag} */,
  {32'h3d23331c, 32'hbd97d7cc} /* (17, 3, 26) {real, imag} */,
  {32'hbbc77178, 32'h3d8bdf7c} /* (17, 3, 25) {real, imag} */,
  {32'h3d90761d, 32'hbdfff03a} /* (17, 3, 24) {real, imag} */,
  {32'hba53b6c0, 32'hbd2bc019} /* (17, 3, 23) {real, imag} */,
  {32'h3b12bb30, 32'hbd97c268} /* (17, 3, 22) {real, imag} */,
  {32'h3c8fac80, 32'hbe237b58} /* (17, 3, 21) {real, imag} */,
  {32'hbcaa46b8, 32'h3c40cacf} /* (17, 3, 20) {real, imag} */,
  {32'hbccdf184, 32'h3c6c31aa} /* (17, 3, 19) {real, imag} */,
  {32'hbdf5c0ca, 32'h3c3e3965} /* (17, 3, 18) {real, imag} */,
  {32'h3d82d3e1, 32'hbcc47176} /* (17, 3, 17) {real, imag} */,
  {32'hbd97cee8, 32'h00000000} /* (17, 3, 16) {real, imag} */,
  {32'h3d82d3e1, 32'h3cc47176} /* (17, 3, 15) {real, imag} */,
  {32'hbdf5c0ca, 32'hbc3e3965} /* (17, 3, 14) {real, imag} */,
  {32'hbccdf184, 32'hbc6c31aa} /* (17, 3, 13) {real, imag} */,
  {32'hbcaa46b8, 32'hbc40cacf} /* (17, 3, 12) {real, imag} */,
  {32'h3c8fac80, 32'h3e237b58} /* (17, 3, 11) {real, imag} */,
  {32'h3b12bb30, 32'h3d97c268} /* (17, 3, 10) {real, imag} */,
  {32'hba53b6c0, 32'h3d2bc019} /* (17, 3, 9) {real, imag} */,
  {32'h3d90761d, 32'h3dfff03a} /* (17, 3, 8) {real, imag} */,
  {32'hbbc77178, 32'hbd8bdf7c} /* (17, 3, 7) {real, imag} */,
  {32'h3d23331c, 32'h3d97d7cc} /* (17, 3, 6) {real, imag} */,
  {32'h3e187c8c, 32'hbe988bda} /* (17, 3, 5) {real, imag} */,
  {32'h3e4ce992, 32'h3e1374fc} /* (17, 3, 4) {real, imag} */,
  {32'h3e512bb7, 32'hbe3a35be} /* (17, 3, 3) {real, imag} */,
  {32'hbead3484, 32'h3f718cae} /* (17, 3, 2) {real, imag} */,
  {32'hbfe0f38d, 32'hc011965f} /* (17, 3, 1) {real, imag} */,
  {32'hc013893a, 32'h00000000} /* (17, 3, 0) {real, imag} */,
  {32'hbfd14def, 32'h40071064} /* (17, 2, 31) {real, imag} */,
  {32'hbeb35f0e, 32'hbf71e9ba} /* (17, 2, 30) {real, imag} */,
  {32'h3e937a69, 32'h3e748ee4} /* (17, 2, 29) {real, imag} */,
  {32'h3c7a4100, 32'hbeb8ec6c} /* (17, 2, 28) {real, imag} */,
  {32'h3d9ecc7e, 32'h3e791de1} /* (17, 2, 27) {real, imag} */,
  {32'h3d7cbdb9, 32'hbdc81c10} /* (17, 2, 26) {real, imag} */,
  {32'hbd8607b5, 32'h3e0f4e9f} /* (17, 2, 25) {real, imag} */,
  {32'h3df93f04, 32'hbe199ea5} /* (17, 2, 24) {real, imag} */,
  {32'hbd64bb9c, 32'hbd945600} /* (17, 2, 23) {real, imag} */,
  {32'h3d17098d, 32'hbcb03a46} /* (17, 2, 22) {real, imag} */,
  {32'hbdbc9ef6, 32'hbdbbe582} /* (17, 2, 21) {real, imag} */,
  {32'h3d9f080e, 32'h3daca09e} /* (17, 2, 20) {real, imag} */,
  {32'hbcc9237e, 32'h3d39a0ec} /* (17, 2, 19) {real, imag} */,
  {32'hbce6254e, 32'hbd113a52} /* (17, 2, 18) {real, imag} */,
  {32'h3da8071e, 32'h3c5efe90} /* (17, 2, 17) {real, imag} */,
  {32'hbdfaf381, 32'h00000000} /* (17, 2, 16) {real, imag} */,
  {32'h3da8071e, 32'hbc5efe90} /* (17, 2, 15) {real, imag} */,
  {32'hbce6254e, 32'h3d113a52} /* (17, 2, 14) {real, imag} */,
  {32'hbcc9237e, 32'hbd39a0ec} /* (17, 2, 13) {real, imag} */,
  {32'h3d9f080e, 32'hbdaca09e} /* (17, 2, 12) {real, imag} */,
  {32'hbdbc9ef6, 32'h3dbbe582} /* (17, 2, 11) {real, imag} */,
  {32'h3d17098d, 32'h3cb03a46} /* (17, 2, 10) {real, imag} */,
  {32'hbd64bb9c, 32'h3d945600} /* (17, 2, 9) {real, imag} */,
  {32'h3df93f04, 32'h3e199ea5} /* (17, 2, 8) {real, imag} */,
  {32'hbd8607b5, 32'hbe0f4e9f} /* (17, 2, 7) {real, imag} */,
  {32'h3d7cbdb9, 32'h3dc81c10} /* (17, 2, 6) {real, imag} */,
  {32'h3d9ecc7e, 32'hbe791de1} /* (17, 2, 5) {real, imag} */,
  {32'h3c7a4100, 32'h3eb8ec6c} /* (17, 2, 4) {real, imag} */,
  {32'h3e937a69, 32'hbe748ee4} /* (17, 2, 3) {real, imag} */,
  {32'hbeb35f0e, 32'h3f71e9ba} /* (17, 2, 2) {real, imag} */,
  {32'hbfd14def, 32'hc0071064} /* (17, 2, 1) {real, imag} */,
  {32'hc01b9977, 32'h00000000} /* (17, 2, 0) {real, imag} */,
  {32'hbfd0e884, 32'h3ff913cb} /* (17, 1, 31) {real, imag} */,
  {32'hbe41b94a, 32'hbf61c57b} /* (17, 1, 30) {real, imag} */,
  {32'h3e60b47e, 32'h3e61d376} /* (17, 1, 29) {real, imag} */,
  {32'h3ceafe4c, 32'hbebe165d} /* (17, 1, 28) {real, imag} */,
  {32'h3dfb813f, 32'h3e78ffef} /* (17, 1, 27) {real, imag} */,
  {32'hbd24a1f1, 32'hbd9e9be4} /* (17, 1, 26) {real, imag} */,
  {32'hbd369183, 32'h3d9eda2a} /* (17, 1, 25) {real, imag} */,
  {32'h3c9a73ad, 32'hbdf4b0d2} /* (17, 1, 24) {real, imag} */,
  {32'h3c60e0d2, 32'hbdd4fb20} /* (17, 1, 23) {real, imag} */,
  {32'hbbaebf30, 32'hbd0113c5} /* (17, 1, 22) {real, imag} */,
  {32'h3c9bec44, 32'hbcc197b6} /* (17, 1, 21) {real, imag} */,
  {32'h3dab70e6, 32'h3d31136e} /* (17, 1, 20) {real, imag} */,
  {32'hbc131816, 32'hbcaabd5c} /* (17, 1, 19) {real, imag} */,
  {32'hbcca334b, 32'h3dc5c9fe} /* (17, 1, 18) {real, imag} */,
  {32'h3cefdf1f, 32'hbca4dca3} /* (17, 1, 17) {real, imag} */,
  {32'h3cd73a1d, 32'h00000000} /* (17, 1, 16) {real, imag} */,
  {32'h3cefdf1f, 32'h3ca4dca3} /* (17, 1, 15) {real, imag} */,
  {32'hbcca334b, 32'hbdc5c9fe} /* (17, 1, 14) {real, imag} */,
  {32'hbc131816, 32'h3caabd5c} /* (17, 1, 13) {real, imag} */,
  {32'h3dab70e6, 32'hbd31136e} /* (17, 1, 12) {real, imag} */,
  {32'h3c9bec44, 32'h3cc197b6} /* (17, 1, 11) {real, imag} */,
  {32'hbbaebf30, 32'h3d0113c5} /* (17, 1, 10) {real, imag} */,
  {32'h3c60e0d2, 32'h3dd4fb20} /* (17, 1, 9) {real, imag} */,
  {32'h3c9a73ad, 32'h3df4b0d2} /* (17, 1, 8) {real, imag} */,
  {32'hbd369183, 32'hbd9eda2a} /* (17, 1, 7) {real, imag} */,
  {32'hbd24a1f1, 32'h3d9e9be4} /* (17, 1, 6) {real, imag} */,
  {32'h3dfb813f, 32'hbe78ffef} /* (17, 1, 5) {real, imag} */,
  {32'h3ceafe4c, 32'h3ebe165d} /* (17, 1, 4) {real, imag} */,
  {32'h3e60b47e, 32'hbe61d376} /* (17, 1, 3) {real, imag} */,
  {32'hbe41b94a, 32'h3f61c57b} /* (17, 1, 2) {real, imag} */,
  {32'hbfd0e884, 32'hbff913cb} /* (17, 1, 1) {real, imag} */,
  {32'hc028b830, 32'h00000000} /* (17, 1, 0) {real, imag} */,
  {32'hbfdfa87c, 32'h3fc76120} /* (17, 0, 31) {real, imag} */,
  {32'h3d625df0, 32'hbf1ba575} /* (17, 0, 30) {real, imag} */,
  {32'h3dbaf1f5, 32'h3e0110fc} /* (17, 0, 29) {real, imag} */,
  {32'h3c42cf00, 32'hbdd01c08} /* (17, 0, 28) {real, imag} */,
  {32'h3d94237f, 32'hbc26b8a8} /* (17, 0, 27) {real, imag} */,
  {32'h3ce6fb1b, 32'h3985f680} /* (17, 0, 26) {real, imag} */,
  {32'hbc9e17c8, 32'h3d8427ae} /* (17, 0, 25) {real, imag} */,
  {32'h3d096f4e, 32'hbc036f94} /* (17, 0, 24) {real, imag} */,
  {32'h3cc69ab2, 32'h3c3fe33c} /* (17, 0, 23) {real, imag} */,
  {32'hbd08d186, 32'h3c88848d} /* (17, 0, 22) {real, imag} */,
  {32'hbc8f24c2, 32'h3cc571a4} /* (17, 0, 21) {real, imag} */,
  {32'h3d283c5c, 32'h3d3c3370} /* (17, 0, 20) {real, imag} */,
  {32'hbc6396c1, 32'h3cf4d766} /* (17, 0, 19) {real, imag} */,
  {32'h3c5158d8, 32'h3d071ebe} /* (17, 0, 18) {real, imag} */,
  {32'hbc59425c, 32'h3aa80050} /* (17, 0, 17) {real, imag} */,
  {32'h3c627f9c, 32'h00000000} /* (17, 0, 16) {real, imag} */,
  {32'hbc59425c, 32'hbaa80050} /* (17, 0, 15) {real, imag} */,
  {32'h3c5158d8, 32'hbd071ebe} /* (17, 0, 14) {real, imag} */,
  {32'hbc6396c1, 32'hbcf4d766} /* (17, 0, 13) {real, imag} */,
  {32'h3d283c5c, 32'hbd3c3370} /* (17, 0, 12) {real, imag} */,
  {32'hbc8f24c2, 32'hbcc571a4} /* (17, 0, 11) {real, imag} */,
  {32'hbd08d186, 32'hbc88848d} /* (17, 0, 10) {real, imag} */,
  {32'h3cc69ab2, 32'hbc3fe33c} /* (17, 0, 9) {real, imag} */,
  {32'h3d096f4e, 32'h3c036f94} /* (17, 0, 8) {real, imag} */,
  {32'hbc9e17c8, 32'hbd8427ae} /* (17, 0, 7) {real, imag} */,
  {32'h3ce6fb1b, 32'hb985f680} /* (17, 0, 6) {real, imag} */,
  {32'h3d94237f, 32'h3c26b8a8} /* (17, 0, 5) {real, imag} */,
  {32'h3c42cf00, 32'h3dd01c08} /* (17, 0, 4) {real, imag} */,
  {32'h3dbaf1f5, 32'hbe0110fc} /* (17, 0, 3) {real, imag} */,
  {32'h3d625df0, 32'h3f1ba575} /* (17, 0, 2) {real, imag} */,
  {32'hbfdfa87c, 32'hbfc76120} /* (17, 0, 1) {real, imag} */,
  {32'hc01fc958, 32'h00000000} /* (17, 0, 0) {real, imag} */,
  {32'hbf4cda95, 32'h3e9cadae} /* (16, 31, 31) {real, imag} */,
  {32'h3e2d539a, 32'hbe7c54be} /* (16, 31, 30) {real, imag} */,
  {32'h3d4da90e, 32'h3da4fe42} /* (16, 31, 29) {real, imag} */,
  {32'hbd9b9a69, 32'h3d795a4e} /* (16, 31, 28) {real, imag} */,
  {32'h3dd4e3ad, 32'hbcc4dff0} /* (16, 31, 27) {real, imag} */,
  {32'h3d21b926, 32'hbc544bd4} /* (16, 31, 26) {real, imag} */,
  {32'hbcaed732, 32'h3b589470} /* (16, 31, 25) {real, imag} */,
  {32'h3b129328, 32'h3d89d4c5} /* (16, 31, 24) {real, imag} */,
  {32'hbc488120, 32'hbc4e57c5} /* (16, 31, 23) {real, imag} */,
  {32'h3b523fdc, 32'hbb188e58} /* (16, 31, 22) {real, imag} */,
  {32'h3c554c0a, 32'h3cfcd610} /* (16, 31, 21) {real, imag} */,
  {32'hbb86c5fe, 32'h3ba12d20} /* (16, 31, 20) {real, imag} */,
  {32'hbdc628ac, 32'hbdb52652} /* (16, 31, 19) {real, imag} */,
  {32'h3d2d493a, 32'hbd211fe3} /* (16, 31, 18) {real, imag} */,
  {32'h3c6efa24, 32'hbcabedb0} /* (16, 31, 17) {real, imag} */,
  {32'h3dab895e, 32'h00000000} /* (16, 31, 16) {real, imag} */,
  {32'h3c6efa24, 32'h3cabedb0} /* (16, 31, 15) {real, imag} */,
  {32'h3d2d493a, 32'h3d211fe3} /* (16, 31, 14) {real, imag} */,
  {32'hbdc628ac, 32'h3db52652} /* (16, 31, 13) {real, imag} */,
  {32'hbb86c5fe, 32'hbba12d20} /* (16, 31, 12) {real, imag} */,
  {32'h3c554c0a, 32'hbcfcd610} /* (16, 31, 11) {real, imag} */,
  {32'h3b523fdc, 32'h3b188e58} /* (16, 31, 10) {real, imag} */,
  {32'hbc488120, 32'h3c4e57c5} /* (16, 31, 9) {real, imag} */,
  {32'h3b129328, 32'hbd89d4c5} /* (16, 31, 8) {real, imag} */,
  {32'hbcaed732, 32'hbb589470} /* (16, 31, 7) {real, imag} */,
  {32'h3d21b926, 32'h3c544bd4} /* (16, 31, 6) {real, imag} */,
  {32'h3dd4e3ad, 32'h3cc4dff0} /* (16, 31, 5) {real, imag} */,
  {32'hbd9b9a69, 32'hbd795a4e} /* (16, 31, 4) {real, imag} */,
  {32'h3d4da90e, 32'hbda4fe42} /* (16, 31, 3) {real, imag} */,
  {32'h3e2d539a, 32'h3e7c54be} /* (16, 31, 2) {real, imag} */,
  {32'hbf4cda95, 32'hbe9cadae} /* (16, 31, 1) {real, imag} */,
  {32'hbf8fd602, 32'h00000000} /* (16, 31, 0) {real, imag} */,
  {32'hbf95eedc, 32'h3e168e68} /* (16, 30, 31) {real, imag} */,
  {32'h3ea675da, 32'hbe27c75e} /* (16, 30, 30) {real, imag} */,
  {32'h3dd17991, 32'h3dedc80e} /* (16, 30, 29) {real, imag} */,
  {32'hbcd8ec1d, 32'h3cc33e10} /* (16, 30, 28) {real, imag} */,
  {32'h3e47428f, 32'hbdef2d26} /* (16, 30, 27) {real, imag} */,
  {32'h3db82066, 32'hbdcdd6b0} /* (16, 30, 26) {real, imag} */,
  {32'hbaa6ff00, 32'h3dfce8ee} /* (16, 30, 25) {real, imag} */,
  {32'hbcdd4c6e, 32'hbaa8e890} /* (16, 30, 24) {real, imag} */,
  {32'hbac76180, 32'hbc88bf60} /* (16, 30, 23) {real, imag} */,
  {32'hbc82faa4, 32'hbd22bac2} /* (16, 30, 22) {real, imag} */,
  {32'h3d39959a, 32'hbc467b70} /* (16, 30, 21) {real, imag} */,
  {32'hbc1b6472, 32'h3cc3532d} /* (16, 30, 20) {real, imag} */,
  {32'hbd1a6ca6, 32'h3d7d0f74} /* (16, 30, 19) {real, imag} */,
  {32'hbda291f3, 32'h3da49903} /* (16, 30, 18) {real, imag} */,
  {32'hbcb2708a, 32'hbc38b857} /* (16, 30, 17) {real, imag} */,
  {32'hbc879631, 32'h00000000} /* (16, 30, 16) {real, imag} */,
  {32'hbcb2708a, 32'h3c38b857} /* (16, 30, 15) {real, imag} */,
  {32'hbda291f3, 32'hbda49903} /* (16, 30, 14) {real, imag} */,
  {32'hbd1a6ca6, 32'hbd7d0f74} /* (16, 30, 13) {real, imag} */,
  {32'hbc1b6472, 32'hbcc3532d} /* (16, 30, 12) {real, imag} */,
  {32'h3d39959a, 32'h3c467b70} /* (16, 30, 11) {real, imag} */,
  {32'hbc82faa4, 32'h3d22bac2} /* (16, 30, 10) {real, imag} */,
  {32'hbac76180, 32'h3c88bf60} /* (16, 30, 9) {real, imag} */,
  {32'hbcdd4c6e, 32'h3aa8e890} /* (16, 30, 8) {real, imag} */,
  {32'hbaa6ff00, 32'hbdfce8ee} /* (16, 30, 7) {real, imag} */,
  {32'h3db82066, 32'h3dcdd6b0} /* (16, 30, 6) {real, imag} */,
  {32'h3e47428f, 32'h3def2d26} /* (16, 30, 5) {real, imag} */,
  {32'hbcd8ec1d, 32'hbcc33e10} /* (16, 30, 4) {real, imag} */,
  {32'h3dd17991, 32'hbdedc80e} /* (16, 30, 3) {real, imag} */,
  {32'h3ea675da, 32'h3e27c75e} /* (16, 30, 2) {real, imag} */,
  {32'hbf95eedc, 32'hbe168e68} /* (16, 30, 1) {real, imag} */,
  {32'hbf908a20, 32'h00000000} /* (16, 30, 0) {real, imag} */,
  {32'hbfc948c1, 32'h3de088a4} /* (16, 29, 31) {real, imag} */,
  {32'h3ed72d76, 32'hbe731e8a} /* (16, 29, 30) {real, imag} */,
  {32'h3da2dbdc, 32'h3c939cdc} /* (16, 29, 29) {real, imag} */,
  {32'hbe2578c0, 32'h3bb4e0e0} /* (16, 29, 28) {real, imag} */,
  {32'h3e1b16f4, 32'hbe012303} /* (16, 29, 27) {real, imag} */,
  {32'h3e3a0d2e, 32'hbe2f76af} /* (16, 29, 26) {real, imag} */,
  {32'hbd7bd6f8, 32'hbd1874b7} /* (16, 29, 25) {real, imag} */,
  {32'hbc34f682, 32'h3a809300} /* (16, 29, 24) {real, imag} */,
  {32'h3dc29442, 32'hbc326142} /* (16, 29, 23) {real, imag} */,
  {32'hbb948e22, 32'h3d33c56a} /* (16, 29, 22) {real, imag} */,
  {32'hbccd283c, 32'hbd856e87} /* (16, 29, 21) {real, imag} */,
  {32'hbd4d840a, 32'h3c22c8cc} /* (16, 29, 20) {real, imag} */,
  {32'h3d913f64, 32'hbcb0156b} /* (16, 29, 19) {real, imag} */,
  {32'hbd8e3966, 32'h3d2d200a} /* (16, 29, 18) {real, imag} */,
  {32'hbc589e56, 32'h3d436710} /* (16, 29, 17) {real, imag} */,
  {32'hbca61850, 32'h00000000} /* (16, 29, 16) {real, imag} */,
  {32'hbc589e56, 32'hbd436710} /* (16, 29, 15) {real, imag} */,
  {32'hbd8e3966, 32'hbd2d200a} /* (16, 29, 14) {real, imag} */,
  {32'h3d913f64, 32'h3cb0156b} /* (16, 29, 13) {real, imag} */,
  {32'hbd4d840a, 32'hbc22c8cc} /* (16, 29, 12) {real, imag} */,
  {32'hbccd283c, 32'h3d856e87} /* (16, 29, 11) {real, imag} */,
  {32'hbb948e22, 32'hbd33c56a} /* (16, 29, 10) {real, imag} */,
  {32'h3dc29442, 32'h3c326142} /* (16, 29, 9) {real, imag} */,
  {32'hbc34f682, 32'hba809300} /* (16, 29, 8) {real, imag} */,
  {32'hbd7bd6f8, 32'h3d1874b7} /* (16, 29, 7) {real, imag} */,
  {32'h3e3a0d2e, 32'h3e2f76af} /* (16, 29, 6) {real, imag} */,
  {32'h3e1b16f4, 32'h3e012303} /* (16, 29, 5) {real, imag} */,
  {32'hbe2578c0, 32'hbbb4e0e0} /* (16, 29, 4) {real, imag} */,
  {32'h3da2dbdc, 32'hbc939cdc} /* (16, 29, 3) {real, imag} */,
  {32'h3ed72d76, 32'h3e731e8a} /* (16, 29, 2) {real, imag} */,
  {32'hbfc948c1, 32'hbde088a4} /* (16, 29, 1) {real, imag} */,
  {32'hbf6a51fc, 32'h00000000} /* (16, 29, 0) {real, imag} */,
  {32'hbfca6a6d, 32'h3e35b078} /* (16, 28, 31) {real, imag} */,
  {32'h3edc085d, 32'hbe9cced3} /* (16, 28, 30) {real, imag} */,
  {32'hbb0235c8, 32'hbc95f5be} /* (16, 28, 29) {real, imag} */,
  {32'hbe6011db, 32'hbde387d4} /* (16, 28, 28) {real, imag} */,
  {32'h3dce9854, 32'hbc2498d6} /* (16, 28, 27) {real, imag} */,
  {32'h3df34626, 32'h3d4f4eb4} /* (16, 28, 26) {real, imag} */,
  {32'h3d005a94, 32'hbd7e4d84} /* (16, 28, 25) {real, imag} */,
  {32'hbd23fe5e, 32'h3dad4b03} /* (16, 28, 24) {real, imag} */,
  {32'h3e45c7e6, 32'h3d658d25} /* (16, 28, 23) {real, imag} */,
  {32'hbd1b2790, 32'hbc926d16} /* (16, 28, 22) {real, imag} */,
  {32'hbcc18860, 32'h3c61b498} /* (16, 28, 21) {real, imag} */,
  {32'h3cefa3ce, 32'hbe197897} /* (16, 28, 20) {real, imag} */,
  {32'h3d46a6da, 32'hbb6f6ee4} /* (16, 28, 19) {real, imag} */,
  {32'h3ced0e2c, 32'hbd98b0d6} /* (16, 28, 18) {real, imag} */,
  {32'h39f1b518, 32'h3d28f16a} /* (16, 28, 17) {real, imag} */,
  {32'h3e05d9d8, 32'h00000000} /* (16, 28, 16) {real, imag} */,
  {32'h39f1b518, 32'hbd28f16a} /* (16, 28, 15) {real, imag} */,
  {32'h3ced0e2c, 32'h3d98b0d6} /* (16, 28, 14) {real, imag} */,
  {32'h3d46a6da, 32'h3b6f6ee4} /* (16, 28, 13) {real, imag} */,
  {32'h3cefa3ce, 32'h3e197897} /* (16, 28, 12) {real, imag} */,
  {32'hbcc18860, 32'hbc61b498} /* (16, 28, 11) {real, imag} */,
  {32'hbd1b2790, 32'h3c926d16} /* (16, 28, 10) {real, imag} */,
  {32'h3e45c7e6, 32'hbd658d25} /* (16, 28, 9) {real, imag} */,
  {32'hbd23fe5e, 32'hbdad4b03} /* (16, 28, 8) {real, imag} */,
  {32'h3d005a94, 32'h3d7e4d84} /* (16, 28, 7) {real, imag} */,
  {32'h3df34626, 32'hbd4f4eb4} /* (16, 28, 6) {real, imag} */,
  {32'h3dce9854, 32'h3c2498d6} /* (16, 28, 5) {real, imag} */,
  {32'hbe6011db, 32'h3de387d4} /* (16, 28, 4) {real, imag} */,
  {32'hbb0235c8, 32'h3c95f5be} /* (16, 28, 3) {real, imag} */,
  {32'h3edc085d, 32'h3e9cced3} /* (16, 28, 2) {real, imag} */,
  {32'hbfca6a6d, 32'hbe35b078} /* (16, 28, 1) {real, imag} */,
  {32'hbf88915a, 32'h00000000} /* (16, 28, 0) {real, imag} */,
  {32'hbfb1f2a3, 32'h3d6199f0} /* (16, 27, 31) {real, imag} */,
  {32'h3eb9beb0, 32'hbe570365} /* (16, 27, 30) {real, imag} */,
  {32'h3d11121b, 32'hbc07c53c} /* (16, 27, 29) {real, imag} */,
  {32'hbe53ff3d, 32'hbd8ad592} /* (16, 27, 28) {real, imag} */,
  {32'h3dded714, 32'h3c8efedc} /* (16, 27, 27) {real, imag} */,
  {32'h3d98a654, 32'hbdb70b71} /* (16, 27, 26) {real, imag} */,
  {32'hbd21cf64, 32'h3cfd346c} /* (16, 27, 25) {real, imag} */,
  {32'hbd416f04, 32'hbd2a26a6} /* (16, 27, 24) {real, imag} */,
  {32'h3cc02bfd, 32'h3d89c4d4} /* (16, 27, 23) {real, imag} */,
  {32'hbd18a514, 32'hbd573e68} /* (16, 27, 22) {real, imag} */,
  {32'h3be38418, 32'hbd4cf186} /* (16, 27, 21) {real, imag} */,
  {32'hbc05916f, 32'hbd34ceb7} /* (16, 27, 20) {real, imag} */,
  {32'h3ca73c94, 32'h3d89e064} /* (16, 27, 19) {real, imag} */,
  {32'h3b4ea2cc, 32'hba3b5bb0} /* (16, 27, 18) {real, imag} */,
  {32'hbb4d5ea8, 32'hbd35d424} /* (16, 27, 17) {real, imag} */,
  {32'hbc853e48, 32'h00000000} /* (16, 27, 16) {real, imag} */,
  {32'hbb4d5ea8, 32'h3d35d424} /* (16, 27, 15) {real, imag} */,
  {32'h3b4ea2cc, 32'h3a3b5bb0} /* (16, 27, 14) {real, imag} */,
  {32'h3ca73c94, 32'hbd89e064} /* (16, 27, 13) {real, imag} */,
  {32'hbc05916f, 32'h3d34ceb7} /* (16, 27, 12) {real, imag} */,
  {32'h3be38418, 32'h3d4cf186} /* (16, 27, 11) {real, imag} */,
  {32'hbd18a514, 32'h3d573e68} /* (16, 27, 10) {real, imag} */,
  {32'h3cc02bfd, 32'hbd89c4d4} /* (16, 27, 9) {real, imag} */,
  {32'hbd416f04, 32'h3d2a26a6} /* (16, 27, 8) {real, imag} */,
  {32'hbd21cf64, 32'hbcfd346c} /* (16, 27, 7) {real, imag} */,
  {32'h3d98a654, 32'h3db70b71} /* (16, 27, 6) {real, imag} */,
  {32'h3dded714, 32'hbc8efedc} /* (16, 27, 5) {real, imag} */,
  {32'hbe53ff3d, 32'h3d8ad592} /* (16, 27, 4) {real, imag} */,
  {32'h3d11121b, 32'h3c07c53c} /* (16, 27, 3) {real, imag} */,
  {32'h3eb9beb0, 32'h3e570365} /* (16, 27, 2) {real, imag} */,
  {32'hbfb1f2a3, 32'hbd6199f0} /* (16, 27, 1) {real, imag} */,
  {32'hbf8cee4c, 32'h00000000} /* (16, 27, 0) {real, imag} */,
  {32'hbfa184df, 32'h3a16a200} /* (16, 26, 31) {real, imag} */,
  {32'h3e9e38cf, 32'hbe0b80a2} /* (16, 26, 30) {real, imag} */,
  {32'h3d1a8528, 32'hbd567f06} /* (16, 26, 29) {real, imag} */,
  {32'hbe6166a5, 32'hbd824484} /* (16, 26, 28) {real, imag} */,
  {32'h3c82896a, 32'hbd7aa0a8} /* (16, 26, 27) {real, imag} */,
  {32'h3d75cd98, 32'hbd7051e1} /* (16, 26, 26) {real, imag} */,
  {32'hbcbba58f, 32'hbceb322f} /* (16, 26, 25) {real, imag} */,
  {32'h3d512c32, 32'hbb8ee860} /* (16, 26, 24) {real, imag} */,
  {32'h3d9e499f, 32'h3b8ffd6e} /* (16, 26, 23) {real, imag} */,
  {32'h3db48160, 32'h3d58de66} /* (16, 26, 22) {real, imag} */,
  {32'h3d6ebc1c, 32'hbde6bed2} /* (16, 26, 21) {real, imag} */,
  {32'hbd8232fe, 32'hbc2135c6} /* (16, 26, 20) {real, imag} */,
  {32'h3cf61c06, 32'h3d3e6844} /* (16, 26, 19) {real, imag} */,
  {32'hbd296d25, 32'h3c8d8b4c} /* (16, 26, 18) {real, imag} */,
  {32'hbd60f90f, 32'hbc3cc277} /* (16, 26, 17) {real, imag} */,
  {32'hbcc2e71e, 32'h00000000} /* (16, 26, 16) {real, imag} */,
  {32'hbd60f90f, 32'h3c3cc277} /* (16, 26, 15) {real, imag} */,
  {32'hbd296d25, 32'hbc8d8b4c} /* (16, 26, 14) {real, imag} */,
  {32'h3cf61c06, 32'hbd3e6844} /* (16, 26, 13) {real, imag} */,
  {32'hbd8232fe, 32'h3c2135c6} /* (16, 26, 12) {real, imag} */,
  {32'h3d6ebc1c, 32'h3de6bed2} /* (16, 26, 11) {real, imag} */,
  {32'h3db48160, 32'hbd58de66} /* (16, 26, 10) {real, imag} */,
  {32'h3d9e499f, 32'hbb8ffd6e} /* (16, 26, 9) {real, imag} */,
  {32'h3d512c32, 32'h3b8ee860} /* (16, 26, 8) {real, imag} */,
  {32'hbcbba58f, 32'h3ceb322f} /* (16, 26, 7) {real, imag} */,
  {32'h3d75cd98, 32'h3d7051e1} /* (16, 26, 6) {real, imag} */,
  {32'h3c82896a, 32'h3d7aa0a8} /* (16, 26, 5) {real, imag} */,
  {32'hbe6166a5, 32'h3d824484} /* (16, 26, 4) {real, imag} */,
  {32'h3d1a8528, 32'h3d567f06} /* (16, 26, 3) {real, imag} */,
  {32'h3e9e38cf, 32'h3e0b80a2} /* (16, 26, 2) {real, imag} */,
  {32'hbfa184df, 32'hba16a200} /* (16, 26, 1) {real, imag} */,
  {32'hbf9e1ac1, 32'h00000000} /* (16, 26, 0) {real, imag} */,
  {32'hbf9c833d, 32'h3d92b61c} /* (16, 25, 31) {real, imag} */,
  {32'h3e9d580b, 32'hbe02f988} /* (16, 25, 30) {real, imag} */,
  {32'hbcb4b334, 32'hbdd95ed9} /* (16, 25, 29) {real, imag} */,
  {32'hbe45402c, 32'hbd7d50e8} /* (16, 25, 28) {real, imag} */,
  {32'h3e2ae79d, 32'hbb70c0c0} /* (16, 25, 27) {real, imag} */,
  {32'h3d81f97c, 32'hbd0eee40} /* (16, 25, 26) {real, imag} */,
  {32'hbd807510, 32'h3ad4ba70} /* (16, 25, 25) {real, imag} */,
  {32'h3dd67009, 32'hbd944dd1} /* (16, 25, 24) {real, imag} */,
  {32'hbb3cda20, 32'hbcf38b22} /* (16, 25, 23) {real, imag} */,
  {32'hbc4a2f87, 32'h3cd16af4} /* (16, 25, 22) {real, imag} */,
  {32'hbd29f6a9, 32'hbd3a6548} /* (16, 25, 21) {real, imag} */,
  {32'h3d2d6068, 32'hbd90f5bd} /* (16, 25, 20) {real, imag} */,
  {32'h3d50a6cc, 32'h3d413074} /* (16, 25, 19) {real, imag} */,
  {32'hbc7cad2c, 32'hbd253eaa} /* (16, 25, 18) {real, imag} */,
  {32'h3da8b1a0, 32'h3d066b34} /* (16, 25, 17) {real, imag} */,
  {32'hbceae242, 32'h00000000} /* (16, 25, 16) {real, imag} */,
  {32'h3da8b1a0, 32'hbd066b34} /* (16, 25, 15) {real, imag} */,
  {32'hbc7cad2c, 32'h3d253eaa} /* (16, 25, 14) {real, imag} */,
  {32'h3d50a6cc, 32'hbd413074} /* (16, 25, 13) {real, imag} */,
  {32'h3d2d6068, 32'h3d90f5bd} /* (16, 25, 12) {real, imag} */,
  {32'hbd29f6a9, 32'h3d3a6548} /* (16, 25, 11) {real, imag} */,
  {32'hbc4a2f87, 32'hbcd16af4} /* (16, 25, 10) {real, imag} */,
  {32'hbb3cda20, 32'h3cf38b22} /* (16, 25, 9) {real, imag} */,
  {32'h3dd67009, 32'h3d944dd1} /* (16, 25, 8) {real, imag} */,
  {32'hbd807510, 32'hbad4ba70} /* (16, 25, 7) {real, imag} */,
  {32'h3d81f97c, 32'h3d0eee40} /* (16, 25, 6) {real, imag} */,
  {32'h3e2ae79d, 32'h3b70c0c0} /* (16, 25, 5) {real, imag} */,
  {32'hbe45402c, 32'h3d7d50e8} /* (16, 25, 4) {real, imag} */,
  {32'hbcb4b334, 32'h3dd95ed9} /* (16, 25, 3) {real, imag} */,
  {32'h3e9d580b, 32'h3e02f988} /* (16, 25, 2) {real, imag} */,
  {32'hbf9c833d, 32'hbd92b61c} /* (16, 25, 1) {real, imag} */,
  {32'hbf9956ac, 32'h00000000} /* (16, 25, 0) {real, imag} */,
  {32'hbf8e3966, 32'h3da58e50} /* (16, 24, 31) {real, imag} */,
  {32'h3edf03d2, 32'hbe4f4914} /* (16, 24, 30) {real, imag} */,
  {32'hbd4e02dc, 32'hbe36c37d} /* (16, 24, 29) {real, imag} */,
  {32'hbe83d40f, 32'hbdbc08b0} /* (16, 24, 28) {real, imag} */,
  {32'h3e1fbac6, 32'hbdff6ca8} /* (16, 24, 27) {real, imag} */,
  {32'h3d6cef47, 32'h3d960c67} /* (16, 24, 26) {real, imag} */,
  {32'hbdbf16ce, 32'hbcd32bba} /* (16, 24, 25) {real, imag} */,
  {32'h3de2485e, 32'hbc676554} /* (16, 24, 24) {real, imag} */,
  {32'h3dcce6e3, 32'h3d9c21fb} /* (16, 24, 23) {real, imag} */,
  {32'h3d5d3fe1, 32'h3d11291c} /* (16, 24, 22) {real, imag} */,
  {32'h3c915964, 32'hbcf29743} /* (16, 24, 21) {real, imag} */,
  {32'h3c714dc0, 32'h3da63bca} /* (16, 24, 20) {real, imag} */,
  {32'hbd42ffc1, 32'hbd06adae} /* (16, 24, 19) {real, imag} */,
  {32'h3d2d1f3e, 32'h3d948f54} /* (16, 24, 18) {real, imag} */,
  {32'h3d0ac37e, 32'hbda7912a} /* (16, 24, 17) {real, imag} */,
  {32'h3d55196c, 32'h00000000} /* (16, 24, 16) {real, imag} */,
  {32'h3d0ac37e, 32'h3da7912a} /* (16, 24, 15) {real, imag} */,
  {32'h3d2d1f3e, 32'hbd948f54} /* (16, 24, 14) {real, imag} */,
  {32'hbd42ffc1, 32'h3d06adae} /* (16, 24, 13) {real, imag} */,
  {32'h3c714dc0, 32'hbda63bca} /* (16, 24, 12) {real, imag} */,
  {32'h3c915964, 32'h3cf29743} /* (16, 24, 11) {real, imag} */,
  {32'h3d5d3fe1, 32'hbd11291c} /* (16, 24, 10) {real, imag} */,
  {32'h3dcce6e3, 32'hbd9c21fb} /* (16, 24, 9) {real, imag} */,
  {32'h3de2485e, 32'h3c676554} /* (16, 24, 8) {real, imag} */,
  {32'hbdbf16ce, 32'h3cd32bba} /* (16, 24, 7) {real, imag} */,
  {32'h3d6cef47, 32'hbd960c67} /* (16, 24, 6) {real, imag} */,
  {32'h3e1fbac6, 32'h3dff6ca8} /* (16, 24, 5) {real, imag} */,
  {32'hbe83d40f, 32'h3dbc08b0} /* (16, 24, 4) {real, imag} */,
  {32'hbd4e02dc, 32'h3e36c37d} /* (16, 24, 3) {real, imag} */,
  {32'h3edf03d2, 32'h3e4f4914} /* (16, 24, 2) {real, imag} */,
  {32'hbf8e3966, 32'hbda58e50} /* (16, 24, 1) {real, imag} */,
  {32'hbf97702b, 32'h00000000} /* (16, 24, 0) {real, imag} */,
  {32'hbf565dea, 32'h3e01d4de} /* (16, 23, 31) {real, imag} */,
  {32'h3efbefd7, 32'hbcd31a21} /* (16, 23, 30) {real, imag} */,
  {32'hbd75cf7b, 32'hbde7c415} /* (16, 23, 29) {real, imag} */,
  {32'hbe469827, 32'hbe00f6b7} /* (16, 23, 28) {real, imag} */,
  {32'h3d9599b2, 32'hbd6bd2d8} /* (16, 23, 27) {real, imag} */,
  {32'hbe03639f, 32'hbd4a62dc} /* (16, 23, 26) {real, imag} */,
  {32'hbe0b5e03, 32'h3bbb09a8} /* (16, 23, 25) {real, imag} */,
  {32'h3e16476d, 32'hbd45650e} /* (16, 23, 24) {real, imag} */,
  {32'h3dd2b543, 32'hbd14449d} /* (16, 23, 23) {real, imag} */,
  {32'h3daa3cbb, 32'hbd3eaffe} /* (16, 23, 22) {real, imag} */,
  {32'h3d2e4734, 32'h3dae8eb7} /* (16, 23, 21) {real, imag} */,
  {32'hbd9474c2, 32'h3dbb0cc4} /* (16, 23, 20) {real, imag} */,
  {32'h3ce8ebec, 32'h3b61d080} /* (16, 23, 19) {real, imag} */,
  {32'hb9bdd700, 32'hbde62c15} /* (16, 23, 18) {real, imag} */,
  {32'hbd2bcd02, 32'h3d37dadd} /* (16, 23, 17) {real, imag} */,
  {32'h3d5c2aaa, 32'h00000000} /* (16, 23, 16) {real, imag} */,
  {32'hbd2bcd02, 32'hbd37dadd} /* (16, 23, 15) {real, imag} */,
  {32'hb9bdd700, 32'h3de62c15} /* (16, 23, 14) {real, imag} */,
  {32'h3ce8ebec, 32'hbb61d080} /* (16, 23, 13) {real, imag} */,
  {32'hbd9474c2, 32'hbdbb0cc4} /* (16, 23, 12) {real, imag} */,
  {32'h3d2e4734, 32'hbdae8eb7} /* (16, 23, 11) {real, imag} */,
  {32'h3daa3cbb, 32'h3d3eaffe} /* (16, 23, 10) {real, imag} */,
  {32'h3dd2b543, 32'h3d14449d} /* (16, 23, 9) {real, imag} */,
  {32'h3e16476d, 32'h3d45650e} /* (16, 23, 8) {real, imag} */,
  {32'hbe0b5e03, 32'hbbbb09a8} /* (16, 23, 7) {real, imag} */,
  {32'hbe03639f, 32'h3d4a62dc} /* (16, 23, 6) {real, imag} */,
  {32'h3d9599b2, 32'h3d6bd2d8} /* (16, 23, 5) {real, imag} */,
  {32'hbe469827, 32'h3e00f6b7} /* (16, 23, 4) {real, imag} */,
  {32'hbd75cf7b, 32'h3de7c415} /* (16, 23, 3) {real, imag} */,
  {32'h3efbefd7, 32'h3cd31a21} /* (16, 23, 2) {real, imag} */,
  {32'hbf565dea, 32'hbe01d4de} /* (16, 23, 1) {real, imag} */,
  {32'hbf89fc32, 32'h00000000} /* (16, 23, 0) {real, imag} */,
  {32'hbf372cca, 32'h3db95010} /* (16, 22, 31) {real, imag} */,
  {32'h3ecb5dfa, 32'hbcc92c7a} /* (16, 22, 30) {real, imag} */,
  {32'hbd846ed6, 32'hbd3adec2} /* (16, 22, 29) {real, imag} */,
  {32'hbe3ec336, 32'hbd7e2b93} /* (16, 22, 28) {real, imag} */,
  {32'h3daedfa6, 32'hbcdda36d} /* (16, 22, 27) {real, imag} */,
  {32'hbbed23c8, 32'hbd906468} /* (16, 22, 26) {real, imag} */,
  {32'h3c9f90e5, 32'h3d7e6dbe} /* (16, 22, 25) {real, imag} */,
  {32'h3d135044, 32'hbcf723cc} /* (16, 22, 24) {real, imag} */,
  {32'hbd3f3062, 32'hbd6d3314} /* (16, 22, 23) {real, imag} */,
  {32'h3d10b2f2, 32'h3da71cae} /* (16, 22, 22) {real, imag} */,
  {32'hbc74f177, 32'hbd9bcfcc} /* (16, 22, 21) {real, imag} */,
  {32'h3d7d2c05, 32'hbd1e6a70} /* (16, 22, 20) {real, imag} */,
  {32'h3d5c6dae, 32'h3d1f680a} /* (16, 22, 19) {real, imag} */,
  {32'h3d802e00, 32'hbd42e1d1} /* (16, 22, 18) {real, imag} */,
  {32'h3d463f2c, 32'h3d5a0fb4} /* (16, 22, 17) {real, imag} */,
  {32'h3c06acd8, 32'h00000000} /* (16, 22, 16) {real, imag} */,
  {32'h3d463f2c, 32'hbd5a0fb4} /* (16, 22, 15) {real, imag} */,
  {32'h3d802e00, 32'h3d42e1d1} /* (16, 22, 14) {real, imag} */,
  {32'h3d5c6dae, 32'hbd1f680a} /* (16, 22, 13) {real, imag} */,
  {32'h3d7d2c05, 32'h3d1e6a70} /* (16, 22, 12) {real, imag} */,
  {32'hbc74f177, 32'h3d9bcfcc} /* (16, 22, 11) {real, imag} */,
  {32'h3d10b2f2, 32'hbda71cae} /* (16, 22, 10) {real, imag} */,
  {32'hbd3f3062, 32'h3d6d3314} /* (16, 22, 9) {real, imag} */,
  {32'h3d135044, 32'h3cf723cc} /* (16, 22, 8) {real, imag} */,
  {32'h3c9f90e5, 32'hbd7e6dbe} /* (16, 22, 7) {real, imag} */,
  {32'hbbed23c8, 32'h3d906468} /* (16, 22, 6) {real, imag} */,
  {32'h3daedfa6, 32'h3cdda36d} /* (16, 22, 5) {real, imag} */,
  {32'hbe3ec336, 32'h3d7e2b93} /* (16, 22, 4) {real, imag} */,
  {32'hbd846ed6, 32'h3d3adec2} /* (16, 22, 3) {real, imag} */,
  {32'h3ecb5dfa, 32'h3cc92c7a} /* (16, 22, 2) {real, imag} */,
  {32'hbf372cca, 32'hbdb95010} /* (16, 22, 1) {real, imag} */,
  {32'hbf6f4ab9, 32'h00000000} /* (16, 22, 0) {real, imag} */,
  {32'hbea7658a, 32'h3d3eace0} /* (16, 21, 31) {real, imag} */,
  {32'h3e7ddfe0, 32'h3da8de70} /* (16, 21, 30) {real, imag} */,
  {32'h3d82a200, 32'hbbea8168} /* (16, 21, 29) {real, imag} */,
  {32'h3d30c732, 32'hbdb4c189} /* (16, 21, 28) {real, imag} */,
  {32'hbccb4ed0, 32'hbcaceee1} /* (16, 21, 27) {real, imag} */,
  {32'h3cb1c8c6, 32'hbd209e7c} /* (16, 21, 26) {real, imag} */,
  {32'h3dbf34c8, 32'h3d826530} /* (16, 21, 25) {real, imag} */,
  {32'hbb9deefc, 32'hbd85c282} /* (16, 21, 24) {real, imag} */,
  {32'h3c990fd1, 32'h3d800618} /* (16, 21, 23) {real, imag} */,
  {32'h3c0954c0, 32'h3d8e46c0} /* (16, 21, 22) {real, imag} */,
  {32'hbdafcdac, 32'h3d0479f0} /* (16, 21, 21) {real, imag} */,
  {32'hbdbbd1e8, 32'h3aed7ae0} /* (16, 21, 20) {real, imag} */,
  {32'hbaada2e0, 32'hbd930e2d} /* (16, 21, 19) {real, imag} */,
  {32'h3c8d04b4, 32'h3d248835} /* (16, 21, 18) {real, imag} */,
  {32'h3cfd1873, 32'hbd677525} /* (16, 21, 17) {real, imag} */,
  {32'hbb6ef940, 32'h00000000} /* (16, 21, 16) {real, imag} */,
  {32'h3cfd1873, 32'h3d677525} /* (16, 21, 15) {real, imag} */,
  {32'h3c8d04b4, 32'hbd248835} /* (16, 21, 14) {real, imag} */,
  {32'hbaada2e0, 32'h3d930e2d} /* (16, 21, 13) {real, imag} */,
  {32'hbdbbd1e8, 32'hbaed7ae0} /* (16, 21, 12) {real, imag} */,
  {32'hbdafcdac, 32'hbd0479f0} /* (16, 21, 11) {real, imag} */,
  {32'h3c0954c0, 32'hbd8e46c0} /* (16, 21, 10) {real, imag} */,
  {32'h3c990fd1, 32'hbd800618} /* (16, 21, 9) {real, imag} */,
  {32'hbb9deefc, 32'h3d85c282} /* (16, 21, 8) {real, imag} */,
  {32'h3dbf34c8, 32'hbd826530} /* (16, 21, 7) {real, imag} */,
  {32'h3cb1c8c6, 32'h3d209e7c} /* (16, 21, 6) {real, imag} */,
  {32'hbccb4ed0, 32'h3caceee1} /* (16, 21, 5) {real, imag} */,
  {32'h3d30c732, 32'h3db4c189} /* (16, 21, 4) {real, imag} */,
  {32'h3d82a200, 32'h3bea8168} /* (16, 21, 3) {real, imag} */,
  {32'h3e7ddfe0, 32'hbda8de70} /* (16, 21, 2) {real, imag} */,
  {32'hbea7658a, 32'hbd3eace0} /* (16, 21, 1) {real, imag} */,
  {32'hbf2bf9d9, 32'h00000000} /* (16, 21, 0) {real, imag} */,
  {32'h3e8408a5, 32'h3d148354} /* (16, 20, 31) {real, imag} */,
  {32'hbc52aeb0, 32'h3e5b1b6e} /* (16, 20, 30) {real, imag} */,
  {32'h3d0fc4dc, 32'h3dde8461} /* (16, 20, 29) {real, imag} */,
  {32'h3e5a4586, 32'hbdf9181f} /* (16, 20, 28) {real, imag} */,
  {32'hbde39916, 32'h3c32ba48} /* (16, 20, 27) {real, imag} */,
  {32'hbe538d6c, 32'hbe0152f2} /* (16, 20, 26) {real, imag} */,
  {32'h3d2b4658, 32'h3cbc11d2} /* (16, 20, 25) {real, imag} */,
  {32'hbde3e9a6, 32'h3b3190e0} /* (16, 20, 24) {real, imag} */,
  {32'h3c4ec188, 32'hbc368010} /* (16, 20, 23) {real, imag} */,
  {32'hbda6af60, 32'hbd14e9e8} /* (16, 20, 22) {real, imag} */,
  {32'h3db50792, 32'hbcd15554} /* (16, 20, 21) {real, imag} */,
  {32'h3d0f4888, 32'h3bcb62c8} /* (16, 20, 20) {real, imag} */,
  {32'hbd1337b2, 32'hbb645ef8} /* (16, 20, 19) {real, imag} */,
  {32'h3cd1117e, 32'hbb9b49c0} /* (16, 20, 18) {real, imag} */,
  {32'h3d83ba0a, 32'h3d448a7c} /* (16, 20, 17) {real, imag} */,
  {32'h3bf02ccc, 32'h00000000} /* (16, 20, 16) {real, imag} */,
  {32'h3d83ba0a, 32'hbd448a7c} /* (16, 20, 15) {real, imag} */,
  {32'h3cd1117e, 32'h3b9b49c0} /* (16, 20, 14) {real, imag} */,
  {32'hbd1337b2, 32'h3b645ef8} /* (16, 20, 13) {real, imag} */,
  {32'h3d0f4888, 32'hbbcb62c8} /* (16, 20, 12) {real, imag} */,
  {32'h3db50792, 32'h3cd15554} /* (16, 20, 11) {real, imag} */,
  {32'hbda6af60, 32'h3d14e9e8} /* (16, 20, 10) {real, imag} */,
  {32'h3c4ec188, 32'h3c368010} /* (16, 20, 9) {real, imag} */,
  {32'hbde3e9a6, 32'hbb3190e0} /* (16, 20, 8) {real, imag} */,
  {32'h3d2b4658, 32'hbcbc11d2} /* (16, 20, 7) {real, imag} */,
  {32'hbe538d6c, 32'h3e0152f2} /* (16, 20, 6) {real, imag} */,
  {32'hbde39916, 32'hbc32ba48} /* (16, 20, 5) {real, imag} */,
  {32'h3e5a4586, 32'h3df9181f} /* (16, 20, 4) {real, imag} */,
  {32'h3d0fc4dc, 32'hbdde8461} /* (16, 20, 3) {real, imag} */,
  {32'hbc52aeb0, 32'hbe5b1b6e} /* (16, 20, 2) {real, imag} */,
  {32'h3e8408a5, 32'hbd148354} /* (16, 20, 1) {real, imag} */,
  {32'hbc0fc120, 32'h00000000} /* (16, 20, 0) {real, imag} */,
  {32'h3f0582e0, 32'h3abb1700} /* (16, 19, 31) {real, imag} */,
  {32'hbe66c1d1, 32'h3e8d33e5} /* (16, 19, 30) {real, imag} */,
  {32'h3e42ebed, 32'h3dc8f931} /* (16, 19, 29) {real, imag} */,
  {32'h3e178a0c, 32'hbc7fde90} /* (16, 19, 28) {real, imag} */,
  {32'hbe2fb97e, 32'h3d237cdc} /* (16, 19, 27) {real, imag} */,
  {32'h3d2b9a48, 32'h3da321b2} /* (16, 19, 26) {real, imag} */,
  {32'h3e05ccab, 32'hbdb80055} /* (16, 19, 25) {real, imag} */,
  {32'hbde112fc, 32'h3e2da6b8} /* (16, 19, 24) {real, imag} */,
  {32'hbbbec778, 32'h3cdf7e08} /* (16, 19, 23) {real, imag} */,
  {32'hbbda0af0, 32'hbc055543} /* (16, 19, 22) {real, imag} */,
  {32'h3ca71f6c, 32'h3ccbd870} /* (16, 19, 21) {real, imag} */,
  {32'hbdc2cb54, 32'hbb460230} /* (16, 19, 20) {real, imag} */,
  {32'h3d1abdb1, 32'h3bb12781} /* (16, 19, 19) {real, imag} */,
  {32'hbd0b3b3c, 32'h3d0a2f9e} /* (16, 19, 18) {real, imag} */,
  {32'hbd1b0cb2, 32'h3ceae296} /* (16, 19, 17) {real, imag} */,
  {32'h3ce549e4, 32'h00000000} /* (16, 19, 16) {real, imag} */,
  {32'hbd1b0cb2, 32'hbceae296} /* (16, 19, 15) {real, imag} */,
  {32'hbd0b3b3c, 32'hbd0a2f9e} /* (16, 19, 14) {real, imag} */,
  {32'h3d1abdb1, 32'hbbb12781} /* (16, 19, 13) {real, imag} */,
  {32'hbdc2cb54, 32'h3b460230} /* (16, 19, 12) {real, imag} */,
  {32'h3ca71f6c, 32'hbccbd870} /* (16, 19, 11) {real, imag} */,
  {32'hbbda0af0, 32'h3c055543} /* (16, 19, 10) {real, imag} */,
  {32'hbbbec778, 32'hbcdf7e08} /* (16, 19, 9) {real, imag} */,
  {32'hbde112fc, 32'hbe2da6b8} /* (16, 19, 8) {real, imag} */,
  {32'h3e05ccab, 32'h3db80055} /* (16, 19, 7) {real, imag} */,
  {32'h3d2b9a48, 32'hbda321b2} /* (16, 19, 6) {real, imag} */,
  {32'hbe2fb97e, 32'hbd237cdc} /* (16, 19, 5) {real, imag} */,
  {32'h3e178a0c, 32'h3c7fde90} /* (16, 19, 4) {real, imag} */,
  {32'h3e42ebed, 32'hbdc8f931} /* (16, 19, 3) {real, imag} */,
  {32'hbe66c1d1, 32'hbe8d33e5} /* (16, 19, 2) {real, imag} */,
  {32'h3f0582e0, 32'hbabb1700} /* (16, 19, 1) {real, imag} */,
  {32'h3ec3540e, 32'h00000000} /* (16, 19, 0) {real, imag} */,
  {32'h3f4aa1e0, 32'hbd887656} /* (16, 18, 31) {real, imag} */,
  {32'hbeefc907, 32'h3dac0464} /* (16, 18, 30) {real, imag} */,
  {32'h3e82d715, 32'h3e0cf94c} /* (16, 18, 29) {real, imag} */,
  {32'h3e183d4a, 32'h3ce336e8} /* (16, 18, 28) {real, imag} */,
  {32'hbd79c3bc, 32'h3d3e6b74} /* (16, 18, 27) {real, imag} */,
  {32'h3d1598ac, 32'hbd903a11} /* (16, 18, 26) {real, imag} */,
  {32'h3dc2ac2a, 32'h3d266f57} /* (16, 18, 25) {real, imag} */,
  {32'h3ca06d8a, 32'hbc9e2e14} /* (16, 18, 24) {real, imag} */,
  {32'hbdb3fb90, 32'h3c4c8b3e} /* (16, 18, 23) {real, imag} */,
  {32'hbd4893b9, 32'h3dc23642} /* (16, 18, 22) {real, imag} */,
  {32'h3d308db5, 32'h3dcf92da} /* (16, 18, 21) {real, imag} */,
  {32'hbd45496e, 32'hbcc7a834} /* (16, 18, 20) {real, imag} */,
  {32'hbdd229dc, 32'hbda3f59a} /* (16, 18, 19) {real, imag} */,
  {32'h3bfc7e4e, 32'h3d5563e0} /* (16, 18, 18) {real, imag} */,
  {32'hbc995f8e, 32'hbd1d4840} /* (16, 18, 17) {real, imag} */,
  {32'h3d5c474c, 32'h00000000} /* (16, 18, 16) {real, imag} */,
  {32'hbc995f8e, 32'h3d1d4840} /* (16, 18, 15) {real, imag} */,
  {32'h3bfc7e4e, 32'hbd5563e0} /* (16, 18, 14) {real, imag} */,
  {32'hbdd229dc, 32'h3da3f59a} /* (16, 18, 13) {real, imag} */,
  {32'hbd45496e, 32'h3cc7a834} /* (16, 18, 12) {real, imag} */,
  {32'h3d308db5, 32'hbdcf92da} /* (16, 18, 11) {real, imag} */,
  {32'hbd4893b9, 32'hbdc23642} /* (16, 18, 10) {real, imag} */,
  {32'hbdb3fb90, 32'hbc4c8b3e} /* (16, 18, 9) {real, imag} */,
  {32'h3ca06d8a, 32'h3c9e2e14} /* (16, 18, 8) {real, imag} */,
  {32'h3dc2ac2a, 32'hbd266f57} /* (16, 18, 7) {real, imag} */,
  {32'h3d1598ac, 32'h3d903a11} /* (16, 18, 6) {real, imag} */,
  {32'hbd79c3bc, 32'hbd3e6b74} /* (16, 18, 5) {real, imag} */,
  {32'h3e183d4a, 32'hbce336e8} /* (16, 18, 4) {real, imag} */,
  {32'h3e82d715, 32'hbe0cf94c} /* (16, 18, 3) {real, imag} */,
  {32'hbeefc907, 32'hbdac0464} /* (16, 18, 2) {real, imag} */,
  {32'h3f4aa1e0, 32'h3d887656} /* (16, 18, 1) {real, imag} */,
  {32'h3f2d92d1, 32'h00000000} /* (16, 18, 0) {real, imag} */,
  {32'h3f6a1dd3, 32'hbde1133c} /* (16, 17, 31) {real, imag} */,
  {32'hbf197ade, 32'h3d7af27a} /* (16, 17, 30) {real, imag} */,
  {32'h3e9262bc, 32'hbda2c4d9} /* (16, 17, 29) {real, imag} */,
  {32'h3e3addec, 32'h3da2e3b7} /* (16, 17, 28) {real, imag} */,
  {32'hbe02bc64, 32'h3c5eeac8} /* (16, 17, 27) {real, imag} */,
  {32'hbbc1fde0, 32'hbde68f96} /* (16, 17, 26) {real, imag} */,
  {32'h3d2a47e5, 32'hbdb2e06d} /* (16, 17, 25) {real, imag} */,
  {32'h3de86a29, 32'h3dae4683} /* (16, 17, 24) {real, imag} */,
  {32'h3dba7213, 32'hbcb2f2e0} /* (16, 17, 23) {real, imag} */,
  {32'hbab855d0, 32'hbe055af8} /* (16, 17, 22) {real, imag} */,
  {32'hbd8d89fe, 32'h3e22673e} /* (16, 17, 21) {real, imag} */,
  {32'h3d33a17f, 32'h3d98e397} /* (16, 17, 20) {real, imag} */,
  {32'hbd305122, 32'hbd3c2f19} /* (16, 17, 19) {real, imag} */,
  {32'hbd20a2f6, 32'h3d462c5d} /* (16, 17, 18) {real, imag} */,
  {32'h3cfb4642, 32'h39d600c0} /* (16, 17, 17) {real, imag} */,
  {32'h3cf80378, 32'h00000000} /* (16, 17, 16) {real, imag} */,
  {32'h3cfb4642, 32'hb9d600c0} /* (16, 17, 15) {real, imag} */,
  {32'hbd20a2f6, 32'hbd462c5d} /* (16, 17, 14) {real, imag} */,
  {32'hbd305122, 32'h3d3c2f19} /* (16, 17, 13) {real, imag} */,
  {32'h3d33a17f, 32'hbd98e397} /* (16, 17, 12) {real, imag} */,
  {32'hbd8d89fe, 32'hbe22673e} /* (16, 17, 11) {real, imag} */,
  {32'hbab855d0, 32'h3e055af8} /* (16, 17, 10) {real, imag} */,
  {32'h3dba7213, 32'h3cb2f2e0} /* (16, 17, 9) {real, imag} */,
  {32'h3de86a29, 32'hbdae4683} /* (16, 17, 8) {real, imag} */,
  {32'h3d2a47e5, 32'h3db2e06d} /* (16, 17, 7) {real, imag} */,
  {32'hbbc1fde0, 32'h3de68f96} /* (16, 17, 6) {real, imag} */,
  {32'hbe02bc64, 32'hbc5eeac8} /* (16, 17, 5) {real, imag} */,
  {32'h3e3addec, 32'hbda2e3b7} /* (16, 17, 4) {real, imag} */,
  {32'h3e9262bc, 32'h3da2c4d9} /* (16, 17, 3) {real, imag} */,
  {32'hbf197ade, 32'hbd7af27a} /* (16, 17, 2) {real, imag} */,
  {32'h3f6a1dd3, 32'h3de1133c} /* (16, 17, 1) {real, imag} */,
  {32'h3f36565e, 32'h00000000} /* (16, 17, 0) {real, imag} */,
  {32'h3f780559, 32'hbd0296a0} /* (16, 16, 31) {real, imag} */,
  {32'hbf01073f, 32'h3dad03ca} /* (16, 16, 30) {real, imag} */,
  {32'h3e0b83d3, 32'hbd8a6e34} /* (16, 16, 29) {real, imag} */,
  {32'h3dddeeb9, 32'h3da13f5b} /* (16, 16, 28) {real, imag} */,
  {32'hbe5c9e1d, 32'h3e21a39e} /* (16, 16, 27) {real, imag} */,
  {32'hbd6a7d40, 32'h3ca5ef96} /* (16, 16, 26) {real, imag} */,
  {32'h3d9b5a23, 32'hbcbba47e} /* (16, 16, 25) {real, imag} */,
  {32'hbbe42a40, 32'h3b05a5c0} /* (16, 16, 24) {real, imag} */,
  {32'h3cfcd110, 32'hbd277a71} /* (16, 16, 23) {real, imag} */,
  {32'hbcceb671, 32'hbd173899} /* (16, 16, 22) {real, imag} */,
  {32'hbdbf7a77, 32'h3cf03dc4} /* (16, 16, 21) {real, imag} */,
  {32'h3d89d87e, 32'hbe164d26} /* (16, 16, 20) {real, imag} */,
  {32'h3d7318ae, 32'h3d3b1f50} /* (16, 16, 19) {real, imag} */,
  {32'hbdbff628, 32'hbd03c9ea} /* (16, 16, 18) {real, imag} */,
  {32'h3c855448, 32'h3ca33db3} /* (16, 16, 17) {real, imag} */,
  {32'hbd221375, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h3c855448, 32'hbca33db3} /* (16, 16, 15) {real, imag} */,
  {32'hbdbff628, 32'h3d03c9ea} /* (16, 16, 14) {real, imag} */,
  {32'h3d7318ae, 32'hbd3b1f50} /* (16, 16, 13) {real, imag} */,
  {32'h3d89d87e, 32'h3e164d26} /* (16, 16, 12) {real, imag} */,
  {32'hbdbf7a77, 32'hbcf03dc4} /* (16, 16, 11) {real, imag} */,
  {32'hbcceb671, 32'h3d173899} /* (16, 16, 10) {real, imag} */,
  {32'h3cfcd110, 32'h3d277a71} /* (16, 16, 9) {real, imag} */,
  {32'hbbe42a40, 32'hbb05a5c0} /* (16, 16, 8) {real, imag} */,
  {32'h3d9b5a23, 32'h3cbba47e} /* (16, 16, 7) {real, imag} */,
  {32'hbd6a7d40, 32'hbca5ef96} /* (16, 16, 6) {real, imag} */,
  {32'hbe5c9e1d, 32'hbe21a39e} /* (16, 16, 5) {real, imag} */,
  {32'h3dddeeb9, 32'hbda13f5b} /* (16, 16, 4) {real, imag} */,
  {32'h3e0b83d3, 32'h3d8a6e34} /* (16, 16, 3) {real, imag} */,
  {32'hbf01073f, 32'hbdad03ca} /* (16, 16, 2) {real, imag} */,
  {32'h3f780559, 32'h3d0296a0} /* (16, 16, 1) {real, imag} */,
  {32'h3f047db0, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h3f4df0f1, 32'h3e2cfd26} /* (16, 15, 31) {real, imag} */,
  {32'hbee9459c, 32'h3d2955b6} /* (16, 15, 30) {real, imag} */,
  {32'h3e17a0aa, 32'hbd8a6d39} /* (16, 15, 29) {real, imag} */,
  {32'hbd467be6, 32'h3e025c90} /* (16, 15, 28) {real, imag} */,
  {32'hbe49b074, 32'h3e07b424} /* (16, 15, 27) {real, imag} */,
  {32'h3cb84f22, 32'h3daaf756} /* (16, 15, 26) {real, imag} */,
  {32'h3c94f55a, 32'hbd9d436b} /* (16, 15, 25) {real, imag} */,
  {32'hbcb2c324, 32'h3c0fef68} /* (16, 15, 24) {real, imag} */,
  {32'h3c9c2ebc, 32'h39eab7a0} /* (16, 15, 23) {real, imag} */,
  {32'h3d6ef5aa, 32'hbd2a047e} /* (16, 15, 22) {real, imag} */,
  {32'hbce3e8df, 32'h3d0dceaa} /* (16, 15, 21) {real, imag} */,
  {32'hbd768e75, 32'h3aee1500} /* (16, 15, 20) {real, imag} */,
  {32'hbc865981, 32'hbc48ca70} /* (16, 15, 19) {real, imag} */,
  {32'h3cd96cc9, 32'hbafc7420} /* (16, 15, 18) {real, imag} */,
  {32'h3c07ab4c, 32'h3d4d19a0} /* (16, 15, 17) {real, imag} */,
  {32'hbc11c2f1, 32'h00000000} /* (16, 15, 16) {real, imag} */,
  {32'h3c07ab4c, 32'hbd4d19a0} /* (16, 15, 15) {real, imag} */,
  {32'h3cd96cc9, 32'h3afc7420} /* (16, 15, 14) {real, imag} */,
  {32'hbc865981, 32'h3c48ca70} /* (16, 15, 13) {real, imag} */,
  {32'hbd768e75, 32'hbaee1500} /* (16, 15, 12) {real, imag} */,
  {32'hbce3e8df, 32'hbd0dceaa} /* (16, 15, 11) {real, imag} */,
  {32'h3d6ef5aa, 32'h3d2a047e} /* (16, 15, 10) {real, imag} */,
  {32'h3c9c2ebc, 32'hb9eab7a0} /* (16, 15, 9) {real, imag} */,
  {32'hbcb2c324, 32'hbc0fef68} /* (16, 15, 8) {real, imag} */,
  {32'h3c94f55a, 32'h3d9d436b} /* (16, 15, 7) {real, imag} */,
  {32'h3cb84f22, 32'hbdaaf756} /* (16, 15, 6) {real, imag} */,
  {32'hbe49b074, 32'hbe07b424} /* (16, 15, 5) {real, imag} */,
  {32'hbd467be6, 32'hbe025c90} /* (16, 15, 4) {real, imag} */,
  {32'h3e17a0aa, 32'h3d8a6d39} /* (16, 15, 3) {real, imag} */,
  {32'hbee9459c, 32'hbd2955b6} /* (16, 15, 2) {real, imag} */,
  {32'h3f4df0f1, 32'hbe2cfd26} /* (16, 15, 1) {real, imag} */,
  {32'h3f22978e, 32'h00000000} /* (16, 15, 0) {real, imag} */,
  {32'h3f24a678, 32'h3e39e65d} /* (16, 14, 31) {real, imag} */,
  {32'hbebf37d1, 32'h3da64b56} /* (16, 14, 30) {real, imag} */,
  {32'h3da13704, 32'h3c014ec0} /* (16, 14, 29) {real, imag} */,
  {32'h3da76594, 32'h3c863b48} /* (16, 14, 28) {real, imag} */,
  {32'hbe86629a, 32'h3d134048} /* (16, 14, 27) {real, imag} */,
  {32'h3d857a2a, 32'h3c984c2f} /* (16, 14, 26) {real, imag} */,
  {32'h3ccd4360, 32'hbe0003e4} /* (16, 14, 25) {real, imag} */,
  {32'hbd8f32ba, 32'h3d36433a} /* (16, 14, 24) {real, imag} */,
  {32'h3cc90014, 32'hbb980a7d} /* (16, 14, 23) {real, imag} */,
  {32'hbba73728, 32'h3c5a7d30} /* (16, 14, 22) {real, imag} */,
  {32'h3d8a500a, 32'h3d13d935} /* (16, 14, 21) {real, imag} */,
  {32'h3b02c1e8, 32'hbb1b72d0} /* (16, 14, 20) {real, imag} */,
  {32'h3d445da4, 32'hbc99e345} /* (16, 14, 19) {real, imag} */,
  {32'hbd01e688, 32'hbcf6b6d0} /* (16, 14, 18) {real, imag} */,
  {32'hbd73f7a3, 32'hbcaf9af3} /* (16, 14, 17) {real, imag} */,
  {32'hbc75fa00, 32'h00000000} /* (16, 14, 16) {real, imag} */,
  {32'hbd73f7a3, 32'h3caf9af3} /* (16, 14, 15) {real, imag} */,
  {32'hbd01e688, 32'h3cf6b6d0} /* (16, 14, 14) {real, imag} */,
  {32'h3d445da4, 32'h3c99e345} /* (16, 14, 13) {real, imag} */,
  {32'h3b02c1e8, 32'h3b1b72d0} /* (16, 14, 12) {real, imag} */,
  {32'h3d8a500a, 32'hbd13d935} /* (16, 14, 11) {real, imag} */,
  {32'hbba73728, 32'hbc5a7d30} /* (16, 14, 10) {real, imag} */,
  {32'h3cc90014, 32'h3b980a7d} /* (16, 14, 9) {real, imag} */,
  {32'hbd8f32ba, 32'hbd36433a} /* (16, 14, 8) {real, imag} */,
  {32'h3ccd4360, 32'h3e0003e4} /* (16, 14, 7) {real, imag} */,
  {32'h3d857a2a, 32'hbc984c2f} /* (16, 14, 6) {real, imag} */,
  {32'hbe86629a, 32'hbd134048} /* (16, 14, 5) {real, imag} */,
  {32'h3da76594, 32'hbc863b48} /* (16, 14, 4) {real, imag} */,
  {32'h3da13704, 32'hbc014ec0} /* (16, 14, 3) {real, imag} */,
  {32'hbebf37d1, 32'hbda64b56} /* (16, 14, 2) {real, imag} */,
  {32'h3f24a678, 32'hbe39e65d} /* (16, 14, 1) {real, imag} */,
  {32'h3f15a1cb, 32'h00000000} /* (16, 14, 0) {real, imag} */,
  {32'h3f2bb184, 32'h3e455032} /* (16, 13, 31) {real, imag} */,
  {32'hbea33508, 32'h3da01623} /* (16, 13, 30) {real, imag} */,
  {32'hbd537f90, 32'h3d418122} /* (16, 13, 29) {real, imag} */,
  {32'h3de219a8, 32'h3dc0a6aa} /* (16, 13, 28) {real, imag} */,
  {32'hbe45b854, 32'h3d00665c} /* (16, 13, 27) {real, imag} */,
  {32'hbdb31e6e, 32'hbcd655fa} /* (16, 13, 26) {real, imag} */,
  {32'hbd90754c, 32'hbdd6a36f} /* (16, 13, 25) {real, imag} */,
  {32'hbd5d9748, 32'hbc23d8e0} /* (16, 13, 24) {real, imag} */,
  {32'h3cd8b0b2, 32'h3d00f784} /* (16, 13, 23) {real, imag} */,
  {32'h3d507656, 32'hba6cd4b0} /* (16, 13, 22) {real, imag} */,
  {32'h3b13f4c4, 32'h3d597132} /* (16, 13, 21) {real, imag} */,
  {32'h3d3e83fc, 32'hbcdbba6e} /* (16, 13, 20) {real, imag} */,
  {32'h3c288294, 32'hbaf536bc} /* (16, 13, 19) {real, imag} */,
  {32'hbd3e86c2, 32'h3d90dd4f} /* (16, 13, 18) {real, imag} */,
  {32'hbd54d5d6, 32'hbc914caa} /* (16, 13, 17) {real, imag} */,
  {32'hbd097b90, 32'h00000000} /* (16, 13, 16) {real, imag} */,
  {32'hbd54d5d6, 32'h3c914caa} /* (16, 13, 15) {real, imag} */,
  {32'hbd3e86c2, 32'hbd90dd4f} /* (16, 13, 14) {real, imag} */,
  {32'h3c288294, 32'h3af536bc} /* (16, 13, 13) {real, imag} */,
  {32'h3d3e83fc, 32'h3cdbba6e} /* (16, 13, 12) {real, imag} */,
  {32'h3b13f4c4, 32'hbd597132} /* (16, 13, 11) {real, imag} */,
  {32'h3d507656, 32'h3a6cd4b0} /* (16, 13, 10) {real, imag} */,
  {32'h3cd8b0b2, 32'hbd00f784} /* (16, 13, 9) {real, imag} */,
  {32'hbd5d9748, 32'h3c23d8e0} /* (16, 13, 8) {real, imag} */,
  {32'hbd90754c, 32'h3dd6a36f} /* (16, 13, 7) {real, imag} */,
  {32'hbdb31e6e, 32'h3cd655fa} /* (16, 13, 6) {real, imag} */,
  {32'hbe45b854, 32'hbd00665c} /* (16, 13, 5) {real, imag} */,
  {32'h3de219a8, 32'hbdc0a6aa} /* (16, 13, 4) {real, imag} */,
  {32'hbd537f90, 32'hbd418122} /* (16, 13, 3) {real, imag} */,
  {32'hbea33508, 32'hbda01623} /* (16, 13, 2) {real, imag} */,
  {32'h3f2bb184, 32'hbe455032} /* (16, 13, 1) {real, imag} */,
  {32'h3f4010bd, 32'h00000000} /* (16, 13, 0) {real, imag} */,
  {32'h3f182680, 32'h3e1bb5c3} /* (16, 12, 31) {real, imag} */,
  {32'hbec138bc, 32'h3dc46d1f} /* (16, 12, 30) {real, imag} */,
  {32'h3daf6a29, 32'h3d9b1f3f} /* (16, 12, 29) {real, imag} */,
  {32'h3beaa480, 32'h3dc22e89} /* (16, 12, 28) {real, imag} */,
  {32'hbda919a2, 32'h3da8ce1f} /* (16, 12, 27) {real, imag} */,
  {32'h3d5ee502, 32'h3d5a9ee2} /* (16, 12, 26) {real, imag} */,
  {32'hbdacd686, 32'hbc8db5b2} /* (16, 12, 25) {real, imag} */,
  {32'hbd2eeee0, 32'h3e0b3c16} /* (16, 12, 24) {real, imag} */,
  {32'h3c7a0858, 32'hbdb155b2} /* (16, 12, 23) {real, imag} */,
  {32'h3c5830b0, 32'h3d3e0582} /* (16, 12, 22) {real, imag} */,
  {32'h3b4cf240, 32'h3d095291} /* (16, 12, 21) {real, imag} */,
  {32'h3c9c35e4, 32'hbd23c2e1} /* (16, 12, 20) {real, imag} */,
  {32'hbd193a68, 32'hbd1b45b4} /* (16, 12, 19) {real, imag} */,
  {32'hb9723bc0, 32'hbda20248} /* (16, 12, 18) {real, imag} */,
  {32'h3d5102ed, 32'hbd810332} /* (16, 12, 17) {real, imag} */,
  {32'hbd2d94bc, 32'h00000000} /* (16, 12, 16) {real, imag} */,
  {32'h3d5102ed, 32'h3d810332} /* (16, 12, 15) {real, imag} */,
  {32'hb9723bc0, 32'h3da20248} /* (16, 12, 14) {real, imag} */,
  {32'hbd193a68, 32'h3d1b45b4} /* (16, 12, 13) {real, imag} */,
  {32'h3c9c35e4, 32'h3d23c2e1} /* (16, 12, 12) {real, imag} */,
  {32'h3b4cf240, 32'hbd095291} /* (16, 12, 11) {real, imag} */,
  {32'h3c5830b0, 32'hbd3e0582} /* (16, 12, 10) {real, imag} */,
  {32'h3c7a0858, 32'h3db155b2} /* (16, 12, 9) {real, imag} */,
  {32'hbd2eeee0, 32'hbe0b3c16} /* (16, 12, 8) {real, imag} */,
  {32'hbdacd686, 32'h3c8db5b2} /* (16, 12, 7) {real, imag} */,
  {32'h3d5ee502, 32'hbd5a9ee2} /* (16, 12, 6) {real, imag} */,
  {32'hbda919a2, 32'hbda8ce1f} /* (16, 12, 5) {real, imag} */,
  {32'h3beaa480, 32'hbdc22e89} /* (16, 12, 4) {real, imag} */,
  {32'h3daf6a29, 32'hbd9b1f3f} /* (16, 12, 3) {real, imag} */,
  {32'hbec138bc, 32'hbdc46d1f} /* (16, 12, 2) {real, imag} */,
  {32'h3f182680, 32'hbe1bb5c3} /* (16, 12, 1) {real, imag} */,
  {32'h3f6a6db6, 32'h00000000} /* (16, 12, 0) {real, imag} */,
  {32'h3ea17cfa, 32'h3ea1fc44} /* (16, 11, 31) {real, imag} */,
  {32'hbe7190ea, 32'h3e090805} /* (16, 11, 30) {real, imag} */,
  {32'h3d4eff25, 32'hbd8bf662} /* (16, 11, 29) {real, imag} */,
  {32'hbcfeeaad, 32'hbe0c9656} /* (16, 11, 28) {real, imag} */,
  {32'hbd989473, 32'h3d13c534} /* (16, 11, 27) {real, imag} */,
  {32'h3dc01bde, 32'h3da4039e} /* (16, 11, 26) {real, imag} */,
  {32'h3d2f02bf, 32'hbdddd486} /* (16, 11, 25) {real, imag} */,
  {32'h3ce3b18f, 32'h3e12878f} /* (16, 11, 24) {real, imag} */,
  {32'hbce89969, 32'hbd5ee5e2} /* (16, 11, 23) {real, imag} */,
  {32'hbe1c6f16, 32'h3ca9e8ae} /* (16, 11, 22) {real, imag} */,
  {32'h3d4a1391, 32'h3aef7a08} /* (16, 11, 21) {real, imag} */,
  {32'h3dfa79a8, 32'h3d5018a7} /* (16, 11, 20) {real, imag} */,
  {32'hbd10d0fd, 32'h3d72a1bd} /* (16, 11, 19) {real, imag} */,
  {32'h3aebc318, 32'h3cf4993e} /* (16, 11, 18) {real, imag} */,
  {32'h3d48e594, 32'hbd3604cb} /* (16, 11, 17) {real, imag} */,
  {32'h3da1be04, 32'h00000000} /* (16, 11, 16) {real, imag} */,
  {32'h3d48e594, 32'h3d3604cb} /* (16, 11, 15) {real, imag} */,
  {32'h3aebc318, 32'hbcf4993e} /* (16, 11, 14) {real, imag} */,
  {32'hbd10d0fd, 32'hbd72a1bd} /* (16, 11, 13) {real, imag} */,
  {32'h3dfa79a8, 32'hbd5018a7} /* (16, 11, 12) {real, imag} */,
  {32'h3d4a1391, 32'hbaef7a08} /* (16, 11, 11) {real, imag} */,
  {32'hbe1c6f16, 32'hbca9e8ae} /* (16, 11, 10) {real, imag} */,
  {32'hbce89969, 32'h3d5ee5e2} /* (16, 11, 9) {real, imag} */,
  {32'h3ce3b18f, 32'hbe12878f} /* (16, 11, 8) {real, imag} */,
  {32'h3d2f02bf, 32'h3dddd486} /* (16, 11, 7) {real, imag} */,
  {32'h3dc01bde, 32'hbda4039e} /* (16, 11, 6) {real, imag} */,
  {32'hbd989473, 32'hbd13c534} /* (16, 11, 5) {real, imag} */,
  {32'hbcfeeaad, 32'h3e0c9656} /* (16, 11, 4) {real, imag} */,
  {32'h3d4eff25, 32'h3d8bf662} /* (16, 11, 3) {real, imag} */,
  {32'hbe7190ea, 32'hbe090805} /* (16, 11, 2) {real, imag} */,
  {32'h3ea17cfa, 32'hbea1fc44} /* (16, 11, 1) {real, imag} */,
  {32'h3f5d321b, 32'h00000000} /* (16, 11, 0) {real, imag} */,
  {32'hbeb2aedd, 32'h3eb4bc28} /* (16, 10, 31) {real, imag} */,
  {32'h3e622238, 32'h3dba361e} /* (16, 10, 30) {real, imag} */,
  {32'hbd9f11c0, 32'hbd33fbe2} /* (16, 10, 29) {real, imag} */,
  {32'hbcd461c0, 32'hbd80ce1c} /* (16, 10, 28) {real, imag} */,
  {32'hbca99512, 32'hbd062650} /* (16, 10, 27) {real, imag} */,
  {32'hbd07671a, 32'h3d1f1426} /* (16, 10, 26) {real, imag} */,
  {32'hbc0f0cfe, 32'h3ddaf137} /* (16, 10, 25) {real, imag} */,
  {32'h3aa27ce0, 32'h3be06f80} /* (16, 10, 24) {real, imag} */,
  {32'hb9fcb8c0, 32'h3d8b68fe} /* (16, 10, 23) {real, imag} */,
  {32'h3d284e9c, 32'hbdbbe15c} /* (16, 10, 22) {real, imag} */,
  {32'h3d1f7240, 32'hba80bb20} /* (16, 10, 21) {real, imag} */,
  {32'h3cdbcec6, 32'hbc6c1ba8} /* (16, 10, 20) {real, imag} */,
  {32'h3d8c4b25, 32'h3dc589bf} /* (16, 10, 19) {real, imag} */,
  {32'hbcf164fe, 32'hbd1d4769} /* (16, 10, 18) {real, imag} */,
  {32'h3d0139ac, 32'hbd0df39a} /* (16, 10, 17) {real, imag} */,
  {32'h3d3397c3, 32'h00000000} /* (16, 10, 16) {real, imag} */,
  {32'h3d0139ac, 32'h3d0df39a} /* (16, 10, 15) {real, imag} */,
  {32'hbcf164fe, 32'h3d1d4769} /* (16, 10, 14) {real, imag} */,
  {32'h3d8c4b25, 32'hbdc589bf} /* (16, 10, 13) {real, imag} */,
  {32'h3cdbcec6, 32'h3c6c1ba8} /* (16, 10, 12) {real, imag} */,
  {32'h3d1f7240, 32'h3a80bb20} /* (16, 10, 11) {real, imag} */,
  {32'h3d284e9c, 32'h3dbbe15c} /* (16, 10, 10) {real, imag} */,
  {32'hb9fcb8c0, 32'hbd8b68fe} /* (16, 10, 9) {real, imag} */,
  {32'h3aa27ce0, 32'hbbe06f80} /* (16, 10, 8) {real, imag} */,
  {32'hbc0f0cfe, 32'hbddaf137} /* (16, 10, 7) {real, imag} */,
  {32'hbd07671a, 32'hbd1f1426} /* (16, 10, 6) {real, imag} */,
  {32'hbca99512, 32'h3d062650} /* (16, 10, 5) {real, imag} */,
  {32'hbcd461c0, 32'h3d80ce1c} /* (16, 10, 4) {real, imag} */,
  {32'hbd9f11c0, 32'h3d33fbe2} /* (16, 10, 3) {real, imag} */,
  {32'h3e622238, 32'hbdba361e} /* (16, 10, 2) {real, imag} */,
  {32'hbeb2aedd, 32'hbeb4bc28} /* (16, 10, 1) {real, imag} */,
  {32'h3e8b907e, 32'h00000000} /* (16, 10, 0) {real, imag} */,
  {32'hbf511574, 32'h3e9baf47} /* (16, 9, 31) {real, imag} */,
  {32'h3eda9751, 32'hbb9cfdbc} /* (16, 9, 30) {real, imag} */,
  {32'hbe188913, 32'h3d847bed} /* (16, 9, 29) {real, imag} */,
  {32'h3ba63480, 32'h3d358a78} /* (16, 9, 28) {real, imag} */,
  {32'h3d75dded, 32'hbc95f2d8} /* (16, 9, 27) {real, imag} */,
  {32'h3c85f858, 32'hbc020ea2} /* (16, 9, 26) {real, imag} */,
  {32'hbdf702f6, 32'h3df831da} /* (16, 9, 25) {real, imag} */,
  {32'h3d337d25, 32'hbd2dbf18} /* (16, 9, 24) {real, imag} */,
  {32'h3da70b15, 32'hbd21fce3} /* (16, 9, 23) {real, imag} */,
  {32'h3d41ff82, 32'hbc89e844} /* (16, 9, 22) {real, imag} */,
  {32'h3d99a9b1, 32'h3c05c4b8} /* (16, 9, 21) {real, imag} */,
  {32'hbd8cdd62, 32'hbc9cdbbc} /* (16, 9, 20) {real, imag} */,
  {32'hbdc07719, 32'hbccc452a} /* (16, 9, 19) {real, imag} */,
  {32'hbd8f0ce7, 32'h3ca12a7c} /* (16, 9, 18) {real, imag} */,
  {32'h3d1f2f44, 32'h3c95b1ce} /* (16, 9, 17) {real, imag} */,
  {32'hbcb93228, 32'h00000000} /* (16, 9, 16) {real, imag} */,
  {32'h3d1f2f44, 32'hbc95b1ce} /* (16, 9, 15) {real, imag} */,
  {32'hbd8f0ce7, 32'hbca12a7c} /* (16, 9, 14) {real, imag} */,
  {32'hbdc07719, 32'h3ccc452a} /* (16, 9, 13) {real, imag} */,
  {32'hbd8cdd62, 32'h3c9cdbbc} /* (16, 9, 12) {real, imag} */,
  {32'h3d99a9b1, 32'hbc05c4b8} /* (16, 9, 11) {real, imag} */,
  {32'h3d41ff82, 32'h3c89e844} /* (16, 9, 10) {real, imag} */,
  {32'h3da70b15, 32'h3d21fce3} /* (16, 9, 9) {real, imag} */,
  {32'h3d337d25, 32'h3d2dbf18} /* (16, 9, 8) {real, imag} */,
  {32'hbdf702f6, 32'hbdf831da} /* (16, 9, 7) {real, imag} */,
  {32'h3c85f858, 32'h3c020ea2} /* (16, 9, 6) {real, imag} */,
  {32'h3d75dded, 32'h3c95f2d8} /* (16, 9, 5) {real, imag} */,
  {32'h3ba63480, 32'hbd358a78} /* (16, 9, 4) {real, imag} */,
  {32'hbe188913, 32'hbd847bed} /* (16, 9, 3) {real, imag} */,
  {32'h3eda9751, 32'h3b9cfdbc} /* (16, 9, 2) {real, imag} */,
  {32'hbf511574, 32'hbe9baf47} /* (16, 9, 1) {real, imag} */,
  {32'hbe09ca3c, 32'h00000000} /* (16, 9, 0) {real, imag} */,
  {32'hbf83e942, 32'h3eaa6950} /* (16, 8, 31) {real, imag} */,
  {32'h3eaccb02, 32'hbe095eae} /* (16, 8, 30) {real, imag} */,
  {32'hbe80556a, 32'hbc278910} /* (16, 8, 29) {real, imag} */,
  {32'hbd8e7eb8, 32'h3c643790} /* (16, 8, 28) {real, imag} */,
  {32'hbbf4ad80, 32'hbc04d8f0} /* (16, 8, 27) {real, imag} */,
  {32'hbdfec4fe, 32'h3d16cfb8} /* (16, 8, 26) {real, imag} */,
  {32'hbda40c96, 32'hbdaacc40} /* (16, 8, 25) {real, imag} */,
  {32'h3d27b3b3, 32'hbdfe5492} /* (16, 8, 24) {real, imag} */,
  {32'hbcc82bd0, 32'hbdbc5081} /* (16, 8, 23) {real, imag} */,
  {32'hbbe3d7d0, 32'hbd4c51ec} /* (16, 8, 22) {real, imag} */,
  {32'hbdd88d8b, 32'hbcd8a415} /* (16, 8, 21) {real, imag} */,
  {32'h3d6e0350, 32'h3d92ef16} /* (16, 8, 20) {real, imag} */,
  {32'hbdb21308, 32'hbd46daca} /* (16, 8, 19) {real, imag} */,
  {32'hbd173112, 32'h3d0030bd} /* (16, 8, 18) {real, imag} */,
  {32'hbb413784, 32'hbd2969a7} /* (16, 8, 17) {real, imag} */,
  {32'h3d048f90, 32'h00000000} /* (16, 8, 16) {real, imag} */,
  {32'hbb413784, 32'h3d2969a7} /* (16, 8, 15) {real, imag} */,
  {32'hbd173112, 32'hbd0030bd} /* (16, 8, 14) {real, imag} */,
  {32'hbdb21308, 32'h3d46daca} /* (16, 8, 13) {real, imag} */,
  {32'h3d6e0350, 32'hbd92ef16} /* (16, 8, 12) {real, imag} */,
  {32'hbdd88d8b, 32'h3cd8a415} /* (16, 8, 11) {real, imag} */,
  {32'hbbe3d7d0, 32'h3d4c51ec} /* (16, 8, 10) {real, imag} */,
  {32'hbcc82bd0, 32'h3dbc5081} /* (16, 8, 9) {real, imag} */,
  {32'h3d27b3b3, 32'h3dfe5492} /* (16, 8, 8) {real, imag} */,
  {32'hbda40c96, 32'h3daacc40} /* (16, 8, 7) {real, imag} */,
  {32'hbdfec4fe, 32'hbd16cfb8} /* (16, 8, 6) {real, imag} */,
  {32'hbbf4ad80, 32'h3c04d8f0} /* (16, 8, 5) {real, imag} */,
  {32'hbd8e7eb8, 32'hbc643790} /* (16, 8, 4) {real, imag} */,
  {32'hbe80556a, 32'h3c278910} /* (16, 8, 3) {real, imag} */,
  {32'h3eaccb02, 32'h3e095eae} /* (16, 8, 2) {real, imag} */,
  {32'hbf83e942, 32'hbeaa6950} /* (16, 8, 1) {real, imag} */,
  {32'hbea6b5d9, 32'h00000000} /* (16, 8, 0) {real, imag} */,
  {32'hbf86f407, 32'h3ef0f183} /* (16, 7, 31) {real, imag} */,
  {32'h3e8b976d, 32'hbe690d8a} /* (16, 7, 30) {real, imag} */,
  {32'hbda04ad0, 32'h3d18221a} /* (16, 7, 29) {real, imag} */,
  {32'hbdc399c1, 32'hbcb4fd38} /* (16, 7, 28) {real, imag} */,
  {32'h3dbff836, 32'hbd19e48c} /* (16, 7, 27) {real, imag} */,
  {32'hbd0c1c7c, 32'h3e1f75bf} /* (16, 7, 26) {real, imag} */,
  {32'hbc114edc, 32'hbcec2e3d} /* (16, 7, 25) {real, imag} */,
  {32'h3c3cd7a0, 32'hbd2947b4} /* (16, 7, 24) {real, imag} */,
  {32'h3d494c98, 32'hbd73e237} /* (16, 7, 23) {real, imag} */,
  {32'hbc86d190, 32'h3e025994} /* (16, 7, 22) {real, imag} */,
  {32'h3d174173, 32'hbe206349} /* (16, 7, 21) {real, imag} */,
  {32'h3ded9cf8, 32'h3cbcfd29} /* (16, 7, 20) {real, imag} */,
  {32'hbc9a41b9, 32'hbc7fdc7e} /* (16, 7, 19) {real, imag} */,
  {32'h3cde0806, 32'h3c96ab49} /* (16, 7, 18) {real, imag} */,
  {32'h3c92a61e, 32'h3da5bd02} /* (16, 7, 17) {real, imag} */,
  {32'hbe10dd18, 32'h00000000} /* (16, 7, 16) {real, imag} */,
  {32'h3c92a61e, 32'hbda5bd02} /* (16, 7, 15) {real, imag} */,
  {32'h3cde0806, 32'hbc96ab49} /* (16, 7, 14) {real, imag} */,
  {32'hbc9a41b9, 32'h3c7fdc7e} /* (16, 7, 13) {real, imag} */,
  {32'h3ded9cf8, 32'hbcbcfd29} /* (16, 7, 12) {real, imag} */,
  {32'h3d174173, 32'h3e206349} /* (16, 7, 11) {real, imag} */,
  {32'hbc86d190, 32'hbe025994} /* (16, 7, 10) {real, imag} */,
  {32'h3d494c98, 32'h3d73e237} /* (16, 7, 9) {real, imag} */,
  {32'h3c3cd7a0, 32'h3d2947b4} /* (16, 7, 8) {real, imag} */,
  {32'hbc114edc, 32'h3cec2e3d} /* (16, 7, 7) {real, imag} */,
  {32'hbd0c1c7c, 32'hbe1f75bf} /* (16, 7, 6) {real, imag} */,
  {32'h3dbff836, 32'h3d19e48c} /* (16, 7, 5) {real, imag} */,
  {32'hbdc399c1, 32'h3cb4fd38} /* (16, 7, 4) {real, imag} */,
  {32'hbda04ad0, 32'hbd18221a} /* (16, 7, 3) {real, imag} */,
  {32'h3e8b976d, 32'h3e690d8a} /* (16, 7, 2) {real, imag} */,
  {32'hbf86f407, 32'hbef0f183} /* (16, 7, 1) {real, imag} */,
  {32'hbf31f69c, 32'h00000000} /* (16, 7, 0) {real, imag} */,
  {32'hbf8a543d, 32'h3f080290} /* (16, 6, 31) {real, imag} */,
  {32'h3e60c70e, 32'hbe31368c} /* (16, 6, 30) {real, imag} */,
  {32'hbdc6d490, 32'hbc113d08} /* (16, 6, 29) {real, imag} */,
  {32'hbd51cabc, 32'hbd0fc19d} /* (16, 6, 28) {real, imag} */,
  {32'h3da95600, 32'hbdee5d04} /* (16, 6, 27) {real, imag} */,
  {32'h3d0ce9c0, 32'hbcbf2ace} /* (16, 6, 26) {real, imag} */,
  {32'h3cc2013d, 32'h3b2ee7b8} /* (16, 6, 25) {real, imag} */,
  {32'h3d3a49ae, 32'hbe1090c5} /* (16, 6, 24) {real, imag} */,
  {32'hbb3bbb20, 32'hbc911724} /* (16, 6, 23) {real, imag} */,
  {32'hbd20a72f, 32'h3db898d1} /* (16, 6, 22) {real, imag} */,
  {32'hbd8f495a, 32'hbd23afe5} /* (16, 6, 21) {real, imag} */,
  {32'h3dd50212, 32'hbd2373aa} /* (16, 6, 20) {real, imag} */,
  {32'h3d761dc9, 32'h3d65719a} /* (16, 6, 19) {real, imag} */,
  {32'h3c4f61d5, 32'hbd4bdab8} /* (16, 6, 18) {real, imag} */,
  {32'h3d34a941, 32'h3cba5d78} /* (16, 6, 17) {real, imag} */,
  {32'hbbe0c320, 32'h00000000} /* (16, 6, 16) {real, imag} */,
  {32'h3d34a941, 32'hbcba5d78} /* (16, 6, 15) {real, imag} */,
  {32'h3c4f61d5, 32'h3d4bdab8} /* (16, 6, 14) {real, imag} */,
  {32'h3d761dc9, 32'hbd65719a} /* (16, 6, 13) {real, imag} */,
  {32'h3dd50212, 32'h3d2373aa} /* (16, 6, 12) {real, imag} */,
  {32'hbd8f495a, 32'h3d23afe5} /* (16, 6, 11) {real, imag} */,
  {32'hbd20a72f, 32'hbdb898d1} /* (16, 6, 10) {real, imag} */,
  {32'hbb3bbb20, 32'h3c911724} /* (16, 6, 9) {real, imag} */,
  {32'h3d3a49ae, 32'h3e1090c5} /* (16, 6, 8) {real, imag} */,
  {32'h3cc2013d, 32'hbb2ee7b8} /* (16, 6, 7) {real, imag} */,
  {32'h3d0ce9c0, 32'h3cbf2ace} /* (16, 6, 6) {real, imag} */,
  {32'h3da95600, 32'h3dee5d04} /* (16, 6, 5) {real, imag} */,
  {32'hbd51cabc, 32'h3d0fc19d} /* (16, 6, 4) {real, imag} */,
  {32'hbdc6d490, 32'h3c113d08} /* (16, 6, 3) {real, imag} */,
  {32'h3e60c70e, 32'h3e31368c} /* (16, 6, 2) {real, imag} */,
  {32'hbf8a543d, 32'hbf080290} /* (16, 6, 1) {real, imag} */,
  {32'hbf3a5c44, 32'h00000000} /* (16, 6, 0) {real, imag} */,
  {32'hbf7f8c66, 32'h3f456861} /* (16, 5, 31) {real, imag} */,
  {32'hbdb7241e, 32'hbe8849ac} /* (16, 5, 30) {real, imag} */,
  {32'hbdb138b0, 32'hbd940ea4} /* (16, 5, 29) {real, imag} */,
  {32'h3df29c62, 32'hbdc99de0} /* (16, 5, 28) {real, imag} */,
  {32'h3e2c694c, 32'hbc9d63ce} /* (16, 5, 27) {real, imag} */,
  {32'hbd00d67e, 32'hbd99e81b} /* (16, 5, 26) {real, imag} */,
  {32'h3e076c07, 32'h3d0ec2b2} /* (16, 5, 25) {real, imag} */,
  {32'h3d9afc66, 32'hbd3254f6} /* (16, 5, 24) {real, imag} */,
  {32'h3cb4f82b, 32'hbc9b306d} /* (16, 5, 23) {real, imag} */,
  {32'h3d5484e4, 32'hbd48d8dc} /* (16, 5, 22) {real, imag} */,
  {32'hbd9088aa, 32'hba7dd180} /* (16, 5, 21) {real, imag} */,
  {32'hbaba1ab8, 32'h3d714521} /* (16, 5, 20) {real, imag} */,
  {32'h3d5be344, 32'hbd7c2070} /* (16, 5, 19) {real, imag} */,
  {32'hbd010bef, 32'hbcd85924} /* (16, 5, 18) {real, imag} */,
  {32'hbd6e16ac, 32'hbd6d7ec4} /* (16, 5, 17) {real, imag} */,
  {32'hbc178f7b, 32'h00000000} /* (16, 5, 16) {real, imag} */,
  {32'hbd6e16ac, 32'h3d6d7ec4} /* (16, 5, 15) {real, imag} */,
  {32'hbd010bef, 32'h3cd85924} /* (16, 5, 14) {real, imag} */,
  {32'h3d5be344, 32'h3d7c2070} /* (16, 5, 13) {real, imag} */,
  {32'hbaba1ab8, 32'hbd714521} /* (16, 5, 12) {real, imag} */,
  {32'hbd9088aa, 32'h3a7dd180} /* (16, 5, 11) {real, imag} */,
  {32'h3d5484e4, 32'h3d48d8dc} /* (16, 5, 10) {real, imag} */,
  {32'h3cb4f82b, 32'h3c9b306d} /* (16, 5, 9) {real, imag} */,
  {32'h3d9afc66, 32'h3d3254f6} /* (16, 5, 8) {real, imag} */,
  {32'h3e076c07, 32'hbd0ec2b2} /* (16, 5, 7) {real, imag} */,
  {32'hbd00d67e, 32'h3d99e81b} /* (16, 5, 6) {real, imag} */,
  {32'h3e2c694c, 32'h3c9d63ce} /* (16, 5, 5) {real, imag} */,
  {32'h3df29c62, 32'h3dc99de0} /* (16, 5, 4) {real, imag} */,
  {32'hbdb138b0, 32'h3d940ea4} /* (16, 5, 3) {real, imag} */,
  {32'hbdb7241e, 32'h3e8849ac} /* (16, 5, 2) {real, imag} */,
  {32'hbf7f8c66, 32'hbf456861} /* (16, 5, 1) {real, imag} */,
  {32'hbf462805, 32'h00000000} /* (16, 5, 0) {real, imag} */,
  {32'hbf333586, 32'h3f69f7ac} /* (16, 4, 31) {real, imag} */,
  {32'hbec84819, 32'hbebc9c3d} /* (16, 4, 30) {real, imag} */,
  {32'h3c640d8a, 32'h3d30bded} /* (16, 4, 29) {real, imag} */,
  {32'h3e0bfe47, 32'hbe3474fa} /* (16, 4, 28) {real, imag} */,
  {32'h3e33d1c0, 32'hbcc6ca6d} /* (16, 4, 27) {real, imag} */,
  {32'h3d02dbc9, 32'h3dbc70d6} /* (16, 4, 26) {real, imag} */,
  {32'h3e3559ec, 32'hbd7cb058} /* (16, 4, 25) {real, imag} */,
  {32'hbe19dcc6, 32'h3c2b15b8} /* (16, 4, 24) {real, imag} */,
  {32'h3c059bb8, 32'h3cf400c6} /* (16, 4, 23) {real, imag} */,
  {32'hbdfb8e5a, 32'hbdb22f08} /* (16, 4, 22) {real, imag} */,
  {32'h3c136ef4, 32'hbd4ef644} /* (16, 4, 21) {real, imag} */,
  {32'h3d094a65, 32'h3dacc0d6} /* (16, 4, 20) {real, imag} */,
  {32'hbda9ba5b, 32'h3cba4324} /* (16, 4, 19) {real, imag} */,
  {32'hbcca78e4, 32'h3d2b9db4} /* (16, 4, 18) {real, imag} */,
  {32'h3b37295d, 32'hbbfbf62c} /* (16, 4, 17) {real, imag} */,
  {32'hbd929778, 32'h00000000} /* (16, 4, 16) {real, imag} */,
  {32'h3b37295d, 32'h3bfbf62c} /* (16, 4, 15) {real, imag} */,
  {32'hbcca78e4, 32'hbd2b9db4} /* (16, 4, 14) {real, imag} */,
  {32'hbda9ba5b, 32'hbcba4324} /* (16, 4, 13) {real, imag} */,
  {32'h3d094a65, 32'hbdacc0d6} /* (16, 4, 12) {real, imag} */,
  {32'h3c136ef4, 32'h3d4ef644} /* (16, 4, 11) {real, imag} */,
  {32'hbdfb8e5a, 32'h3db22f08} /* (16, 4, 10) {real, imag} */,
  {32'h3c059bb8, 32'hbcf400c6} /* (16, 4, 9) {real, imag} */,
  {32'hbe19dcc6, 32'hbc2b15b8} /* (16, 4, 8) {real, imag} */,
  {32'h3e3559ec, 32'h3d7cb058} /* (16, 4, 7) {real, imag} */,
  {32'h3d02dbc9, 32'hbdbc70d6} /* (16, 4, 6) {real, imag} */,
  {32'h3e33d1c0, 32'h3cc6ca6d} /* (16, 4, 5) {real, imag} */,
  {32'h3e0bfe47, 32'h3e3474fa} /* (16, 4, 4) {real, imag} */,
  {32'h3c640d8a, 32'hbd30bded} /* (16, 4, 3) {real, imag} */,
  {32'hbec84819, 32'h3ebc9c3d} /* (16, 4, 2) {real, imag} */,
  {32'hbf333586, 32'hbf69f7ac} /* (16, 4, 1) {real, imag} */,
  {32'hbf3c66b5, 32'h00000000} /* (16, 4, 0) {real, imag} */,
  {32'hbf1443ea, 32'h3f77b4e0} /* (16, 3, 31) {real, imag} */,
  {32'hbe75c364, 32'hbeabea61} /* (16, 3, 30) {real, imag} */,
  {32'h3d2b77ec, 32'h3df9ea53} /* (16, 3, 29) {real, imag} */,
  {32'h3d502202, 32'hbd6f1d7c} /* (16, 3, 28) {real, imag} */,
  {32'h3dcc67bc, 32'h3e044137} /* (16, 3, 27) {real, imag} */,
  {32'h3caa4c0c, 32'hbc8a7228} /* (16, 3, 26) {real, imag} */,
  {32'h3d33f1d4, 32'h3d8d2366} /* (16, 3, 25) {real, imag} */,
  {32'h3a946210, 32'hbdc47998} /* (16, 3, 24) {real, imag} */,
  {32'h3cc0a94a, 32'hbd1857da} /* (16, 3, 23) {real, imag} */,
  {32'h3caa3508, 32'hbd3b6d42} /* (16, 3, 22) {real, imag} */,
  {32'h3ca07df0, 32'hbdbaebb5} /* (16, 3, 21) {real, imag} */,
  {32'h3b1a99e0, 32'h3daf9026} /* (16, 3, 20) {real, imag} */,
  {32'hbd7aa943, 32'h3c7bcf4a} /* (16, 3, 19) {real, imag} */,
  {32'hbd2304ce, 32'h3d67bfca} /* (16, 3, 18) {real, imag} */,
  {32'h3d17228e, 32'hbd7aeb6c} /* (16, 3, 17) {real, imag} */,
  {32'hbbd5e44e, 32'h00000000} /* (16, 3, 16) {real, imag} */,
  {32'h3d17228e, 32'h3d7aeb6c} /* (16, 3, 15) {real, imag} */,
  {32'hbd2304ce, 32'hbd67bfca} /* (16, 3, 14) {real, imag} */,
  {32'hbd7aa943, 32'hbc7bcf4a} /* (16, 3, 13) {real, imag} */,
  {32'h3b1a99e0, 32'hbdaf9026} /* (16, 3, 12) {real, imag} */,
  {32'h3ca07df0, 32'h3dbaebb5} /* (16, 3, 11) {real, imag} */,
  {32'h3caa3508, 32'h3d3b6d42} /* (16, 3, 10) {real, imag} */,
  {32'h3cc0a94a, 32'h3d1857da} /* (16, 3, 9) {real, imag} */,
  {32'h3a946210, 32'h3dc47998} /* (16, 3, 8) {real, imag} */,
  {32'h3d33f1d4, 32'hbd8d2366} /* (16, 3, 7) {real, imag} */,
  {32'h3caa4c0c, 32'h3c8a7228} /* (16, 3, 6) {real, imag} */,
  {32'h3dcc67bc, 32'hbe044137} /* (16, 3, 5) {real, imag} */,
  {32'h3d502202, 32'h3d6f1d7c} /* (16, 3, 4) {real, imag} */,
  {32'h3d2b77ec, 32'hbdf9ea53} /* (16, 3, 3) {real, imag} */,
  {32'hbe75c364, 32'h3eabea61} /* (16, 3, 2) {real, imag} */,
  {32'hbf1443ea, 32'hbf77b4e0} /* (16, 3, 1) {real, imag} */,
  {32'hbf3aa1b4, 32'h00000000} /* (16, 3, 0) {real, imag} */,
  {32'hbf212180, 32'h3f731b40} /* (16, 2, 31) {real, imag} */,
  {32'hbe1e6b83, 32'hbeeabbf9} /* (16, 2, 30) {real, imag} */,
  {32'h3e1622a4, 32'h3d97cd92} /* (16, 2, 29) {real, imag} */,
  {32'h3cc9a9ed, 32'hbe6909f4} /* (16, 2, 28) {real, imag} */,
  {32'hbc4cd510, 32'h3deb3a54} /* (16, 2, 27) {real, imag} */,
  {32'hbcaaf558, 32'hbd8ed7ea} /* (16, 2, 26) {real, imag} */,
  {32'h3d2749ab, 32'h3d13a2e4} /* (16, 2, 25) {real, imag} */,
  {32'h3ddcd4a4, 32'hbd2ae740} /* (16, 2, 24) {real, imag} */,
  {32'hbdb6cda1, 32'h3c594ca3} /* (16, 2, 23) {real, imag} */,
  {32'h3da2a951, 32'h3ce6f7ad} /* (16, 2, 22) {real, imag} */,
  {32'hbceef948, 32'h3d1eb472} /* (16, 2, 21) {real, imag} */,
  {32'h3c1ecd3a, 32'h3c6a833a} /* (16, 2, 20) {real, imag} */,
  {32'h3ce715fc, 32'h3af35fd0} /* (16, 2, 19) {real, imag} */,
  {32'h3c9649b0, 32'hbd06fb3a} /* (16, 2, 18) {real, imag} */,
  {32'hbd64abe9, 32'h3d085c12} /* (16, 2, 17) {real, imag} */,
  {32'hbbd2f05c, 32'h00000000} /* (16, 2, 16) {real, imag} */,
  {32'hbd64abe9, 32'hbd085c12} /* (16, 2, 15) {real, imag} */,
  {32'h3c9649b0, 32'h3d06fb3a} /* (16, 2, 14) {real, imag} */,
  {32'h3ce715fc, 32'hbaf35fd0} /* (16, 2, 13) {real, imag} */,
  {32'h3c1ecd3a, 32'hbc6a833a} /* (16, 2, 12) {real, imag} */,
  {32'hbceef948, 32'hbd1eb472} /* (16, 2, 11) {real, imag} */,
  {32'h3da2a951, 32'hbce6f7ad} /* (16, 2, 10) {real, imag} */,
  {32'hbdb6cda1, 32'hbc594ca3} /* (16, 2, 9) {real, imag} */,
  {32'h3ddcd4a4, 32'h3d2ae740} /* (16, 2, 8) {real, imag} */,
  {32'h3d2749ab, 32'hbd13a2e4} /* (16, 2, 7) {real, imag} */,
  {32'hbcaaf558, 32'h3d8ed7ea} /* (16, 2, 6) {real, imag} */,
  {32'hbc4cd510, 32'hbdeb3a54} /* (16, 2, 5) {real, imag} */,
  {32'h3cc9a9ed, 32'h3e6909f4} /* (16, 2, 4) {real, imag} */,
  {32'h3e1622a4, 32'hbd97cd92} /* (16, 2, 3) {real, imag} */,
  {32'hbe1e6b83, 32'h3eeabbf9} /* (16, 2, 2) {real, imag} */,
  {32'hbf212180, 32'hbf731b40} /* (16, 2, 1) {real, imag} */,
  {32'hbf51706c, 32'h00000000} /* (16, 2, 0) {real, imag} */,
  {32'hbf323fe7, 32'h3f489173} /* (16, 1, 31) {real, imag} */,
  {32'hbd481eb0, 32'hbee22563} /* (16, 1, 30) {real, imag} */,
  {32'h3dca7525, 32'h3e046cf0} /* (16, 1, 29) {real, imag} */,
  {32'h3c076248, 32'hbe045d46} /* (16, 1, 28) {real, imag} */,
  {32'h3d8f581b, 32'h3d3bb758} /* (16, 1, 27) {real, imag} */,
  {32'h3bd2e0f8, 32'hbd6d0b3b} /* (16, 1, 26) {real, imag} */,
  {32'hbd26c86d, 32'hbd0df0f5} /* (16, 1, 25) {real, imag} */,
  {32'h3bb6a8d4, 32'hbc950d0b} /* (16, 1, 24) {real, imag} */,
  {32'hbe0a9e65, 32'h3d22cb54} /* (16, 1, 23) {real, imag} */,
  {32'hbcc448a2, 32'h3ca6780b} /* (16, 1, 22) {real, imag} */,
  {32'h3d6264ce, 32'hbd25511c} /* (16, 1, 21) {real, imag} */,
  {32'hbc7209a3, 32'hbd902c57} /* (16, 1, 20) {real, imag} */,
  {32'h3d02d6e0, 32'h3c9fcc30} /* (16, 1, 19) {real, imag} */,
  {32'hbcedd279, 32'hbb9abe28} /* (16, 1, 18) {real, imag} */,
  {32'hbdb94654, 32'hbdec1208} /* (16, 1, 17) {real, imag} */,
  {32'hbd88ed0c, 32'h00000000} /* (16, 1, 16) {real, imag} */,
  {32'hbdb94654, 32'h3dec1208} /* (16, 1, 15) {real, imag} */,
  {32'hbcedd279, 32'h3b9abe28} /* (16, 1, 14) {real, imag} */,
  {32'h3d02d6e0, 32'hbc9fcc30} /* (16, 1, 13) {real, imag} */,
  {32'hbc7209a3, 32'h3d902c57} /* (16, 1, 12) {real, imag} */,
  {32'h3d6264ce, 32'h3d25511c} /* (16, 1, 11) {real, imag} */,
  {32'hbcc448a2, 32'hbca6780b} /* (16, 1, 10) {real, imag} */,
  {32'hbe0a9e65, 32'hbd22cb54} /* (16, 1, 9) {real, imag} */,
  {32'h3bb6a8d4, 32'h3c950d0b} /* (16, 1, 8) {real, imag} */,
  {32'hbd26c86d, 32'h3d0df0f5} /* (16, 1, 7) {real, imag} */,
  {32'h3bd2e0f8, 32'h3d6d0b3b} /* (16, 1, 6) {real, imag} */,
  {32'h3d8f581b, 32'hbd3bb758} /* (16, 1, 5) {real, imag} */,
  {32'h3c076248, 32'h3e045d46} /* (16, 1, 4) {real, imag} */,
  {32'h3dca7525, 32'hbe046cf0} /* (16, 1, 3) {real, imag} */,
  {32'hbd481eb0, 32'h3ee22563} /* (16, 1, 2) {real, imag} */,
  {32'hbf323fe7, 32'hbf489173} /* (16, 1, 1) {real, imag} */,
  {32'hbf68cd18, 32'h00000000} /* (16, 1, 0) {real, imag} */,
  {32'hbf2f29f7, 32'h3f1c302c} /* (16, 0, 31) {real, imag} */,
  {32'h3d9ab908, 32'hbeb0f986} /* (16, 0, 30) {real, imag} */,
  {32'h3d3c11c4, 32'h3d6f9ef0} /* (16, 0, 29) {real, imag} */,
  {32'hbd29325a, 32'hbc1d8c88} /* (16, 0, 28) {real, imag} */,
  {32'h3d31a3cc, 32'h3c77aa78} /* (16, 0, 27) {real, imag} */,
  {32'h3d1bbb52, 32'h3c49270c} /* (16, 0, 26) {real, imag} */,
  {32'hbd37701e, 32'h3d62ada1} /* (16, 0, 25) {real, imag} */,
  {32'hbd240ed6, 32'hbd9c7a95} /* (16, 0, 24) {real, imag} */,
  {32'h3b2118e0, 32'hbd0c3e9f} /* (16, 0, 23) {real, imag} */,
  {32'hbcb9ba11, 32'h3c947290} /* (16, 0, 22) {real, imag} */,
  {32'h3cdce3c4, 32'hbd6fb152} /* (16, 0, 21) {real, imag} */,
  {32'hbd1a2289, 32'h3cf1c670} /* (16, 0, 20) {real, imag} */,
  {32'hbd038c2e, 32'h3c6fb30a} /* (16, 0, 19) {real, imag} */,
  {32'h3c1e4ff4, 32'h3bb853e4} /* (16, 0, 18) {real, imag} */,
  {32'h3c2107ee, 32'hbcb18401} /* (16, 0, 17) {real, imag} */,
  {32'hbdbbd458, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h3c2107ee, 32'h3cb18401} /* (16, 0, 15) {real, imag} */,
  {32'h3c1e4ff4, 32'hbbb853e4} /* (16, 0, 14) {real, imag} */,
  {32'hbd038c2e, 32'hbc6fb30a} /* (16, 0, 13) {real, imag} */,
  {32'hbd1a2289, 32'hbcf1c670} /* (16, 0, 12) {real, imag} */,
  {32'h3cdce3c4, 32'h3d6fb152} /* (16, 0, 11) {real, imag} */,
  {32'hbcb9ba11, 32'hbc947290} /* (16, 0, 10) {real, imag} */,
  {32'h3b2118e0, 32'h3d0c3e9f} /* (16, 0, 9) {real, imag} */,
  {32'hbd240ed6, 32'h3d9c7a95} /* (16, 0, 8) {real, imag} */,
  {32'hbd37701e, 32'hbd62ada1} /* (16, 0, 7) {real, imag} */,
  {32'h3d1bbb52, 32'hbc49270c} /* (16, 0, 6) {real, imag} */,
  {32'h3d31a3cc, 32'hbc77aa78} /* (16, 0, 5) {real, imag} */,
  {32'hbd29325a, 32'h3c1d8c88} /* (16, 0, 4) {real, imag} */,
  {32'h3d3c11c4, 32'hbd6f9ef0} /* (16, 0, 3) {real, imag} */,
  {32'h3d9ab908, 32'h3eb0f986} /* (16, 0, 2) {real, imag} */,
  {32'hbf2f29f7, 32'hbf1c302c} /* (16, 0, 1) {real, imag} */,
  {32'hbf71de8c, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h3f52e9ad, 32'hbf02e741} /* (15, 31, 31) {real, imag} */,
  {32'hbe5cdbb9, 32'h3e222470} /* (15, 31, 30) {real, imag} */,
  {32'hbcae8646, 32'h3c0293b4} /* (15, 31, 29) {real, imag} */,
  {32'h3c24effc, 32'hbd4286f6} /* (15, 31, 28) {real, imag} */,
  {32'hbd885437, 32'h3bb9595c} /* (15, 31, 27) {real, imag} */,
  {32'hbc6256fc, 32'h3d5488e3} /* (15, 31, 26) {real, imag} */,
  {32'h3ce4f83d, 32'h3d47d328} /* (15, 31, 25) {real, imag} */,
  {32'hbdef4b80, 32'h3c150808} /* (15, 31, 24) {real, imag} */,
  {32'hbd605cae, 32'h3d13469e} /* (15, 31, 23) {real, imag} */,
  {32'h3cb38bce, 32'hbd1e2b9e} /* (15, 31, 22) {real, imag} */,
  {32'h3c1394b0, 32'h3cf50feb} /* (15, 31, 21) {real, imag} */,
  {32'h3d47db7d, 32'h3ce916d9} /* (15, 31, 20) {real, imag} */,
  {32'hbd4d1283, 32'h3d36af9e} /* (15, 31, 19) {real, imag} */,
  {32'h3cdc577e, 32'hbccf9428} /* (15, 31, 18) {real, imag} */,
  {32'hbd2ec514, 32'hbd03e11e} /* (15, 31, 17) {real, imag} */,
  {32'h3d017e18, 32'h00000000} /* (15, 31, 16) {real, imag} */,
  {32'hbd2ec514, 32'h3d03e11e} /* (15, 31, 15) {real, imag} */,
  {32'h3cdc577e, 32'h3ccf9428} /* (15, 31, 14) {real, imag} */,
  {32'hbd4d1283, 32'hbd36af9e} /* (15, 31, 13) {real, imag} */,
  {32'h3d47db7d, 32'hbce916d9} /* (15, 31, 12) {real, imag} */,
  {32'h3c1394b0, 32'hbcf50feb} /* (15, 31, 11) {real, imag} */,
  {32'h3cb38bce, 32'h3d1e2b9e} /* (15, 31, 10) {real, imag} */,
  {32'hbd605cae, 32'hbd13469e} /* (15, 31, 9) {real, imag} */,
  {32'hbdef4b80, 32'hbc150808} /* (15, 31, 8) {real, imag} */,
  {32'h3ce4f83d, 32'hbd47d328} /* (15, 31, 7) {real, imag} */,
  {32'hbc6256fc, 32'hbd5488e3} /* (15, 31, 6) {real, imag} */,
  {32'hbd885437, 32'hbbb9595c} /* (15, 31, 5) {real, imag} */,
  {32'h3c24effc, 32'h3d4286f6} /* (15, 31, 4) {real, imag} */,
  {32'hbcae8646, 32'hbc0293b4} /* (15, 31, 3) {real, imag} */,
  {32'hbe5cdbb9, 32'hbe222470} /* (15, 31, 2) {real, imag} */,
  {32'h3f52e9ad, 32'h3f02e741} /* (15, 31, 1) {real, imag} */,
  {32'h3f47a1e3, 32'h00000000} /* (15, 31, 0) {real, imag} */,
  {32'h3f52e489, 32'hbed68802} /* (15, 30, 31) {real, imag} */,
  {32'hbeafaaea, 32'h3e320c0d} /* (15, 30, 30) {real, imag} */,
  {32'h3d9356d5, 32'h3dac446a} /* (15, 30, 29) {real, imag} */,
  {32'h3debead8, 32'hbdc3fb12} /* (15, 30, 28) {real, imag} */,
  {32'h3c69c438, 32'h3d7aa1c8} /* (15, 30, 27) {real, imag} */,
  {32'h3db5bed3, 32'hbbf529e4} /* (15, 30, 26) {real, imag} */,
  {32'h3e1ea5da, 32'h3e2e5d56} /* (15, 30, 25) {real, imag} */,
  {32'hbdbc30fc, 32'h3d2683a0} /* (15, 30, 24) {real, imag} */,
  {32'hbb8f8870, 32'h3dbc4e8e} /* (15, 30, 23) {real, imag} */,
  {32'hbd941d70, 32'hbcf1b2f4} /* (15, 30, 22) {real, imag} */,
  {32'hbd346182, 32'hbd63d68e} /* (15, 30, 21) {real, imag} */,
  {32'h3dad7a51, 32'h3d962f4b} /* (15, 30, 20) {real, imag} */,
  {32'h3d037776, 32'h3e11b916} /* (15, 30, 19) {real, imag} */,
  {32'hbc2cd632, 32'h3c3c53d8} /* (15, 30, 18) {real, imag} */,
  {32'h3bc83b76, 32'h3c97f926} /* (15, 30, 17) {real, imag} */,
  {32'hbd6a68dc, 32'h00000000} /* (15, 30, 16) {real, imag} */,
  {32'h3bc83b76, 32'hbc97f926} /* (15, 30, 15) {real, imag} */,
  {32'hbc2cd632, 32'hbc3c53d8} /* (15, 30, 14) {real, imag} */,
  {32'h3d037776, 32'hbe11b916} /* (15, 30, 13) {real, imag} */,
  {32'h3dad7a51, 32'hbd962f4b} /* (15, 30, 12) {real, imag} */,
  {32'hbd346182, 32'h3d63d68e} /* (15, 30, 11) {real, imag} */,
  {32'hbd941d70, 32'h3cf1b2f4} /* (15, 30, 10) {real, imag} */,
  {32'hbb8f8870, 32'hbdbc4e8e} /* (15, 30, 9) {real, imag} */,
  {32'hbdbc30fc, 32'hbd2683a0} /* (15, 30, 8) {real, imag} */,
  {32'h3e1ea5da, 32'hbe2e5d56} /* (15, 30, 7) {real, imag} */,
  {32'h3db5bed3, 32'h3bf529e4} /* (15, 30, 6) {real, imag} */,
  {32'h3c69c438, 32'hbd7aa1c8} /* (15, 30, 5) {real, imag} */,
  {32'h3debead8, 32'h3dc3fb12} /* (15, 30, 4) {real, imag} */,
  {32'h3d9356d5, 32'hbdac446a} /* (15, 30, 3) {real, imag} */,
  {32'hbeafaaea, 32'hbe320c0d} /* (15, 30, 2) {real, imag} */,
  {32'h3f52e489, 32'h3ed68802} /* (15, 30, 1) {real, imag} */,
  {32'h3f6f2e4e, 32'h00000000} /* (15, 30, 0) {real, imag} */,
  {32'h3f219be3, 32'hbec580ec} /* (15, 29, 31) {real, imag} */,
  {32'hbee7a030, 32'h3db40424} /* (15, 29, 30) {real, imag} */,
  {32'h3d81fea0, 32'h3cb511fe} /* (15, 29, 29) {real, imag} */,
  {32'hbd8b0580, 32'hbdaf756a} /* (15, 29, 28) {real, imag} */,
  {32'h3d31fac5, 32'hbb993e60} /* (15, 29, 27) {real, imag} */,
  {32'h3e0a0b8d, 32'h3cac0c91} /* (15, 29, 26) {real, imag} */,
  {32'h3e118b01, 32'hbc85ad22} /* (15, 29, 25) {real, imag} */,
  {32'h3d514f38, 32'h3d8c4416} /* (15, 29, 24) {real, imag} */,
  {32'h3b7e79c0, 32'hbd0a505f} /* (15, 29, 23) {real, imag} */,
  {32'hbdc8a1e1, 32'hbce85d80} /* (15, 29, 22) {real, imag} */,
  {32'hbd8b4c81, 32'h3d85e3a8} /* (15, 29, 21) {real, imag} */,
  {32'hbcbdf1d8, 32'h3c7d1fe4} /* (15, 29, 20) {real, imag} */,
  {32'h3db431ca, 32'hbbd4ade8} /* (15, 29, 19) {real, imag} */,
  {32'h3d18a650, 32'h3d1d6c95} /* (15, 29, 18) {real, imag} */,
  {32'h3d7f7364, 32'h3d58fe91} /* (15, 29, 17) {real, imag} */,
  {32'hbd131adf, 32'h00000000} /* (15, 29, 16) {real, imag} */,
  {32'h3d7f7364, 32'hbd58fe91} /* (15, 29, 15) {real, imag} */,
  {32'h3d18a650, 32'hbd1d6c95} /* (15, 29, 14) {real, imag} */,
  {32'h3db431ca, 32'h3bd4ade8} /* (15, 29, 13) {real, imag} */,
  {32'hbcbdf1d8, 32'hbc7d1fe4} /* (15, 29, 12) {real, imag} */,
  {32'hbd8b4c81, 32'hbd85e3a8} /* (15, 29, 11) {real, imag} */,
  {32'hbdc8a1e1, 32'h3ce85d80} /* (15, 29, 10) {real, imag} */,
  {32'h3b7e79c0, 32'h3d0a505f} /* (15, 29, 9) {real, imag} */,
  {32'h3d514f38, 32'hbd8c4416} /* (15, 29, 8) {real, imag} */,
  {32'h3e118b01, 32'h3c85ad22} /* (15, 29, 7) {real, imag} */,
  {32'h3e0a0b8d, 32'hbcac0c91} /* (15, 29, 6) {real, imag} */,
  {32'h3d31fac5, 32'h3b993e60} /* (15, 29, 5) {real, imag} */,
  {32'hbd8b0580, 32'h3daf756a} /* (15, 29, 4) {real, imag} */,
  {32'h3d81fea0, 32'hbcb511fe} /* (15, 29, 3) {real, imag} */,
  {32'hbee7a030, 32'hbdb40424} /* (15, 29, 2) {real, imag} */,
  {32'h3f219be3, 32'h3ec580ec} /* (15, 29, 1) {real, imag} */,
  {32'h3f8139eb, 32'h00000000} /* (15, 29, 0) {real, imag} */,
  {32'h3efb7a4e, 32'hbeb3ddfa} /* (15, 28, 31) {real, imag} */,
  {32'hbef731fd, 32'hbda57706} /* (15, 28, 30) {real, imag} */,
  {32'h3d6cd4b7, 32'h39087400} /* (15, 28, 29) {real, imag} */,
  {32'h3cabf5ee, 32'hbe0f4b4e} /* (15, 28, 28) {real, imag} */,
  {32'hbdcb0493, 32'h3d2ec338} /* (15, 28, 27) {real, imag} */,
  {32'h3dd27ad8, 32'h3d0ac7ca} /* (15, 28, 26) {real, imag} */,
  {32'h3dfcd1cf, 32'hbdc9dd50} /* (15, 28, 25) {real, imag} */,
  {32'hbcffbf3e, 32'hbc53d634} /* (15, 28, 24) {real, imag} */,
  {32'h3d8f6232, 32'h3d66a617} /* (15, 28, 23) {real, imag} */,
  {32'h3c39e718, 32'hbb0ead36} /* (15, 28, 22) {real, imag} */,
  {32'hbb456d2c, 32'hbc08a324} /* (15, 28, 21) {real, imag} */,
  {32'h3d1bba95, 32'hbc2a68f8} /* (15, 28, 20) {real, imag} */,
  {32'h3cb1c2ec, 32'h3de51528} /* (15, 28, 19) {real, imag} */,
  {32'hbd6a0bf8, 32'h3d3321cc} /* (15, 28, 18) {real, imag} */,
  {32'hbbac8588, 32'hbc911792} /* (15, 28, 17) {real, imag} */,
  {32'h3d06e4a5, 32'h00000000} /* (15, 28, 16) {real, imag} */,
  {32'hbbac8588, 32'h3c911792} /* (15, 28, 15) {real, imag} */,
  {32'hbd6a0bf8, 32'hbd3321cc} /* (15, 28, 14) {real, imag} */,
  {32'h3cb1c2ec, 32'hbde51528} /* (15, 28, 13) {real, imag} */,
  {32'h3d1bba95, 32'h3c2a68f8} /* (15, 28, 12) {real, imag} */,
  {32'hbb456d2c, 32'h3c08a324} /* (15, 28, 11) {real, imag} */,
  {32'h3c39e718, 32'h3b0ead36} /* (15, 28, 10) {real, imag} */,
  {32'h3d8f6232, 32'hbd66a617} /* (15, 28, 9) {real, imag} */,
  {32'hbcffbf3e, 32'h3c53d634} /* (15, 28, 8) {real, imag} */,
  {32'h3dfcd1cf, 32'h3dc9dd50} /* (15, 28, 7) {real, imag} */,
  {32'h3dd27ad8, 32'hbd0ac7ca} /* (15, 28, 6) {real, imag} */,
  {32'hbdcb0493, 32'hbd2ec338} /* (15, 28, 5) {real, imag} */,
  {32'h3cabf5ee, 32'h3e0f4b4e} /* (15, 28, 4) {real, imag} */,
  {32'h3d6cd4b7, 32'hb9087400} /* (15, 28, 3) {real, imag} */,
  {32'hbef731fd, 32'h3da57706} /* (15, 28, 2) {real, imag} */,
  {32'h3efb7a4e, 32'h3eb3ddfa} /* (15, 28, 1) {real, imag} */,
  {32'h3f8c8bf4, 32'h00000000} /* (15, 28, 0) {real, imag} */,
  {32'h3f2b0ecd, 32'hbe88243c} /* (15, 27, 31) {real, imag} */,
  {32'hbf13b8b3, 32'hbc550fa8} /* (15, 27, 30) {real, imag} */,
  {32'h3dd17999, 32'hbb0a74e0} /* (15, 27, 29) {real, imag} */,
  {32'hbd0cebda, 32'hbdf5ea5f} /* (15, 27, 28) {real, imag} */,
  {32'hba0ebc00, 32'hbcb8e924} /* (15, 27, 27) {real, imag} */,
  {32'h3da6033d, 32'hbdb42f29} /* (15, 27, 26) {real, imag} */,
  {32'hbc73e900, 32'hbd2600ff} /* (15, 27, 25) {real, imag} */,
  {32'hbe105b01, 32'h3e500dbc} /* (15, 27, 24) {real, imag} */,
  {32'h3da1081c, 32'hbcc10168} /* (15, 27, 23) {real, imag} */,
  {32'hbd983985, 32'hbd74b499} /* (15, 27, 22) {real, imag} */,
  {32'hbc8c6746, 32'h3c27a234} /* (15, 27, 21) {real, imag} */,
  {32'h3d3a0b3f, 32'hbce82b58} /* (15, 27, 20) {real, imag} */,
  {32'hbd229878, 32'h3c8ce1f4} /* (15, 27, 19) {real, imag} */,
  {32'h3da6cf78, 32'h3dd9914d} /* (15, 27, 18) {real, imag} */,
  {32'hbb32de70, 32'hbd4c73a8} /* (15, 27, 17) {real, imag} */,
  {32'hbc0cd290, 32'h00000000} /* (15, 27, 16) {real, imag} */,
  {32'hbb32de70, 32'h3d4c73a8} /* (15, 27, 15) {real, imag} */,
  {32'h3da6cf78, 32'hbdd9914d} /* (15, 27, 14) {real, imag} */,
  {32'hbd229878, 32'hbc8ce1f4} /* (15, 27, 13) {real, imag} */,
  {32'h3d3a0b3f, 32'h3ce82b58} /* (15, 27, 12) {real, imag} */,
  {32'hbc8c6746, 32'hbc27a234} /* (15, 27, 11) {real, imag} */,
  {32'hbd983985, 32'h3d74b499} /* (15, 27, 10) {real, imag} */,
  {32'h3da1081c, 32'h3cc10168} /* (15, 27, 9) {real, imag} */,
  {32'hbe105b01, 32'hbe500dbc} /* (15, 27, 8) {real, imag} */,
  {32'hbc73e900, 32'h3d2600ff} /* (15, 27, 7) {real, imag} */,
  {32'h3da6033d, 32'h3db42f29} /* (15, 27, 6) {real, imag} */,
  {32'hba0ebc00, 32'h3cb8e924} /* (15, 27, 5) {real, imag} */,
  {32'hbd0cebda, 32'h3df5ea5f} /* (15, 27, 4) {real, imag} */,
  {32'h3dd17999, 32'h3b0a74e0} /* (15, 27, 3) {real, imag} */,
  {32'hbf13b8b3, 32'h3c550fa8} /* (15, 27, 2) {real, imag} */,
  {32'h3f2b0ecd, 32'h3e88243c} /* (15, 27, 1) {real, imag} */,
  {32'h3f6ee5d8, 32'h00000000} /* (15, 27, 0) {real, imag} */,
  {32'h3f5d5fe5, 32'hbe38feec} /* (15, 26, 31) {real, imag} */,
  {32'hbf01f138, 32'h3cf121fc} /* (15, 26, 30) {real, imag} */,
  {32'h3d1e87b8, 32'h3b198370} /* (15, 26, 29) {real, imag} */,
  {32'hbdf11124, 32'hbde6279a} /* (15, 26, 28) {real, imag} */,
  {32'hbd9385e7, 32'h3e3592d1} /* (15, 26, 27) {real, imag} */,
  {32'hbbbe2c58, 32'hbd8bb38c} /* (15, 26, 26) {real, imag} */,
  {32'hbce06000, 32'h3ce856f5} /* (15, 26, 25) {real, imag} */,
  {32'hbe1aeb51, 32'hbccbab42} /* (15, 26, 24) {real, imag} */,
  {32'h3daf823f, 32'hbca8415a} /* (15, 26, 23) {real, imag} */,
  {32'h3d9b233e, 32'hbde601e8} /* (15, 26, 22) {real, imag} */,
  {32'h3bd0cccc, 32'h3dd00388} /* (15, 26, 21) {real, imag} */,
  {32'hbbe8ccd4, 32'hbd887d42} /* (15, 26, 20) {real, imag} */,
  {32'h3d095504, 32'h3c92903a} /* (15, 26, 19) {real, imag} */,
  {32'h3db9dbc0, 32'h3d816d5f} /* (15, 26, 18) {real, imag} */,
  {32'h3d0039c6, 32'hbcc97be6} /* (15, 26, 17) {real, imag} */,
  {32'hbcd45a26, 32'h00000000} /* (15, 26, 16) {real, imag} */,
  {32'h3d0039c6, 32'h3cc97be6} /* (15, 26, 15) {real, imag} */,
  {32'h3db9dbc0, 32'hbd816d5f} /* (15, 26, 14) {real, imag} */,
  {32'h3d095504, 32'hbc92903a} /* (15, 26, 13) {real, imag} */,
  {32'hbbe8ccd4, 32'h3d887d42} /* (15, 26, 12) {real, imag} */,
  {32'h3bd0cccc, 32'hbdd00388} /* (15, 26, 11) {real, imag} */,
  {32'h3d9b233e, 32'h3de601e8} /* (15, 26, 10) {real, imag} */,
  {32'h3daf823f, 32'h3ca8415a} /* (15, 26, 9) {real, imag} */,
  {32'hbe1aeb51, 32'h3ccbab42} /* (15, 26, 8) {real, imag} */,
  {32'hbce06000, 32'hbce856f5} /* (15, 26, 7) {real, imag} */,
  {32'hbbbe2c58, 32'h3d8bb38c} /* (15, 26, 6) {real, imag} */,
  {32'hbd9385e7, 32'hbe3592d1} /* (15, 26, 5) {real, imag} */,
  {32'hbdf11124, 32'h3de6279a} /* (15, 26, 4) {real, imag} */,
  {32'h3d1e87b8, 32'hbb198370} /* (15, 26, 3) {real, imag} */,
  {32'hbf01f138, 32'hbcf121fc} /* (15, 26, 2) {real, imag} */,
  {32'h3f5d5fe5, 32'h3e38feec} /* (15, 26, 1) {real, imag} */,
  {32'h3f3204a4, 32'h00000000} /* (15, 26, 0) {real, imag} */,
  {32'h3f673852, 32'hbe1b54ae} /* (15, 25, 31) {real, imag} */,
  {32'hbf01c6d3, 32'h3dd34958} /* (15, 25, 30) {real, imag} */,
  {32'h3da23f34, 32'hbdae5d63} /* (15, 25, 29) {real, imag} */,
  {32'h3bc8b8d8, 32'hbcf722f4} /* (15, 25, 28) {real, imag} */,
  {32'hbd72da65, 32'h3e0a163e} /* (15, 25, 27) {real, imag} */,
  {32'h3da90978, 32'h3cc43edb} /* (15, 25, 26) {real, imag} */,
  {32'h3d1e3894, 32'h3d6e4250} /* (15, 25, 25) {real, imag} */,
  {32'hbbbf1c14, 32'h3c244ba4} /* (15, 25, 24) {real, imag} */,
  {32'h3da5253a, 32'h3d688a4e} /* (15, 25, 23) {real, imag} */,
  {32'hbd3eac7c, 32'h3d940fe2} /* (15, 25, 22) {real, imag} */,
  {32'h3cc1a147, 32'hbd20e0f0} /* (15, 25, 21) {real, imag} */,
  {32'hbc046faa, 32'h3d49e11b} /* (15, 25, 20) {real, imag} */,
  {32'hbd2b9808, 32'h3c192d48} /* (15, 25, 19) {real, imag} */,
  {32'hbd62412a, 32'h3d805ecd} /* (15, 25, 18) {real, imag} */,
  {32'hbc4c269f, 32'hbca2dc87} /* (15, 25, 17) {real, imag} */,
  {32'hba4a1d20, 32'h00000000} /* (15, 25, 16) {real, imag} */,
  {32'hbc4c269f, 32'h3ca2dc87} /* (15, 25, 15) {real, imag} */,
  {32'hbd62412a, 32'hbd805ecd} /* (15, 25, 14) {real, imag} */,
  {32'hbd2b9808, 32'hbc192d48} /* (15, 25, 13) {real, imag} */,
  {32'hbc046faa, 32'hbd49e11b} /* (15, 25, 12) {real, imag} */,
  {32'h3cc1a147, 32'h3d20e0f0} /* (15, 25, 11) {real, imag} */,
  {32'hbd3eac7c, 32'hbd940fe2} /* (15, 25, 10) {real, imag} */,
  {32'h3da5253a, 32'hbd688a4e} /* (15, 25, 9) {real, imag} */,
  {32'hbbbf1c14, 32'hbc244ba4} /* (15, 25, 8) {real, imag} */,
  {32'h3d1e3894, 32'hbd6e4250} /* (15, 25, 7) {real, imag} */,
  {32'h3da90978, 32'hbcc43edb} /* (15, 25, 6) {real, imag} */,
  {32'hbd72da65, 32'hbe0a163e} /* (15, 25, 5) {real, imag} */,
  {32'h3bc8b8d8, 32'h3cf722f4} /* (15, 25, 4) {real, imag} */,
  {32'h3da23f34, 32'h3dae5d63} /* (15, 25, 3) {real, imag} */,
  {32'hbf01c6d3, 32'hbdd34958} /* (15, 25, 2) {real, imag} */,
  {32'h3f673852, 32'h3e1b54ae} /* (15, 25, 1) {real, imag} */,
  {32'h3f33a4de, 32'h00000000} /* (15, 25, 0) {real, imag} */,
  {32'h3f592fe9, 32'hbe43af4f} /* (15, 24, 31) {real, imag} */,
  {32'hbedce43d, 32'h3e103cb2} /* (15, 24, 30) {real, imag} */,
  {32'h3d8c1ced, 32'hbe1e20ce} /* (15, 24, 29) {real, imag} */,
  {32'h3b73dfa8, 32'hbe135650} /* (15, 24, 28) {real, imag} */,
  {32'hbdb9b116, 32'h3cda2f94} /* (15, 24, 27) {real, imag} */,
  {32'hbd9ed456, 32'h3e118c05} /* (15, 24, 26) {real, imag} */,
  {32'h3d9103cc, 32'hbcfd96bc} /* (15, 24, 25) {real, imag} */,
  {32'h3d15d722, 32'h3d4de0dd} /* (15, 24, 24) {real, imag} */,
  {32'hbd8571fa, 32'hbc18eb8c} /* (15, 24, 23) {real, imag} */,
  {32'hbbe34d78, 32'hbd61776e} /* (15, 24, 22) {real, imag} */,
  {32'h3d30716b, 32'h3d77e8da} /* (15, 24, 21) {real, imag} */,
  {32'hbd4bf9d9, 32'hbc5e2040} /* (15, 24, 20) {real, imag} */,
  {32'h3d42669e, 32'h3ce7eecc} /* (15, 24, 19) {real, imag} */,
  {32'hbcb8fd05, 32'h3d3be2d0} /* (15, 24, 18) {real, imag} */,
  {32'hbc82ef72, 32'hbcdd99ad} /* (15, 24, 17) {real, imag} */,
  {32'h3d61ad94, 32'h00000000} /* (15, 24, 16) {real, imag} */,
  {32'hbc82ef72, 32'h3cdd99ad} /* (15, 24, 15) {real, imag} */,
  {32'hbcb8fd05, 32'hbd3be2d0} /* (15, 24, 14) {real, imag} */,
  {32'h3d42669e, 32'hbce7eecc} /* (15, 24, 13) {real, imag} */,
  {32'hbd4bf9d9, 32'h3c5e2040} /* (15, 24, 12) {real, imag} */,
  {32'h3d30716b, 32'hbd77e8da} /* (15, 24, 11) {real, imag} */,
  {32'hbbe34d78, 32'h3d61776e} /* (15, 24, 10) {real, imag} */,
  {32'hbd8571fa, 32'h3c18eb8c} /* (15, 24, 9) {real, imag} */,
  {32'h3d15d722, 32'hbd4de0dd} /* (15, 24, 8) {real, imag} */,
  {32'h3d9103cc, 32'h3cfd96bc} /* (15, 24, 7) {real, imag} */,
  {32'hbd9ed456, 32'hbe118c05} /* (15, 24, 6) {real, imag} */,
  {32'hbdb9b116, 32'hbcda2f94} /* (15, 24, 5) {real, imag} */,
  {32'h3b73dfa8, 32'h3e135650} /* (15, 24, 4) {real, imag} */,
  {32'h3d8c1ced, 32'h3e1e20ce} /* (15, 24, 3) {real, imag} */,
  {32'hbedce43d, 32'hbe103cb2} /* (15, 24, 2) {real, imag} */,
  {32'h3f592fe9, 32'h3e43af4f} /* (15, 24, 1) {real, imag} */,
  {32'h3f10f00c, 32'h00000000} /* (15, 24, 0) {real, imag} */,
  {32'h3f431bac, 32'hbdcdeec1} /* (15, 23, 31) {real, imag} */,
  {32'hbecdfb6a, 32'h3de7a984} /* (15, 23, 30) {real, imag} */,
  {32'hbd7b7788, 32'hbe7ff318} /* (15, 23, 29) {real, imag} */,
  {32'hbda625d8, 32'hbe7f923a} /* (15, 23, 28) {real, imag} */,
  {32'hbe075132, 32'hbc04575e} /* (15, 23, 27) {real, imag} */,
  {32'hbde5f91c, 32'hbd95428b} /* (15, 23, 26) {real, imag} */,
  {32'h3d92ac85, 32'h3d1cf9b6} /* (15, 23, 25) {real, imag} */,
  {32'hbd128cc2, 32'h3dc4c0f0} /* (15, 23, 24) {real, imag} */,
  {32'h3d4fbac5, 32'h3b8d384d} /* (15, 23, 23) {real, imag} */,
  {32'hbcad8ec8, 32'h3d388505} /* (15, 23, 22) {real, imag} */,
  {32'h3b8abc28, 32'h3caf2405} /* (15, 23, 21) {real, imag} */,
  {32'h3d002238, 32'hbdad5abd} /* (15, 23, 20) {real, imag} */,
  {32'h3a9649a0, 32'hbd88e62f} /* (15, 23, 19) {real, imag} */,
  {32'h3d806b38, 32'h3cc7db25} /* (15, 23, 18) {real, imag} */,
  {32'hbcbf50ea, 32'h3dba8019} /* (15, 23, 17) {real, imag} */,
  {32'hbe027801, 32'h00000000} /* (15, 23, 16) {real, imag} */,
  {32'hbcbf50ea, 32'hbdba8019} /* (15, 23, 15) {real, imag} */,
  {32'h3d806b38, 32'hbcc7db25} /* (15, 23, 14) {real, imag} */,
  {32'h3a9649a0, 32'h3d88e62f} /* (15, 23, 13) {real, imag} */,
  {32'h3d002238, 32'h3dad5abd} /* (15, 23, 12) {real, imag} */,
  {32'h3b8abc28, 32'hbcaf2405} /* (15, 23, 11) {real, imag} */,
  {32'hbcad8ec8, 32'hbd388505} /* (15, 23, 10) {real, imag} */,
  {32'h3d4fbac5, 32'hbb8d384d} /* (15, 23, 9) {real, imag} */,
  {32'hbd128cc2, 32'hbdc4c0f0} /* (15, 23, 8) {real, imag} */,
  {32'h3d92ac85, 32'hbd1cf9b6} /* (15, 23, 7) {real, imag} */,
  {32'hbde5f91c, 32'h3d95428b} /* (15, 23, 6) {real, imag} */,
  {32'hbe075132, 32'h3c04575e} /* (15, 23, 5) {real, imag} */,
  {32'hbda625d8, 32'h3e7f923a} /* (15, 23, 4) {real, imag} */,
  {32'hbd7b7788, 32'h3e7ff318} /* (15, 23, 3) {real, imag} */,
  {32'hbecdfb6a, 32'hbde7a984} /* (15, 23, 2) {real, imag} */,
  {32'h3f431bac, 32'h3dcdeec1} /* (15, 23, 1) {real, imag} */,
  {32'h3eb0aa4d, 32'h00000000} /* (15, 23, 0) {real, imag} */,
  {32'h3f28c32a, 32'hbd925339} /* (15, 22, 31) {real, imag} */,
  {32'hbe81815a, 32'h3dcec0c2} /* (15, 22, 30) {real, imag} */,
  {32'h3d4029de, 32'hbe46ccb4} /* (15, 22, 29) {real, imag} */,
  {32'hbd5925eb, 32'hbe3db051} /* (15, 22, 28) {real, imag} */,
  {32'hbd95f181, 32'h3c928705} /* (15, 22, 27) {real, imag} */,
  {32'hbe26517e, 32'hbd96ea08} /* (15, 22, 26) {real, imag} */,
  {32'h3df16736, 32'h3c7e5e08} /* (15, 22, 25) {real, imag} */,
  {32'hbbef4e40, 32'h3d0c27ba} /* (15, 22, 24) {real, imag} */,
  {32'hbc2ca4ee, 32'h3a0e7570} /* (15, 22, 23) {real, imag} */,
  {32'hbdddb5fe, 32'hbc2fed48} /* (15, 22, 22) {real, imag} */,
  {32'hbd0bb33f, 32'hbd051386} /* (15, 22, 21) {real, imag} */,
  {32'hbd45d0de, 32'hbd4a28ba} /* (15, 22, 20) {real, imag} */,
  {32'h3ba02c20, 32'h3cfd3214} /* (15, 22, 19) {real, imag} */,
  {32'hbd9d165b, 32'h3b2be7b4} /* (15, 22, 18) {real, imag} */,
  {32'hba645e80, 32'hbd3672fb} /* (15, 22, 17) {real, imag} */,
  {32'h3d5aa288, 32'h00000000} /* (15, 22, 16) {real, imag} */,
  {32'hba645e80, 32'h3d3672fb} /* (15, 22, 15) {real, imag} */,
  {32'hbd9d165b, 32'hbb2be7b4} /* (15, 22, 14) {real, imag} */,
  {32'h3ba02c20, 32'hbcfd3214} /* (15, 22, 13) {real, imag} */,
  {32'hbd45d0de, 32'h3d4a28ba} /* (15, 22, 12) {real, imag} */,
  {32'hbd0bb33f, 32'h3d051386} /* (15, 22, 11) {real, imag} */,
  {32'hbdddb5fe, 32'h3c2fed48} /* (15, 22, 10) {real, imag} */,
  {32'hbc2ca4ee, 32'hba0e7570} /* (15, 22, 9) {real, imag} */,
  {32'hbbef4e40, 32'hbd0c27ba} /* (15, 22, 8) {real, imag} */,
  {32'h3df16736, 32'hbc7e5e08} /* (15, 22, 7) {real, imag} */,
  {32'hbe26517e, 32'h3d96ea08} /* (15, 22, 6) {real, imag} */,
  {32'hbd95f181, 32'hbc928705} /* (15, 22, 5) {real, imag} */,
  {32'hbd5925eb, 32'h3e3db051} /* (15, 22, 4) {real, imag} */,
  {32'h3d4029de, 32'h3e46ccb4} /* (15, 22, 3) {real, imag} */,
  {32'hbe81815a, 32'hbdcec0c2} /* (15, 22, 2) {real, imag} */,
  {32'h3f28c32a, 32'h3d925339} /* (15, 22, 1) {real, imag} */,
  {32'h3e72ccf4, 32'h00000000} /* (15, 22, 0) {real, imag} */,
  {32'h3e41400a, 32'hbd83f426} /* (15, 21, 31) {real, imag} */,
  {32'hbda0ee8c, 32'h3e01c91c} /* (15, 21, 30) {real, imag} */,
  {32'h3d8338b0, 32'hbde8fede} /* (15, 21, 29) {real, imag} */,
  {32'h3c98d1a0, 32'hbe27a81b} /* (15, 21, 28) {real, imag} */,
  {32'hbda0159b, 32'hbc139c40} /* (15, 21, 27) {real, imag} */,
  {32'h3d1a29d8, 32'hbd0532a4} /* (15, 21, 26) {real, imag} */,
  {32'h3d74e7e8, 32'h3c46572c} /* (15, 21, 25) {real, imag} */,
  {32'hbd4c2998, 32'hbd1fd2e4} /* (15, 21, 24) {real, imag} */,
  {32'h3c8de962, 32'hbcc4289e} /* (15, 21, 23) {real, imag} */,
  {32'h3c4b04e8, 32'h3c20c264} /* (15, 21, 22) {real, imag} */,
  {32'h3d0306c3, 32'h3e08d8ff} /* (15, 21, 21) {real, imag} */,
  {32'hbc4e3c18, 32'h3d991cd5} /* (15, 21, 20) {real, imag} */,
  {32'h3ad190c0, 32'hbc5579c4} /* (15, 21, 19) {real, imag} */,
  {32'hbbe1fdd2, 32'h3c57d9b4} /* (15, 21, 18) {real, imag} */,
  {32'h3dad825e, 32'h3cd3738a} /* (15, 21, 17) {real, imag} */,
  {32'hbc4b8c78, 32'h00000000} /* (15, 21, 16) {real, imag} */,
  {32'h3dad825e, 32'hbcd3738a} /* (15, 21, 15) {real, imag} */,
  {32'hbbe1fdd2, 32'hbc57d9b4} /* (15, 21, 14) {real, imag} */,
  {32'h3ad190c0, 32'h3c5579c4} /* (15, 21, 13) {real, imag} */,
  {32'hbc4e3c18, 32'hbd991cd5} /* (15, 21, 12) {real, imag} */,
  {32'h3d0306c3, 32'hbe08d8ff} /* (15, 21, 11) {real, imag} */,
  {32'h3c4b04e8, 32'hbc20c264} /* (15, 21, 10) {real, imag} */,
  {32'h3c8de962, 32'h3cc4289e} /* (15, 21, 9) {real, imag} */,
  {32'hbd4c2998, 32'h3d1fd2e4} /* (15, 21, 8) {real, imag} */,
  {32'h3d74e7e8, 32'hbc46572c} /* (15, 21, 7) {real, imag} */,
  {32'h3d1a29d8, 32'h3d0532a4} /* (15, 21, 6) {real, imag} */,
  {32'hbda0159b, 32'h3c139c40} /* (15, 21, 5) {real, imag} */,
  {32'h3c98d1a0, 32'h3e27a81b} /* (15, 21, 4) {real, imag} */,
  {32'h3d8338b0, 32'h3de8fede} /* (15, 21, 3) {real, imag} */,
  {32'hbda0ee8c, 32'hbe01c91c} /* (15, 21, 2) {real, imag} */,
  {32'h3e41400a, 32'h3d83f426} /* (15, 21, 1) {real, imag} */,
  {32'hbc190d70, 32'h00000000} /* (15, 21, 0) {real, imag} */,
  {32'hbefe2f3a, 32'h3e3d83b2} /* (15, 20, 31) {real, imag} */,
  {32'h3e86ae06, 32'hbb705eb0} /* (15, 20, 30) {real, imag} */,
  {32'h3e077f14, 32'hbc831678} /* (15, 20, 29) {real, imag} */,
  {32'h3b7a8b00, 32'hbd7edd4a} /* (15, 20, 28) {real, imag} */,
  {32'h3ccf1f03, 32'h3a512f80} /* (15, 20, 27) {real, imag} */,
  {32'hbc78af2c, 32'hbd9325ca} /* (15, 20, 26) {real, imag} */,
  {32'hbe0c6aa2, 32'hbd2d2df5} /* (15, 20, 25) {real, imag} */,
  {32'h3db05210, 32'hbe05a20f} /* (15, 20, 24) {real, imag} */,
  {32'h3cdb45c2, 32'h3d0c7d26} /* (15, 20, 23) {real, imag} */,
  {32'h3c802615, 32'hbc4626c4} /* (15, 20, 22) {real, imag} */,
  {32'hbd108b43, 32'hbcd13ca0} /* (15, 20, 21) {real, imag} */,
  {32'hbd5a6054, 32'h3d072aba} /* (15, 20, 20) {real, imag} */,
  {32'hbd1b196a, 32'hbd50e24d} /* (15, 20, 19) {real, imag} */,
  {32'hbc2fc2b2, 32'hbcd29695} /* (15, 20, 18) {real, imag} */,
  {32'h3c2c5c15, 32'hbaf10470} /* (15, 20, 17) {real, imag} */,
  {32'h3cd41e39, 32'h00000000} /* (15, 20, 16) {real, imag} */,
  {32'h3c2c5c15, 32'h3af10470} /* (15, 20, 15) {real, imag} */,
  {32'hbc2fc2b2, 32'h3cd29695} /* (15, 20, 14) {real, imag} */,
  {32'hbd1b196a, 32'h3d50e24d} /* (15, 20, 13) {real, imag} */,
  {32'hbd5a6054, 32'hbd072aba} /* (15, 20, 12) {real, imag} */,
  {32'hbd108b43, 32'h3cd13ca0} /* (15, 20, 11) {real, imag} */,
  {32'h3c802615, 32'h3c4626c4} /* (15, 20, 10) {real, imag} */,
  {32'h3cdb45c2, 32'hbd0c7d26} /* (15, 20, 9) {real, imag} */,
  {32'h3db05210, 32'h3e05a20f} /* (15, 20, 8) {real, imag} */,
  {32'hbe0c6aa2, 32'h3d2d2df5} /* (15, 20, 7) {real, imag} */,
  {32'hbc78af2c, 32'h3d9325ca} /* (15, 20, 6) {real, imag} */,
  {32'h3ccf1f03, 32'hba512f80} /* (15, 20, 5) {real, imag} */,
  {32'h3b7a8b00, 32'h3d7edd4a} /* (15, 20, 4) {real, imag} */,
  {32'h3e077f14, 32'h3c831678} /* (15, 20, 3) {real, imag} */,
  {32'h3e86ae06, 32'h3b705eb0} /* (15, 20, 2) {real, imag} */,
  {32'hbefe2f3a, 32'hbe3d83b2} /* (15, 20, 1) {real, imag} */,
  {32'hbeaf4937, 32'h00000000} /* (15, 20, 0) {real, imag} */,
  {32'hbf46a411, 32'h3e56fe53} /* (15, 19, 31) {real, imag} */,
  {32'h3ec305e4, 32'hbd24f326} /* (15, 19, 30) {real, imag} */,
  {32'h3e23f84c, 32'h3d132e34} /* (15, 19, 29) {real, imag} */,
  {32'h3d0aa5ca, 32'hbdee9eb8} /* (15, 19, 28) {real, imag} */,
  {32'h3d9bbe62, 32'h3d077249} /* (15, 19, 27) {real, imag} */,
  {32'hbdb251c2, 32'hbc8299ce} /* (15, 19, 26) {real, imag} */,
  {32'hbdb49dac, 32'h3cdacf6a} /* (15, 19, 25) {real, imag} */,
  {32'h3d107490, 32'hbd1441e5} /* (15, 19, 24) {real, imag} */,
  {32'hbde7a634, 32'h3c01d840} /* (15, 19, 23) {real, imag} */,
  {32'h3bf10770, 32'hbd8cba73} /* (15, 19, 22) {real, imag} */,
  {32'h3c236f72, 32'hbdac8390} /* (15, 19, 21) {real, imag} */,
  {32'h3d793aa1, 32'hbd9311da} /* (15, 19, 20) {real, imag} */,
  {32'hbcaab737, 32'h3ce30b34} /* (15, 19, 19) {real, imag} */,
  {32'hbc8a9b26, 32'h3db534fc} /* (15, 19, 18) {real, imag} */,
  {32'h3c47f7b4, 32'h3d871996} /* (15, 19, 17) {real, imag} */,
  {32'hbb7bc984, 32'h00000000} /* (15, 19, 16) {real, imag} */,
  {32'h3c47f7b4, 32'hbd871996} /* (15, 19, 15) {real, imag} */,
  {32'hbc8a9b26, 32'hbdb534fc} /* (15, 19, 14) {real, imag} */,
  {32'hbcaab737, 32'hbce30b34} /* (15, 19, 13) {real, imag} */,
  {32'h3d793aa1, 32'h3d9311da} /* (15, 19, 12) {real, imag} */,
  {32'h3c236f72, 32'h3dac8390} /* (15, 19, 11) {real, imag} */,
  {32'h3bf10770, 32'h3d8cba73} /* (15, 19, 10) {real, imag} */,
  {32'hbde7a634, 32'hbc01d840} /* (15, 19, 9) {real, imag} */,
  {32'h3d107490, 32'h3d1441e5} /* (15, 19, 8) {real, imag} */,
  {32'hbdb49dac, 32'hbcdacf6a} /* (15, 19, 7) {real, imag} */,
  {32'hbdb251c2, 32'h3c8299ce} /* (15, 19, 6) {real, imag} */,
  {32'h3d9bbe62, 32'hbd077249} /* (15, 19, 5) {real, imag} */,
  {32'h3d0aa5ca, 32'h3dee9eb8} /* (15, 19, 4) {real, imag} */,
  {32'h3e23f84c, 32'hbd132e34} /* (15, 19, 3) {real, imag} */,
  {32'h3ec305e4, 32'h3d24f326} /* (15, 19, 2) {real, imag} */,
  {32'hbf46a411, 32'hbe56fe53} /* (15, 19, 1) {real, imag} */,
  {32'hbec64828, 32'h00000000} /* (15, 19, 0) {real, imag} */,
  {32'hbf54672b, 32'h3d2481a8} /* (15, 18, 31) {real, imag} */,
  {32'h3ed0d966, 32'hbd10af02} /* (15, 18, 30) {real, imag} */,
  {32'h3e0f1c6e, 32'h3d981aae} /* (15, 18, 29) {real, imag} */,
  {32'hbe055fb3, 32'h3e38c1e2} /* (15, 18, 28) {real, imag} */,
  {32'h3daee1ba, 32'hbe0d160f} /* (15, 18, 27) {real, imag} */,
  {32'hbcff0174, 32'hbd0a85fa} /* (15, 18, 26) {real, imag} */,
  {32'h3c5db750, 32'hbcc2c01a} /* (15, 18, 25) {real, imag} */,
  {32'h3dd11bfd, 32'h3db5aa63} /* (15, 18, 24) {real, imag} */,
  {32'h3c8ca675, 32'hbc3ef9ce} /* (15, 18, 23) {real, imag} */,
  {32'hbdc69bf1, 32'h3cb60afc} /* (15, 18, 22) {real, imag} */,
  {32'hbb920bb4, 32'h3db38f5a} /* (15, 18, 21) {real, imag} */,
  {32'h3d5774fc, 32'hbd385dce} /* (15, 18, 20) {real, imag} */,
  {32'hbd9e4911, 32'hbd01a46c} /* (15, 18, 19) {real, imag} */,
  {32'hbd7b66f9, 32'hbd6b3cb4} /* (15, 18, 18) {real, imag} */,
  {32'hbce38901, 32'hbc8612db} /* (15, 18, 17) {real, imag} */,
  {32'hbcb1e30f, 32'h00000000} /* (15, 18, 16) {real, imag} */,
  {32'hbce38901, 32'h3c8612db} /* (15, 18, 15) {real, imag} */,
  {32'hbd7b66f9, 32'h3d6b3cb4} /* (15, 18, 14) {real, imag} */,
  {32'hbd9e4911, 32'h3d01a46c} /* (15, 18, 13) {real, imag} */,
  {32'h3d5774fc, 32'h3d385dce} /* (15, 18, 12) {real, imag} */,
  {32'hbb920bb4, 32'hbdb38f5a} /* (15, 18, 11) {real, imag} */,
  {32'hbdc69bf1, 32'hbcb60afc} /* (15, 18, 10) {real, imag} */,
  {32'h3c8ca675, 32'h3c3ef9ce} /* (15, 18, 9) {real, imag} */,
  {32'h3dd11bfd, 32'hbdb5aa63} /* (15, 18, 8) {real, imag} */,
  {32'h3c5db750, 32'h3cc2c01a} /* (15, 18, 7) {real, imag} */,
  {32'hbcff0174, 32'h3d0a85fa} /* (15, 18, 6) {real, imag} */,
  {32'h3daee1ba, 32'h3e0d160f} /* (15, 18, 5) {real, imag} */,
  {32'hbe055fb3, 32'hbe38c1e2} /* (15, 18, 4) {real, imag} */,
  {32'h3e0f1c6e, 32'hbd981aae} /* (15, 18, 3) {real, imag} */,
  {32'h3ed0d966, 32'h3d10af02} /* (15, 18, 2) {real, imag} */,
  {32'hbf54672b, 32'hbd2481a8} /* (15, 18, 1) {real, imag} */,
  {32'hbef5b7dc, 32'h00000000} /* (15, 18, 0) {real, imag} */,
  {32'hbf6a0e51, 32'h3d053c50} /* (15, 17, 31) {real, imag} */,
  {32'h3ef270dd, 32'hbaf31620} /* (15, 17, 30) {real, imag} */,
  {32'h3db9067e, 32'hbd07b67a} /* (15, 17, 29) {real, imag} */,
  {32'hbcc936fe, 32'h3e363b93} /* (15, 17, 28) {real, imag} */,
  {32'h3c8be5be, 32'hbd94f4ba} /* (15, 17, 27) {real, imag} */,
  {32'hbdd8ef95, 32'h3d81df82} /* (15, 17, 26) {real, imag} */,
  {32'hbddb05d0, 32'hbd0bd1b3} /* (15, 17, 25) {real, imag} */,
  {32'h3e07a58b, 32'hbd94abe8} /* (15, 17, 24) {real, imag} */,
  {32'h3c8065bc, 32'h3c5268a2} /* (15, 17, 23) {real, imag} */,
  {32'hbdb6a4c8, 32'hbc39ba76} /* (15, 17, 22) {real, imag} */,
  {32'h3d258172, 32'hbd74ce8e} /* (15, 17, 21) {real, imag} */,
  {32'hbd86d39e, 32'hbd867952} /* (15, 17, 20) {real, imag} */,
  {32'hbc9f4e52, 32'hbd103a6e} /* (15, 17, 19) {real, imag} */,
  {32'hbc6cdfd4, 32'h3c6db26c} /* (15, 17, 18) {real, imag} */,
  {32'h3b915aa8, 32'h3d04245d} /* (15, 17, 17) {real, imag} */,
  {32'hbd4b82c8, 32'h00000000} /* (15, 17, 16) {real, imag} */,
  {32'h3b915aa8, 32'hbd04245d} /* (15, 17, 15) {real, imag} */,
  {32'hbc6cdfd4, 32'hbc6db26c} /* (15, 17, 14) {real, imag} */,
  {32'hbc9f4e52, 32'h3d103a6e} /* (15, 17, 13) {real, imag} */,
  {32'hbd86d39e, 32'h3d867952} /* (15, 17, 12) {real, imag} */,
  {32'h3d258172, 32'h3d74ce8e} /* (15, 17, 11) {real, imag} */,
  {32'hbdb6a4c8, 32'h3c39ba76} /* (15, 17, 10) {real, imag} */,
  {32'h3c8065bc, 32'hbc5268a2} /* (15, 17, 9) {real, imag} */,
  {32'h3e07a58b, 32'h3d94abe8} /* (15, 17, 8) {real, imag} */,
  {32'hbddb05d0, 32'h3d0bd1b3} /* (15, 17, 7) {real, imag} */,
  {32'hbdd8ef95, 32'hbd81df82} /* (15, 17, 6) {real, imag} */,
  {32'h3c8be5be, 32'h3d94f4ba} /* (15, 17, 5) {real, imag} */,
  {32'hbcc936fe, 32'hbe363b93} /* (15, 17, 4) {real, imag} */,
  {32'h3db9067e, 32'h3d07b67a} /* (15, 17, 3) {real, imag} */,
  {32'h3ef270dd, 32'h3af31620} /* (15, 17, 2) {real, imag} */,
  {32'hbf6a0e51, 32'hbd053c50} /* (15, 17, 1) {real, imag} */,
  {32'hbf439a26, 32'h00000000} /* (15, 17, 0) {real, imag} */,
  {32'hbf801cb5, 32'h3e4e78f5} /* (15, 16, 31) {real, imag} */,
  {32'h3f0b1472, 32'h3c01f5c0} /* (15, 16, 30) {real, imag} */,
  {32'h3e4658f0, 32'hbddd41af} /* (15, 16, 29) {real, imag} */,
  {32'hbe1134f6, 32'h3e4cb82d} /* (15, 16, 28) {real, imag} */,
  {32'hbc6be700, 32'hbd8e0496} /* (15, 16, 27) {real, imag} */,
  {32'hbdba2096, 32'h3c427c90} /* (15, 16, 26) {real, imag} */,
  {32'h3dcced87, 32'h3c50d0b5} /* (15, 16, 25) {real, imag} */,
  {32'h3d93cbcc, 32'hbd0caf2b} /* (15, 16, 24) {real, imag} */,
  {32'h3d3b2579, 32'hbd4da6a5} /* (15, 16, 23) {real, imag} */,
  {32'h3cbc2deb, 32'hbc23f363} /* (15, 16, 22) {real, imag} */,
  {32'h3d281104, 32'hbd29ede4} /* (15, 16, 21) {real, imag} */,
  {32'hbd2e6dba, 32'hbd630a9d} /* (15, 16, 20) {real, imag} */,
  {32'hbd1739f3, 32'h3d3f56b3} /* (15, 16, 19) {real, imag} */,
  {32'h3cb6b077, 32'h3d0d5739} /* (15, 16, 18) {real, imag} */,
  {32'h3d1839c4, 32'hbc30370e} /* (15, 16, 17) {real, imag} */,
  {32'h3c3201ca, 32'h00000000} /* (15, 16, 16) {real, imag} */,
  {32'h3d1839c4, 32'h3c30370e} /* (15, 16, 15) {real, imag} */,
  {32'h3cb6b077, 32'hbd0d5739} /* (15, 16, 14) {real, imag} */,
  {32'hbd1739f3, 32'hbd3f56b3} /* (15, 16, 13) {real, imag} */,
  {32'hbd2e6dba, 32'h3d630a9d} /* (15, 16, 12) {real, imag} */,
  {32'h3d281104, 32'h3d29ede4} /* (15, 16, 11) {real, imag} */,
  {32'h3cbc2deb, 32'h3c23f363} /* (15, 16, 10) {real, imag} */,
  {32'h3d3b2579, 32'h3d4da6a5} /* (15, 16, 9) {real, imag} */,
  {32'h3d93cbcc, 32'h3d0caf2b} /* (15, 16, 8) {real, imag} */,
  {32'h3dcced87, 32'hbc50d0b5} /* (15, 16, 7) {real, imag} */,
  {32'hbdba2096, 32'hbc427c90} /* (15, 16, 6) {real, imag} */,
  {32'hbc6be700, 32'h3d8e0496} /* (15, 16, 5) {real, imag} */,
  {32'hbe1134f6, 32'hbe4cb82d} /* (15, 16, 4) {real, imag} */,
  {32'h3e4658f0, 32'h3ddd41af} /* (15, 16, 3) {real, imag} */,
  {32'h3f0b1472, 32'hbc01f5c0} /* (15, 16, 2) {real, imag} */,
  {32'hbf801cb5, 32'hbe4e78f5} /* (15, 16, 1) {real, imag} */,
  {32'hbf58b48d, 32'h00000000} /* (15, 16, 0) {real, imag} */,
  {32'hbf93541e, 32'h3e86a81a} /* (15, 15, 31) {real, imag} */,
  {32'h3f0f65ad, 32'h3b96bae8} /* (15, 15, 30) {real, imag} */,
  {32'h3e03d352, 32'hbdc7d28f} /* (15, 15, 29) {real, imag} */,
  {32'hbe00caf7, 32'h3db2c5aa} /* (15, 15, 28) {real, imag} */,
  {32'hbd664d59, 32'hbd248938} /* (15, 15, 27) {real, imag} */,
  {32'hbd696dee, 32'h3e011453} /* (15, 15, 26) {real, imag} */,
  {32'h3d0c1d0c, 32'hbd09f29d} /* (15, 15, 25) {real, imag} */,
  {32'h3d85951e, 32'hbd1fea6d} /* (15, 15, 24) {real, imag} */,
  {32'h3d983181, 32'hbcd03659} /* (15, 15, 23) {real, imag} */,
  {32'hbc894f30, 32'h3b8ea6ec} /* (15, 15, 22) {real, imag} */,
  {32'hbb2e0a18, 32'h3d5114a6} /* (15, 15, 21) {real, imag} */,
  {32'h3dae2112, 32'hbd769e44} /* (15, 15, 20) {real, imag} */,
  {32'hbdd9982a, 32'h3d2b70a8} /* (15, 15, 19) {real, imag} */,
  {32'h3d5e7269, 32'hbcc36260} /* (15, 15, 18) {real, imag} */,
  {32'hbd11d0c1, 32'hbd0da55b} /* (15, 15, 17) {real, imag} */,
  {32'h3c45b216, 32'h00000000} /* (15, 15, 16) {real, imag} */,
  {32'hbd11d0c1, 32'h3d0da55b} /* (15, 15, 15) {real, imag} */,
  {32'h3d5e7269, 32'h3cc36260} /* (15, 15, 14) {real, imag} */,
  {32'hbdd9982a, 32'hbd2b70a8} /* (15, 15, 13) {real, imag} */,
  {32'h3dae2112, 32'h3d769e44} /* (15, 15, 12) {real, imag} */,
  {32'hbb2e0a18, 32'hbd5114a6} /* (15, 15, 11) {real, imag} */,
  {32'hbc894f30, 32'hbb8ea6ec} /* (15, 15, 10) {real, imag} */,
  {32'h3d983181, 32'h3cd03659} /* (15, 15, 9) {real, imag} */,
  {32'h3d85951e, 32'h3d1fea6d} /* (15, 15, 8) {real, imag} */,
  {32'h3d0c1d0c, 32'h3d09f29d} /* (15, 15, 7) {real, imag} */,
  {32'hbd696dee, 32'hbe011453} /* (15, 15, 6) {real, imag} */,
  {32'hbd664d59, 32'h3d248938} /* (15, 15, 5) {real, imag} */,
  {32'hbe00caf7, 32'hbdb2c5aa} /* (15, 15, 4) {real, imag} */,
  {32'h3e03d352, 32'h3dc7d28f} /* (15, 15, 3) {real, imag} */,
  {32'h3f0f65ad, 32'hbb96bae8} /* (15, 15, 2) {real, imag} */,
  {32'hbf93541e, 32'hbe86a81a} /* (15, 15, 1) {real, imag} */,
  {32'hbf31085a, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hbfa31fed, 32'h3ee1bec1} /* (15, 14, 31) {real, imag} */,
  {32'h3f023bfd, 32'h3db83523} /* (15, 14, 30) {real, imag} */,
  {32'h3e274f4e, 32'hbc8a35fa} /* (15, 14, 29) {real, imag} */,
  {32'hbd17590c, 32'h3e21be90} /* (15, 14, 28) {real, imag} */,
  {32'h3b35dc90, 32'hbe128fed} /* (15, 14, 27) {real, imag} */,
  {32'h3cb8cdc8, 32'hbd188bc8} /* (15, 14, 26) {real, imag} */,
  {32'h3d36942c, 32'hbdc27fb2} /* (15, 14, 25) {real, imag} */,
  {32'hbc5abdb0, 32'hbe1f4ca8} /* (15, 14, 24) {real, imag} */,
  {32'hbd37dc8e, 32'hbbb8ce1c} /* (15, 14, 23) {real, imag} */,
  {32'hbda54941, 32'h3dc35fd3} /* (15, 14, 22) {real, imag} */,
  {32'h3d236602, 32'h3c99661e} /* (15, 14, 21) {real, imag} */,
  {32'h3d222ae0, 32'hbbf29704} /* (15, 14, 20) {real, imag} */,
  {32'h3d8505c9, 32'h3d5927b2} /* (15, 14, 19) {real, imag} */,
  {32'hbd3751b7, 32'hbceaf0a8} /* (15, 14, 18) {real, imag} */,
  {32'h3d4b9a7e, 32'h3d9a049d} /* (15, 14, 17) {real, imag} */,
  {32'h3d043880, 32'h00000000} /* (15, 14, 16) {real, imag} */,
  {32'h3d4b9a7e, 32'hbd9a049d} /* (15, 14, 15) {real, imag} */,
  {32'hbd3751b7, 32'h3ceaf0a8} /* (15, 14, 14) {real, imag} */,
  {32'h3d8505c9, 32'hbd5927b2} /* (15, 14, 13) {real, imag} */,
  {32'h3d222ae0, 32'h3bf29704} /* (15, 14, 12) {real, imag} */,
  {32'h3d236602, 32'hbc99661e} /* (15, 14, 11) {real, imag} */,
  {32'hbda54941, 32'hbdc35fd3} /* (15, 14, 10) {real, imag} */,
  {32'hbd37dc8e, 32'h3bb8ce1c} /* (15, 14, 9) {real, imag} */,
  {32'hbc5abdb0, 32'h3e1f4ca8} /* (15, 14, 8) {real, imag} */,
  {32'h3d36942c, 32'h3dc27fb2} /* (15, 14, 7) {real, imag} */,
  {32'h3cb8cdc8, 32'h3d188bc8} /* (15, 14, 6) {real, imag} */,
  {32'h3b35dc90, 32'h3e128fed} /* (15, 14, 5) {real, imag} */,
  {32'hbd17590c, 32'hbe21be90} /* (15, 14, 4) {real, imag} */,
  {32'h3e274f4e, 32'h3c8a35fa} /* (15, 14, 3) {real, imag} */,
  {32'h3f023bfd, 32'hbdb83523} /* (15, 14, 2) {real, imag} */,
  {32'hbfa31fed, 32'hbee1bec1} /* (15, 14, 1) {real, imag} */,
  {32'hbf289f06, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'hbf766b5b, 32'h3ec22016} /* (15, 13, 31) {real, imag} */,
  {32'h3ee35c20, 32'hbd96d9af} /* (15, 13, 30) {real, imag} */,
  {32'h3d3aab92, 32'hbb9b3f8c} /* (15, 13, 29) {real, imag} */,
  {32'hbd97fdfb, 32'h3e45e610} /* (15, 13, 28) {real, imag} */,
  {32'h3d3c4446, 32'hbc72edfc} /* (15, 13, 27) {real, imag} */,
  {32'hbd7c66eb, 32'hbd873398} /* (15, 13, 26) {real, imag} */,
  {32'h3db574e8, 32'hbd361449} /* (15, 13, 25) {real, imag} */,
  {32'hbb7f8958, 32'hbc5e0dc0} /* (15, 13, 24) {real, imag} */,
  {32'hbd15359f, 32'h3d9d4ffa} /* (15, 13, 23) {real, imag} */,
  {32'hbdcc31b2, 32'hbd8cedad} /* (15, 13, 22) {real, imag} */,
  {32'hbd5aaa24, 32'hbd69541c} /* (15, 13, 21) {real, imag} */,
  {32'h3b3f67d0, 32'h3c0444ec} /* (15, 13, 20) {real, imag} */,
  {32'hbd0451ac, 32'h3bdcd2d0} /* (15, 13, 19) {real, imag} */,
  {32'h3bcb809a, 32'h3d0c73e3} /* (15, 13, 18) {real, imag} */,
  {32'hbdab9034, 32'h3c9c6b72} /* (15, 13, 17) {real, imag} */,
  {32'hbcb8cfee, 32'h00000000} /* (15, 13, 16) {real, imag} */,
  {32'hbdab9034, 32'hbc9c6b72} /* (15, 13, 15) {real, imag} */,
  {32'h3bcb809a, 32'hbd0c73e3} /* (15, 13, 14) {real, imag} */,
  {32'hbd0451ac, 32'hbbdcd2d0} /* (15, 13, 13) {real, imag} */,
  {32'h3b3f67d0, 32'hbc0444ec} /* (15, 13, 12) {real, imag} */,
  {32'hbd5aaa24, 32'h3d69541c} /* (15, 13, 11) {real, imag} */,
  {32'hbdcc31b2, 32'h3d8cedad} /* (15, 13, 10) {real, imag} */,
  {32'hbd15359f, 32'hbd9d4ffa} /* (15, 13, 9) {real, imag} */,
  {32'hbb7f8958, 32'h3c5e0dc0} /* (15, 13, 8) {real, imag} */,
  {32'h3db574e8, 32'h3d361449} /* (15, 13, 7) {real, imag} */,
  {32'hbd7c66eb, 32'h3d873398} /* (15, 13, 6) {real, imag} */,
  {32'h3d3c4446, 32'h3c72edfc} /* (15, 13, 5) {real, imag} */,
  {32'hbd97fdfb, 32'hbe45e610} /* (15, 13, 4) {real, imag} */,
  {32'h3d3aab92, 32'h3b9b3f8c} /* (15, 13, 3) {real, imag} */,
  {32'h3ee35c20, 32'h3d96d9af} /* (15, 13, 2) {real, imag} */,
  {32'hbf766b5b, 32'hbec22016} /* (15, 13, 1) {real, imag} */,
  {32'hbef487ac, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'hbf51fcc1, 32'h3e7ebcdc} /* (15, 12, 31) {real, imag} */,
  {32'h3eb28bbe, 32'h3b3c3690} /* (15, 12, 30) {real, imag} */,
  {32'h3d529a5a, 32'h3c47cb48} /* (15, 12, 29) {real, imag} */,
  {32'hbe41a85a, 32'h3e10c1cc} /* (15, 12, 28) {real, imag} */,
  {32'h3d9f17e1, 32'hbddbc7eb} /* (15, 12, 27) {real, imag} */,
  {32'h3e03a618, 32'h3e2bc639} /* (15, 12, 26) {real, imag} */,
  {32'hbdbe1398, 32'hbbb276c0} /* (15, 12, 25) {real, imag} */,
  {32'h3dd17254, 32'h3c47911c} /* (15, 12, 24) {real, imag} */,
  {32'hbda771b0, 32'hbd158670} /* (15, 12, 23) {real, imag} */,
  {32'h3d15e302, 32'hbb1df4ee} /* (15, 12, 22) {real, imag} */,
  {32'h3c34c3f7, 32'hbce4db50} /* (15, 12, 21) {real, imag} */,
  {32'hbd9a8674, 32'h3ba6bc02} /* (15, 12, 20) {real, imag} */,
  {32'hbda79299, 32'hbd802386} /* (15, 12, 19) {real, imag} */,
  {32'h3d92be4e, 32'h3d0f1136} /* (15, 12, 18) {real, imag} */,
  {32'h3c74c267, 32'h3d0bb792} /* (15, 12, 17) {real, imag} */,
  {32'h3b3db4a8, 32'h00000000} /* (15, 12, 16) {real, imag} */,
  {32'h3c74c267, 32'hbd0bb792} /* (15, 12, 15) {real, imag} */,
  {32'h3d92be4e, 32'hbd0f1136} /* (15, 12, 14) {real, imag} */,
  {32'hbda79299, 32'h3d802386} /* (15, 12, 13) {real, imag} */,
  {32'hbd9a8674, 32'hbba6bc02} /* (15, 12, 12) {real, imag} */,
  {32'h3c34c3f7, 32'h3ce4db50} /* (15, 12, 11) {real, imag} */,
  {32'h3d15e302, 32'h3b1df4ee} /* (15, 12, 10) {real, imag} */,
  {32'hbda771b0, 32'h3d158670} /* (15, 12, 9) {real, imag} */,
  {32'h3dd17254, 32'hbc47911c} /* (15, 12, 8) {real, imag} */,
  {32'hbdbe1398, 32'h3bb276c0} /* (15, 12, 7) {real, imag} */,
  {32'h3e03a618, 32'hbe2bc639} /* (15, 12, 6) {real, imag} */,
  {32'h3d9f17e1, 32'h3ddbc7eb} /* (15, 12, 5) {real, imag} */,
  {32'hbe41a85a, 32'hbe10c1cc} /* (15, 12, 4) {real, imag} */,
  {32'h3d529a5a, 32'hbc47cb48} /* (15, 12, 3) {real, imag} */,
  {32'h3eb28bbe, 32'hbb3c3690} /* (15, 12, 2) {real, imag} */,
  {32'hbf51fcc1, 32'hbe7ebcdc} /* (15, 12, 1) {real, imag} */,
  {32'h3c67c160, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'hbf0f5e10, 32'h3e1d23a7} /* (15, 11, 31) {real, imag} */,
  {32'h3eb9b12e, 32'h3dace6e6} /* (15, 11, 30) {real, imag} */,
  {32'h3d03712c, 32'hbcbae330} /* (15, 11, 29) {real, imag} */,
  {32'hbe0dad72, 32'h3dd87d82} /* (15, 11, 28) {real, imag} */,
  {32'h3ddadd33, 32'hbda2bc13} /* (15, 11, 27) {real, imag} */,
  {32'h3d8b1397, 32'hbd94ce8c} /* (15, 11, 26) {real, imag} */,
  {32'hbe19677d, 32'h3c6a1158} /* (15, 11, 25) {real, imag} */,
  {32'hbc87d3b8, 32'hbd16c68c} /* (15, 11, 24) {real, imag} */,
  {32'h3d6b72cb, 32'hbdb1ffd6} /* (15, 11, 23) {real, imag} */,
  {32'hbdc8cd01, 32'hbd3c3087} /* (15, 11, 22) {real, imag} */,
  {32'hbca11f72, 32'h3d1e4c4c} /* (15, 11, 21) {real, imag} */,
  {32'h3db8bd20, 32'h3d96e12d} /* (15, 11, 20) {real, imag} */,
  {32'hbda320db, 32'hbd64de8b} /* (15, 11, 19) {real, imag} */,
  {32'hbcc26082, 32'hbd862c5c} /* (15, 11, 18) {real, imag} */,
  {32'h3c464444, 32'h3dd11a84} /* (15, 11, 17) {real, imag} */,
  {32'h3cdabfa0, 32'h00000000} /* (15, 11, 16) {real, imag} */,
  {32'h3c464444, 32'hbdd11a84} /* (15, 11, 15) {real, imag} */,
  {32'hbcc26082, 32'h3d862c5c} /* (15, 11, 14) {real, imag} */,
  {32'hbda320db, 32'h3d64de8b} /* (15, 11, 13) {real, imag} */,
  {32'h3db8bd20, 32'hbd96e12d} /* (15, 11, 12) {real, imag} */,
  {32'hbca11f72, 32'hbd1e4c4c} /* (15, 11, 11) {real, imag} */,
  {32'hbdc8cd01, 32'h3d3c3087} /* (15, 11, 10) {real, imag} */,
  {32'h3d6b72cb, 32'h3db1ffd6} /* (15, 11, 9) {real, imag} */,
  {32'hbc87d3b8, 32'h3d16c68c} /* (15, 11, 8) {real, imag} */,
  {32'hbe19677d, 32'hbc6a1158} /* (15, 11, 7) {real, imag} */,
  {32'h3d8b1397, 32'h3d94ce8c} /* (15, 11, 6) {real, imag} */,
  {32'h3ddadd33, 32'h3da2bc13} /* (15, 11, 5) {real, imag} */,
  {32'hbe0dad72, 32'hbdd87d82} /* (15, 11, 4) {real, imag} */,
  {32'h3d03712c, 32'h3cbae330} /* (15, 11, 3) {real, imag} */,
  {32'h3eb9b12e, 32'hbdace6e6} /* (15, 11, 2) {real, imag} */,
  {32'hbf0f5e10, 32'hbe1d23a7} /* (15, 11, 1) {real, imag} */,
  {32'h3ecaf990, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h3e163062, 32'h3dc5dec9} /* (15, 10, 31) {real, imag} */,
  {32'h3de017a2, 32'h3e0bf050} /* (15, 10, 30) {real, imag} */,
  {32'hbd1be906, 32'hbda76b74} /* (15, 10, 29) {real, imag} */,
  {32'hbd787f8f, 32'hbcc015b8} /* (15, 10, 28) {real, imag} */,
  {32'hbd4dbeaa, 32'h3d902aa8} /* (15, 10, 27) {real, imag} */,
  {32'h3cb13544, 32'h3d12ad5d} /* (15, 10, 26) {real, imag} */,
  {32'hbd810f4e, 32'hbda89853} /* (15, 10, 25) {real, imag} */,
  {32'hbe0d4e1f, 32'h3e2e2746} /* (15, 10, 24) {real, imag} */,
  {32'h3d81574c, 32'h3cb596dc} /* (15, 10, 23) {real, imag} */,
  {32'hbd61fa1c, 32'hbd13b9dc} /* (15, 10, 22) {real, imag} */,
  {32'hbc5e7ea9, 32'hbd9594ac} /* (15, 10, 21) {real, imag} */,
  {32'h3d8d9ed0, 32'h3ce4b978} /* (15, 10, 20) {real, imag} */,
  {32'h3e053681, 32'hbd437082} /* (15, 10, 19) {real, imag} */,
  {32'h3ce7ff9b, 32'hbc82a06e} /* (15, 10, 18) {real, imag} */,
  {32'hbd496850, 32'h3e10693f} /* (15, 10, 17) {real, imag} */,
  {32'h3d973f44, 32'h00000000} /* (15, 10, 16) {real, imag} */,
  {32'hbd496850, 32'hbe10693f} /* (15, 10, 15) {real, imag} */,
  {32'h3ce7ff9b, 32'h3c82a06e} /* (15, 10, 14) {real, imag} */,
  {32'h3e053681, 32'h3d437082} /* (15, 10, 13) {real, imag} */,
  {32'h3d8d9ed0, 32'hbce4b978} /* (15, 10, 12) {real, imag} */,
  {32'hbc5e7ea9, 32'h3d9594ac} /* (15, 10, 11) {real, imag} */,
  {32'hbd61fa1c, 32'h3d13b9dc} /* (15, 10, 10) {real, imag} */,
  {32'h3d81574c, 32'hbcb596dc} /* (15, 10, 9) {real, imag} */,
  {32'hbe0d4e1f, 32'hbe2e2746} /* (15, 10, 8) {real, imag} */,
  {32'hbd810f4e, 32'h3da89853} /* (15, 10, 7) {real, imag} */,
  {32'h3cb13544, 32'hbd12ad5d} /* (15, 10, 6) {real, imag} */,
  {32'hbd4dbeaa, 32'hbd902aa8} /* (15, 10, 5) {real, imag} */,
  {32'hbd787f8f, 32'h3cc015b8} /* (15, 10, 4) {real, imag} */,
  {32'hbd1be906, 32'h3da76b74} /* (15, 10, 3) {real, imag} */,
  {32'h3de017a2, 32'hbe0bf050} /* (15, 10, 2) {real, imag} */,
  {32'h3e163062, 32'hbdc5dec9} /* (15, 10, 1) {real, imag} */,
  {32'h3f45c425, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'h3ed0f1d8, 32'hbd3af246} /* (15, 9, 31) {real, imag} */,
  {32'hbdd17a6a, 32'h3e3ae886} /* (15, 9, 30) {real, imag} */,
  {32'hbdf7c778, 32'h3d5282a0} /* (15, 9, 29) {real, imag} */,
  {32'hbd6ec624, 32'hbcae48fc} /* (15, 9, 28) {real, imag} */,
  {32'hbdfa9e31, 32'hbc6c9bc6} /* (15, 9, 27) {real, imag} */,
  {32'h3d91fc58, 32'h3e11d05a} /* (15, 9, 26) {real, imag} */,
  {32'h3d4304fc, 32'hbd99b97d} /* (15, 9, 25) {real, imag} */,
  {32'hbb4892e8, 32'h3d6ead09} /* (15, 9, 24) {real, imag} */,
  {32'hbd7ad7df, 32'hbbd2d0ad} /* (15, 9, 23) {real, imag} */,
  {32'h3ddff422, 32'hbd9a8e7a} /* (15, 9, 22) {real, imag} */,
  {32'hbcd24988, 32'hbd710b9a} /* (15, 9, 21) {real, imag} */,
  {32'hbb0f6cb8, 32'h3da16a9f} /* (15, 9, 20) {real, imag} */,
  {32'hbdfdc688, 32'hbc849f40} /* (15, 9, 19) {real, imag} */,
  {32'h3ce07239, 32'h3d0c52b7} /* (15, 9, 18) {real, imag} */,
  {32'hbd922756, 32'h3ce11d5c} /* (15, 9, 17) {real, imag} */,
  {32'h3dd920fe, 32'h00000000} /* (15, 9, 16) {real, imag} */,
  {32'hbd922756, 32'hbce11d5c} /* (15, 9, 15) {real, imag} */,
  {32'h3ce07239, 32'hbd0c52b7} /* (15, 9, 14) {real, imag} */,
  {32'hbdfdc688, 32'h3c849f40} /* (15, 9, 13) {real, imag} */,
  {32'hbb0f6cb8, 32'hbda16a9f} /* (15, 9, 12) {real, imag} */,
  {32'hbcd24988, 32'h3d710b9a} /* (15, 9, 11) {real, imag} */,
  {32'h3ddff422, 32'h3d9a8e7a} /* (15, 9, 10) {real, imag} */,
  {32'hbd7ad7df, 32'h3bd2d0ad} /* (15, 9, 9) {real, imag} */,
  {32'hbb4892e8, 32'hbd6ead09} /* (15, 9, 8) {real, imag} */,
  {32'h3d4304fc, 32'h3d99b97d} /* (15, 9, 7) {real, imag} */,
  {32'h3d91fc58, 32'hbe11d05a} /* (15, 9, 6) {real, imag} */,
  {32'hbdfa9e31, 32'h3c6c9bc6} /* (15, 9, 5) {real, imag} */,
  {32'hbd6ec624, 32'h3cae48fc} /* (15, 9, 4) {real, imag} */,
  {32'hbdf7c778, 32'hbd5282a0} /* (15, 9, 3) {real, imag} */,
  {32'hbdd17a6a, 32'hbe3ae886} /* (15, 9, 2) {real, imag} */,
  {32'h3ed0f1d8, 32'h3d3af246} /* (15, 9, 1) {real, imag} */,
  {32'h3f7aac80, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'h3eea8a56, 32'hbe2f7f8f} /* (15, 8, 31) {real, imag} */,
  {32'hbe937051, 32'h3e65a604} /* (15, 8, 30) {real, imag} */,
  {32'hbe27e8ee, 32'hbca5f018} /* (15, 8, 29) {real, imag} */,
  {32'hbc7c60ba, 32'hbdd9b348} /* (15, 8, 28) {real, imag} */,
  {32'hbde45732, 32'h3db4d965} /* (15, 8, 27) {real, imag} */,
  {32'h3dc06e56, 32'hbcbba3ba} /* (15, 8, 26) {real, imag} */,
  {32'hbcfe6ff9, 32'hbcd90afc} /* (15, 8, 25) {real, imag} */,
  {32'hbdc510a1, 32'h3dcf688e} /* (15, 8, 24) {real, imag} */,
  {32'hbd2189cd, 32'hbd99e2e8} /* (15, 8, 23) {real, imag} */,
  {32'h3da1ba26, 32'h3d21442a} /* (15, 8, 22) {real, imag} */,
  {32'h3d91ed3a, 32'h3deb50af} /* (15, 8, 21) {real, imag} */,
  {32'h3e02d50e, 32'h3dacda66} /* (15, 8, 20) {real, imag} */,
  {32'hbdae1991, 32'hbb0ca80c} /* (15, 8, 19) {real, imag} */,
  {32'hbc87b383, 32'h3c8b87b9} /* (15, 8, 18) {real, imag} */,
  {32'h3db922fa, 32'hbdae0075} /* (15, 8, 17) {real, imag} */,
  {32'h3d6eec10, 32'h00000000} /* (15, 8, 16) {real, imag} */,
  {32'h3db922fa, 32'h3dae0075} /* (15, 8, 15) {real, imag} */,
  {32'hbc87b383, 32'hbc8b87b9} /* (15, 8, 14) {real, imag} */,
  {32'hbdae1991, 32'h3b0ca80c} /* (15, 8, 13) {real, imag} */,
  {32'h3e02d50e, 32'hbdacda66} /* (15, 8, 12) {real, imag} */,
  {32'h3d91ed3a, 32'hbdeb50af} /* (15, 8, 11) {real, imag} */,
  {32'h3da1ba26, 32'hbd21442a} /* (15, 8, 10) {real, imag} */,
  {32'hbd2189cd, 32'h3d99e2e8} /* (15, 8, 9) {real, imag} */,
  {32'hbdc510a1, 32'hbdcf688e} /* (15, 8, 8) {real, imag} */,
  {32'hbcfe6ff9, 32'h3cd90afc} /* (15, 8, 7) {real, imag} */,
  {32'h3dc06e56, 32'h3cbba3ba} /* (15, 8, 6) {real, imag} */,
  {32'hbde45732, 32'hbdb4d965} /* (15, 8, 5) {real, imag} */,
  {32'hbc7c60ba, 32'h3dd9b348} /* (15, 8, 4) {real, imag} */,
  {32'hbe27e8ee, 32'h3ca5f018} /* (15, 8, 3) {real, imag} */,
  {32'hbe937051, 32'hbe65a604} /* (15, 8, 2) {real, imag} */,
  {32'h3eea8a56, 32'h3e2f7f8f} /* (15, 8, 1) {real, imag} */,
  {32'h3f81d877, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h3f137dd2, 32'hbe035fe4} /* (15, 7, 31) {real, imag} */,
  {32'hbea0f27e, 32'h3e3455dc} /* (15, 7, 30) {real, imag} */,
  {32'hbd7e14a8, 32'hbd6efbda} /* (15, 7, 29) {real, imag} */,
  {32'h3d61afb4, 32'hbe034f0c} /* (15, 7, 28) {real, imag} */,
  {32'hbe1ca6c5, 32'hbca0dc54} /* (15, 7, 27) {real, imag} */,
  {32'h3d63490f, 32'h3a4ef7e0} /* (15, 7, 26) {real, imag} */,
  {32'hbbeb5e30, 32'hbd362e38} /* (15, 7, 25) {real, imag} */,
  {32'hbd3ea9ec, 32'h3d576d4f} /* (15, 7, 24) {real, imag} */,
  {32'h3dbae2b6, 32'h3d180c82} /* (15, 7, 23) {real, imag} */,
  {32'hbc8170b7, 32'h3d96fe9e} /* (15, 7, 22) {real, imag} */,
  {32'hbd284fa0, 32'hbd4536c0} /* (15, 7, 21) {real, imag} */,
  {32'h3ce66beb, 32'hbc7d5d1c} /* (15, 7, 20) {real, imag} */,
  {32'h3d7663de, 32'h3ce4d6f0} /* (15, 7, 19) {real, imag} */,
  {32'hbd8762ef, 32'h3d495775} /* (15, 7, 18) {real, imag} */,
  {32'hbcaab788, 32'hbcaa1479} /* (15, 7, 17) {real, imag} */,
  {32'hbd606c24, 32'h00000000} /* (15, 7, 16) {real, imag} */,
  {32'hbcaab788, 32'h3caa1479} /* (15, 7, 15) {real, imag} */,
  {32'hbd8762ef, 32'hbd495775} /* (15, 7, 14) {real, imag} */,
  {32'h3d7663de, 32'hbce4d6f0} /* (15, 7, 13) {real, imag} */,
  {32'h3ce66beb, 32'h3c7d5d1c} /* (15, 7, 12) {real, imag} */,
  {32'hbd284fa0, 32'h3d4536c0} /* (15, 7, 11) {real, imag} */,
  {32'hbc8170b7, 32'hbd96fe9e} /* (15, 7, 10) {real, imag} */,
  {32'h3dbae2b6, 32'hbd180c82} /* (15, 7, 9) {real, imag} */,
  {32'hbd3ea9ec, 32'hbd576d4f} /* (15, 7, 8) {real, imag} */,
  {32'hbbeb5e30, 32'h3d362e38} /* (15, 7, 7) {real, imag} */,
  {32'h3d63490f, 32'hba4ef7e0} /* (15, 7, 6) {real, imag} */,
  {32'hbe1ca6c5, 32'h3ca0dc54} /* (15, 7, 5) {real, imag} */,
  {32'h3d61afb4, 32'h3e034f0c} /* (15, 7, 4) {real, imag} */,
  {32'hbd7e14a8, 32'h3d6efbda} /* (15, 7, 3) {real, imag} */,
  {32'hbea0f27e, 32'hbe3455dc} /* (15, 7, 2) {real, imag} */,
  {32'h3f137dd2, 32'h3e035fe4} /* (15, 7, 1) {real, imag} */,
  {32'h3f8fe642, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'h3f060ce9, 32'hbe7057ec} /* (15, 6, 31) {real, imag} */,
  {32'hbeb1347e, 32'h3e5852ba} /* (15, 6, 30) {real, imag} */,
  {32'hbac980b0, 32'h3dffa988} /* (15, 6, 29) {real, imag} */,
  {32'h3cb4af7a, 32'hbdb5d246} /* (15, 6, 28) {real, imag} */,
  {32'hbd89fbfb, 32'h3c7dba70} /* (15, 6, 27) {real, imag} */,
  {32'h3d774781, 32'hbd8ae9f4} /* (15, 6, 26) {real, imag} */,
  {32'h3ce45b5c, 32'hbd06ea9a} /* (15, 6, 25) {real, imag} */,
  {32'hbd16b851, 32'h3c957ade} /* (15, 6, 24) {real, imag} */,
  {32'hbc4695c8, 32'h3d25ae11} /* (15, 6, 23) {real, imag} */,
  {32'hbd50111c, 32'h3ca19f42} /* (15, 6, 22) {real, imag} */,
  {32'hbce9ad49, 32'h3c434d28} /* (15, 6, 21) {real, imag} */,
  {32'h3d13c718, 32'hbd825eaa} /* (15, 6, 20) {real, imag} */,
  {32'hbd25cc6e, 32'h3d300829} /* (15, 6, 19) {real, imag} */,
  {32'hbd08073c, 32'h3d7645b1} /* (15, 6, 18) {real, imag} */,
  {32'h3d3acaec, 32'h3c3fb2b4} /* (15, 6, 17) {real, imag} */,
  {32'h3d27adfd, 32'h00000000} /* (15, 6, 16) {real, imag} */,
  {32'h3d3acaec, 32'hbc3fb2b4} /* (15, 6, 15) {real, imag} */,
  {32'hbd08073c, 32'hbd7645b1} /* (15, 6, 14) {real, imag} */,
  {32'hbd25cc6e, 32'hbd300829} /* (15, 6, 13) {real, imag} */,
  {32'h3d13c718, 32'h3d825eaa} /* (15, 6, 12) {real, imag} */,
  {32'hbce9ad49, 32'hbc434d28} /* (15, 6, 11) {real, imag} */,
  {32'hbd50111c, 32'hbca19f42} /* (15, 6, 10) {real, imag} */,
  {32'hbc4695c8, 32'hbd25ae11} /* (15, 6, 9) {real, imag} */,
  {32'hbd16b851, 32'hbc957ade} /* (15, 6, 8) {real, imag} */,
  {32'h3ce45b5c, 32'h3d06ea9a} /* (15, 6, 7) {real, imag} */,
  {32'h3d774781, 32'h3d8ae9f4} /* (15, 6, 6) {real, imag} */,
  {32'hbd89fbfb, 32'hbc7dba70} /* (15, 6, 5) {real, imag} */,
  {32'h3cb4af7a, 32'h3db5d246} /* (15, 6, 4) {real, imag} */,
  {32'hbac980b0, 32'hbdffa988} /* (15, 6, 3) {real, imag} */,
  {32'hbeb1347e, 32'hbe5852ba} /* (15, 6, 2) {real, imag} */,
  {32'h3f060ce9, 32'h3e7057ec} /* (15, 6, 1) {real, imag} */,
  {32'h3f8a4351, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h3f24e6d7, 32'hbf141149} /* (15, 5, 31) {real, imag} */,
  {32'hbe37133d, 32'h3e84f25b} /* (15, 5, 30) {real, imag} */,
  {32'hbe25f50c, 32'h3debef97} /* (15, 5, 29) {real, imag} */,
  {32'hbda4c2fd, 32'hbdd99c5d} /* (15, 5, 28) {real, imag} */,
  {32'hbda447d6, 32'hbaec4080} /* (15, 5, 27) {real, imag} */,
  {32'hbd096878, 32'hbda30369} /* (15, 5, 26) {real, imag} */,
  {32'h3ddc91c2, 32'hbc252fe0} /* (15, 5, 25) {real, imag} */,
  {32'h3dd32b94, 32'h3d3b2ec8} /* (15, 5, 24) {real, imag} */,
  {32'hbdefb6cc, 32'hbcb6148c} /* (15, 5, 23) {real, imag} */,
  {32'hbd46c526, 32'h3cc288a6} /* (15, 5, 22) {real, imag} */,
  {32'hbce7b32e, 32'h3dabbae6} /* (15, 5, 21) {real, imag} */,
  {32'hbcb3c7f6, 32'h3d6ad658} /* (15, 5, 20) {real, imag} */,
  {32'hbde5034a, 32'h3d84d6fb} /* (15, 5, 19) {real, imag} */,
  {32'hbbd5fa80, 32'hbde99f8f} /* (15, 5, 18) {real, imag} */,
  {32'h3da44032, 32'h3d826ab7} /* (15, 5, 17) {real, imag} */,
  {32'h3de5db73, 32'h00000000} /* (15, 5, 16) {real, imag} */,
  {32'h3da44032, 32'hbd826ab7} /* (15, 5, 15) {real, imag} */,
  {32'hbbd5fa80, 32'h3de99f8f} /* (15, 5, 14) {real, imag} */,
  {32'hbde5034a, 32'hbd84d6fb} /* (15, 5, 13) {real, imag} */,
  {32'hbcb3c7f6, 32'hbd6ad658} /* (15, 5, 12) {real, imag} */,
  {32'hbce7b32e, 32'hbdabbae6} /* (15, 5, 11) {real, imag} */,
  {32'hbd46c526, 32'hbcc288a6} /* (15, 5, 10) {real, imag} */,
  {32'hbdefb6cc, 32'h3cb6148c} /* (15, 5, 9) {real, imag} */,
  {32'h3dd32b94, 32'hbd3b2ec8} /* (15, 5, 8) {real, imag} */,
  {32'h3ddc91c2, 32'h3c252fe0} /* (15, 5, 7) {real, imag} */,
  {32'hbd096878, 32'h3da30369} /* (15, 5, 6) {real, imag} */,
  {32'hbda447d6, 32'h3aec4080} /* (15, 5, 5) {real, imag} */,
  {32'hbda4c2fd, 32'h3dd99c5d} /* (15, 5, 4) {real, imag} */,
  {32'hbe25f50c, 32'hbdebef97} /* (15, 5, 3) {real, imag} */,
  {32'hbe37133d, 32'hbe84f25b} /* (15, 5, 2) {real, imag} */,
  {32'h3f24e6d7, 32'h3f141149} /* (15, 5, 1) {real, imag} */,
  {32'h3f85f083, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'h3f10ca53, 32'hbf4eab07} /* (15, 4, 31) {real, imag} */,
  {32'hbd0ee558, 32'h3e921ca6} /* (15, 4, 30) {real, imag} */,
  {32'hbd547fc9, 32'h3e08b5e3} /* (15, 4, 29) {real, imag} */,
  {32'hbdd688c0, 32'h3d079968} /* (15, 4, 28) {real, imag} */,
  {32'hbe005005, 32'hbc350222} /* (15, 4, 27) {real, imag} */,
  {32'h3bdc2770, 32'hbbc7a684} /* (15, 4, 26) {real, imag} */,
  {32'h3cd00a84, 32'hbc9a8278} /* (15, 4, 25) {real, imag} */,
  {32'h3d2739f1, 32'h3d6931eb} /* (15, 4, 24) {real, imag} */,
  {32'hbc6e6130, 32'hbdc39890} /* (15, 4, 23) {real, imag} */,
  {32'h3cf685be, 32'h3c850cd8} /* (15, 4, 22) {real, imag} */,
  {32'h3cee019c, 32'h3db64972} /* (15, 4, 21) {real, imag} */,
  {32'hbc8d19ba, 32'h3c908a67} /* (15, 4, 20) {real, imag} */,
  {32'h3d6944de, 32'hbd8854b8} /* (15, 4, 19) {real, imag} */,
  {32'h3b176938, 32'h3d999764} /* (15, 4, 18) {real, imag} */,
  {32'hbd7b7d3b, 32'hbb08f426} /* (15, 4, 17) {real, imag} */,
  {32'h3dc8a3b2, 32'h00000000} /* (15, 4, 16) {real, imag} */,
  {32'hbd7b7d3b, 32'h3b08f426} /* (15, 4, 15) {real, imag} */,
  {32'h3b176938, 32'hbd999764} /* (15, 4, 14) {real, imag} */,
  {32'h3d6944de, 32'h3d8854b8} /* (15, 4, 13) {real, imag} */,
  {32'hbc8d19ba, 32'hbc908a67} /* (15, 4, 12) {real, imag} */,
  {32'h3cee019c, 32'hbdb64972} /* (15, 4, 11) {real, imag} */,
  {32'h3cf685be, 32'hbc850cd8} /* (15, 4, 10) {real, imag} */,
  {32'hbc6e6130, 32'h3dc39890} /* (15, 4, 9) {real, imag} */,
  {32'h3d2739f1, 32'hbd6931eb} /* (15, 4, 8) {real, imag} */,
  {32'h3cd00a84, 32'h3c9a8278} /* (15, 4, 7) {real, imag} */,
  {32'h3bdc2770, 32'h3bc7a684} /* (15, 4, 6) {real, imag} */,
  {32'hbe005005, 32'h3c350222} /* (15, 4, 5) {real, imag} */,
  {32'hbdd688c0, 32'hbd079968} /* (15, 4, 4) {real, imag} */,
  {32'hbd547fc9, 32'hbe08b5e3} /* (15, 4, 3) {real, imag} */,
  {32'hbd0ee558, 32'hbe921ca6} /* (15, 4, 2) {real, imag} */,
  {32'h3f10ca53, 32'h3f4eab07} /* (15, 4, 1) {real, imag} */,
  {32'h3f94a8bc, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'h3f28cb0d, 32'hbf3f1f3a} /* (15, 3, 31) {real, imag} */,
  {32'hbd5af77c, 32'h3ebc6983} /* (15, 3, 30) {real, imag} */,
  {32'hbd62d89c, 32'h3d927d4c} /* (15, 3, 29) {real, imag} */,
  {32'hbe2bb559, 32'h3d81c4ae} /* (15, 3, 28) {real, imag} */,
  {32'hbde39dda, 32'hbe0390f3} /* (15, 3, 27) {real, imag} */,
  {32'h3d5bd4dd, 32'hbcf9232b} /* (15, 3, 26) {real, imag} */,
  {32'h3d1a738d, 32'hbe030a95} /* (15, 3, 25) {real, imag} */,
  {32'h3d083604, 32'hbbefa084} /* (15, 3, 24) {real, imag} */,
  {32'h3d58fa06, 32'h3c9b7aae} /* (15, 3, 23) {real, imag} */,
  {32'h3d88ba3f, 32'h3d45a270} /* (15, 3, 22) {real, imag} */,
  {32'hbcf50ca4, 32'hbc14222e} /* (15, 3, 21) {real, imag} */,
  {32'h3d678990, 32'hbc875a32} /* (15, 3, 20) {real, imag} */,
  {32'hbd2777b0, 32'h3d256761} /* (15, 3, 19) {real, imag} */,
  {32'hbc70ebc0, 32'h3cb3fda2} /* (15, 3, 18) {real, imag} */,
  {32'hbd901ea2, 32'h3d946184} /* (15, 3, 17) {real, imag} */,
  {32'h3da2185c, 32'h00000000} /* (15, 3, 16) {real, imag} */,
  {32'hbd901ea2, 32'hbd946184} /* (15, 3, 15) {real, imag} */,
  {32'hbc70ebc0, 32'hbcb3fda2} /* (15, 3, 14) {real, imag} */,
  {32'hbd2777b0, 32'hbd256761} /* (15, 3, 13) {real, imag} */,
  {32'h3d678990, 32'h3c875a32} /* (15, 3, 12) {real, imag} */,
  {32'hbcf50ca4, 32'h3c14222e} /* (15, 3, 11) {real, imag} */,
  {32'h3d88ba3f, 32'hbd45a270} /* (15, 3, 10) {real, imag} */,
  {32'h3d58fa06, 32'hbc9b7aae} /* (15, 3, 9) {real, imag} */,
  {32'h3d083604, 32'h3befa084} /* (15, 3, 8) {real, imag} */,
  {32'h3d1a738d, 32'h3e030a95} /* (15, 3, 7) {real, imag} */,
  {32'h3d5bd4dd, 32'h3cf9232b} /* (15, 3, 6) {real, imag} */,
  {32'hbde39dda, 32'h3e0390f3} /* (15, 3, 5) {real, imag} */,
  {32'hbe2bb559, 32'hbd81c4ae} /* (15, 3, 4) {real, imag} */,
  {32'hbd62d89c, 32'hbd927d4c} /* (15, 3, 3) {real, imag} */,
  {32'hbd5af77c, 32'hbebc6983} /* (15, 3, 2) {real, imag} */,
  {32'h3f28cb0d, 32'h3f3f1f3a} /* (15, 3, 1) {real, imag} */,
  {32'h3fa3c3dd, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'h3f22520b, 32'hbf421e5b} /* (15, 2, 31) {real, imag} */,
  {32'h3d9756b6, 32'h3e9c73a6} /* (15, 2, 30) {real, imag} */,
  {32'hbe17081e, 32'h3c085654} /* (15, 2, 29) {real, imag} */,
  {32'hbcd6b132, 32'h3d473dfc} /* (15, 2, 28) {real, imag} */,
  {32'hbe22c92e, 32'hbdbf9454} /* (15, 2, 27) {real, imag} */,
  {32'hbba0b520, 32'hbaadc9f0} /* (15, 2, 26) {real, imag} */,
  {32'hbcb596c4, 32'hbd22d230} /* (15, 2, 25) {real, imag} */,
  {32'h3d784639, 32'h3c164fe6} /* (15, 2, 24) {real, imag} */,
  {32'hbdfffa53, 32'h3c7ef31c} /* (15, 2, 23) {real, imag} */,
  {32'h3aef9380, 32'h3c9fd42c} /* (15, 2, 22) {real, imag} */,
  {32'hbda0503d, 32'h3b9a5884} /* (15, 2, 21) {real, imag} */,
  {32'h3d733742, 32'hbcd29489} /* (15, 2, 20) {real, imag} */,
  {32'h3a9f7270, 32'h3b56fe00} /* (15, 2, 19) {real, imag} */,
  {32'h3d6326e0, 32'h3dd22cc1} /* (15, 2, 18) {real, imag} */,
  {32'h3d0ef6c0, 32'h3bff9da0} /* (15, 2, 17) {real, imag} */,
  {32'h3db04fd6, 32'h00000000} /* (15, 2, 16) {real, imag} */,
  {32'h3d0ef6c0, 32'hbbff9da0} /* (15, 2, 15) {real, imag} */,
  {32'h3d6326e0, 32'hbdd22cc1} /* (15, 2, 14) {real, imag} */,
  {32'h3a9f7270, 32'hbb56fe00} /* (15, 2, 13) {real, imag} */,
  {32'h3d733742, 32'h3cd29489} /* (15, 2, 12) {real, imag} */,
  {32'hbda0503d, 32'hbb9a5884} /* (15, 2, 11) {real, imag} */,
  {32'h3aef9380, 32'hbc9fd42c} /* (15, 2, 10) {real, imag} */,
  {32'hbdfffa53, 32'hbc7ef31c} /* (15, 2, 9) {real, imag} */,
  {32'h3d784639, 32'hbc164fe6} /* (15, 2, 8) {real, imag} */,
  {32'hbcb596c4, 32'h3d22d230} /* (15, 2, 7) {real, imag} */,
  {32'hbba0b520, 32'h3aadc9f0} /* (15, 2, 6) {real, imag} */,
  {32'hbe22c92e, 32'h3dbf9454} /* (15, 2, 5) {real, imag} */,
  {32'hbcd6b132, 32'hbd473dfc} /* (15, 2, 4) {real, imag} */,
  {32'hbe17081e, 32'hbc085654} /* (15, 2, 3) {real, imag} */,
  {32'h3d9756b6, 32'hbe9c73a6} /* (15, 2, 2) {real, imag} */,
  {32'h3f22520b, 32'h3f421e5b} /* (15, 2, 1) {real, imag} */,
  {32'h3f9b8f6d, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'h3f08c6f7, 32'hbf6a3331} /* (15, 1, 31) {real, imag} */,
  {32'h3da58a96, 32'h3e447fc8} /* (15, 1, 30) {real, imag} */,
  {32'h3d00682f, 32'h3d643695} /* (15, 1, 29) {real, imag} */,
  {32'hbd9068c2, 32'h3db01261} /* (15, 1, 28) {real, imag} */,
  {32'hbdd37c65, 32'h3d1677e2} /* (15, 1, 27) {real, imag} */,
  {32'hbd36310b, 32'h3dbb7822} /* (15, 1, 26) {real, imag} */,
  {32'hbd9373e8, 32'hbda725a4} /* (15, 1, 25) {real, imag} */,
  {32'h3d28fe27, 32'hbca03e8a} /* (15, 1, 24) {real, imag} */,
  {32'hbd858cb3, 32'h3b89adfc} /* (15, 1, 23) {real, imag} */,
  {32'h3d09faca, 32'h3d801ea7} /* (15, 1, 22) {real, imag} */,
  {32'hbdd97192, 32'hbcae0db7} /* (15, 1, 21) {real, imag} */,
  {32'hbd2d726f, 32'h3d834c56} /* (15, 1, 20) {real, imag} */,
  {32'h3c9afe26, 32'hbcc20579} /* (15, 1, 19) {real, imag} */,
  {32'h3a9048a8, 32'hbd0ef7dd} /* (15, 1, 18) {real, imag} */,
  {32'h3d024cdc, 32'h3c17a3e1} /* (15, 1, 17) {real, imag} */,
  {32'hbd602828, 32'h00000000} /* (15, 1, 16) {real, imag} */,
  {32'h3d024cdc, 32'hbc17a3e1} /* (15, 1, 15) {real, imag} */,
  {32'h3a9048a8, 32'h3d0ef7dd} /* (15, 1, 14) {real, imag} */,
  {32'h3c9afe26, 32'h3cc20579} /* (15, 1, 13) {real, imag} */,
  {32'hbd2d726f, 32'hbd834c56} /* (15, 1, 12) {real, imag} */,
  {32'hbdd97192, 32'h3cae0db7} /* (15, 1, 11) {real, imag} */,
  {32'h3d09faca, 32'hbd801ea7} /* (15, 1, 10) {real, imag} */,
  {32'hbd858cb3, 32'hbb89adfc} /* (15, 1, 9) {real, imag} */,
  {32'h3d28fe27, 32'h3ca03e8a} /* (15, 1, 8) {real, imag} */,
  {32'hbd9373e8, 32'h3da725a4} /* (15, 1, 7) {real, imag} */,
  {32'hbd36310b, 32'hbdbb7822} /* (15, 1, 6) {real, imag} */,
  {32'hbdd37c65, 32'hbd1677e2} /* (15, 1, 5) {real, imag} */,
  {32'hbd9068c2, 32'hbdb01261} /* (15, 1, 4) {real, imag} */,
  {32'h3d00682f, 32'hbd643695} /* (15, 1, 3) {real, imag} */,
  {32'h3da58a96, 32'hbe447fc8} /* (15, 1, 2) {real, imag} */,
  {32'h3f08c6f7, 32'h3f6a3331} /* (15, 1, 1) {real, imag} */,
  {32'h3f4ec941, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'h3f15afcb, 32'hbf2b896b} /* (15, 0, 31) {real, imag} */,
  {32'hbcf9e1d0, 32'h3e238fde} /* (15, 0, 30) {real, imag} */,
  {32'hbc363970, 32'h3dc3a941} /* (15, 0, 29) {real, imag} */,
  {32'hbcf757ba, 32'h3d913e16} /* (15, 0, 28) {real, imag} */,
  {32'hbddf31fc, 32'hbc4dea82} /* (15, 0, 27) {real, imag} */,
  {32'h3b22ef10, 32'h3d98c1df} /* (15, 0, 26) {real, imag} */,
  {32'hbd8d10d7, 32'hbd0e30e3} /* (15, 0, 25) {real, imag} */,
  {32'h3d0dc387, 32'hbd19860f} /* (15, 0, 24) {real, imag} */,
  {32'hbd853214, 32'h3c7eefc4} /* (15, 0, 23) {real, imag} */,
  {32'hb999e340, 32'hbd160fef} /* (15, 0, 22) {real, imag} */,
  {32'hbc0fdaf2, 32'hbd7b9c7e} /* (15, 0, 21) {real, imag} */,
  {32'hbd29049c, 32'hbcf0c92e} /* (15, 0, 20) {real, imag} */,
  {32'h3c158728, 32'hbc7f065b} /* (15, 0, 19) {real, imag} */,
  {32'h3ccb3ef5, 32'h3d22f87b} /* (15, 0, 18) {real, imag} */,
  {32'h3bcea744, 32'hbc5d8c4e} /* (15, 0, 17) {real, imag} */,
  {32'h3c832fd1, 32'h00000000} /* (15, 0, 16) {real, imag} */,
  {32'h3bcea744, 32'h3c5d8c4e} /* (15, 0, 15) {real, imag} */,
  {32'h3ccb3ef5, 32'hbd22f87b} /* (15, 0, 14) {real, imag} */,
  {32'h3c158728, 32'h3c7f065b} /* (15, 0, 13) {real, imag} */,
  {32'hbd29049c, 32'h3cf0c92e} /* (15, 0, 12) {real, imag} */,
  {32'hbc0fdaf2, 32'h3d7b9c7e} /* (15, 0, 11) {real, imag} */,
  {32'hb999e340, 32'h3d160fef} /* (15, 0, 10) {real, imag} */,
  {32'hbd853214, 32'hbc7eefc4} /* (15, 0, 9) {real, imag} */,
  {32'h3d0dc387, 32'h3d19860f} /* (15, 0, 8) {real, imag} */,
  {32'hbd8d10d7, 32'h3d0e30e3} /* (15, 0, 7) {real, imag} */,
  {32'h3b22ef10, 32'hbd98c1df} /* (15, 0, 6) {real, imag} */,
  {32'hbddf31fc, 32'h3c4dea82} /* (15, 0, 5) {real, imag} */,
  {32'hbcf757ba, 32'hbd913e16} /* (15, 0, 4) {real, imag} */,
  {32'hbc363970, 32'hbdc3a941} /* (15, 0, 3) {real, imag} */,
  {32'hbcf9e1d0, 32'hbe238fde} /* (15, 0, 2) {real, imag} */,
  {32'h3f15afcb, 32'h3f2b896b} /* (15, 0, 1) {real, imag} */,
  {32'h3f3277c3, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h3ff3120e, 32'hbfa1e9ca} /* (14, 31, 31) {real, imag} */,
  {32'hbee6e8f9, 32'h3e90bc8c} /* (14, 31, 30) {real, imag} */,
  {32'hbc9c3b90, 32'h3dc3c85c} /* (14, 31, 29) {real, imag} */,
  {32'h3d237202, 32'hbcc661b4} /* (14, 31, 28) {real, imag} */,
  {32'hbcac1590, 32'h3c585746} /* (14, 31, 27) {real, imag} */,
  {32'hbcc924a8, 32'h3cd04472} /* (14, 31, 26) {real, imag} */,
  {32'hbb8b2f70, 32'h3d224089} /* (14, 31, 25) {real, imag} */,
  {32'h3c4c55b8, 32'h3ca60edb} /* (14, 31, 24) {real, imag} */,
  {32'hbd08378b, 32'h3cc32a29} /* (14, 31, 23) {real, imag} */,
  {32'h398fcf80, 32'hbd62eb90} /* (14, 31, 22) {real, imag} */,
  {32'hbd32eb28, 32'h3c61f31f} /* (14, 31, 21) {real, imag} */,
  {32'h3ccd5c36, 32'hbc46a7a8} /* (14, 31, 20) {real, imag} */,
  {32'h3c7765ed, 32'hbd794f6e} /* (14, 31, 19) {real, imag} */,
  {32'hbd6dedfa, 32'h3a52ad30} /* (14, 31, 18) {real, imag} */,
  {32'hbca0f109, 32'h3d0ea118} /* (14, 31, 17) {real, imag} */,
  {32'h3d681c11, 32'h00000000} /* (14, 31, 16) {real, imag} */,
  {32'hbca0f109, 32'hbd0ea118} /* (14, 31, 15) {real, imag} */,
  {32'hbd6dedfa, 32'hba52ad30} /* (14, 31, 14) {real, imag} */,
  {32'h3c7765ed, 32'h3d794f6e} /* (14, 31, 13) {real, imag} */,
  {32'h3ccd5c36, 32'h3c46a7a8} /* (14, 31, 12) {real, imag} */,
  {32'hbd32eb28, 32'hbc61f31f} /* (14, 31, 11) {real, imag} */,
  {32'h398fcf80, 32'h3d62eb90} /* (14, 31, 10) {real, imag} */,
  {32'hbd08378b, 32'hbcc32a29} /* (14, 31, 9) {real, imag} */,
  {32'h3c4c55b8, 32'hbca60edb} /* (14, 31, 8) {real, imag} */,
  {32'hbb8b2f70, 32'hbd224089} /* (14, 31, 7) {real, imag} */,
  {32'hbcc924a8, 32'hbcd04472} /* (14, 31, 6) {real, imag} */,
  {32'hbcac1590, 32'hbc585746} /* (14, 31, 5) {real, imag} */,
  {32'h3d237202, 32'h3cc661b4} /* (14, 31, 4) {real, imag} */,
  {32'hbc9c3b90, 32'hbdc3c85c} /* (14, 31, 3) {real, imag} */,
  {32'hbee6e8f9, 32'hbe90bc8c} /* (14, 31, 2) {real, imag} */,
  {32'h3ff3120e, 32'h3fa1e9ca} /* (14, 31, 1) {real, imag} */,
  {32'h401a6f8e, 32'h00000000} /* (14, 31, 0) {real, imag} */,
  {32'h40157487, 32'hbf93bace} /* (14, 30, 31) {real, imag} */,
  {32'hbf6858c5, 32'h3e37a81f} /* (14, 30, 30) {real, imag} */,
  {32'h3d6c9417, 32'h3e03f189} /* (14, 30, 29) {real, imag} */,
  {32'h3e4a2995, 32'h3be6df50} /* (14, 30, 28) {real, imag} */,
  {32'hbd081c6c, 32'h3c0d0d2a} /* (14, 30, 27) {real, imag} */,
  {32'h3d27e94a, 32'hbdd9ebef} /* (14, 30, 26) {real, imag} */,
  {32'hbbdb5be8, 32'h3d831f14} /* (14, 30, 25) {real, imag} */,
  {32'h3d2c7be5, 32'h3db593ee} /* (14, 30, 24) {real, imag} */,
  {32'hbd9dd30a, 32'hbc1e4494} /* (14, 30, 23) {real, imag} */,
  {32'h3e030f37, 32'h3d89f147} /* (14, 30, 22) {real, imag} */,
  {32'hbb68d368, 32'h3d637e56} /* (14, 30, 21) {real, imag} */,
  {32'h3d8b9e29, 32'h3b6c4430} /* (14, 30, 20) {real, imag} */,
  {32'hbd675ba0, 32'hbd117978} /* (14, 30, 19) {real, imag} */,
  {32'h3b0eb058, 32'h3d5fc270} /* (14, 30, 18) {real, imag} */,
  {32'h3cb9c76c, 32'h3d6a8110} /* (14, 30, 17) {real, imag} */,
  {32'h3d450735, 32'h00000000} /* (14, 30, 16) {real, imag} */,
  {32'h3cb9c76c, 32'hbd6a8110} /* (14, 30, 15) {real, imag} */,
  {32'h3b0eb058, 32'hbd5fc270} /* (14, 30, 14) {real, imag} */,
  {32'hbd675ba0, 32'h3d117978} /* (14, 30, 13) {real, imag} */,
  {32'h3d8b9e29, 32'hbb6c4430} /* (14, 30, 12) {real, imag} */,
  {32'hbb68d368, 32'hbd637e56} /* (14, 30, 11) {real, imag} */,
  {32'h3e030f37, 32'hbd89f147} /* (14, 30, 10) {real, imag} */,
  {32'hbd9dd30a, 32'h3c1e4494} /* (14, 30, 9) {real, imag} */,
  {32'h3d2c7be5, 32'hbdb593ee} /* (14, 30, 8) {real, imag} */,
  {32'hbbdb5be8, 32'hbd831f14} /* (14, 30, 7) {real, imag} */,
  {32'h3d27e94a, 32'h3dd9ebef} /* (14, 30, 6) {real, imag} */,
  {32'hbd081c6c, 32'hbc0d0d2a} /* (14, 30, 5) {real, imag} */,
  {32'h3e4a2995, 32'hbbe6df50} /* (14, 30, 4) {real, imag} */,
  {32'h3d6c9417, 32'hbe03f189} /* (14, 30, 3) {real, imag} */,
  {32'hbf6858c5, 32'hbe37a81f} /* (14, 30, 2) {real, imag} */,
  {32'h40157487, 32'h3f93bace} /* (14, 30, 1) {real, imag} */,
  {32'h401ebfd6, 32'h00000000} /* (14, 30, 0) {real, imag} */,
  {32'h401a9d66, 32'hbf3ff838} /* (14, 29, 31) {real, imag} */,
  {32'hbf5c8030, 32'h3e109618} /* (14, 29, 30) {real, imag} */,
  {32'h3d7a3e93, 32'h3d8c97f8} /* (14, 29, 29) {real, imag} */,
  {32'h3daa35d8, 32'hbd1efe4f} /* (14, 29, 28) {real, imag} */,
  {32'hbcc04220, 32'hbb5c4cb0} /* (14, 29, 27) {real, imag} */,
  {32'h3d9c3d9a, 32'h3bafbba2} /* (14, 29, 26) {real, imag} */,
  {32'h3e1b73bb, 32'h3d84a81c} /* (14, 29, 25) {real, imag} */,
  {32'h3bdac28a, 32'h3db5978d} /* (14, 29, 24) {real, imag} */,
  {32'hbd4ec9ae, 32'h3cfb5852} /* (14, 29, 23) {real, imag} */,
  {32'hbc8c4af4, 32'h3de3f65c} /* (14, 29, 22) {real, imag} */,
  {32'hbd0ab5d8, 32'h3d46279d} /* (14, 29, 21) {real, imag} */,
  {32'h3c0694a8, 32'h3c83d635} /* (14, 29, 20) {real, imag} */,
  {32'h3c49e7c4, 32'h3db19d8a} /* (14, 29, 19) {real, imag} */,
  {32'hbbff5c20, 32'h3db2cadd} /* (14, 29, 18) {real, imag} */,
  {32'h37829000, 32'hbd0d2efe} /* (14, 29, 17) {real, imag} */,
  {32'hbdb5a5f6, 32'h00000000} /* (14, 29, 16) {real, imag} */,
  {32'h37829000, 32'h3d0d2efe} /* (14, 29, 15) {real, imag} */,
  {32'hbbff5c20, 32'hbdb2cadd} /* (14, 29, 14) {real, imag} */,
  {32'h3c49e7c4, 32'hbdb19d8a} /* (14, 29, 13) {real, imag} */,
  {32'h3c0694a8, 32'hbc83d635} /* (14, 29, 12) {real, imag} */,
  {32'hbd0ab5d8, 32'hbd46279d} /* (14, 29, 11) {real, imag} */,
  {32'hbc8c4af4, 32'hbde3f65c} /* (14, 29, 10) {real, imag} */,
  {32'hbd4ec9ae, 32'hbcfb5852} /* (14, 29, 9) {real, imag} */,
  {32'h3bdac28a, 32'hbdb5978d} /* (14, 29, 8) {real, imag} */,
  {32'h3e1b73bb, 32'hbd84a81c} /* (14, 29, 7) {real, imag} */,
  {32'h3d9c3d9a, 32'hbbafbba2} /* (14, 29, 6) {real, imag} */,
  {32'hbcc04220, 32'h3b5c4cb0} /* (14, 29, 5) {real, imag} */,
  {32'h3daa35d8, 32'h3d1efe4f} /* (14, 29, 4) {real, imag} */,
  {32'h3d7a3e93, 32'hbd8c97f8} /* (14, 29, 3) {real, imag} */,
  {32'hbf5c8030, 32'hbe109618} /* (14, 29, 2) {real, imag} */,
  {32'h401a9d66, 32'h3f3ff838} /* (14, 29, 1) {real, imag} */,
  {32'h402149c2, 32'h00000000} /* (14, 29, 0) {real, imag} */,
  {32'h40181b21, 32'hbf11fa9b} /* (14, 28, 31) {real, imag} */,
  {32'hbf839fd8, 32'h3df5e508} /* (14, 28, 30) {real, imag} */,
  {32'h3db183bd, 32'hbd27ed10} /* (14, 28, 29) {real, imag} */,
  {32'hbc8657ac, 32'hbdfaf042} /* (14, 28, 28) {real, imag} */,
  {32'hbd4e8b36, 32'h3e1825a0} /* (14, 28, 27) {real, imag} */,
  {32'h3b202460, 32'hbcb8453e} /* (14, 28, 26) {real, imag} */,
  {32'h3dfc849b, 32'hba918180} /* (14, 28, 25) {real, imag} */,
  {32'h3af06758, 32'h3d83eb76} /* (14, 28, 24) {real, imag} */,
  {32'hbdb06890, 32'h3cb4bc44} /* (14, 28, 23) {real, imag} */,
  {32'hbc4eece0, 32'hbdcd8d08} /* (14, 28, 22) {real, imag} */,
  {32'h3d3e1224, 32'h3d64a7de} /* (14, 28, 21) {real, imag} */,
  {32'hbcd4a852, 32'h3ce3ed07} /* (14, 28, 20) {real, imag} */,
  {32'h3cbae2df, 32'hbc59e710} /* (14, 28, 19) {real, imag} */,
  {32'hbcafddd4, 32'h3d1eb019} /* (14, 28, 18) {real, imag} */,
  {32'h3d11e41f, 32'h3b92c938} /* (14, 28, 17) {real, imag} */,
  {32'hbc9f87c1, 32'h00000000} /* (14, 28, 16) {real, imag} */,
  {32'h3d11e41f, 32'hbb92c938} /* (14, 28, 15) {real, imag} */,
  {32'hbcafddd4, 32'hbd1eb019} /* (14, 28, 14) {real, imag} */,
  {32'h3cbae2df, 32'h3c59e710} /* (14, 28, 13) {real, imag} */,
  {32'hbcd4a852, 32'hbce3ed07} /* (14, 28, 12) {real, imag} */,
  {32'h3d3e1224, 32'hbd64a7de} /* (14, 28, 11) {real, imag} */,
  {32'hbc4eece0, 32'h3dcd8d08} /* (14, 28, 10) {real, imag} */,
  {32'hbdb06890, 32'hbcb4bc44} /* (14, 28, 9) {real, imag} */,
  {32'h3af06758, 32'hbd83eb76} /* (14, 28, 8) {real, imag} */,
  {32'h3dfc849b, 32'h3a918180} /* (14, 28, 7) {real, imag} */,
  {32'h3b202460, 32'h3cb8453e} /* (14, 28, 6) {real, imag} */,
  {32'hbd4e8b36, 32'hbe1825a0} /* (14, 28, 5) {real, imag} */,
  {32'hbc8657ac, 32'h3dfaf042} /* (14, 28, 4) {real, imag} */,
  {32'h3db183bd, 32'h3d27ed10} /* (14, 28, 3) {real, imag} */,
  {32'hbf839fd8, 32'hbdf5e508} /* (14, 28, 2) {real, imag} */,
  {32'h40181b21, 32'h3f11fa9b} /* (14, 28, 1) {real, imag} */,
  {32'h4023b8b1, 32'h00000000} /* (14, 28, 0) {real, imag} */,
  {32'h4019c6cf, 32'hbf1d6277} /* (14, 27, 31) {real, imag} */,
  {32'hbf887f53, 32'h3e686a51} /* (14, 27, 30) {real, imag} */,
  {32'hbd0255af, 32'hbe011b4c} /* (14, 27, 29) {real, imag} */,
  {32'h3d795972, 32'hbea38308} /* (14, 27, 28) {real, imag} */,
  {32'hbe0d4274, 32'h3e3428b2} /* (14, 27, 27) {real, imag} */,
  {32'hbdaa4c00, 32'hba8988a0} /* (14, 27, 26) {real, imag} */,
  {32'hbc744134, 32'hbd55d29e} /* (14, 27, 25) {real, imag} */,
  {32'hbd9e4f78, 32'h3e40f148} /* (14, 27, 24) {real, imag} */,
  {32'hbde827b5, 32'h3bc2be64} /* (14, 27, 23) {real, imag} */,
  {32'h3d1153d7, 32'hbdfc2cfa} /* (14, 27, 22) {real, imag} */,
  {32'h3cb5921f, 32'h3e0db24a} /* (14, 27, 21) {real, imag} */,
  {32'hbcab20de, 32'hbd6b03c8} /* (14, 27, 20) {real, imag} */,
  {32'h3d8ded5a, 32'hbd2973b8} /* (14, 27, 19) {real, imag} */,
  {32'hbdaca7ed, 32'h3d4fe81e} /* (14, 27, 18) {real, imag} */,
  {32'h3d51d5d9, 32'hbd049f3e} /* (14, 27, 17) {real, imag} */,
  {32'h3dcb09b2, 32'h00000000} /* (14, 27, 16) {real, imag} */,
  {32'h3d51d5d9, 32'h3d049f3e} /* (14, 27, 15) {real, imag} */,
  {32'hbdaca7ed, 32'hbd4fe81e} /* (14, 27, 14) {real, imag} */,
  {32'h3d8ded5a, 32'h3d2973b8} /* (14, 27, 13) {real, imag} */,
  {32'hbcab20de, 32'h3d6b03c8} /* (14, 27, 12) {real, imag} */,
  {32'h3cb5921f, 32'hbe0db24a} /* (14, 27, 11) {real, imag} */,
  {32'h3d1153d7, 32'h3dfc2cfa} /* (14, 27, 10) {real, imag} */,
  {32'hbde827b5, 32'hbbc2be64} /* (14, 27, 9) {real, imag} */,
  {32'hbd9e4f78, 32'hbe40f148} /* (14, 27, 8) {real, imag} */,
  {32'hbc744134, 32'h3d55d29e} /* (14, 27, 7) {real, imag} */,
  {32'hbdaa4c00, 32'h3a8988a0} /* (14, 27, 6) {real, imag} */,
  {32'hbe0d4274, 32'hbe3428b2} /* (14, 27, 5) {real, imag} */,
  {32'h3d795972, 32'h3ea38308} /* (14, 27, 4) {real, imag} */,
  {32'hbd0255af, 32'h3e011b4c} /* (14, 27, 3) {real, imag} */,
  {32'hbf887f53, 32'hbe686a51} /* (14, 27, 2) {real, imag} */,
  {32'h4019c6cf, 32'h3f1d6277} /* (14, 27, 1) {real, imag} */,
  {32'h40249dc7, 32'h00000000} /* (14, 27, 0) {real, imag} */,
  {32'h40229fee, 32'hbeeaa004} /* (14, 26, 31) {real, imag} */,
  {32'hbf9036d2, 32'h3e808881} /* (14, 26, 30) {real, imag} */,
  {32'hbdfc3c81, 32'hbdab8fe4} /* (14, 26, 29) {real, imag} */,
  {32'h3d208ee0, 32'hbe0e861c} /* (14, 26, 28) {real, imag} */,
  {32'hbd1805be, 32'h3e2d708f} /* (14, 26, 27) {real, imag} */,
  {32'hbd2ee8cc, 32'h3dd2ad62} /* (14, 26, 26) {real, imag} */,
  {32'hbd38168e, 32'h3d84b0b9} /* (14, 26, 25) {real, imag} */,
  {32'hbd304444, 32'h3d414ca6} /* (14, 26, 24) {real, imag} */,
  {32'h3e060d30, 32'hbd48b4b2} /* (14, 26, 23) {real, imag} */,
  {32'h3ba5f618, 32'hbd9bb1b4} /* (14, 26, 22) {real, imag} */,
  {32'hbc8cb7fe, 32'h3d12f57e} /* (14, 26, 21) {real, imag} */,
  {32'hbd0b4417, 32'h3beffa20} /* (14, 26, 20) {real, imag} */,
  {32'h3dd01edf, 32'hbac571b0} /* (14, 26, 19) {real, imag} */,
  {32'hbd7966c2, 32'h3d38b0f3} /* (14, 26, 18) {real, imag} */,
  {32'h3d7ba604, 32'hbd8365f0} /* (14, 26, 17) {real, imag} */,
  {32'hbb8281c0, 32'h00000000} /* (14, 26, 16) {real, imag} */,
  {32'h3d7ba604, 32'h3d8365f0} /* (14, 26, 15) {real, imag} */,
  {32'hbd7966c2, 32'hbd38b0f3} /* (14, 26, 14) {real, imag} */,
  {32'h3dd01edf, 32'h3ac571b0} /* (14, 26, 13) {real, imag} */,
  {32'hbd0b4417, 32'hbbeffa20} /* (14, 26, 12) {real, imag} */,
  {32'hbc8cb7fe, 32'hbd12f57e} /* (14, 26, 11) {real, imag} */,
  {32'h3ba5f618, 32'h3d9bb1b4} /* (14, 26, 10) {real, imag} */,
  {32'h3e060d30, 32'h3d48b4b2} /* (14, 26, 9) {real, imag} */,
  {32'hbd304444, 32'hbd414ca6} /* (14, 26, 8) {real, imag} */,
  {32'hbd38168e, 32'hbd84b0b9} /* (14, 26, 7) {real, imag} */,
  {32'hbd2ee8cc, 32'hbdd2ad62} /* (14, 26, 6) {real, imag} */,
  {32'hbd1805be, 32'hbe2d708f} /* (14, 26, 5) {real, imag} */,
  {32'h3d208ee0, 32'h3e0e861c} /* (14, 26, 4) {real, imag} */,
  {32'hbdfc3c81, 32'h3dab8fe4} /* (14, 26, 3) {real, imag} */,
  {32'hbf9036d2, 32'hbe808881} /* (14, 26, 2) {real, imag} */,
  {32'h40229fee, 32'h3eeaa004} /* (14, 26, 1) {real, imag} */,
  {32'h401693d3, 32'h00000000} /* (14, 26, 0) {real, imag} */,
  {32'h40257c8b, 32'hbef087fc} /* (14, 25, 31) {real, imag} */,
  {32'hbf984704, 32'h3e682560} /* (14, 25, 30) {real, imag} */,
  {32'h3cc6ec0a, 32'hbd283eb8} /* (14, 25, 29) {real, imag} */,
  {32'h3dbf6a38, 32'hbdd60a41} /* (14, 25, 28) {real, imag} */,
  {32'hbe611ef6, 32'h3de88991} /* (14, 25, 27) {real, imag} */,
  {32'h3d75da5a, 32'hbb054c10} /* (14, 25, 26) {real, imag} */,
  {32'h3ca78410, 32'h3da31e89} /* (14, 25, 25) {real, imag} */,
  {32'hbde25446, 32'h3d7e5442} /* (14, 25, 24) {real, imag} */,
  {32'h3da78ea1, 32'hbd0d765e} /* (14, 25, 23) {real, imag} */,
  {32'hbdf89de0, 32'hbc8fd3ca} /* (14, 25, 22) {real, imag} */,
  {32'hbd15f34b, 32'h3d7750da} /* (14, 25, 21) {real, imag} */,
  {32'h3bcce074, 32'h3d8fb8ec} /* (14, 25, 20) {real, imag} */,
  {32'h3b159d68, 32'h3d742eb3} /* (14, 25, 19) {real, imag} */,
  {32'h3cd1daf6, 32'h3b7c9850} /* (14, 25, 18) {real, imag} */,
  {32'hbc39dfe5, 32'h3d5f1efc} /* (14, 25, 17) {real, imag} */,
  {32'hbd82a708, 32'h00000000} /* (14, 25, 16) {real, imag} */,
  {32'hbc39dfe5, 32'hbd5f1efc} /* (14, 25, 15) {real, imag} */,
  {32'h3cd1daf6, 32'hbb7c9850} /* (14, 25, 14) {real, imag} */,
  {32'h3b159d68, 32'hbd742eb3} /* (14, 25, 13) {real, imag} */,
  {32'h3bcce074, 32'hbd8fb8ec} /* (14, 25, 12) {real, imag} */,
  {32'hbd15f34b, 32'hbd7750da} /* (14, 25, 11) {real, imag} */,
  {32'hbdf89de0, 32'h3c8fd3ca} /* (14, 25, 10) {real, imag} */,
  {32'h3da78ea1, 32'h3d0d765e} /* (14, 25, 9) {real, imag} */,
  {32'hbde25446, 32'hbd7e5442} /* (14, 25, 8) {real, imag} */,
  {32'h3ca78410, 32'hbda31e89} /* (14, 25, 7) {real, imag} */,
  {32'h3d75da5a, 32'h3b054c10} /* (14, 25, 6) {real, imag} */,
  {32'hbe611ef6, 32'hbde88991} /* (14, 25, 5) {real, imag} */,
  {32'h3dbf6a38, 32'h3dd60a41} /* (14, 25, 4) {real, imag} */,
  {32'h3cc6ec0a, 32'h3d283eb8} /* (14, 25, 3) {real, imag} */,
  {32'hbf984704, 32'hbe682560} /* (14, 25, 2) {real, imag} */,
  {32'h40257c8b, 32'h3ef087fc} /* (14, 25, 1) {real, imag} */,
  {32'h40063682, 32'h00000000} /* (14, 25, 0) {real, imag} */,
  {32'h4019b710, 32'hbecf621a} /* (14, 24, 31) {real, imag} */,
  {32'hbf898d34, 32'h3eba2558} /* (14, 24, 30) {real, imag} */,
  {32'h3cc46cde, 32'hbe3b7c8f} /* (14, 24, 29) {real, imag} */,
  {32'h3e222fde, 32'hbe3f4b6b} /* (14, 24, 28) {real, imag} */,
  {32'hbe816bb6, 32'h3e322795} /* (14, 24, 27) {real, imag} */,
  {32'hbe0e5f6a, 32'h3ae89e00} /* (14, 24, 26) {real, imag} */,
  {32'h3e1bc801, 32'hbd8576df} /* (14, 24, 25) {real, imag} */,
  {32'h3d21ed74, 32'hbcad5092} /* (14, 24, 24) {real, imag} */,
  {32'h3d643858, 32'hbcaf07e0} /* (14, 24, 23) {real, imag} */,
  {32'hbd521334, 32'hbd836a68} /* (14, 24, 22) {real, imag} */,
  {32'hbd5624bc, 32'h3d0684ec} /* (14, 24, 21) {real, imag} */,
  {32'hbd8774d2, 32'h3d341d3e} /* (14, 24, 20) {real, imag} */,
  {32'hbd428e0c, 32'hbad880f0} /* (14, 24, 19) {real, imag} */,
  {32'hbdee75a9, 32'h3b9be9a0} /* (14, 24, 18) {real, imag} */,
  {32'hbdc1b31c, 32'h3d777724} /* (14, 24, 17) {real, imag} */,
  {32'hbc718c32, 32'h00000000} /* (14, 24, 16) {real, imag} */,
  {32'hbdc1b31c, 32'hbd777724} /* (14, 24, 15) {real, imag} */,
  {32'hbdee75a9, 32'hbb9be9a0} /* (14, 24, 14) {real, imag} */,
  {32'hbd428e0c, 32'h3ad880f0} /* (14, 24, 13) {real, imag} */,
  {32'hbd8774d2, 32'hbd341d3e} /* (14, 24, 12) {real, imag} */,
  {32'hbd5624bc, 32'hbd0684ec} /* (14, 24, 11) {real, imag} */,
  {32'hbd521334, 32'h3d836a68} /* (14, 24, 10) {real, imag} */,
  {32'h3d643858, 32'h3caf07e0} /* (14, 24, 9) {real, imag} */,
  {32'h3d21ed74, 32'h3cad5092} /* (14, 24, 8) {real, imag} */,
  {32'h3e1bc801, 32'h3d8576df} /* (14, 24, 7) {real, imag} */,
  {32'hbe0e5f6a, 32'hbae89e00} /* (14, 24, 6) {real, imag} */,
  {32'hbe816bb6, 32'hbe322795} /* (14, 24, 5) {real, imag} */,
  {32'h3e222fde, 32'h3e3f4b6b} /* (14, 24, 4) {real, imag} */,
  {32'h3cc46cde, 32'h3e3b7c8f} /* (14, 24, 3) {real, imag} */,
  {32'hbf898d34, 32'hbeba2558} /* (14, 24, 2) {real, imag} */,
  {32'h4019b710, 32'h3ecf621a} /* (14, 24, 1) {real, imag} */,
  {32'h3fe49fb3, 32'h00000000} /* (14, 24, 0) {real, imag} */,
  {32'h3ffe9254, 32'hbe88e780} /* (14, 23, 31) {real, imag} */,
  {32'hbf67c811, 32'h3e73f35c} /* (14, 23, 30) {real, imag} */,
  {32'h3d6d37a9, 32'hbe26bfc2} /* (14, 23, 29) {real, imag} */,
  {32'h3e03c72e, 32'hbe249cd6} /* (14, 23, 28) {real, imag} */,
  {32'hbe352074, 32'h3d952570} /* (14, 23, 27) {real, imag} */,
  {32'hbbfb8580, 32'hbc4d421a} /* (14, 23, 26) {real, imag} */,
  {32'h3dfdd4f1, 32'h3cdda000} /* (14, 23, 25) {real, imag} */,
  {32'hbd0aebc5, 32'h3c91762a} /* (14, 23, 24) {real, imag} */,
  {32'hbc1c1d80, 32'h3de64c16} /* (14, 23, 23) {real, imag} */,
  {32'hbcf876a4, 32'hbddb8856} /* (14, 23, 22) {real, imag} */,
  {32'h3d4d8cee, 32'hbd0e0b06} /* (14, 23, 21) {real, imag} */,
  {32'h3d105eac, 32'h3d107313} /* (14, 23, 20) {real, imag} */,
  {32'h3c496bc2, 32'h3d3eb35a} /* (14, 23, 19) {real, imag} */,
  {32'hbac36e68, 32'h3d8aa58f} /* (14, 23, 18) {real, imag} */,
  {32'h3d3a87b2, 32'h3d213bd6} /* (14, 23, 17) {real, imag} */,
  {32'hbc49cc16, 32'h00000000} /* (14, 23, 16) {real, imag} */,
  {32'h3d3a87b2, 32'hbd213bd6} /* (14, 23, 15) {real, imag} */,
  {32'hbac36e68, 32'hbd8aa58f} /* (14, 23, 14) {real, imag} */,
  {32'h3c496bc2, 32'hbd3eb35a} /* (14, 23, 13) {real, imag} */,
  {32'h3d105eac, 32'hbd107313} /* (14, 23, 12) {real, imag} */,
  {32'h3d4d8cee, 32'h3d0e0b06} /* (14, 23, 11) {real, imag} */,
  {32'hbcf876a4, 32'h3ddb8856} /* (14, 23, 10) {real, imag} */,
  {32'hbc1c1d80, 32'hbde64c16} /* (14, 23, 9) {real, imag} */,
  {32'hbd0aebc5, 32'hbc91762a} /* (14, 23, 8) {real, imag} */,
  {32'h3dfdd4f1, 32'hbcdda000} /* (14, 23, 7) {real, imag} */,
  {32'hbbfb8580, 32'h3c4d421a} /* (14, 23, 6) {real, imag} */,
  {32'hbe352074, 32'hbd952570} /* (14, 23, 5) {real, imag} */,
  {32'h3e03c72e, 32'h3e249cd6} /* (14, 23, 4) {real, imag} */,
  {32'h3d6d37a9, 32'h3e26bfc2} /* (14, 23, 3) {real, imag} */,
  {32'hbf67c811, 32'hbe73f35c} /* (14, 23, 2) {real, imag} */,
  {32'h3ffe9254, 32'h3e88e780} /* (14, 23, 1) {real, imag} */,
  {32'h3faa08e2, 32'h00000000} /* (14, 23, 0) {real, imag} */,
  {32'h3fb4b1a7, 32'hbe300817} /* (14, 22, 31) {real, imag} */,
  {32'hbf21733d, 32'h3e2ab9d6} /* (14, 22, 30) {real, imag} */,
  {32'h3c3a4670, 32'hbe2d93a4} /* (14, 22, 29) {real, imag} */,
  {32'h3e159aa6, 32'hbe65557e} /* (14, 22, 28) {real, imag} */,
  {32'hbe3e53a0, 32'h3dcb2c7a} /* (14, 22, 27) {real, imag} */,
  {32'hbd8efbd0, 32'h3d809522} /* (14, 22, 26) {real, imag} */,
  {32'h3df92e79, 32'h3cce29c9} /* (14, 22, 25) {real, imag} */,
  {32'hbd237ddc, 32'h3db5ed98} /* (14, 22, 24) {real, imag} */,
  {32'hbdd127de, 32'h3e186f21} /* (14, 22, 23) {real, imag} */,
  {32'hbd1cd015, 32'h3d1876ae} /* (14, 22, 22) {real, imag} */,
  {32'hbdd7be15, 32'hbda1f628} /* (14, 22, 21) {real, imag} */,
  {32'h3d8259da, 32'hbd9c7d36} /* (14, 22, 20) {real, imag} */,
  {32'h3cd7db8f, 32'hbbbfd830} /* (14, 22, 19) {real, imag} */,
  {32'hbd26cd0e, 32'h3d438c8c} /* (14, 22, 18) {real, imag} */,
  {32'hbcb46e6a, 32'hbde52132} /* (14, 22, 17) {real, imag} */,
  {32'h3d804c96, 32'h00000000} /* (14, 22, 16) {real, imag} */,
  {32'hbcb46e6a, 32'h3de52132} /* (14, 22, 15) {real, imag} */,
  {32'hbd26cd0e, 32'hbd438c8c} /* (14, 22, 14) {real, imag} */,
  {32'h3cd7db8f, 32'h3bbfd830} /* (14, 22, 13) {real, imag} */,
  {32'h3d8259da, 32'h3d9c7d36} /* (14, 22, 12) {real, imag} */,
  {32'hbdd7be15, 32'h3da1f628} /* (14, 22, 11) {real, imag} */,
  {32'hbd1cd015, 32'hbd1876ae} /* (14, 22, 10) {real, imag} */,
  {32'hbdd127de, 32'hbe186f21} /* (14, 22, 9) {real, imag} */,
  {32'hbd237ddc, 32'hbdb5ed98} /* (14, 22, 8) {real, imag} */,
  {32'h3df92e79, 32'hbcce29c9} /* (14, 22, 7) {real, imag} */,
  {32'hbd8efbd0, 32'hbd809522} /* (14, 22, 6) {real, imag} */,
  {32'hbe3e53a0, 32'hbdcb2c7a} /* (14, 22, 5) {real, imag} */,
  {32'h3e159aa6, 32'h3e65557e} /* (14, 22, 4) {real, imag} */,
  {32'h3c3a4670, 32'h3e2d93a4} /* (14, 22, 3) {real, imag} */,
  {32'hbf21733d, 32'hbe2ab9d6} /* (14, 22, 2) {real, imag} */,
  {32'h3fb4b1a7, 32'h3e300817} /* (14, 22, 1) {real, imag} */,
  {32'h3f983438, 32'h00000000} /* (14, 22, 0) {real, imag} */,
  {32'h3ec06862, 32'h3da054c0} /* (14, 21, 31) {real, imag} */,
  {32'hbe4af16d, 32'h3e22a25f} /* (14, 21, 30) {real, imag} */,
  {32'h3dec9d13, 32'hbdf0fef9} /* (14, 21, 29) {real, imag} */,
  {32'h3dff8134, 32'hbdfdd604} /* (14, 21, 28) {real, imag} */,
  {32'hbe085644, 32'h3dc35fe7} /* (14, 21, 27) {real, imag} */,
  {32'hbdcc8c9c, 32'h3b354378} /* (14, 21, 26) {real, imag} */,
  {32'h3cb46217, 32'hbde2926d} /* (14, 21, 25) {real, imag} */,
  {32'h3d9206b5, 32'hbcb956c3} /* (14, 21, 24) {real, imag} */,
  {32'hba83c7e0, 32'h3d4db68a} /* (14, 21, 23) {real, imag} */,
  {32'h3c2de2c8, 32'hbd30d216} /* (14, 21, 22) {real, imag} */,
  {32'hbc3fbb4c, 32'h3bea3cc4} /* (14, 21, 21) {real, imag} */,
  {32'hbc35954b, 32'h3e0a888e} /* (14, 21, 20) {real, imag} */,
  {32'h3d0315d6, 32'h3b6a33a8} /* (14, 21, 19) {real, imag} */,
  {32'hbd884641, 32'hbd5e1aac} /* (14, 21, 18) {real, imag} */,
  {32'hbd04071a, 32'h3c7a60d4} /* (14, 21, 17) {real, imag} */,
  {32'hbd2eb2b1, 32'h00000000} /* (14, 21, 16) {real, imag} */,
  {32'hbd04071a, 32'hbc7a60d4} /* (14, 21, 15) {real, imag} */,
  {32'hbd884641, 32'h3d5e1aac} /* (14, 21, 14) {real, imag} */,
  {32'h3d0315d6, 32'hbb6a33a8} /* (14, 21, 13) {real, imag} */,
  {32'hbc35954b, 32'hbe0a888e} /* (14, 21, 12) {real, imag} */,
  {32'hbc3fbb4c, 32'hbbea3cc4} /* (14, 21, 11) {real, imag} */,
  {32'h3c2de2c8, 32'h3d30d216} /* (14, 21, 10) {real, imag} */,
  {32'hba83c7e0, 32'hbd4db68a} /* (14, 21, 9) {real, imag} */,
  {32'h3d9206b5, 32'h3cb956c3} /* (14, 21, 8) {real, imag} */,
  {32'h3cb46217, 32'h3de2926d} /* (14, 21, 7) {real, imag} */,
  {32'hbdcc8c9c, 32'hbb354378} /* (14, 21, 6) {real, imag} */,
  {32'hbe085644, 32'hbdc35fe7} /* (14, 21, 5) {real, imag} */,
  {32'h3dff8134, 32'h3dfdd604} /* (14, 21, 4) {real, imag} */,
  {32'h3dec9d13, 32'h3df0fef9} /* (14, 21, 3) {real, imag} */,
  {32'hbe4af16d, 32'hbe22a25f} /* (14, 21, 2) {real, imag} */,
  {32'h3ec06862, 32'hbda054c0} /* (14, 21, 1) {real, imag} */,
  {32'h3f152456, 32'h00000000} /* (14, 21, 0) {real, imag} */,
  {32'hbf7477ed, 32'h3e674b40} /* (14, 20, 31) {real, imag} */,
  {32'h3eddeb3e, 32'h3c41e300} /* (14, 20, 30) {real, imag} */,
  {32'h3df8d476, 32'hbc020434} /* (14, 20, 29) {real, imag} */,
  {32'hbbf606f0, 32'hbd0ebf04} /* (14, 20, 28) {real, imag} */,
  {32'h3ce55b10, 32'hbe067566} /* (14, 20, 27) {real, imag} */,
  {32'h3d0b2d90, 32'hbdfbf2c5} /* (14, 20, 26) {real, imag} */,
  {32'hbbcd1ad8, 32'hbd18eacf} /* (14, 20, 25) {real, imag} */,
  {32'h3d1cfb38, 32'hbd901da6} /* (14, 20, 24) {real, imag} */,
  {32'hbd9bf326, 32'hbb3492cc} /* (14, 20, 23) {real, imag} */,
  {32'hbdd5bb9f, 32'h3dbc5f00} /* (14, 20, 22) {real, imag} */,
  {32'h3dbb628d, 32'h3d13d66e} /* (14, 20, 21) {real, imag} */,
  {32'h3d987bec, 32'h3d9a16df} /* (14, 20, 20) {real, imag} */,
  {32'hbdaef105, 32'h3d2df589} /* (14, 20, 19) {real, imag} */,
  {32'h3d81b9da, 32'hbde5cf5c} /* (14, 20, 18) {real, imag} */,
  {32'hbc91a1ca, 32'h3d7c0db4} /* (14, 20, 17) {real, imag} */,
  {32'hbd21fee5, 32'h00000000} /* (14, 20, 16) {real, imag} */,
  {32'hbc91a1ca, 32'hbd7c0db4} /* (14, 20, 15) {real, imag} */,
  {32'h3d81b9da, 32'h3de5cf5c} /* (14, 20, 14) {real, imag} */,
  {32'hbdaef105, 32'hbd2df589} /* (14, 20, 13) {real, imag} */,
  {32'h3d987bec, 32'hbd9a16df} /* (14, 20, 12) {real, imag} */,
  {32'h3dbb628d, 32'hbd13d66e} /* (14, 20, 11) {real, imag} */,
  {32'hbdd5bb9f, 32'hbdbc5f00} /* (14, 20, 10) {real, imag} */,
  {32'hbd9bf326, 32'h3b3492cc} /* (14, 20, 9) {real, imag} */,
  {32'h3d1cfb38, 32'h3d901da6} /* (14, 20, 8) {real, imag} */,
  {32'hbbcd1ad8, 32'h3d18eacf} /* (14, 20, 7) {real, imag} */,
  {32'h3d0b2d90, 32'h3dfbf2c5} /* (14, 20, 6) {real, imag} */,
  {32'h3ce55b10, 32'h3e067566} /* (14, 20, 5) {real, imag} */,
  {32'hbbf606f0, 32'h3d0ebf04} /* (14, 20, 4) {real, imag} */,
  {32'h3df8d476, 32'h3c020434} /* (14, 20, 3) {real, imag} */,
  {32'h3eddeb3e, 32'hbc41e300} /* (14, 20, 2) {real, imag} */,
  {32'hbf7477ed, 32'hbe674b40} /* (14, 20, 1) {real, imag} */,
  {32'hbf1197b0, 32'h00000000} /* (14, 20, 0) {real, imag} */,
  {32'hbfc6b476, 32'h3e86b0c7} /* (14, 19, 31) {real, imag} */,
  {32'h3f42fd8a, 32'hbde0645a} /* (14, 19, 30) {real, imag} */,
  {32'h3e62faab, 32'h3c38ac20} /* (14, 19, 29) {real, imag} */,
  {32'hbe171922, 32'h3d9565ef} /* (14, 19, 28) {real, imag} */,
  {32'h3de2d35b, 32'hbe10b76c} /* (14, 19, 27) {real, imag} */,
  {32'hbda60bb6, 32'hbd29b170} /* (14, 19, 26) {real, imag} */,
  {32'hbc8bc170, 32'h3dae58cc} /* (14, 19, 25) {real, imag} */,
  {32'h3dcacbcf, 32'h3d431044} /* (14, 19, 24) {real, imag} */,
  {32'hbcb7b0b2, 32'h3d150708} /* (14, 19, 23) {real, imag} */,
  {32'hbdadfd48, 32'hbd9936a8} /* (14, 19, 22) {real, imag} */,
  {32'h3d017e38, 32'hbda8767b} /* (14, 19, 21) {real, imag} */,
  {32'h3c7eeb72, 32'hbca8eb22} /* (14, 19, 20) {real, imag} */,
  {32'hbd63e32e, 32'h3d96dcc0} /* (14, 19, 19) {real, imag} */,
  {32'hbbeb6e10, 32'h3cf6e2ec} /* (14, 19, 18) {real, imag} */,
  {32'h3c154c40, 32'hbd48dd78} /* (14, 19, 17) {real, imag} */,
  {32'h3b522b00, 32'h00000000} /* (14, 19, 16) {real, imag} */,
  {32'h3c154c40, 32'h3d48dd78} /* (14, 19, 15) {real, imag} */,
  {32'hbbeb6e10, 32'hbcf6e2ec} /* (14, 19, 14) {real, imag} */,
  {32'hbd63e32e, 32'hbd96dcc0} /* (14, 19, 13) {real, imag} */,
  {32'h3c7eeb72, 32'h3ca8eb22} /* (14, 19, 12) {real, imag} */,
  {32'h3d017e38, 32'h3da8767b} /* (14, 19, 11) {real, imag} */,
  {32'hbdadfd48, 32'h3d9936a8} /* (14, 19, 10) {real, imag} */,
  {32'hbcb7b0b2, 32'hbd150708} /* (14, 19, 9) {real, imag} */,
  {32'h3dcacbcf, 32'hbd431044} /* (14, 19, 8) {real, imag} */,
  {32'hbc8bc170, 32'hbdae58cc} /* (14, 19, 7) {real, imag} */,
  {32'hbda60bb6, 32'h3d29b170} /* (14, 19, 6) {real, imag} */,
  {32'h3de2d35b, 32'h3e10b76c} /* (14, 19, 5) {real, imag} */,
  {32'hbe171922, 32'hbd9565ef} /* (14, 19, 4) {real, imag} */,
  {32'h3e62faab, 32'hbc38ac20} /* (14, 19, 3) {real, imag} */,
  {32'h3f42fd8a, 32'h3de0645a} /* (14, 19, 2) {real, imag} */,
  {32'hbfc6b476, 32'hbe86b0c7} /* (14, 19, 1) {real, imag} */,
  {32'hbf75c510, 32'h00000000} /* (14, 19, 0) {real, imag} */,
  {32'hbff6d3dc, 32'h3e921bed} /* (14, 18, 31) {real, imag} */,
  {32'h3f55d7f0, 32'hbe81e218} /* (14, 18, 30) {real, imag} */,
  {32'h3e08cccc, 32'hbd6c5253} /* (14, 18, 29) {real, imag} */,
  {32'hbe11d9f3, 32'h3e025cd5} /* (14, 18, 28) {real, imag} */,
  {32'h3d5e36ee, 32'hbc81602e} /* (14, 18, 27) {real, imag} */,
  {32'hbda35503, 32'hbd07bcee} /* (14, 18, 26) {real, imag} */,
  {32'hbde38beb, 32'h3cf82068} /* (14, 18, 25) {real, imag} */,
  {32'h3d52a9d9, 32'hbd1ca296} /* (14, 18, 24) {real, imag} */,
  {32'hbd08dca2, 32'hbcd338c4} /* (14, 18, 23) {real, imag} */,
  {32'h3c2af075, 32'hbd47f048} /* (14, 18, 22) {real, imag} */,
  {32'hbdcb8484, 32'hbd8aec35} /* (14, 18, 21) {real, imag} */,
  {32'h3d248e3a, 32'hbd6340bd} /* (14, 18, 20) {real, imag} */,
  {32'h3cbdb0ee, 32'hbd0f5cba} /* (14, 18, 19) {real, imag} */,
  {32'h3dc5ff14, 32'hbda2a4d1} /* (14, 18, 18) {real, imag} */,
  {32'h3db14f5d, 32'h3b89d500} /* (14, 18, 17) {real, imag} */,
  {32'h3bff6460, 32'h00000000} /* (14, 18, 16) {real, imag} */,
  {32'h3db14f5d, 32'hbb89d500} /* (14, 18, 15) {real, imag} */,
  {32'h3dc5ff14, 32'h3da2a4d1} /* (14, 18, 14) {real, imag} */,
  {32'h3cbdb0ee, 32'h3d0f5cba} /* (14, 18, 13) {real, imag} */,
  {32'h3d248e3a, 32'h3d6340bd} /* (14, 18, 12) {real, imag} */,
  {32'hbdcb8484, 32'h3d8aec35} /* (14, 18, 11) {real, imag} */,
  {32'h3c2af075, 32'h3d47f048} /* (14, 18, 10) {real, imag} */,
  {32'hbd08dca2, 32'h3cd338c4} /* (14, 18, 9) {real, imag} */,
  {32'h3d52a9d9, 32'h3d1ca296} /* (14, 18, 8) {real, imag} */,
  {32'hbde38beb, 32'hbcf82068} /* (14, 18, 7) {real, imag} */,
  {32'hbda35503, 32'h3d07bcee} /* (14, 18, 6) {real, imag} */,
  {32'h3d5e36ee, 32'h3c81602e} /* (14, 18, 5) {real, imag} */,
  {32'hbe11d9f3, 32'hbe025cd5} /* (14, 18, 4) {real, imag} */,
  {32'h3e08cccc, 32'h3d6c5253} /* (14, 18, 3) {real, imag} */,
  {32'h3f55d7f0, 32'h3e81e218} /* (14, 18, 2) {real, imag} */,
  {32'hbff6d3dc, 32'hbe921bed} /* (14, 18, 1) {real, imag} */,
  {32'hbfa6ce38, 32'h00000000} /* (14, 18, 0) {real, imag} */,
  {32'hc00b6eb6, 32'h3e5a8902} /* (14, 17, 31) {real, imag} */,
  {32'h3f83c118, 32'hbe4f7e2a} /* (14, 17, 30) {real, imag} */,
  {32'h3e11d72d, 32'hbe20246b} /* (14, 17, 29) {real, imag} */,
  {32'hbe18e79c, 32'h3e18d274} /* (14, 17, 28) {real, imag} */,
  {32'h3df69eb2, 32'h3c82c4f5} /* (14, 17, 27) {real, imag} */,
  {32'hbe550d82, 32'hbcfa8060} /* (14, 17, 26) {real, imag} */,
  {32'hbd917e57, 32'hbd651a2a} /* (14, 17, 25) {real, imag} */,
  {32'h3dd880e9, 32'hbddbe528} /* (14, 17, 24) {real, imag} */,
  {32'h3bffdec0, 32'hbcd15d6f} /* (14, 17, 23) {real, imag} */,
  {32'h3d655940, 32'hbd064c16} /* (14, 17, 22) {real, imag} */,
  {32'h3d031f65, 32'hbbc64230} /* (14, 17, 21) {real, imag} */,
  {32'h3cefe528, 32'hbd371ff1} /* (14, 17, 20) {real, imag} */,
  {32'hbd8539d2, 32'hbd54be30} /* (14, 17, 19) {real, imag} */,
  {32'hbcdb872a, 32'hbb6c0aa4} /* (14, 17, 18) {real, imag} */,
  {32'hbc0fb39a, 32'h3d922c44} /* (14, 17, 17) {real, imag} */,
  {32'h3d279b7c, 32'h00000000} /* (14, 17, 16) {real, imag} */,
  {32'hbc0fb39a, 32'hbd922c44} /* (14, 17, 15) {real, imag} */,
  {32'hbcdb872a, 32'h3b6c0aa4} /* (14, 17, 14) {real, imag} */,
  {32'hbd8539d2, 32'h3d54be30} /* (14, 17, 13) {real, imag} */,
  {32'h3cefe528, 32'h3d371ff1} /* (14, 17, 12) {real, imag} */,
  {32'h3d031f65, 32'h3bc64230} /* (14, 17, 11) {real, imag} */,
  {32'h3d655940, 32'h3d064c16} /* (14, 17, 10) {real, imag} */,
  {32'h3bffdec0, 32'h3cd15d6f} /* (14, 17, 9) {real, imag} */,
  {32'h3dd880e9, 32'h3ddbe528} /* (14, 17, 8) {real, imag} */,
  {32'hbd917e57, 32'h3d651a2a} /* (14, 17, 7) {real, imag} */,
  {32'hbe550d82, 32'h3cfa8060} /* (14, 17, 6) {real, imag} */,
  {32'h3df69eb2, 32'hbc82c4f5} /* (14, 17, 5) {real, imag} */,
  {32'hbe18e79c, 32'hbe18d274} /* (14, 17, 4) {real, imag} */,
  {32'h3e11d72d, 32'h3e20246b} /* (14, 17, 3) {real, imag} */,
  {32'h3f83c118, 32'h3e4f7e2a} /* (14, 17, 2) {real, imag} */,
  {32'hc00b6eb6, 32'hbe5a8902} /* (14, 17, 1) {real, imag} */,
  {32'hbfe53322, 32'h00000000} /* (14, 17, 0) {real, imag} */,
  {32'hc01badd4, 32'h3ec0a560} /* (14, 16, 31) {real, imag} */,
  {32'h3f8dfabd, 32'hbe86087f} /* (14, 16, 30) {real, imag} */,
  {32'h3d932dca, 32'hbe2e91c5} /* (14, 16, 29) {real, imag} */,
  {32'hbe1528a2, 32'h3e8e612c} /* (14, 16, 28) {real, imag} */,
  {32'h3e1ce952, 32'hbdae9e2c} /* (14, 16, 27) {real, imag} */,
  {32'h3cda6c7a, 32'hbd891eec} /* (14, 16, 26) {real, imag} */,
  {32'hbd81ebf7, 32'h3c87d08c} /* (14, 16, 25) {real, imag} */,
  {32'h3d859c07, 32'h3d79fd17} /* (14, 16, 24) {real, imag} */,
  {32'h3d464378, 32'hbd13c785} /* (14, 16, 23) {real, imag} */,
  {32'hba51ab38, 32'hbd774f2e} /* (14, 16, 22) {real, imag} */,
  {32'h3da46a18, 32'hbdb8aebc} /* (14, 16, 21) {real, imag} */,
  {32'hbc4049d5, 32'h3dc0102e} /* (14, 16, 20) {real, imag} */,
  {32'hbdb2b8aa, 32'h3d9abefd} /* (14, 16, 19) {real, imag} */,
  {32'h3c05702a, 32'h3ca36260} /* (14, 16, 18) {real, imag} */,
  {32'h3b82c780, 32'h3cac232e} /* (14, 16, 17) {real, imag} */,
  {32'hbc4fa25c, 32'h00000000} /* (14, 16, 16) {real, imag} */,
  {32'h3b82c780, 32'hbcac232e} /* (14, 16, 15) {real, imag} */,
  {32'h3c05702a, 32'hbca36260} /* (14, 16, 14) {real, imag} */,
  {32'hbdb2b8aa, 32'hbd9abefd} /* (14, 16, 13) {real, imag} */,
  {32'hbc4049d5, 32'hbdc0102e} /* (14, 16, 12) {real, imag} */,
  {32'h3da46a18, 32'h3db8aebc} /* (14, 16, 11) {real, imag} */,
  {32'hba51ab38, 32'h3d774f2e} /* (14, 16, 10) {real, imag} */,
  {32'h3d464378, 32'h3d13c785} /* (14, 16, 9) {real, imag} */,
  {32'h3d859c07, 32'hbd79fd17} /* (14, 16, 8) {real, imag} */,
  {32'hbd81ebf7, 32'hbc87d08c} /* (14, 16, 7) {real, imag} */,
  {32'h3cda6c7a, 32'h3d891eec} /* (14, 16, 6) {real, imag} */,
  {32'h3e1ce952, 32'h3dae9e2c} /* (14, 16, 5) {real, imag} */,
  {32'hbe1528a2, 32'hbe8e612c} /* (14, 16, 4) {real, imag} */,
  {32'h3d932dca, 32'h3e2e91c5} /* (14, 16, 3) {real, imag} */,
  {32'h3f8dfabd, 32'h3e86087f} /* (14, 16, 2) {real, imag} */,
  {32'hc01badd4, 32'hbec0a560} /* (14, 16, 1) {real, imag} */,
  {32'hbfdb99c9, 32'h00000000} /* (14, 16, 0) {real, imag} */,
  {32'hc0249cee, 32'h3ef758f3} /* (14, 15, 31) {real, imag} */,
  {32'h3f87af84, 32'hbe697dae} /* (14, 15, 30) {real, imag} */,
  {32'h3d9035da, 32'hbdbffce6} /* (14, 15, 29) {real, imag} */,
  {32'hbe0995f8, 32'h3e935d28} /* (14, 15, 28) {real, imag} */,
  {32'h3d8f1cb2, 32'hbd70318c} /* (14, 15, 27) {real, imag} */,
  {32'h3cb87100, 32'hbe89f6be} /* (14, 15, 26) {real, imag} */,
  {32'hbd98e41f, 32'h3d344c92} /* (14, 15, 25) {real, imag} */,
  {32'h3e4997a4, 32'hbcec7738} /* (14, 15, 24) {real, imag} */,
  {32'h3e027f5b, 32'hbd2e7e80} /* (14, 15, 23) {real, imag} */,
  {32'hbd8b8535, 32'hbd406f12} /* (14, 15, 22) {real, imag} */,
  {32'hbda69dc0, 32'h3d934561} /* (14, 15, 21) {real, imag} */,
  {32'h3d256170, 32'h3d888ca2} /* (14, 15, 20) {real, imag} */,
  {32'hbde5e440, 32'hbde8195c} /* (14, 15, 19) {real, imag} */,
  {32'hbd1a1b0f, 32'hbc50d3e9} /* (14, 15, 18) {real, imag} */,
  {32'hbd2b7dfa, 32'h3cb793a8} /* (14, 15, 17) {real, imag} */,
  {32'hbd0ec7dc, 32'h00000000} /* (14, 15, 16) {real, imag} */,
  {32'hbd2b7dfa, 32'hbcb793a8} /* (14, 15, 15) {real, imag} */,
  {32'hbd1a1b0f, 32'h3c50d3e9} /* (14, 15, 14) {real, imag} */,
  {32'hbde5e440, 32'h3de8195c} /* (14, 15, 13) {real, imag} */,
  {32'h3d256170, 32'hbd888ca2} /* (14, 15, 12) {real, imag} */,
  {32'hbda69dc0, 32'hbd934561} /* (14, 15, 11) {real, imag} */,
  {32'hbd8b8535, 32'h3d406f12} /* (14, 15, 10) {real, imag} */,
  {32'h3e027f5b, 32'h3d2e7e80} /* (14, 15, 9) {real, imag} */,
  {32'h3e4997a4, 32'h3cec7738} /* (14, 15, 8) {real, imag} */,
  {32'hbd98e41f, 32'hbd344c92} /* (14, 15, 7) {real, imag} */,
  {32'h3cb87100, 32'h3e89f6be} /* (14, 15, 6) {real, imag} */,
  {32'h3d8f1cb2, 32'h3d70318c} /* (14, 15, 5) {real, imag} */,
  {32'hbe0995f8, 32'hbe935d28} /* (14, 15, 4) {real, imag} */,
  {32'h3d9035da, 32'h3dbffce6} /* (14, 15, 3) {real, imag} */,
  {32'h3f87af84, 32'h3e697dae} /* (14, 15, 2) {real, imag} */,
  {32'hc0249cee, 32'hbef758f3} /* (14, 15, 1) {real, imag} */,
  {32'hbfed1ec4, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'hc020b3cc, 32'h3ec886ff} /* (14, 14, 31) {real, imag} */,
  {32'h3f57b00e, 32'hbe356b77} /* (14, 14, 30) {real, imag} */,
  {32'h3d71a97e, 32'h3cd29922} /* (14, 14, 29) {real, imag} */,
  {32'hbbcdde60, 32'h3e3aa18f} /* (14, 14, 28) {real, imag} */,
  {32'h3e1b1020, 32'hbdc0ebbc} /* (14, 14, 27) {real, imag} */,
  {32'h3cfac247, 32'hbdd02ab9} /* (14, 14, 26) {real, imag} */,
  {32'hbdbad88d, 32'hbc99b2d8} /* (14, 14, 25) {real, imag} */,
  {32'h3dfe50d2, 32'h3c8430eb} /* (14, 14, 24) {real, imag} */,
  {32'h3c62be36, 32'h3942c400} /* (14, 14, 23) {real, imag} */,
  {32'hbccbb10a, 32'h3bc77564} /* (14, 14, 22) {real, imag} */,
  {32'hbc271d64, 32'hbdc32775} /* (14, 14, 21) {real, imag} */,
  {32'h3c25e482, 32'hbcf95e42} /* (14, 14, 20) {real, imag} */,
  {32'hbc08cbdc, 32'h3d2e9206} /* (14, 14, 19) {real, imag} */,
  {32'h3c1d4fcc, 32'hbc05bab8} /* (14, 14, 18) {real, imag} */,
  {32'h3d7addde, 32'h3d8ec286} /* (14, 14, 17) {real, imag} */,
  {32'h3c82cd1e, 32'h00000000} /* (14, 14, 16) {real, imag} */,
  {32'h3d7addde, 32'hbd8ec286} /* (14, 14, 15) {real, imag} */,
  {32'h3c1d4fcc, 32'h3c05bab8} /* (14, 14, 14) {real, imag} */,
  {32'hbc08cbdc, 32'hbd2e9206} /* (14, 14, 13) {real, imag} */,
  {32'h3c25e482, 32'h3cf95e42} /* (14, 14, 12) {real, imag} */,
  {32'hbc271d64, 32'h3dc32775} /* (14, 14, 11) {real, imag} */,
  {32'hbccbb10a, 32'hbbc77564} /* (14, 14, 10) {real, imag} */,
  {32'h3c62be36, 32'hb942c400} /* (14, 14, 9) {real, imag} */,
  {32'h3dfe50d2, 32'hbc8430eb} /* (14, 14, 8) {real, imag} */,
  {32'hbdbad88d, 32'h3c99b2d8} /* (14, 14, 7) {real, imag} */,
  {32'h3cfac247, 32'h3dd02ab9} /* (14, 14, 6) {real, imag} */,
  {32'h3e1b1020, 32'h3dc0ebbc} /* (14, 14, 5) {real, imag} */,
  {32'hbbcdde60, 32'hbe3aa18f} /* (14, 14, 4) {real, imag} */,
  {32'h3d71a97e, 32'hbcd29922} /* (14, 14, 3) {real, imag} */,
  {32'h3f57b00e, 32'h3e356b77} /* (14, 14, 2) {real, imag} */,
  {32'hc020b3cc, 32'hbec886ff} /* (14, 14, 1) {real, imag} */,
  {32'hbfc9ba90, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'hc00c7100, 32'h3e56be92} /* (14, 13, 31) {real, imag} */,
  {32'h3f393126, 32'hbdaf20d6} /* (14, 13, 30) {real, imag} */,
  {32'h3decfbd2, 32'h3d36ec18} /* (14, 13, 29) {real, imag} */,
  {32'hbdf5cd9f, 32'h3e497a28} /* (14, 13, 28) {real, imag} */,
  {32'h3ddca137, 32'hbe1f0dc0} /* (14, 13, 27) {real, imag} */,
  {32'h3d466eb3, 32'hbd9e0a90} /* (14, 13, 26) {real, imag} */,
  {32'hbc0f6bb8, 32'h3c28ae5c} /* (14, 13, 25) {real, imag} */,
  {32'h3d8f7371, 32'h3ce0f2dd} /* (14, 13, 24) {real, imag} */,
  {32'hbd0f4eef, 32'h3d9d5259} /* (14, 13, 23) {real, imag} */,
  {32'h3d3c330f, 32'h3bf6a368} /* (14, 13, 22) {real, imag} */,
  {32'h3d501ad6, 32'hbe1ebb0e} /* (14, 13, 21) {real, imag} */,
  {32'hbd651ea2, 32'hbdb359aa} /* (14, 13, 20) {real, imag} */,
  {32'h3cb0012b, 32'hbcb048c2} /* (14, 13, 19) {real, imag} */,
  {32'hbd1d72f4, 32'hbda9aca4} /* (14, 13, 18) {real, imag} */,
  {32'hbc3777b0, 32'h3b2ee158} /* (14, 13, 17) {real, imag} */,
  {32'h3d1cd716, 32'h00000000} /* (14, 13, 16) {real, imag} */,
  {32'hbc3777b0, 32'hbb2ee158} /* (14, 13, 15) {real, imag} */,
  {32'hbd1d72f4, 32'h3da9aca4} /* (14, 13, 14) {real, imag} */,
  {32'h3cb0012b, 32'h3cb048c2} /* (14, 13, 13) {real, imag} */,
  {32'hbd651ea2, 32'h3db359aa} /* (14, 13, 12) {real, imag} */,
  {32'h3d501ad6, 32'h3e1ebb0e} /* (14, 13, 11) {real, imag} */,
  {32'h3d3c330f, 32'hbbf6a368} /* (14, 13, 10) {real, imag} */,
  {32'hbd0f4eef, 32'hbd9d5259} /* (14, 13, 9) {real, imag} */,
  {32'h3d8f7371, 32'hbce0f2dd} /* (14, 13, 8) {real, imag} */,
  {32'hbc0f6bb8, 32'hbc28ae5c} /* (14, 13, 7) {real, imag} */,
  {32'h3d466eb3, 32'h3d9e0a90} /* (14, 13, 6) {real, imag} */,
  {32'h3ddca137, 32'h3e1f0dc0} /* (14, 13, 5) {real, imag} */,
  {32'hbdf5cd9f, 32'hbe497a28} /* (14, 13, 4) {real, imag} */,
  {32'h3decfbd2, 32'hbd36ec18} /* (14, 13, 3) {real, imag} */,
  {32'h3f393126, 32'h3daf20d6} /* (14, 13, 2) {real, imag} */,
  {32'hc00c7100, 32'hbe56be92} /* (14, 13, 1) {real, imag} */,
  {32'hbf8fc6f2, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'hbfe09d72, 32'h3e5ab408} /* (14, 12, 31) {real, imag} */,
  {32'h3f1d5295, 32'hbb8f8c40} /* (14, 12, 30) {real, imag} */,
  {32'h3d0fff30, 32'hbba3fe78} /* (14, 12, 29) {real, imag} */,
  {32'hbe368df8, 32'h3e5ded6f} /* (14, 12, 28) {real, imag} */,
  {32'h3e6b0b42, 32'hbe34201e} /* (14, 12, 27) {real, imag} */,
  {32'h3d3ff080, 32'hbb7647a0} /* (14, 12, 26) {real, imag} */,
  {32'h3db62d54, 32'hbd827786} /* (14, 12, 25) {real, imag} */,
  {32'h3d9b0696, 32'hbc2b286c} /* (14, 12, 24) {real, imag} */,
  {32'hbb3fa6f0, 32'h3cb25f66} /* (14, 12, 23) {real, imag} */,
  {32'h3c300410, 32'hbd4c06d3} /* (14, 12, 22) {real, imag} */,
  {32'h3d6293a6, 32'hbd96cd13} /* (14, 12, 21) {real, imag} */,
  {32'hbc9e270a, 32'hbd752baa} /* (14, 12, 20) {real, imag} */,
  {32'h3d3b815e, 32'h3d06b4af} /* (14, 12, 19) {real, imag} */,
  {32'h3cf64df0, 32'h3b96a140} /* (14, 12, 18) {real, imag} */,
  {32'h3cb43c5a, 32'hbd626c14} /* (14, 12, 17) {real, imag} */,
  {32'hbdb13818, 32'h00000000} /* (14, 12, 16) {real, imag} */,
  {32'h3cb43c5a, 32'h3d626c14} /* (14, 12, 15) {real, imag} */,
  {32'h3cf64df0, 32'hbb96a140} /* (14, 12, 14) {real, imag} */,
  {32'h3d3b815e, 32'hbd06b4af} /* (14, 12, 13) {real, imag} */,
  {32'hbc9e270a, 32'h3d752baa} /* (14, 12, 12) {real, imag} */,
  {32'h3d6293a6, 32'h3d96cd13} /* (14, 12, 11) {real, imag} */,
  {32'h3c300410, 32'h3d4c06d3} /* (14, 12, 10) {real, imag} */,
  {32'hbb3fa6f0, 32'hbcb25f66} /* (14, 12, 9) {real, imag} */,
  {32'h3d9b0696, 32'h3c2b286c} /* (14, 12, 8) {real, imag} */,
  {32'h3db62d54, 32'h3d827786} /* (14, 12, 7) {real, imag} */,
  {32'h3d3ff080, 32'h3b7647a0} /* (14, 12, 6) {real, imag} */,
  {32'h3e6b0b42, 32'h3e34201e} /* (14, 12, 5) {real, imag} */,
  {32'hbe368df8, 32'hbe5ded6f} /* (14, 12, 4) {real, imag} */,
  {32'h3d0fff30, 32'h3ba3fe78} /* (14, 12, 3) {real, imag} */,
  {32'h3f1d5295, 32'h3b8f8c40} /* (14, 12, 2) {real, imag} */,
  {32'hbfe09d72, 32'hbe5ab408} /* (14, 12, 1) {real, imag} */,
  {32'hbf14aa94, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'hbf6d4421, 32'h3dfaf5f0} /* (14, 11, 31) {real, imag} */,
  {32'h3f0dd2ef, 32'h3da52262} /* (14, 11, 30) {real, imag} */,
  {32'h3d4b0bda, 32'h3d626dce} /* (14, 11, 29) {real, imag} */,
  {32'hbd857418, 32'h3daf0d4a} /* (14, 11, 28) {real, imag} */,
  {32'h3dd2d22f, 32'hbe1f544c} /* (14, 11, 27) {real, imag} */,
  {32'h3d9a83ac, 32'h3ce74e43} /* (14, 11, 26) {real, imag} */,
  {32'hbd8b99bd, 32'hbddac313} /* (14, 11, 25) {real, imag} */,
  {32'h3d3fcbde, 32'hbcf83e0f} /* (14, 11, 24) {real, imag} */,
  {32'hbdedfb2e, 32'hbdd7caaf} /* (14, 11, 23) {real, imag} */,
  {32'hbdc22a4a, 32'hbd35f358} /* (14, 11, 22) {real, imag} */,
  {32'hbd9dc13e, 32'hbd11af48} /* (14, 11, 21) {real, imag} */,
  {32'hbb0b293c, 32'h3e29155c} /* (14, 11, 20) {real, imag} */,
  {32'h3de1ed59, 32'h3d223fa0} /* (14, 11, 19) {real, imag} */,
  {32'h3d7ad0ca, 32'h3c31c800} /* (14, 11, 18) {real, imag} */,
  {32'h3d5e0d28, 32'h3b397cc0} /* (14, 11, 17) {real, imag} */,
  {32'hbcb6b172, 32'h00000000} /* (14, 11, 16) {real, imag} */,
  {32'h3d5e0d28, 32'hbb397cc0} /* (14, 11, 15) {real, imag} */,
  {32'h3d7ad0ca, 32'hbc31c800} /* (14, 11, 14) {real, imag} */,
  {32'h3de1ed59, 32'hbd223fa0} /* (14, 11, 13) {real, imag} */,
  {32'hbb0b293c, 32'hbe29155c} /* (14, 11, 12) {real, imag} */,
  {32'hbd9dc13e, 32'h3d11af48} /* (14, 11, 11) {real, imag} */,
  {32'hbdc22a4a, 32'h3d35f358} /* (14, 11, 10) {real, imag} */,
  {32'hbdedfb2e, 32'h3dd7caaf} /* (14, 11, 9) {real, imag} */,
  {32'h3d3fcbde, 32'h3cf83e0f} /* (14, 11, 8) {real, imag} */,
  {32'hbd8b99bd, 32'h3ddac313} /* (14, 11, 7) {real, imag} */,
  {32'h3d9a83ac, 32'hbce74e43} /* (14, 11, 6) {real, imag} */,
  {32'h3dd2d22f, 32'h3e1f544c} /* (14, 11, 5) {real, imag} */,
  {32'hbd857418, 32'hbdaf0d4a} /* (14, 11, 4) {real, imag} */,
  {32'h3d4b0bda, 32'hbd626dce} /* (14, 11, 3) {real, imag} */,
  {32'h3f0dd2ef, 32'hbda52262} /* (14, 11, 2) {real, imag} */,
  {32'hbf6d4421, 32'hbdfaf5f0} /* (14, 11, 1) {real, imag} */,
  {32'h3b0f9e00, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h3f03599a, 32'hbe7ad559} /* (14, 10, 31) {real, imag} */,
  {32'h3d8a6928, 32'h3dee1b4c} /* (14, 10, 30) {real, imag} */,
  {32'h3d1ef388, 32'h3d665443} /* (14, 10, 29) {real, imag} */,
  {32'hbd3a6c80, 32'hbbc2a070} /* (14, 10, 28) {real, imag} */,
  {32'hbe47ac70, 32'h3d73c50b} /* (14, 10, 27) {real, imag} */,
  {32'hbd2420fc, 32'h3d893e8c} /* (14, 10, 26) {real, imag} */,
  {32'hbdafe03b, 32'h3cf93aed} /* (14, 10, 25) {real, imag} */,
  {32'h3ccc75af, 32'h3d0df6d0} /* (14, 10, 24) {real, imag} */,
  {32'h3c1a8ba0, 32'h3df26aba} /* (14, 10, 23) {real, imag} */,
  {32'h3ce793e2, 32'hbc343a3c} /* (14, 10, 22) {real, imag} */,
  {32'h3beaf9f0, 32'hbd901522} /* (14, 10, 21) {real, imag} */,
  {32'h3d6a1244, 32'hbd01fbac} /* (14, 10, 20) {real, imag} */,
  {32'hbc7845fa, 32'hbdfcaa9d} /* (14, 10, 19) {real, imag} */,
  {32'hbdf70479, 32'hbcd6fa10} /* (14, 10, 18) {real, imag} */,
  {32'hbdd7a252, 32'hbd3f3dc0} /* (14, 10, 17) {real, imag} */,
  {32'hbc8e3884, 32'h00000000} /* (14, 10, 16) {real, imag} */,
  {32'hbdd7a252, 32'h3d3f3dc0} /* (14, 10, 15) {real, imag} */,
  {32'hbdf70479, 32'h3cd6fa10} /* (14, 10, 14) {real, imag} */,
  {32'hbc7845fa, 32'h3dfcaa9d} /* (14, 10, 13) {real, imag} */,
  {32'h3d6a1244, 32'h3d01fbac} /* (14, 10, 12) {real, imag} */,
  {32'h3beaf9f0, 32'h3d901522} /* (14, 10, 11) {real, imag} */,
  {32'h3ce793e2, 32'h3c343a3c} /* (14, 10, 10) {real, imag} */,
  {32'h3c1a8ba0, 32'hbdf26aba} /* (14, 10, 9) {real, imag} */,
  {32'h3ccc75af, 32'hbd0df6d0} /* (14, 10, 8) {real, imag} */,
  {32'hbdafe03b, 32'hbcf93aed} /* (14, 10, 7) {real, imag} */,
  {32'hbd2420fc, 32'hbd893e8c} /* (14, 10, 6) {real, imag} */,
  {32'hbe47ac70, 32'hbd73c50b} /* (14, 10, 5) {real, imag} */,
  {32'hbd3a6c80, 32'h3bc2a070} /* (14, 10, 4) {real, imag} */,
  {32'h3d1ef388, 32'hbd665443} /* (14, 10, 3) {real, imag} */,
  {32'h3d8a6928, 32'hbdee1b4c} /* (14, 10, 2) {real, imag} */,
  {32'h3f03599a, 32'h3e7ad559} /* (14, 10, 1) {real, imag} */,
  {32'h3f7a318d, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'h3f9e886a, 32'hbee28374} /* (14, 9, 31) {real, imag} */,
  {32'hbef0dde2, 32'h3e49d9ac} /* (14, 9, 30) {real, imag} */,
  {32'hbcafbbfa, 32'h3e21b840} /* (14, 9, 29) {real, imag} */,
  {32'hbd0afe17, 32'hbb7f2720} /* (14, 9, 28) {real, imag} */,
  {32'hbe372b78, 32'h3e71d200} /* (14, 9, 27) {real, imag} */,
  {32'h3d8a7a96, 32'hbcbdea17} /* (14, 9, 26) {real, imag} */,
  {32'hbdea040f, 32'hbbebb558} /* (14, 9, 25) {real, imag} */,
  {32'h3c9a98d6, 32'h3de55cfa} /* (14, 9, 24) {real, imag} */,
  {32'hbab7df40, 32'h3cbecc8a} /* (14, 9, 23) {real, imag} */,
  {32'h3c9865b4, 32'h3d93d302} /* (14, 9, 22) {real, imag} */,
  {32'hbc9b3667, 32'h3dae5b31} /* (14, 9, 21) {real, imag} */,
  {32'h3defff5a, 32'hbd4f89c3} /* (14, 9, 20) {real, imag} */,
  {32'hbcd3a997, 32'hbd886278} /* (14, 9, 19) {real, imag} */,
  {32'hbcd4cf1e, 32'h3db0bfff} /* (14, 9, 18) {real, imag} */,
  {32'h3d8ca143, 32'hbd57fc94} /* (14, 9, 17) {real, imag} */,
  {32'h3ceb7177, 32'h00000000} /* (14, 9, 16) {real, imag} */,
  {32'h3d8ca143, 32'h3d57fc94} /* (14, 9, 15) {real, imag} */,
  {32'hbcd4cf1e, 32'hbdb0bfff} /* (14, 9, 14) {real, imag} */,
  {32'hbcd3a997, 32'h3d886278} /* (14, 9, 13) {real, imag} */,
  {32'h3defff5a, 32'h3d4f89c3} /* (14, 9, 12) {real, imag} */,
  {32'hbc9b3667, 32'hbdae5b31} /* (14, 9, 11) {real, imag} */,
  {32'h3c9865b4, 32'hbd93d302} /* (14, 9, 10) {real, imag} */,
  {32'hbab7df40, 32'hbcbecc8a} /* (14, 9, 9) {real, imag} */,
  {32'h3c9a98d6, 32'hbde55cfa} /* (14, 9, 8) {real, imag} */,
  {32'hbdea040f, 32'h3bebb558} /* (14, 9, 7) {real, imag} */,
  {32'h3d8a7a96, 32'h3cbdea17} /* (14, 9, 6) {real, imag} */,
  {32'hbe372b78, 32'hbe71d200} /* (14, 9, 5) {real, imag} */,
  {32'hbd0afe17, 32'h3b7f2720} /* (14, 9, 4) {real, imag} */,
  {32'hbcafbbfa, 32'hbe21b840} /* (14, 9, 3) {real, imag} */,
  {32'hbef0dde2, 32'hbe49d9ac} /* (14, 9, 2) {real, imag} */,
  {32'h3f9e886a, 32'h3ee28374} /* (14, 9, 1) {real, imag} */,
  {32'h3fdb576a, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'h3fc06eed, 32'hbf08687f} /* (14, 8, 31) {real, imag} */,
  {32'hbf2836ce, 32'h3ec824d8} /* (14, 8, 30) {real, imag} */,
  {32'hbd32e6fd, 32'h3dfede0a} /* (14, 8, 29) {real, imag} */,
  {32'h3e0faa86, 32'hbd7f856b} /* (14, 8, 28) {real, imag} */,
  {32'hbdabe6b2, 32'h3bb39e60} /* (14, 8, 27) {real, imag} */,
  {32'h3c5966e8, 32'h3de50d74} /* (14, 8, 26) {real, imag} */,
  {32'hbd5734cc, 32'h3dc0bca1} /* (14, 8, 25) {real, imag} */,
  {32'hbdaf2586, 32'h3dd209e0} /* (14, 8, 24) {real, imag} */,
  {32'hbd8abefe, 32'hbd6f2a16} /* (14, 8, 23) {real, imag} */,
  {32'hbd4d49ce, 32'hbdb2ff1a} /* (14, 8, 22) {real, imag} */,
  {32'hbd4a0bce, 32'hbccf3890} /* (14, 8, 21) {real, imag} */,
  {32'hbd4dcb82, 32'h3c995ce4} /* (14, 8, 20) {real, imag} */,
  {32'h3d8d5b78, 32'hbcd6a109} /* (14, 8, 19) {real, imag} */,
  {32'hbd662a72, 32'h3d9bf8b8} /* (14, 8, 18) {real, imag} */,
  {32'hbdae477e, 32'h3dd6a18a} /* (14, 8, 17) {real, imag} */,
  {32'h3bdac844, 32'h00000000} /* (14, 8, 16) {real, imag} */,
  {32'hbdae477e, 32'hbdd6a18a} /* (14, 8, 15) {real, imag} */,
  {32'hbd662a72, 32'hbd9bf8b8} /* (14, 8, 14) {real, imag} */,
  {32'h3d8d5b78, 32'h3cd6a109} /* (14, 8, 13) {real, imag} */,
  {32'hbd4dcb82, 32'hbc995ce4} /* (14, 8, 12) {real, imag} */,
  {32'hbd4a0bce, 32'h3ccf3890} /* (14, 8, 11) {real, imag} */,
  {32'hbd4d49ce, 32'h3db2ff1a} /* (14, 8, 10) {real, imag} */,
  {32'hbd8abefe, 32'h3d6f2a16} /* (14, 8, 9) {real, imag} */,
  {32'hbdaf2586, 32'hbdd209e0} /* (14, 8, 8) {real, imag} */,
  {32'hbd5734cc, 32'hbdc0bca1} /* (14, 8, 7) {real, imag} */,
  {32'h3c5966e8, 32'hbde50d74} /* (14, 8, 6) {real, imag} */,
  {32'hbdabe6b2, 32'hbbb39e60} /* (14, 8, 5) {real, imag} */,
  {32'h3e0faa86, 32'h3d7f856b} /* (14, 8, 4) {real, imag} */,
  {32'hbd32e6fd, 32'hbdfede0a} /* (14, 8, 3) {real, imag} */,
  {32'hbf2836ce, 32'hbec824d8} /* (14, 8, 2) {real, imag} */,
  {32'h3fc06eed, 32'h3f08687f} /* (14, 8, 1) {real, imag} */,
  {32'h40025d86, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'h3fdac22e, 32'hbf2ce0dc} /* (14, 7, 31) {real, imag} */,
  {32'hbf3d8a21, 32'h3ed09a10} /* (14, 7, 30) {real, imag} */,
  {32'hbd7d79b9, 32'h3d7bc146} /* (14, 7, 29) {real, imag} */,
  {32'h3e1e7320, 32'hbda33d59} /* (14, 7, 28) {real, imag} */,
  {32'hbdf87f3b, 32'h3cc52d24} /* (14, 7, 27) {real, imag} */,
  {32'h3d4ca9ca, 32'h3dc65d18} /* (14, 7, 26) {real, imag} */,
  {32'hbd308158, 32'h3c160ef8} /* (14, 7, 25) {real, imag} */,
  {32'hbdef662a, 32'hbce13010} /* (14, 7, 24) {real, imag} */,
  {32'hbcc20a0c, 32'h3d84587a} /* (14, 7, 23) {real, imag} */,
  {32'h3d33457d, 32'hbdd10b04} /* (14, 7, 22) {real, imag} */,
  {32'hbd9feb72, 32'h3cba1fb4} /* (14, 7, 21) {real, imag} */,
  {32'h3cec90a1, 32'hbd1e08d2} /* (14, 7, 20) {real, imag} */,
  {32'h3d432c82, 32'hbd92cdee} /* (14, 7, 19) {real, imag} */,
  {32'hbc9034ce, 32'h3da9f644} /* (14, 7, 18) {real, imag} */,
  {32'h3c185129, 32'h3d1ec9e6} /* (14, 7, 17) {real, imag} */,
  {32'h3dc48baa, 32'h00000000} /* (14, 7, 16) {real, imag} */,
  {32'h3c185129, 32'hbd1ec9e6} /* (14, 7, 15) {real, imag} */,
  {32'hbc9034ce, 32'hbda9f644} /* (14, 7, 14) {real, imag} */,
  {32'h3d432c82, 32'h3d92cdee} /* (14, 7, 13) {real, imag} */,
  {32'h3cec90a1, 32'h3d1e08d2} /* (14, 7, 12) {real, imag} */,
  {32'hbd9feb72, 32'hbcba1fb4} /* (14, 7, 11) {real, imag} */,
  {32'h3d33457d, 32'h3dd10b04} /* (14, 7, 10) {real, imag} */,
  {32'hbcc20a0c, 32'hbd84587a} /* (14, 7, 9) {real, imag} */,
  {32'hbdef662a, 32'h3ce13010} /* (14, 7, 8) {real, imag} */,
  {32'hbd308158, 32'hbc160ef8} /* (14, 7, 7) {real, imag} */,
  {32'h3d4ca9ca, 32'hbdc65d18} /* (14, 7, 6) {real, imag} */,
  {32'hbdf87f3b, 32'hbcc52d24} /* (14, 7, 5) {real, imag} */,
  {32'h3e1e7320, 32'h3da33d59} /* (14, 7, 4) {real, imag} */,
  {32'hbd7d79b9, 32'hbd7bc146} /* (14, 7, 3) {real, imag} */,
  {32'hbf3d8a21, 32'hbed09a10} /* (14, 7, 2) {real, imag} */,
  {32'h3fdac22e, 32'h3f2ce0dc} /* (14, 7, 1) {real, imag} */,
  {32'h401048ba, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'h3feda8a1, 32'hbf7e9606} /* (14, 6, 31) {real, imag} */,
  {32'hbf211a33, 32'h3f0561f6} /* (14, 6, 30) {real, imag} */,
  {32'hbde5971d, 32'h3ddfb66a} /* (14, 6, 29) {real, imag} */,
  {32'h3ddf21a4, 32'h3bf10030} /* (14, 6, 28) {real, imag} */,
  {32'hbe298158, 32'h3e2bdf27} /* (14, 6, 27) {real, imag} */,
  {32'h3db020ac, 32'h3c460510} /* (14, 6, 26) {real, imag} */,
  {32'h3d4da6f0, 32'hbe09a9f4} /* (14, 6, 25) {real, imag} */,
  {32'h3c7e1684, 32'h3c398c02} /* (14, 6, 24) {real, imag} */,
  {32'hbaa09f80, 32'h3dda7bcd} /* (14, 6, 23) {real, imag} */,
  {32'h3d9e5e76, 32'h3d543b9c} /* (14, 6, 22) {real, imag} */,
  {32'hbcb83994, 32'h3de6096f} /* (14, 6, 21) {real, imag} */,
  {32'h3cb1b446, 32'h3d5f9f6c} /* (14, 6, 20) {real, imag} */,
  {32'hbdb2b89d, 32'h3c6b60be} /* (14, 6, 19) {real, imag} */,
  {32'hbd4181c4, 32'hbd161255} /* (14, 6, 18) {real, imag} */,
  {32'hbd52aace, 32'hbd9db1f6} /* (14, 6, 17) {real, imag} */,
  {32'hbd8a7e99, 32'h00000000} /* (14, 6, 16) {real, imag} */,
  {32'hbd52aace, 32'h3d9db1f6} /* (14, 6, 15) {real, imag} */,
  {32'hbd4181c4, 32'h3d161255} /* (14, 6, 14) {real, imag} */,
  {32'hbdb2b89d, 32'hbc6b60be} /* (14, 6, 13) {real, imag} */,
  {32'h3cb1b446, 32'hbd5f9f6c} /* (14, 6, 12) {real, imag} */,
  {32'hbcb83994, 32'hbde6096f} /* (14, 6, 11) {real, imag} */,
  {32'h3d9e5e76, 32'hbd543b9c} /* (14, 6, 10) {real, imag} */,
  {32'hbaa09f80, 32'hbdda7bcd} /* (14, 6, 9) {real, imag} */,
  {32'h3c7e1684, 32'hbc398c02} /* (14, 6, 8) {real, imag} */,
  {32'h3d4da6f0, 32'h3e09a9f4} /* (14, 6, 7) {real, imag} */,
  {32'h3db020ac, 32'hbc460510} /* (14, 6, 6) {real, imag} */,
  {32'hbe298158, 32'hbe2bdf27} /* (14, 6, 5) {real, imag} */,
  {32'h3ddf21a4, 32'hbbf10030} /* (14, 6, 4) {real, imag} */,
  {32'hbde5971d, 32'hbddfb66a} /* (14, 6, 3) {real, imag} */,
  {32'hbf211a33, 32'hbf0561f6} /* (14, 6, 2) {real, imag} */,
  {32'h3feda8a1, 32'h3f7e9606} /* (14, 6, 1) {real, imag} */,
  {32'h401cdc75, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h3fdfb27e, 32'hbfd1b090} /* (14, 5, 31) {real, imag} */,
  {32'hbe479b68, 32'h3f28d9a4} /* (14, 5, 30) {real, imag} */,
  {32'hbdb9cbd8, 32'h3e11dee0} /* (14, 5, 29) {real, imag} */,
  {32'hbe1009a2, 32'hbc01b930} /* (14, 5, 28) {real, imag} */,
  {32'hbe428f38, 32'h3d1708a6} /* (14, 5, 27) {real, imag} */,
  {32'h3dc2df88, 32'h3de4e47c} /* (14, 5, 26) {real, imag} */,
  {32'hbdc38458, 32'hbd5046ca} /* (14, 5, 25) {real, imag} */,
  {32'h3d6b4070, 32'hbc52bf00} /* (14, 5, 24) {real, imag} */,
  {32'hbd705a16, 32'hbd186c1c} /* (14, 5, 23) {real, imag} */,
  {32'hbbc94938, 32'hbd7b4933} /* (14, 5, 22) {real, imag} */,
  {32'hbcae2e09, 32'h3d0d2f50} /* (14, 5, 21) {real, imag} */,
  {32'h3d969e64, 32'h3b47c7e8} /* (14, 5, 20) {real, imag} */,
  {32'h3cccb077, 32'h3bf2613c} /* (14, 5, 19) {real, imag} */,
  {32'hbc72ceb8, 32'h3c9e443c} /* (14, 5, 18) {real, imag} */,
  {32'h3c4d447c, 32'h3d8c892f} /* (14, 5, 17) {real, imag} */,
  {32'h3d2b1444, 32'h00000000} /* (14, 5, 16) {real, imag} */,
  {32'h3c4d447c, 32'hbd8c892f} /* (14, 5, 15) {real, imag} */,
  {32'hbc72ceb8, 32'hbc9e443c} /* (14, 5, 14) {real, imag} */,
  {32'h3cccb077, 32'hbbf2613c} /* (14, 5, 13) {real, imag} */,
  {32'h3d969e64, 32'hbb47c7e8} /* (14, 5, 12) {real, imag} */,
  {32'hbcae2e09, 32'hbd0d2f50} /* (14, 5, 11) {real, imag} */,
  {32'hbbc94938, 32'h3d7b4933} /* (14, 5, 10) {real, imag} */,
  {32'hbd705a16, 32'h3d186c1c} /* (14, 5, 9) {real, imag} */,
  {32'h3d6b4070, 32'h3c52bf00} /* (14, 5, 8) {real, imag} */,
  {32'hbdc38458, 32'h3d5046ca} /* (14, 5, 7) {real, imag} */,
  {32'h3dc2df88, 32'hbde4e47c} /* (14, 5, 6) {real, imag} */,
  {32'hbe428f38, 32'hbd1708a6} /* (14, 5, 5) {real, imag} */,
  {32'hbe1009a2, 32'h3c01b930} /* (14, 5, 4) {real, imag} */,
  {32'hbdb9cbd8, 32'hbe11dee0} /* (14, 5, 3) {real, imag} */,
  {32'hbe479b68, 32'hbf28d9a4} /* (14, 5, 2) {real, imag} */,
  {32'h3fdfb27e, 32'h3fd1b090} /* (14, 5, 1) {real, imag} */,
  {32'h401d2969, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'h3fc8f5de, 32'hc0040571} /* (14, 4, 31) {real, imag} */,
  {32'h3d6d3e18, 32'h3f377415} /* (14, 4, 30) {real, imag} */,
  {32'hbda543b5, 32'h3e43dbb2} /* (14, 4, 29) {real, imag} */,
  {32'hbe534e22, 32'h3ab23b20} /* (14, 4, 28) {real, imag} */,
  {32'hbe459586, 32'h3cc9647c} /* (14, 4, 27) {real, imag} */,
  {32'h3db73499, 32'h3db96754} /* (14, 4, 26) {real, imag} */,
  {32'hbe1c706b, 32'hbca69350} /* (14, 4, 25) {real, imag} */,
  {32'h3c345489, 32'hbc836e42} /* (14, 4, 24) {real, imag} */,
  {32'h3bf40c78, 32'hbc8d2958} /* (14, 4, 23) {real, imag} */,
  {32'hbd24fc52, 32'h3c8c299a} /* (14, 4, 22) {real, imag} */,
  {32'hbd143a9c, 32'hbce5cd5b} /* (14, 4, 21) {real, imag} */,
  {32'h3cc36ac2, 32'hbc74fe4a} /* (14, 4, 20) {real, imag} */,
  {32'h3d14524a, 32'h3c077ee0} /* (14, 4, 19) {real, imag} */,
  {32'hbcab4774, 32'h3c9f87c0} /* (14, 4, 18) {real, imag} */,
  {32'h3b815148, 32'hbc4b6e30} /* (14, 4, 17) {real, imag} */,
  {32'h3d8163af, 32'h00000000} /* (14, 4, 16) {real, imag} */,
  {32'h3b815148, 32'h3c4b6e30} /* (14, 4, 15) {real, imag} */,
  {32'hbcab4774, 32'hbc9f87c0} /* (14, 4, 14) {real, imag} */,
  {32'h3d14524a, 32'hbc077ee0} /* (14, 4, 13) {real, imag} */,
  {32'h3cc36ac2, 32'h3c74fe4a} /* (14, 4, 12) {real, imag} */,
  {32'hbd143a9c, 32'h3ce5cd5b} /* (14, 4, 11) {real, imag} */,
  {32'hbd24fc52, 32'hbc8c299a} /* (14, 4, 10) {real, imag} */,
  {32'h3bf40c78, 32'h3c8d2958} /* (14, 4, 9) {real, imag} */,
  {32'h3c345489, 32'h3c836e42} /* (14, 4, 8) {real, imag} */,
  {32'hbe1c706b, 32'h3ca69350} /* (14, 4, 7) {real, imag} */,
  {32'h3db73499, 32'hbdb96754} /* (14, 4, 6) {real, imag} */,
  {32'hbe459586, 32'hbcc9647c} /* (14, 4, 5) {real, imag} */,
  {32'hbe534e22, 32'hbab23b20} /* (14, 4, 4) {real, imag} */,
  {32'hbda543b5, 32'hbe43dbb2} /* (14, 4, 3) {real, imag} */,
  {32'h3d6d3e18, 32'hbf377415} /* (14, 4, 2) {real, imag} */,
  {32'h3fc8f5de, 32'h40040571} /* (14, 4, 1) {real, imag} */,
  {32'h40355c83, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'h3fc4a16e, 32'hc007d3bd} /* (14, 3, 31) {real, imag} */,
  {32'h3db1c7c0, 32'h3f3fc5b2} /* (14, 3, 30) {real, imag} */,
  {32'hbe270b19, 32'h3d8da4a8} /* (14, 3, 29) {real, imag} */,
  {32'hbe049aba, 32'h3da92cb4} /* (14, 3, 28) {real, imag} */,
  {32'hbdfc6796, 32'hbd8562de} /* (14, 3, 27) {real, imag} */,
  {32'h3db61db6, 32'hbc375401} /* (14, 3, 26) {real, imag} */,
  {32'h3db03496, 32'hbe01f9f0} /* (14, 3, 25) {real, imag} */,
  {32'h3c68fd13, 32'hbd47012a} /* (14, 3, 24) {real, imag} */,
  {32'hbc31e2c8, 32'hbd740987} /* (14, 3, 23) {real, imag} */,
  {32'hbd9caf82, 32'hbcbed3de} /* (14, 3, 22) {real, imag} */,
  {32'hbd2b96ea, 32'h3d3c0677} /* (14, 3, 21) {real, imag} */,
  {32'h3bb7bbc0, 32'hbcec4857} /* (14, 3, 20) {real, imag} */,
  {32'h3caf3d94, 32'hbc654424} /* (14, 3, 19) {real, imag} */,
  {32'h3d6fc812, 32'hbdb02cad} /* (14, 3, 18) {real, imag} */,
  {32'hbe071082, 32'h3d65ebd8} /* (14, 3, 17) {real, imag} */,
  {32'h3c0658bc, 32'h00000000} /* (14, 3, 16) {real, imag} */,
  {32'hbe071082, 32'hbd65ebd8} /* (14, 3, 15) {real, imag} */,
  {32'h3d6fc812, 32'h3db02cad} /* (14, 3, 14) {real, imag} */,
  {32'h3caf3d94, 32'h3c654424} /* (14, 3, 13) {real, imag} */,
  {32'h3bb7bbc0, 32'h3cec4857} /* (14, 3, 12) {real, imag} */,
  {32'hbd2b96ea, 32'hbd3c0677} /* (14, 3, 11) {real, imag} */,
  {32'hbd9caf82, 32'h3cbed3de} /* (14, 3, 10) {real, imag} */,
  {32'hbc31e2c8, 32'h3d740987} /* (14, 3, 9) {real, imag} */,
  {32'h3c68fd13, 32'h3d47012a} /* (14, 3, 8) {real, imag} */,
  {32'h3db03496, 32'h3e01f9f0} /* (14, 3, 7) {real, imag} */,
  {32'h3db61db6, 32'h3c375401} /* (14, 3, 6) {real, imag} */,
  {32'hbdfc6796, 32'h3d8562de} /* (14, 3, 5) {real, imag} */,
  {32'hbe049aba, 32'hbda92cb4} /* (14, 3, 4) {real, imag} */,
  {32'hbe270b19, 32'hbd8da4a8} /* (14, 3, 3) {real, imag} */,
  {32'h3db1c7c0, 32'hbf3fc5b2} /* (14, 3, 2) {real, imag} */,
  {32'h3fc4a16e, 32'h4007d3bd} /* (14, 3, 1) {real, imag} */,
  {32'h4041208e, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h3fc9cfd6, 32'hc0020043} /* (14, 2, 31) {real, imag} */,
  {32'h3e32b0cc, 32'h3f29c3ce} /* (14, 2, 30) {real, imag} */,
  {32'hbdaf7afe, 32'h3df53f8e} /* (14, 2, 29) {real, imag} */,
  {32'hbdaf48ee, 32'h3e16ea52} /* (14, 2, 28) {real, imag} */,
  {32'hbe68f1f9, 32'hbd8f14d2} /* (14, 2, 27) {real, imag} */,
  {32'hbd8879c2, 32'hbd055982} /* (14, 2, 26) {real, imag} */,
  {32'hbd4d95b9, 32'hbdf4e82c} /* (14, 2, 25) {real, imag} */,
  {32'hbd017459, 32'hbd9e04d4} /* (14, 2, 24) {real, imag} */,
  {32'h3cfffc18, 32'hbdf63932} /* (14, 2, 23) {real, imag} */,
  {32'hbd824dd6, 32'h3d921c43} /* (14, 2, 22) {real, imag} */,
  {32'hbd6f0c84, 32'hbd1945ca} /* (14, 2, 21) {real, imag} */,
  {32'h3d6ebd4e, 32'h3d70a07f} /* (14, 2, 20) {real, imag} */,
  {32'hbd8a6c88, 32'h3d154fa8} /* (14, 2, 19) {real, imag} */,
  {32'h3c571d22, 32'h3dc832b4} /* (14, 2, 18) {real, imag} */,
  {32'hbc4fa020, 32'hbd10795c} /* (14, 2, 17) {real, imag} */,
  {32'h3d00a05f, 32'h00000000} /* (14, 2, 16) {real, imag} */,
  {32'hbc4fa020, 32'h3d10795c} /* (14, 2, 15) {real, imag} */,
  {32'h3c571d22, 32'hbdc832b4} /* (14, 2, 14) {real, imag} */,
  {32'hbd8a6c88, 32'hbd154fa8} /* (14, 2, 13) {real, imag} */,
  {32'h3d6ebd4e, 32'hbd70a07f} /* (14, 2, 12) {real, imag} */,
  {32'hbd6f0c84, 32'h3d1945ca} /* (14, 2, 11) {real, imag} */,
  {32'hbd824dd6, 32'hbd921c43} /* (14, 2, 10) {real, imag} */,
  {32'h3cfffc18, 32'h3df63932} /* (14, 2, 9) {real, imag} */,
  {32'hbd017459, 32'h3d9e04d4} /* (14, 2, 8) {real, imag} */,
  {32'hbd4d95b9, 32'h3df4e82c} /* (14, 2, 7) {real, imag} */,
  {32'hbd8879c2, 32'h3d055982} /* (14, 2, 6) {real, imag} */,
  {32'hbe68f1f9, 32'h3d8f14d2} /* (14, 2, 5) {real, imag} */,
  {32'hbdaf48ee, 32'hbe16ea52} /* (14, 2, 4) {real, imag} */,
  {32'hbdaf7afe, 32'hbdf53f8e} /* (14, 2, 3) {real, imag} */,
  {32'h3e32b0cc, 32'hbf29c3ce} /* (14, 2, 2) {real, imag} */,
  {32'h3fc9cfd6, 32'h40020043} /* (14, 2, 1) {real, imag} */,
  {32'h4032c1de, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h3fce41bc, 32'hc0018ebb} /* (14, 1, 31) {real, imag} */,
  {32'h3dd31b54, 32'h3f098264} /* (14, 1, 30) {real, imag} */,
  {32'hbe4dd37e, 32'h3dadc47e} /* (14, 1, 29) {real, imag} */,
  {32'hbe0b5042, 32'h3dc5e3a7} /* (14, 1, 28) {real, imag} */,
  {32'hbe1eb710, 32'hbd89b560} /* (14, 1, 27) {real, imag} */,
  {32'hbd29b154, 32'h3c36a75c} /* (14, 1, 26) {real, imag} */,
  {32'hbdaa6b25, 32'h3d63d979} /* (14, 1, 25) {real, imag} */,
  {32'h3c9c20bc, 32'h3b894a34} /* (14, 1, 24) {real, imag} */,
  {32'h3c4e8518, 32'h3bda920c} /* (14, 1, 23) {real, imag} */,
  {32'hbd984894, 32'hbda82c32} /* (14, 1, 22) {real, imag} */,
  {32'hbd51808e, 32'hbc619c5f} /* (14, 1, 21) {real, imag} */,
  {32'h3d4a32e9, 32'h3d73bb48} /* (14, 1, 20) {real, imag} */,
  {32'h3d08b679, 32'hbdc4ae75} /* (14, 1, 19) {real, imag} */,
  {32'h3c4f8b78, 32'h3cc64800} /* (14, 1, 18) {real, imag} */,
  {32'h3ce0dd57, 32'h3d928cb8} /* (14, 1, 17) {real, imag} */,
  {32'h3d047007, 32'h00000000} /* (14, 1, 16) {real, imag} */,
  {32'h3ce0dd57, 32'hbd928cb8} /* (14, 1, 15) {real, imag} */,
  {32'h3c4f8b78, 32'hbcc64800} /* (14, 1, 14) {real, imag} */,
  {32'h3d08b679, 32'h3dc4ae75} /* (14, 1, 13) {real, imag} */,
  {32'h3d4a32e9, 32'hbd73bb48} /* (14, 1, 12) {real, imag} */,
  {32'hbd51808e, 32'h3c619c5f} /* (14, 1, 11) {real, imag} */,
  {32'hbd984894, 32'h3da82c32} /* (14, 1, 10) {real, imag} */,
  {32'h3c4e8518, 32'hbbda920c} /* (14, 1, 9) {real, imag} */,
  {32'h3c9c20bc, 32'hbb894a34} /* (14, 1, 8) {real, imag} */,
  {32'hbdaa6b25, 32'hbd63d979} /* (14, 1, 7) {real, imag} */,
  {32'hbd29b154, 32'hbc36a75c} /* (14, 1, 6) {real, imag} */,
  {32'hbe1eb710, 32'h3d89b560} /* (14, 1, 5) {real, imag} */,
  {32'hbe0b5042, 32'hbdc5e3a7} /* (14, 1, 4) {real, imag} */,
  {32'hbe4dd37e, 32'hbdadc47e} /* (14, 1, 3) {real, imag} */,
  {32'h3dd31b54, 32'hbf098264} /* (14, 1, 2) {real, imag} */,
  {32'h3fce41bc, 32'h40018ebb} /* (14, 1, 1) {real, imag} */,
  {32'h4022cb82, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h3fd3fa4d, 32'hbfd42970} /* (14, 0, 31) {real, imag} */,
  {32'hbe073970, 32'h3ebe42ef} /* (14, 0, 30) {real, imag} */,
  {32'hbe097bba, 32'h3c162d70} /* (14, 0, 29) {real, imag} */,
  {32'hbde7c704, 32'h3e077f51} /* (14, 0, 28) {real, imag} */,
  {32'hbdffa789, 32'hbd326b57} /* (14, 0, 27) {real, imag} */,
  {32'h3d300d59, 32'hbc953d26} /* (14, 0, 26) {real, imag} */,
  {32'h3cda6579, 32'hbc1552f1} /* (14, 0, 25) {real, imag} */,
  {32'hbc33bee6, 32'hbd245811} /* (14, 0, 24) {real, imag} */,
  {32'hbd60688e, 32'h3c02426c} /* (14, 0, 23) {real, imag} */,
  {32'h3c4bb42c, 32'hbcfa18d4} /* (14, 0, 22) {real, imag} */,
  {32'h3d2b6e2d, 32'h3d4acfc9} /* (14, 0, 21) {real, imag} */,
  {32'hbbd3f4c6, 32'h3c22cb10} /* (14, 0, 20) {real, imag} */,
  {32'h3b8b3bf8, 32'h3cf94e1c} /* (14, 0, 19) {real, imag} */,
  {32'h3d52c632, 32'hbd591080} /* (14, 0, 18) {real, imag} */,
  {32'hbd30546c, 32'h3c64105c} /* (14, 0, 17) {real, imag} */,
  {32'hbd0b1247, 32'h00000000} /* (14, 0, 16) {real, imag} */,
  {32'hbd30546c, 32'hbc64105c} /* (14, 0, 15) {real, imag} */,
  {32'h3d52c632, 32'h3d591080} /* (14, 0, 14) {real, imag} */,
  {32'h3b8b3bf8, 32'hbcf94e1c} /* (14, 0, 13) {real, imag} */,
  {32'hbbd3f4c6, 32'hbc22cb10} /* (14, 0, 12) {real, imag} */,
  {32'h3d2b6e2d, 32'hbd4acfc9} /* (14, 0, 11) {real, imag} */,
  {32'h3c4bb42c, 32'h3cfa18d4} /* (14, 0, 10) {real, imag} */,
  {32'hbd60688e, 32'hbc02426c} /* (14, 0, 9) {real, imag} */,
  {32'hbc33bee6, 32'h3d245811} /* (14, 0, 8) {real, imag} */,
  {32'h3cda6579, 32'h3c1552f1} /* (14, 0, 7) {real, imag} */,
  {32'h3d300d59, 32'h3c953d26} /* (14, 0, 6) {real, imag} */,
  {32'hbdffa789, 32'h3d326b57} /* (14, 0, 5) {real, imag} */,
  {32'hbde7c704, 32'hbe077f51} /* (14, 0, 4) {real, imag} */,
  {32'hbe097bba, 32'hbc162d70} /* (14, 0, 3) {real, imag} */,
  {32'hbe073970, 32'hbebe42ef} /* (14, 0, 2) {real, imag} */,
  {32'h3fd3fa4d, 32'h3fd42970} /* (14, 0, 1) {real, imag} */,
  {32'h40126baa, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h403a3993, 32'hbfdc5cca} /* (13, 31, 31) {real, imag} */,
  {32'hbf2e461c, 32'h3eb3c684} /* (13, 31, 30) {real, imag} */,
  {32'hbdc73438, 32'h3ca9777c} /* (13, 31, 29) {real, imag} */,
  {32'hbce864d4, 32'hbcad0c28} /* (13, 31, 28) {real, imag} */,
  {32'hbde31f01, 32'hbe0bf3d8} /* (13, 31, 27) {real, imag} */,
  {32'h3d84e654, 32'hbdcdb984} /* (13, 31, 26) {real, imag} */,
  {32'hbcb513b2, 32'h3d3a7baa} /* (13, 31, 25) {real, imag} */,
  {32'hbd9db974, 32'h3cf60137} /* (13, 31, 24) {real, imag} */,
  {32'hbdc3b318, 32'h3dbdd816} /* (13, 31, 23) {real, imag} */,
  {32'h3a4e1e20, 32'h3d37fc3c} /* (13, 31, 22) {real, imag} */,
  {32'h3bd13d94, 32'h3d3d02ab} /* (13, 31, 21) {real, imag} */,
  {32'hbb9ed370, 32'hbc8dddf2} /* (13, 31, 20) {real, imag} */,
  {32'hbd0ca99c, 32'hbcaf6db4} /* (13, 31, 19) {real, imag} */,
  {32'h3d1516be, 32'h3d6e6ce6} /* (13, 31, 18) {real, imag} */,
  {32'h3ca8c7a0, 32'h3d18a27e} /* (13, 31, 17) {real, imag} */,
  {32'h3d392964, 32'h00000000} /* (13, 31, 16) {real, imag} */,
  {32'h3ca8c7a0, 32'hbd18a27e} /* (13, 31, 15) {real, imag} */,
  {32'h3d1516be, 32'hbd6e6ce6} /* (13, 31, 14) {real, imag} */,
  {32'hbd0ca99c, 32'h3caf6db4} /* (13, 31, 13) {real, imag} */,
  {32'hbb9ed370, 32'h3c8dddf2} /* (13, 31, 12) {real, imag} */,
  {32'h3bd13d94, 32'hbd3d02ab} /* (13, 31, 11) {real, imag} */,
  {32'h3a4e1e20, 32'hbd37fc3c} /* (13, 31, 10) {real, imag} */,
  {32'hbdc3b318, 32'hbdbdd816} /* (13, 31, 9) {real, imag} */,
  {32'hbd9db974, 32'hbcf60137} /* (13, 31, 8) {real, imag} */,
  {32'hbcb513b2, 32'hbd3a7baa} /* (13, 31, 7) {real, imag} */,
  {32'h3d84e654, 32'h3dcdb984} /* (13, 31, 6) {real, imag} */,
  {32'hbde31f01, 32'h3e0bf3d8} /* (13, 31, 5) {real, imag} */,
  {32'hbce864d4, 32'h3cad0c28} /* (13, 31, 4) {real, imag} */,
  {32'hbdc73438, 32'hbca9777c} /* (13, 31, 3) {real, imag} */,
  {32'hbf2e461c, 32'hbeb3c684} /* (13, 31, 2) {real, imag} */,
  {32'h403a3993, 32'h3fdc5cca} /* (13, 31, 1) {real, imag} */,
  {32'h40708aa0, 32'h00000000} /* (13, 31, 0) {real, imag} */,
  {32'h4054571a, 32'hbfabdc7e} /* (13, 30, 31) {real, imag} */,
  {32'hbf944aa7, 32'h3eb1d5a4} /* (13, 30, 30) {real, imag} */,
  {32'hbcd7f900, 32'h3dc4c2f2} /* (13, 30, 29) {real, imag} */,
  {32'h3e26cde5, 32'hbdb97aac} /* (13, 30, 28) {real, imag} */,
  {32'hbe4110e9, 32'hbdebc80c} /* (13, 30, 27) {real, imag} */,
  {32'h3d026cf1, 32'hbc1628d0} /* (13, 30, 26) {real, imag} */,
  {32'h3caec43e, 32'hbcd381d0} /* (13, 30, 25) {real, imag} */,
  {32'hbd8599e0, 32'h3d9c9582} /* (13, 30, 24) {real, imag} */,
  {32'hbd4de024, 32'hbb3f6a50} /* (13, 30, 23) {real, imag} */,
  {32'h3dcfd1a5, 32'hbe1b9266} /* (13, 30, 22) {real, imag} */,
  {32'hbae328c0, 32'h3c7308fc} /* (13, 30, 21) {real, imag} */,
  {32'hbd0fb1f8, 32'h3e2aec93} /* (13, 30, 20) {real, imag} */,
  {32'hbd1d69d8, 32'hbd76ad62} /* (13, 30, 19) {real, imag} */,
  {32'hbcbde2a3, 32'hbd263deb} /* (13, 30, 18) {real, imag} */,
  {32'hbb84283c, 32'hbd2ec59e} /* (13, 30, 17) {real, imag} */,
  {32'h3c15d758, 32'h00000000} /* (13, 30, 16) {real, imag} */,
  {32'hbb84283c, 32'h3d2ec59e} /* (13, 30, 15) {real, imag} */,
  {32'hbcbde2a3, 32'h3d263deb} /* (13, 30, 14) {real, imag} */,
  {32'hbd1d69d8, 32'h3d76ad62} /* (13, 30, 13) {real, imag} */,
  {32'hbd0fb1f8, 32'hbe2aec93} /* (13, 30, 12) {real, imag} */,
  {32'hbae328c0, 32'hbc7308fc} /* (13, 30, 11) {real, imag} */,
  {32'h3dcfd1a5, 32'h3e1b9266} /* (13, 30, 10) {real, imag} */,
  {32'hbd4de024, 32'h3b3f6a50} /* (13, 30, 9) {real, imag} */,
  {32'hbd8599e0, 32'hbd9c9582} /* (13, 30, 8) {real, imag} */,
  {32'h3caec43e, 32'h3cd381d0} /* (13, 30, 7) {real, imag} */,
  {32'h3d026cf1, 32'h3c1628d0} /* (13, 30, 6) {real, imag} */,
  {32'hbe4110e9, 32'h3debc80c} /* (13, 30, 5) {real, imag} */,
  {32'h3e26cde5, 32'h3db97aac} /* (13, 30, 4) {real, imag} */,
  {32'hbcd7f900, 32'hbdc4c2f2} /* (13, 30, 3) {real, imag} */,
  {32'hbf944aa7, 32'hbeb1d5a4} /* (13, 30, 2) {real, imag} */,
  {32'h4054571a, 32'h3fabdc7e} /* (13, 30, 1) {real, imag} */,
  {32'h40789434, 32'h00000000} /* (13, 30, 0) {real, imag} */,
  {32'h40671dcf, 32'hbf7f0678} /* (13, 29, 31) {real, imag} */,
  {32'hbfa04b8a, 32'h3ea1fffe} /* (13, 29, 30) {real, imag} */,
  {32'h3e258a0f, 32'h3dd638ce} /* (13, 29, 29) {real, imag} */,
  {32'h3e1155ed, 32'hbd9d3845} /* (13, 29, 28) {real, imag} */,
  {32'hbe0dd511, 32'hbb32f510} /* (13, 29, 27) {real, imag} */,
  {32'h3b625bcc, 32'hbcf090ac} /* (13, 29, 26) {real, imag} */,
  {32'hbb295948, 32'hbd05c89f} /* (13, 29, 25) {real, imag} */,
  {32'hbe554480, 32'h3e298d62} /* (13, 29, 24) {real, imag} */,
  {32'hbda3ff15, 32'h3e02d5f7} /* (13, 29, 23) {real, imag} */,
  {32'h3d42cacf, 32'hbc3b9a5a} /* (13, 29, 22) {real, imag} */,
  {32'hbc50c70a, 32'h3cdcc9c8} /* (13, 29, 21) {real, imag} */,
  {32'hbd830fd2, 32'h3c80add6} /* (13, 29, 20) {real, imag} */,
  {32'hbda6f722, 32'hbc43fb54} /* (13, 29, 19) {real, imag} */,
  {32'h3cb22a4a, 32'hbd4c5fb5} /* (13, 29, 18) {real, imag} */,
  {32'hbd9e59d4, 32'hbc170ce2} /* (13, 29, 17) {real, imag} */,
  {32'hbd0ba8f7, 32'h00000000} /* (13, 29, 16) {real, imag} */,
  {32'hbd9e59d4, 32'h3c170ce2} /* (13, 29, 15) {real, imag} */,
  {32'h3cb22a4a, 32'h3d4c5fb5} /* (13, 29, 14) {real, imag} */,
  {32'hbda6f722, 32'h3c43fb54} /* (13, 29, 13) {real, imag} */,
  {32'hbd830fd2, 32'hbc80add6} /* (13, 29, 12) {real, imag} */,
  {32'hbc50c70a, 32'hbcdcc9c8} /* (13, 29, 11) {real, imag} */,
  {32'h3d42cacf, 32'h3c3b9a5a} /* (13, 29, 10) {real, imag} */,
  {32'hbda3ff15, 32'hbe02d5f7} /* (13, 29, 9) {real, imag} */,
  {32'hbe554480, 32'hbe298d62} /* (13, 29, 8) {real, imag} */,
  {32'hbb295948, 32'h3d05c89f} /* (13, 29, 7) {real, imag} */,
  {32'h3b625bcc, 32'h3cf090ac} /* (13, 29, 6) {real, imag} */,
  {32'hbe0dd511, 32'h3b32f510} /* (13, 29, 5) {real, imag} */,
  {32'h3e1155ed, 32'h3d9d3845} /* (13, 29, 4) {real, imag} */,
  {32'h3e258a0f, 32'hbdd638ce} /* (13, 29, 3) {real, imag} */,
  {32'hbfa04b8a, 32'hbea1fffe} /* (13, 29, 2) {real, imag} */,
  {32'h40671dcf, 32'h3f7f0678} /* (13, 29, 1) {real, imag} */,
  {32'h407c6bc2, 32'h00000000} /* (13, 29, 0) {real, imag} */,
  {32'h406d3b6c, 32'hbf638032} /* (13, 28, 31) {real, imag} */,
  {32'hbfaecae2, 32'h3e826f26} /* (13, 28, 30) {real, imag} */,
  {32'hbb8dc15c, 32'hbc87b0f6} /* (13, 28, 29) {real, imag} */,
  {32'h3d678c54, 32'hbe4226f3} /* (13, 28, 28) {real, imag} */,
  {32'hbd3351a6, 32'h3d79e24c} /* (13, 28, 27) {real, imag} */,
  {32'h3d295226, 32'h3c32863c} /* (13, 28, 26) {real, imag} */,
  {32'h3d337aa7, 32'h3d04a6ff} /* (13, 28, 25) {real, imag} */,
  {32'hbcf8c841, 32'h3df2c819} /* (13, 28, 24) {real, imag} */,
  {32'hbdd6c8c1, 32'h3b35ce98} /* (13, 28, 23) {real, imag} */,
  {32'hbdd30a0e, 32'h3ca35150} /* (13, 28, 22) {real, imag} */,
  {32'hbc808339, 32'h3b816bc8} /* (13, 28, 21) {real, imag} */,
  {32'h3d264821, 32'hbd9f1d6d} /* (13, 28, 20) {real, imag} */,
  {32'h3d86bfa4, 32'hbc296497} /* (13, 28, 19) {real, imag} */,
  {32'h3d0cfa14, 32'h3d6d6668} /* (13, 28, 18) {real, imag} */,
  {32'h3d15c4e2, 32'h3ca6fa94} /* (13, 28, 17) {real, imag} */,
  {32'hbd56ce0a, 32'h00000000} /* (13, 28, 16) {real, imag} */,
  {32'h3d15c4e2, 32'hbca6fa94} /* (13, 28, 15) {real, imag} */,
  {32'h3d0cfa14, 32'hbd6d6668} /* (13, 28, 14) {real, imag} */,
  {32'h3d86bfa4, 32'h3c296497} /* (13, 28, 13) {real, imag} */,
  {32'h3d264821, 32'h3d9f1d6d} /* (13, 28, 12) {real, imag} */,
  {32'hbc808339, 32'hbb816bc8} /* (13, 28, 11) {real, imag} */,
  {32'hbdd30a0e, 32'hbca35150} /* (13, 28, 10) {real, imag} */,
  {32'hbdd6c8c1, 32'hbb35ce98} /* (13, 28, 9) {real, imag} */,
  {32'hbcf8c841, 32'hbdf2c819} /* (13, 28, 8) {real, imag} */,
  {32'h3d337aa7, 32'hbd04a6ff} /* (13, 28, 7) {real, imag} */,
  {32'h3d295226, 32'hbc32863c} /* (13, 28, 6) {real, imag} */,
  {32'hbd3351a6, 32'hbd79e24c} /* (13, 28, 5) {real, imag} */,
  {32'h3d678c54, 32'h3e4226f3} /* (13, 28, 4) {real, imag} */,
  {32'hbb8dc15c, 32'h3c87b0f6} /* (13, 28, 3) {real, imag} */,
  {32'hbfaecae2, 32'hbe826f26} /* (13, 28, 2) {real, imag} */,
  {32'h406d3b6c, 32'h3f638032} /* (13, 28, 1) {real, imag} */,
  {32'h4074286a, 32'h00000000} /* (13, 28, 0) {real, imag} */,
  {32'h407069b0, 32'hbf5d5c91} /* (13, 27, 31) {real, imag} */,
  {32'hbfbbdd31, 32'h3e4e3804} /* (13, 27, 30) {real, imag} */,
  {32'h3cbca0c0, 32'hbe025356} /* (13, 27, 29) {real, imag} */,
  {32'h3d588a80, 32'hbe375fa6} /* (13, 27, 28) {real, imag} */,
  {32'hbdf25d0a, 32'h3e2e7522} /* (13, 27, 27) {real, imag} */,
  {32'hbd33f0c4, 32'h3d25a00b} /* (13, 27, 26) {real, imag} */,
  {32'h3dae90b4, 32'hbcda6f8a} /* (13, 27, 25) {real, imag} */,
  {32'h3c9e0cde, 32'h3d6d2dd7} /* (13, 27, 24) {real, imag} */,
  {32'h3c9ea78e, 32'hbdb5d36b} /* (13, 27, 23) {real, imag} */,
  {32'h3dc533da, 32'hbc370094} /* (13, 27, 22) {real, imag} */,
  {32'hbda6fa04, 32'h3d09470c} /* (13, 27, 21) {real, imag} */,
  {32'h3da54166, 32'h3e18f85e} /* (13, 27, 20) {real, imag} */,
  {32'h3d2a8f18, 32'hbc42d820} /* (13, 27, 19) {real, imag} */,
  {32'h3d4dbd5f, 32'h3c256713} /* (13, 27, 18) {real, imag} */,
  {32'hbda29b71, 32'h3b048c68} /* (13, 27, 17) {real, imag} */,
  {32'h3d26d8b2, 32'h00000000} /* (13, 27, 16) {real, imag} */,
  {32'hbda29b71, 32'hbb048c68} /* (13, 27, 15) {real, imag} */,
  {32'h3d4dbd5f, 32'hbc256713} /* (13, 27, 14) {real, imag} */,
  {32'h3d2a8f18, 32'h3c42d820} /* (13, 27, 13) {real, imag} */,
  {32'h3da54166, 32'hbe18f85e} /* (13, 27, 12) {real, imag} */,
  {32'hbda6fa04, 32'hbd09470c} /* (13, 27, 11) {real, imag} */,
  {32'h3dc533da, 32'h3c370094} /* (13, 27, 10) {real, imag} */,
  {32'h3c9ea78e, 32'h3db5d36b} /* (13, 27, 9) {real, imag} */,
  {32'h3c9e0cde, 32'hbd6d2dd7} /* (13, 27, 8) {real, imag} */,
  {32'h3dae90b4, 32'h3cda6f8a} /* (13, 27, 7) {real, imag} */,
  {32'hbd33f0c4, 32'hbd25a00b} /* (13, 27, 6) {real, imag} */,
  {32'hbdf25d0a, 32'hbe2e7522} /* (13, 27, 5) {real, imag} */,
  {32'h3d588a80, 32'h3e375fa6} /* (13, 27, 4) {real, imag} */,
  {32'h3cbca0c0, 32'h3e025356} /* (13, 27, 3) {real, imag} */,
  {32'hbfbbdd31, 32'hbe4e3804} /* (13, 27, 2) {real, imag} */,
  {32'h407069b0, 32'h3f5d5c91} /* (13, 27, 1) {real, imag} */,
  {32'h40760581, 32'h00000000} /* (13, 27, 0) {real, imag} */,
  {32'h406fb89a, 32'hbf307fa5} /* (13, 26, 31) {real, imag} */,
  {32'hbfc6962a, 32'h3e33078e} /* (13, 26, 30) {real, imag} */,
  {32'hbdace63a, 32'hbd93c3c6} /* (13, 26, 29) {real, imag} */,
  {32'h3e056ad7, 32'hbe3ec25f} /* (13, 26, 28) {real, imag} */,
  {32'hbd756067, 32'h3deff9be} /* (13, 26, 27) {real, imag} */,
  {32'hbdbddc62, 32'hbd308716} /* (13, 26, 26) {real, imag} */,
  {32'hbd07b8f0, 32'hbd4e71bb} /* (13, 26, 25) {real, imag} */,
  {32'hbe263c5e, 32'h3dae3535} /* (13, 26, 24) {real, imag} */,
  {32'h3d01e583, 32'h3d8938da} /* (13, 26, 23) {real, imag} */,
  {32'h3d9cfda6, 32'h3d8d87e3} /* (13, 26, 22) {real, imag} */,
  {32'hbd9b5c22, 32'hbe4750b4} /* (13, 26, 21) {real, imag} */,
  {32'hbd536dc8, 32'h3c75fa96} /* (13, 26, 20) {real, imag} */,
  {32'hbb927834, 32'h3c40eeb8} /* (13, 26, 19) {real, imag} */,
  {32'h3c99e129, 32'hbc1cc34a} /* (13, 26, 18) {real, imag} */,
  {32'h3d00b408, 32'h3cf444bb} /* (13, 26, 17) {real, imag} */,
  {32'hbd9886fa, 32'h00000000} /* (13, 26, 16) {real, imag} */,
  {32'h3d00b408, 32'hbcf444bb} /* (13, 26, 15) {real, imag} */,
  {32'h3c99e129, 32'h3c1cc34a} /* (13, 26, 14) {real, imag} */,
  {32'hbb927834, 32'hbc40eeb8} /* (13, 26, 13) {real, imag} */,
  {32'hbd536dc8, 32'hbc75fa96} /* (13, 26, 12) {real, imag} */,
  {32'hbd9b5c22, 32'h3e4750b4} /* (13, 26, 11) {real, imag} */,
  {32'h3d9cfda6, 32'hbd8d87e3} /* (13, 26, 10) {real, imag} */,
  {32'h3d01e583, 32'hbd8938da} /* (13, 26, 9) {real, imag} */,
  {32'hbe263c5e, 32'hbdae3535} /* (13, 26, 8) {real, imag} */,
  {32'hbd07b8f0, 32'h3d4e71bb} /* (13, 26, 7) {real, imag} */,
  {32'hbdbddc62, 32'h3d308716} /* (13, 26, 6) {real, imag} */,
  {32'hbd756067, 32'hbdeff9be} /* (13, 26, 5) {real, imag} */,
  {32'h3e056ad7, 32'h3e3ec25f} /* (13, 26, 4) {real, imag} */,
  {32'hbdace63a, 32'h3d93c3c6} /* (13, 26, 3) {real, imag} */,
  {32'hbfc6962a, 32'hbe33078e} /* (13, 26, 2) {real, imag} */,
  {32'h406fb89a, 32'h3f307fa5} /* (13, 26, 1) {real, imag} */,
  {32'h4068a0c4, 32'h00000000} /* (13, 26, 0) {real, imag} */,
  {32'h4068c330, 32'hbf2aee1b} /* (13, 25, 31) {real, imag} */,
  {32'hbfc36562, 32'h3e748719} /* (13, 25, 30) {real, imag} */,
  {32'hbd4880fe, 32'hbde349e0} /* (13, 25, 29) {real, imag} */,
  {32'h3e6c7139, 32'hbddf8180} /* (13, 25, 28) {real, imag} */,
  {32'hbe4bce94, 32'h3db25794} /* (13, 25, 27) {real, imag} */,
  {32'hbce83300, 32'hbdf3ad08} /* (13, 25, 26) {real, imag} */,
  {32'h3c48a408, 32'hbc84c29c} /* (13, 25, 25) {real, imag} */,
  {32'hbbe80850, 32'h3e015cfb} /* (13, 25, 24) {real, imag} */,
  {32'h3d99563a, 32'h3dd39d42} /* (13, 25, 23) {real, imag} */,
  {32'hbdbd6f96, 32'hbd7798a3} /* (13, 25, 22) {real, imag} */,
  {32'h3d9f039a, 32'hbc94f9b0} /* (13, 25, 21) {real, imag} */,
  {32'h3c1f037a, 32'h3ba5ae58} /* (13, 25, 20) {real, imag} */,
  {32'h3d41c991, 32'hbd06889a} /* (13, 25, 19) {real, imag} */,
  {32'hba67db60, 32'h3d495192} /* (13, 25, 18) {real, imag} */,
  {32'hbd8d7883, 32'hbd8bc598} /* (13, 25, 17) {real, imag} */,
  {32'hbd91057a, 32'h00000000} /* (13, 25, 16) {real, imag} */,
  {32'hbd8d7883, 32'h3d8bc598} /* (13, 25, 15) {real, imag} */,
  {32'hba67db60, 32'hbd495192} /* (13, 25, 14) {real, imag} */,
  {32'h3d41c991, 32'h3d06889a} /* (13, 25, 13) {real, imag} */,
  {32'h3c1f037a, 32'hbba5ae58} /* (13, 25, 12) {real, imag} */,
  {32'h3d9f039a, 32'h3c94f9b0} /* (13, 25, 11) {real, imag} */,
  {32'hbdbd6f96, 32'h3d7798a3} /* (13, 25, 10) {real, imag} */,
  {32'h3d99563a, 32'hbdd39d42} /* (13, 25, 9) {real, imag} */,
  {32'hbbe80850, 32'hbe015cfb} /* (13, 25, 8) {real, imag} */,
  {32'h3c48a408, 32'h3c84c29c} /* (13, 25, 7) {real, imag} */,
  {32'hbce83300, 32'h3df3ad08} /* (13, 25, 6) {real, imag} */,
  {32'hbe4bce94, 32'hbdb25794} /* (13, 25, 5) {real, imag} */,
  {32'h3e6c7139, 32'h3ddf8180} /* (13, 25, 4) {real, imag} */,
  {32'hbd4880fe, 32'h3de349e0} /* (13, 25, 3) {real, imag} */,
  {32'hbfc36562, 32'hbe748719} /* (13, 25, 2) {real, imag} */,
  {32'h4068c330, 32'h3f2aee1b} /* (13, 25, 1) {real, imag} */,
  {32'h405378e4, 32'h00000000} /* (13, 25, 0) {real, imag} */,
  {32'h4054d23d, 32'hbf2b1978} /* (13, 24, 31) {real, imag} */,
  {32'hbfbc5d71, 32'h3eb74457} /* (13, 24, 30) {real, imag} */,
  {32'h3c7abfec, 32'hbe56ca8e} /* (13, 24, 29) {real, imag} */,
  {32'h3e849e7c, 32'hbd8dac74} /* (13, 24, 28) {real, imag} */,
  {32'hbe62045e, 32'h3e2c8c35} /* (13, 24, 27) {real, imag} */,
  {32'hbd326f5f, 32'hbe4bed18} /* (13, 24, 26) {real, imag} */,
  {32'h3d42e1db, 32'h3d96f9e1} /* (13, 24, 25) {real, imag} */,
  {32'h3d125b14, 32'h3d7a24ee} /* (13, 24, 24) {real, imag} */,
  {32'h3e1ef564, 32'h3d1c0cc4} /* (13, 24, 23) {real, imag} */,
  {32'hbd6d0132, 32'hbd1b975d} /* (13, 24, 22) {real, imag} */,
  {32'h3d6e6cea, 32'h3d28e994} /* (13, 24, 21) {real, imag} */,
  {32'hbd097840, 32'h3c63a864} /* (13, 24, 20) {real, imag} */,
  {32'h3d158132, 32'hbdf9223e} /* (13, 24, 19) {real, imag} */,
  {32'hbd23750c, 32'h3d14b87e} /* (13, 24, 18) {real, imag} */,
  {32'hbb0bf3e0, 32'h3c4942c2} /* (13, 24, 17) {real, imag} */,
  {32'h3ce3f4ea, 32'h00000000} /* (13, 24, 16) {real, imag} */,
  {32'hbb0bf3e0, 32'hbc4942c2} /* (13, 24, 15) {real, imag} */,
  {32'hbd23750c, 32'hbd14b87e} /* (13, 24, 14) {real, imag} */,
  {32'h3d158132, 32'h3df9223e} /* (13, 24, 13) {real, imag} */,
  {32'hbd097840, 32'hbc63a864} /* (13, 24, 12) {real, imag} */,
  {32'h3d6e6cea, 32'hbd28e994} /* (13, 24, 11) {real, imag} */,
  {32'hbd6d0132, 32'h3d1b975d} /* (13, 24, 10) {real, imag} */,
  {32'h3e1ef564, 32'hbd1c0cc4} /* (13, 24, 9) {real, imag} */,
  {32'h3d125b14, 32'hbd7a24ee} /* (13, 24, 8) {real, imag} */,
  {32'h3d42e1db, 32'hbd96f9e1} /* (13, 24, 7) {real, imag} */,
  {32'hbd326f5f, 32'h3e4bed18} /* (13, 24, 6) {real, imag} */,
  {32'hbe62045e, 32'hbe2c8c35} /* (13, 24, 5) {real, imag} */,
  {32'h3e849e7c, 32'h3d8dac74} /* (13, 24, 4) {real, imag} */,
  {32'h3c7abfec, 32'h3e56ca8e} /* (13, 24, 3) {real, imag} */,
  {32'hbfbc5d71, 32'hbeb74457} /* (13, 24, 2) {real, imag} */,
  {32'h4054d23d, 32'h3f2b1978} /* (13, 24, 1) {real, imag} */,
  {32'h40266250, 32'h00000000} /* (13, 24, 0) {real, imag} */,
  {32'h40320657, 32'hbee5cbde} /* (13, 23, 31) {real, imag} */,
  {32'hbf9083ed, 32'h3eb9a7bc} /* (13, 23, 30) {real, imag} */,
  {32'hbd83cba6, 32'hbe327d54} /* (13, 23, 29) {real, imag} */,
  {32'h3e8007d2, 32'hbe15ef53} /* (13, 23, 28) {real, imag} */,
  {32'hbe2639c9, 32'h3db59888} /* (13, 23, 27) {real, imag} */,
  {32'hbdace850, 32'h3b7307f8} /* (13, 23, 26) {real, imag} */,
  {32'h3cd68292, 32'hbd843a43} /* (13, 23, 25) {real, imag} */,
  {32'hbd56b61b, 32'h3cc1ab04} /* (13, 23, 24) {real, imag} */,
  {32'h3d1c0529, 32'h3d43ce59} /* (13, 23, 23) {real, imag} */,
  {32'hbd5dacd3, 32'h3c95c762} /* (13, 23, 22) {real, imag} */,
  {32'hbd2f048f, 32'h3c03cab0} /* (13, 23, 21) {real, imag} */,
  {32'h3d4158a6, 32'h3c8b7bfa} /* (13, 23, 20) {real, imag} */,
  {32'hbd11d11c, 32'h3ca49524} /* (13, 23, 19) {real, imag} */,
  {32'hbc3378b8, 32'h3dc66907} /* (13, 23, 18) {real, imag} */,
  {32'h3d6814dc, 32'hbcd6ec17} /* (13, 23, 17) {real, imag} */,
  {32'h3d2ae316, 32'h00000000} /* (13, 23, 16) {real, imag} */,
  {32'h3d6814dc, 32'h3cd6ec17} /* (13, 23, 15) {real, imag} */,
  {32'hbc3378b8, 32'hbdc66907} /* (13, 23, 14) {real, imag} */,
  {32'hbd11d11c, 32'hbca49524} /* (13, 23, 13) {real, imag} */,
  {32'h3d4158a6, 32'hbc8b7bfa} /* (13, 23, 12) {real, imag} */,
  {32'hbd2f048f, 32'hbc03cab0} /* (13, 23, 11) {real, imag} */,
  {32'hbd5dacd3, 32'hbc95c762} /* (13, 23, 10) {real, imag} */,
  {32'h3d1c0529, 32'hbd43ce59} /* (13, 23, 9) {real, imag} */,
  {32'hbd56b61b, 32'hbcc1ab04} /* (13, 23, 8) {real, imag} */,
  {32'h3cd68292, 32'h3d843a43} /* (13, 23, 7) {real, imag} */,
  {32'hbdace850, 32'hbb7307f8} /* (13, 23, 6) {real, imag} */,
  {32'hbe2639c9, 32'hbdb59888} /* (13, 23, 5) {real, imag} */,
  {32'h3e8007d2, 32'h3e15ef53} /* (13, 23, 4) {real, imag} */,
  {32'hbd83cba6, 32'h3e327d54} /* (13, 23, 3) {real, imag} */,
  {32'hbf9083ed, 32'hbeb9a7bc} /* (13, 23, 2) {real, imag} */,
  {32'h40320657, 32'h3ee5cbde} /* (13, 23, 1) {real, imag} */,
  {32'h4002e690, 32'h00000000} /* (13, 23, 0) {real, imag} */,
  {32'h3ff6c0ec, 32'hbe811890} /* (13, 22, 31) {real, imag} */,
  {32'hbf317d09, 32'h3e1eb5ca} /* (13, 22, 30) {real, imag} */,
  {32'hbe008c1f, 32'hbdeef69c} /* (13, 22, 29) {real, imag} */,
  {32'h3e77b5eb, 32'hbe755a27} /* (13, 22, 28) {real, imag} */,
  {32'hbe54683b, 32'h3dec3032} /* (13, 22, 27) {real, imag} */,
  {32'hbd9e26ea, 32'h3d4ec6cc} /* (13, 22, 26) {real, imag} */,
  {32'h3b4357e8, 32'hbce58824} /* (13, 22, 25) {real, imag} */,
  {32'hbdb24034, 32'h3c68b7c0} /* (13, 22, 24) {real, imag} */,
  {32'hbd00df10, 32'h3cbc50f0} /* (13, 22, 23) {real, imag} */,
  {32'h3af4edd0, 32'hbd6e44d4} /* (13, 22, 22) {real, imag} */,
  {32'hbd695f02, 32'h3b0cbc30} /* (13, 22, 21) {real, imag} */,
  {32'hbd74e2cc, 32'hbcc1e116} /* (13, 22, 20) {real, imag} */,
  {32'hbd5185c8, 32'hbdbb204a} /* (13, 22, 19) {real, imag} */,
  {32'h3d16c0e6, 32'h3d13f586} /* (13, 22, 18) {real, imag} */,
  {32'h3d070778, 32'h3d85d717} /* (13, 22, 17) {real, imag} */,
  {32'hbc5bd7e6, 32'h00000000} /* (13, 22, 16) {real, imag} */,
  {32'h3d070778, 32'hbd85d717} /* (13, 22, 15) {real, imag} */,
  {32'h3d16c0e6, 32'hbd13f586} /* (13, 22, 14) {real, imag} */,
  {32'hbd5185c8, 32'h3dbb204a} /* (13, 22, 13) {real, imag} */,
  {32'hbd74e2cc, 32'h3cc1e116} /* (13, 22, 12) {real, imag} */,
  {32'hbd695f02, 32'hbb0cbc30} /* (13, 22, 11) {real, imag} */,
  {32'h3af4edd0, 32'h3d6e44d4} /* (13, 22, 10) {real, imag} */,
  {32'hbd00df10, 32'hbcbc50f0} /* (13, 22, 9) {real, imag} */,
  {32'hbdb24034, 32'hbc68b7c0} /* (13, 22, 8) {real, imag} */,
  {32'h3b4357e8, 32'h3ce58824} /* (13, 22, 7) {real, imag} */,
  {32'hbd9e26ea, 32'hbd4ec6cc} /* (13, 22, 6) {real, imag} */,
  {32'hbe54683b, 32'hbdec3032} /* (13, 22, 5) {real, imag} */,
  {32'h3e77b5eb, 32'h3e755a27} /* (13, 22, 4) {real, imag} */,
  {32'hbe008c1f, 32'h3deef69c} /* (13, 22, 3) {real, imag} */,
  {32'hbf317d09, 32'hbe1eb5ca} /* (13, 22, 2) {real, imag} */,
  {32'h3ff6c0ec, 32'h3e811890} /* (13, 22, 1) {real, imag} */,
  {32'h3fbf6c7d, 32'h00000000} /* (13, 22, 0) {real, imag} */,
  {32'h3f00e193, 32'h3d14c690} /* (13, 21, 31) {real, imag} */,
  {32'hbe4c8ffa, 32'h3d9c0b56} /* (13, 21, 30) {real, imag} */,
  {32'h3d80f310, 32'hbd929b34} /* (13, 21, 29) {real, imag} */,
  {32'h3e070504, 32'hbe081042} /* (13, 21, 28) {real, imag} */,
  {32'hbdb6e35e, 32'h3e1ebc2e} /* (13, 21, 27) {real, imag} */,
  {32'hbe011425, 32'hbcf7c973} /* (13, 21, 26) {real, imag} */,
  {32'h3d9f8a1d, 32'hbd840796} /* (13, 21, 25) {real, imag} */,
  {32'h3e2dddf4, 32'h3d01fd1f} /* (13, 21, 24) {real, imag} */,
  {32'hbda794de, 32'h3d3d7e70} /* (13, 21, 23) {real, imag} */,
  {32'hbd256dc2, 32'h3d1e84f7} /* (13, 21, 22) {real, imag} */,
  {32'h3cfa1087, 32'h3d1193f4} /* (13, 21, 21) {real, imag} */,
  {32'h3cd812a2, 32'hbd80beeb} /* (13, 21, 20) {real, imag} */,
  {32'h3d874389, 32'hbdaaf772} /* (13, 21, 19) {real, imag} */,
  {32'h3c8d453c, 32'hbd11c38f} /* (13, 21, 18) {real, imag} */,
  {32'hbcf50bf5, 32'h3de4e644} /* (13, 21, 17) {real, imag} */,
  {32'h3d771ea2, 32'h00000000} /* (13, 21, 16) {real, imag} */,
  {32'hbcf50bf5, 32'hbde4e644} /* (13, 21, 15) {real, imag} */,
  {32'h3c8d453c, 32'h3d11c38f} /* (13, 21, 14) {real, imag} */,
  {32'h3d874389, 32'h3daaf772} /* (13, 21, 13) {real, imag} */,
  {32'h3cd812a2, 32'h3d80beeb} /* (13, 21, 12) {real, imag} */,
  {32'h3cfa1087, 32'hbd1193f4} /* (13, 21, 11) {real, imag} */,
  {32'hbd256dc2, 32'hbd1e84f7} /* (13, 21, 10) {real, imag} */,
  {32'hbda794de, 32'hbd3d7e70} /* (13, 21, 9) {real, imag} */,
  {32'h3e2dddf4, 32'hbd01fd1f} /* (13, 21, 8) {real, imag} */,
  {32'h3d9f8a1d, 32'h3d840796} /* (13, 21, 7) {real, imag} */,
  {32'hbe011425, 32'h3cf7c973} /* (13, 21, 6) {real, imag} */,
  {32'hbdb6e35e, 32'hbe1ebc2e} /* (13, 21, 5) {real, imag} */,
  {32'h3e070504, 32'h3e081042} /* (13, 21, 4) {real, imag} */,
  {32'h3d80f310, 32'h3d929b34} /* (13, 21, 3) {real, imag} */,
  {32'hbe4c8ffa, 32'hbd9c0b56} /* (13, 21, 2) {real, imag} */,
  {32'h3f00e193, 32'hbd14c690} /* (13, 21, 1) {real, imag} */,
  {32'h3f1c3f21, 32'h00000000} /* (13, 21, 0) {real, imag} */,
  {32'hbf966038, 32'h3e1eabec} /* (13, 20, 31) {real, imag} */,
  {32'h3efaf4d0, 32'hbdc64c9a} /* (13, 20, 30) {real, imag} */,
  {32'h3d529b22, 32'hbd59efb3} /* (13, 20, 29) {real, imag} */,
  {32'h3cd3bf44, 32'h3c51e390} /* (13, 20, 28) {real, imag} */,
  {32'h3df31331, 32'hbdec32d0} /* (13, 20, 27) {real, imag} */,
  {32'hbdc617d4, 32'hbd36dcd9} /* (13, 20, 26) {real, imag} */,
  {32'h3ca90b80, 32'hbd5a1db7} /* (13, 20, 25) {real, imag} */,
  {32'h3d820d34, 32'hbc80045c} /* (13, 20, 24) {real, imag} */,
  {32'h3c9fe4c1, 32'h3d03d9a6} /* (13, 20, 23) {real, imag} */,
  {32'hbd16da4e, 32'h3c86eab4} /* (13, 20, 22) {real, imag} */,
  {32'h3dfc40b8, 32'h3a616b60} /* (13, 20, 21) {real, imag} */,
  {32'h3c39733d, 32'h3d66e60f} /* (13, 20, 20) {real, imag} */,
  {32'hbd380564, 32'hbd0bac25} /* (13, 20, 19) {real, imag} */,
  {32'h3c6dda82, 32'h3c644472} /* (13, 20, 18) {real, imag} */,
  {32'hbd7ced3b, 32'h3d725aff} /* (13, 20, 17) {real, imag} */,
  {32'hbd513a42, 32'h00000000} /* (13, 20, 16) {real, imag} */,
  {32'hbd7ced3b, 32'hbd725aff} /* (13, 20, 15) {real, imag} */,
  {32'h3c6dda82, 32'hbc644472} /* (13, 20, 14) {real, imag} */,
  {32'hbd380564, 32'h3d0bac25} /* (13, 20, 13) {real, imag} */,
  {32'h3c39733d, 32'hbd66e60f} /* (13, 20, 12) {real, imag} */,
  {32'h3dfc40b8, 32'hba616b60} /* (13, 20, 11) {real, imag} */,
  {32'hbd16da4e, 32'hbc86eab4} /* (13, 20, 10) {real, imag} */,
  {32'h3c9fe4c1, 32'hbd03d9a6} /* (13, 20, 9) {real, imag} */,
  {32'h3d820d34, 32'h3c80045c} /* (13, 20, 8) {real, imag} */,
  {32'h3ca90b80, 32'h3d5a1db7} /* (13, 20, 7) {real, imag} */,
  {32'hbdc617d4, 32'h3d36dcd9} /* (13, 20, 6) {real, imag} */,
  {32'h3df31331, 32'h3dec32d0} /* (13, 20, 5) {real, imag} */,
  {32'h3cd3bf44, 32'hbc51e390} /* (13, 20, 4) {real, imag} */,
  {32'h3d529b22, 32'h3d59efb3} /* (13, 20, 3) {real, imag} */,
  {32'h3efaf4d0, 32'h3dc64c9a} /* (13, 20, 2) {real, imag} */,
  {32'hbf966038, 32'hbe1eabec} /* (13, 20, 1) {real, imag} */,
  {32'hbf33eae2, 32'h00000000} /* (13, 20, 0) {real, imag} */,
  {32'hc0065280, 32'h3e8e7cc2} /* (13, 19, 31) {real, imag} */,
  {32'h3f71bcd4, 32'hbe0ed1c3} /* (13, 19, 30) {real, imag} */,
  {32'h3d0054a8, 32'hbc33cbec} /* (13, 19, 29) {real, imag} */,
  {32'hbd935e99, 32'h3e16cdaf} /* (13, 19, 28) {real, imag} */,
  {32'h3e5b5159, 32'hbe2d488a} /* (13, 19, 27) {real, imag} */,
  {32'h3c40f5a6, 32'hbe062c89} /* (13, 19, 26) {real, imag} */,
  {32'h3ba509e4, 32'h3cd02ab2} /* (13, 19, 25) {real, imag} */,
  {32'h3d4d7931, 32'hbd9793a8} /* (13, 19, 24) {real, imag} */,
  {32'h3b828e38, 32'h3de49cb8} /* (13, 19, 23) {real, imag} */,
  {32'hbd4c6bac, 32'hbdbd0a7f} /* (13, 19, 22) {real, imag} */,
  {32'h3d36d62a, 32'hbc1485c0} /* (13, 19, 21) {real, imag} */,
  {32'hbd13279e, 32'h3da3918e} /* (13, 19, 20) {real, imag} */,
  {32'hbd766db6, 32'h3c8be880} /* (13, 19, 19) {real, imag} */,
  {32'hbd05dc3d, 32'h3c83dd92} /* (13, 19, 18) {real, imag} */,
  {32'h3c84f8de, 32'hbba17b54} /* (13, 19, 17) {real, imag} */,
  {32'h3df0c498, 32'h00000000} /* (13, 19, 16) {real, imag} */,
  {32'h3c84f8de, 32'h3ba17b54} /* (13, 19, 15) {real, imag} */,
  {32'hbd05dc3d, 32'hbc83dd92} /* (13, 19, 14) {real, imag} */,
  {32'hbd766db6, 32'hbc8be880} /* (13, 19, 13) {real, imag} */,
  {32'hbd13279e, 32'hbda3918e} /* (13, 19, 12) {real, imag} */,
  {32'h3d36d62a, 32'h3c1485c0} /* (13, 19, 11) {real, imag} */,
  {32'hbd4c6bac, 32'h3dbd0a7f} /* (13, 19, 10) {real, imag} */,
  {32'h3b828e38, 32'hbde49cb8} /* (13, 19, 9) {real, imag} */,
  {32'h3d4d7931, 32'h3d9793a8} /* (13, 19, 8) {real, imag} */,
  {32'h3ba509e4, 32'hbcd02ab2} /* (13, 19, 7) {real, imag} */,
  {32'h3c40f5a6, 32'h3e062c89} /* (13, 19, 6) {real, imag} */,
  {32'h3e5b5159, 32'h3e2d488a} /* (13, 19, 5) {real, imag} */,
  {32'hbd935e99, 32'hbe16cdaf} /* (13, 19, 4) {real, imag} */,
  {32'h3d0054a8, 32'h3c33cbec} /* (13, 19, 3) {real, imag} */,
  {32'h3f71bcd4, 32'h3e0ed1c3} /* (13, 19, 2) {real, imag} */,
  {32'hc0065280, 32'hbe8e7cc2} /* (13, 19, 1) {real, imag} */,
  {32'hbfb4d430, 32'h00000000} /* (13, 19, 0) {real, imag} */,
  {32'hc028d5da, 32'h3eb9f0f8} /* (13, 18, 31) {real, imag} */,
  {32'h3f964f49, 32'hbeacde47} /* (13, 18, 30) {real, imag} */,
  {32'h3dc31369, 32'hbd8218d4} /* (13, 18, 29) {real, imag} */,
  {32'hbe133b25, 32'h3e2f01a8} /* (13, 18, 28) {real, imag} */,
  {32'h3e6b1034, 32'hbd23afa3} /* (13, 18, 27) {real, imag} */,
  {32'h3c189864, 32'hbcead3a8} /* (13, 18, 26) {real, imag} */,
  {32'hbd635674, 32'h3cc2ddd2} /* (13, 18, 25) {real, imag} */,
  {32'h3d357f70, 32'hbd9a3967} /* (13, 18, 24) {real, imag} */,
  {32'h3d6a2e8c, 32'hbb8173ae} /* (13, 18, 23) {real, imag} */,
  {32'h3da37dca, 32'hbbe86d50} /* (13, 18, 22) {real, imag} */,
  {32'hbd7d0868, 32'hbd8ab974} /* (13, 18, 21) {real, imag} */,
  {32'h3c1c9acc, 32'h3d8fef06} /* (13, 18, 20) {real, imag} */,
  {32'hbd6bfffc, 32'hbd4795d8} /* (13, 18, 19) {real, imag} */,
  {32'h3ca724a3, 32'hbd60189a} /* (13, 18, 18) {real, imag} */,
  {32'hbc932242, 32'h3d188ef3} /* (13, 18, 17) {real, imag} */,
  {32'hbdc6ed9e, 32'h00000000} /* (13, 18, 16) {real, imag} */,
  {32'hbc932242, 32'hbd188ef3} /* (13, 18, 15) {real, imag} */,
  {32'h3ca724a3, 32'h3d60189a} /* (13, 18, 14) {real, imag} */,
  {32'hbd6bfffc, 32'h3d4795d8} /* (13, 18, 13) {real, imag} */,
  {32'h3c1c9acc, 32'hbd8fef06} /* (13, 18, 12) {real, imag} */,
  {32'hbd7d0868, 32'h3d8ab974} /* (13, 18, 11) {real, imag} */,
  {32'h3da37dca, 32'h3be86d50} /* (13, 18, 10) {real, imag} */,
  {32'h3d6a2e8c, 32'h3b8173ae} /* (13, 18, 9) {real, imag} */,
  {32'h3d357f70, 32'h3d9a3967} /* (13, 18, 8) {real, imag} */,
  {32'hbd635674, 32'hbcc2ddd2} /* (13, 18, 7) {real, imag} */,
  {32'h3c189864, 32'h3cead3a8} /* (13, 18, 6) {real, imag} */,
  {32'h3e6b1034, 32'h3d23afa3} /* (13, 18, 5) {real, imag} */,
  {32'hbe133b25, 32'hbe2f01a8} /* (13, 18, 4) {real, imag} */,
  {32'h3dc31369, 32'h3d8218d4} /* (13, 18, 3) {real, imag} */,
  {32'h3f964f49, 32'h3eacde47} /* (13, 18, 2) {real, imag} */,
  {32'hc028d5da, 32'hbeb9f0f8} /* (13, 18, 1) {real, imag} */,
  {32'hc00392bc, 32'h00000000} /* (13, 18, 0) {real, imag} */,
  {32'hc042bccb, 32'h3ed1b05e} /* (13, 17, 31) {real, imag} */,
  {32'h3fad2e9e, 32'hbea89e34} /* (13, 17, 30) {real, imag} */,
  {32'h3de91d5e, 32'hbd7a0d72} /* (13, 17, 29) {real, imag} */,
  {32'hbe169be6, 32'h3e78a459} /* (13, 17, 28) {real, imag} */,
  {32'h3e659f9e, 32'hbd1c2f5e} /* (13, 17, 27) {real, imag} */,
  {32'h3d6efcc4, 32'hbdd778cf} /* (13, 17, 26) {real, imag} */,
  {32'hbdf66f89, 32'h3cb268d3} /* (13, 17, 25) {real, imag} */,
  {32'h3da56258, 32'hbd7ef44c} /* (13, 17, 24) {real, imag} */,
  {32'h3cc3d3a4, 32'hbd4b55e5} /* (13, 17, 23) {real, imag} */,
  {32'hbd9fbdeb, 32'hbda40ba8} /* (13, 17, 22) {real, imag} */,
  {32'hbd8b866c, 32'hbd5c348f} /* (13, 17, 21) {real, imag} */,
  {32'hbd52bea0, 32'hbd5e7f54} /* (13, 17, 20) {real, imag} */,
  {32'h3cc8da66, 32'hb9b0d9c0} /* (13, 17, 19) {real, imag} */,
  {32'h3dfdca50, 32'h3de9cb1b} /* (13, 17, 18) {real, imag} */,
  {32'h3d965c44, 32'hbc785234} /* (13, 17, 17) {real, imag} */,
  {32'hbd89af40, 32'h00000000} /* (13, 17, 16) {real, imag} */,
  {32'h3d965c44, 32'h3c785234} /* (13, 17, 15) {real, imag} */,
  {32'h3dfdca50, 32'hbde9cb1b} /* (13, 17, 14) {real, imag} */,
  {32'h3cc8da66, 32'h39b0d9c0} /* (13, 17, 13) {real, imag} */,
  {32'hbd52bea0, 32'h3d5e7f54} /* (13, 17, 12) {real, imag} */,
  {32'hbd8b866c, 32'h3d5c348f} /* (13, 17, 11) {real, imag} */,
  {32'hbd9fbdeb, 32'h3da40ba8} /* (13, 17, 10) {real, imag} */,
  {32'h3cc3d3a4, 32'h3d4b55e5} /* (13, 17, 9) {real, imag} */,
  {32'h3da56258, 32'h3d7ef44c} /* (13, 17, 8) {real, imag} */,
  {32'hbdf66f89, 32'hbcb268d3} /* (13, 17, 7) {real, imag} */,
  {32'h3d6efcc4, 32'h3dd778cf} /* (13, 17, 6) {real, imag} */,
  {32'h3e659f9e, 32'h3d1c2f5e} /* (13, 17, 5) {real, imag} */,
  {32'hbe169be6, 32'hbe78a459} /* (13, 17, 4) {real, imag} */,
  {32'h3de91d5e, 32'h3d7a0d72} /* (13, 17, 3) {real, imag} */,
  {32'h3fad2e9e, 32'h3ea89e34} /* (13, 17, 2) {real, imag} */,
  {32'hc042bccb, 32'hbed1b05e} /* (13, 17, 1) {real, imag} */,
  {32'hc0231140, 32'h00000000} /* (13, 17, 0) {real, imag} */,
  {32'hc0571582, 32'h3f132e0a} /* (13, 16, 31) {real, imag} */,
  {32'h3fb0a2e2, 32'hbe8bd41a} /* (13, 16, 30) {real, imag} */,
  {32'h3daa4e0b, 32'hbe00dec2} /* (13, 16, 29) {real, imag} */,
  {32'hbe2634ed, 32'h3e3d9ad6} /* (13, 16, 28) {real, imag} */,
  {32'h3e053d12, 32'hbde11dbe} /* (13, 16, 27) {real, imag} */,
  {32'h3d18473c, 32'hbd930017} /* (13, 16, 26) {real, imag} */,
  {32'hbe2e64d8, 32'h3bbd00d8} /* (13, 16, 25) {real, imag} */,
  {32'h3e1669ae, 32'hbd6244a9} /* (13, 16, 24) {real, imag} */,
  {32'hbb457690, 32'hbd35b6d2} /* (13, 16, 23) {real, imag} */,
  {32'hbd12b0c3, 32'h3cd06a02} /* (13, 16, 22) {real, imag} */,
  {32'h3db0372b, 32'hbbd7fd94} /* (13, 16, 21) {real, imag} */,
  {32'hbdc48528, 32'hbd9009e8} /* (13, 16, 20) {real, imag} */,
  {32'h3d140281, 32'h3cbcb255} /* (13, 16, 19) {real, imag} */,
  {32'hbc8f5cf4, 32'h3cd752b4} /* (13, 16, 18) {real, imag} */,
  {32'h3d372db8, 32'hbd998222} /* (13, 16, 17) {real, imag} */,
  {32'h3d082bce, 32'h00000000} /* (13, 16, 16) {real, imag} */,
  {32'h3d372db8, 32'h3d998222} /* (13, 16, 15) {real, imag} */,
  {32'hbc8f5cf4, 32'hbcd752b4} /* (13, 16, 14) {real, imag} */,
  {32'h3d140281, 32'hbcbcb255} /* (13, 16, 13) {real, imag} */,
  {32'hbdc48528, 32'h3d9009e8} /* (13, 16, 12) {real, imag} */,
  {32'h3db0372b, 32'h3bd7fd94} /* (13, 16, 11) {real, imag} */,
  {32'hbd12b0c3, 32'hbcd06a02} /* (13, 16, 10) {real, imag} */,
  {32'hbb457690, 32'h3d35b6d2} /* (13, 16, 9) {real, imag} */,
  {32'h3e1669ae, 32'h3d6244a9} /* (13, 16, 8) {real, imag} */,
  {32'hbe2e64d8, 32'hbbbd00d8} /* (13, 16, 7) {real, imag} */,
  {32'h3d18473c, 32'h3d930017} /* (13, 16, 6) {real, imag} */,
  {32'h3e053d12, 32'h3de11dbe} /* (13, 16, 5) {real, imag} */,
  {32'hbe2634ed, 32'hbe3d9ad6} /* (13, 16, 4) {real, imag} */,
  {32'h3daa4e0b, 32'h3e00dec2} /* (13, 16, 3) {real, imag} */,
  {32'h3fb0a2e2, 32'h3e8bd41a} /* (13, 16, 2) {real, imag} */,
  {32'hc0571582, 32'hbf132e0a} /* (13, 16, 1) {real, imag} */,
  {32'hc019f5e5, 32'h00000000} /* (13, 16, 0) {real, imag} */,
  {32'hc0600e19, 32'h3f0145df} /* (13, 15, 31) {real, imag} */,
  {32'h3f9b6bf8, 32'hbe6afe11} /* (13, 15, 30) {real, imag} */,
  {32'h3c8522e0, 32'h3c0efa58} /* (13, 15, 29) {real, imag} */,
  {32'hbe4934a6, 32'h3e60c6fb} /* (13, 15, 28) {real, imag} */,
  {32'h3dce1b44, 32'hbe81ef06} /* (13, 15, 27) {real, imag} */,
  {32'hbcd27a20, 32'hbe0c67d6} /* (13, 15, 26) {real, imag} */,
  {32'hbdaa65f1, 32'hbcc603cb} /* (13, 15, 25) {real, imag} */,
  {32'h3d377113, 32'hbd8fe7a2} /* (13, 15, 24) {real, imag} */,
  {32'hbcf295a8, 32'hbd09bc63} /* (13, 15, 23) {real, imag} */,
  {32'hbda18eab, 32'hba3d7dc0} /* (13, 15, 22) {real, imag} */,
  {32'h3c94fb46, 32'hbd4ec647} /* (13, 15, 21) {real, imag} */,
  {32'h3d2f911a, 32'h3bceb640} /* (13, 15, 20) {real, imag} */,
  {32'h3ddaeeb2, 32'hbbda1e24} /* (13, 15, 19) {real, imag} */,
  {32'hbd07d7a7, 32'h3c24b348} /* (13, 15, 18) {real, imag} */,
  {32'h3cc1cc18, 32'h3d6ea5cb} /* (13, 15, 17) {real, imag} */,
  {32'h3d431d18, 32'h00000000} /* (13, 15, 16) {real, imag} */,
  {32'h3cc1cc18, 32'hbd6ea5cb} /* (13, 15, 15) {real, imag} */,
  {32'hbd07d7a7, 32'hbc24b348} /* (13, 15, 14) {real, imag} */,
  {32'h3ddaeeb2, 32'h3bda1e24} /* (13, 15, 13) {real, imag} */,
  {32'h3d2f911a, 32'hbbceb640} /* (13, 15, 12) {real, imag} */,
  {32'h3c94fb46, 32'h3d4ec647} /* (13, 15, 11) {real, imag} */,
  {32'hbda18eab, 32'h3a3d7dc0} /* (13, 15, 10) {real, imag} */,
  {32'hbcf295a8, 32'h3d09bc63} /* (13, 15, 9) {real, imag} */,
  {32'h3d377113, 32'h3d8fe7a2} /* (13, 15, 8) {real, imag} */,
  {32'hbdaa65f1, 32'h3cc603cb} /* (13, 15, 7) {real, imag} */,
  {32'hbcd27a20, 32'h3e0c67d6} /* (13, 15, 6) {real, imag} */,
  {32'h3dce1b44, 32'h3e81ef06} /* (13, 15, 5) {real, imag} */,
  {32'hbe4934a6, 32'hbe60c6fb} /* (13, 15, 4) {real, imag} */,
  {32'h3c8522e0, 32'hbc0efa58} /* (13, 15, 3) {real, imag} */,
  {32'h3f9b6bf8, 32'h3e6afe11} /* (13, 15, 2) {real, imag} */,
  {32'hc0600e19, 32'hbf0145df} /* (13, 15, 1) {real, imag} */,
  {32'hc0201d42, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'hc051ba7e, 32'h3e813898} /* (13, 14, 31) {real, imag} */,
  {32'h3f839641, 32'hbe457762} /* (13, 14, 30) {real, imag} */,
  {32'h3c3c3e48, 32'hbce4a0ea} /* (13, 14, 29) {real, imag} */,
  {32'hbe14b843, 32'h3d807fd0} /* (13, 14, 28) {real, imag} */,
  {32'h3da6d26c, 32'hbdf14d76} /* (13, 14, 27) {real, imag} */,
  {32'h3b34c520, 32'hbe3bb03f} /* (13, 14, 26) {real, imag} */,
  {32'hbdfacc9e, 32'hbdaacad4} /* (13, 14, 25) {real, imag} */,
  {32'h3b57b9a0, 32'hbcc6fae8} /* (13, 14, 24) {real, imag} */,
  {32'hbd20d328, 32'h3c485a27} /* (13, 14, 23) {real, imag} */,
  {32'hbd6dfe05, 32'hbd97bd1d} /* (13, 14, 22) {real, imag} */,
  {32'hbdaa5e58, 32'h3c1a432c} /* (13, 14, 21) {real, imag} */,
  {32'h3dc633ac, 32'hbcb8b4ec} /* (13, 14, 20) {real, imag} */,
  {32'hbd83eff7, 32'hbcf7104c} /* (13, 14, 19) {real, imag} */,
  {32'hbbc02acc, 32'h3bd97790} /* (13, 14, 18) {real, imag} */,
  {32'hbca7668c, 32'h3cd67262} /* (13, 14, 17) {real, imag} */,
  {32'hbd6fa718, 32'h00000000} /* (13, 14, 16) {real, imag} */,
  {32'hbca7668c, 32'hbcd67262} /* (13, 14, 15) {real, imag} */,
  {32'hbbc02acc, 32'hbbd97790} /* (13, 14, 14) {real, imag} */,
  {32'hbd83eff7, 32'h3cf7104c} /* (13, 14, 13) {real, imag} */,
  {32'h3dc633ac, 32'h3cb8b4ec} /* (13, 14, 12) {real, imag} */,
  {32'hbdaa5e58, 32'hbc1a432c} /* (13, 14, 11) {real, imag} */,
  {32'hbd6dfe05, 32'h3d97bd1d} /* (13, 14, 10) {real, imag} */,
  {32'hbd20d328, 32'hbc485a27} /* (13, 14, 9) {real, imag} */,
  {32'h3b57b9a0, 32'h3cc6fae8} /* (13, 14, 8) {real, imag} */,
  {32'hbdfacc9e, 32'h3daacad4} /* (13, 14, 7) {real, imag} */,
  {32'h3b34c520, 32'h3e3bb03f} /* (13, 14, 6) {real, imag} */,
  {32'h3da6d26c, 32'h3df14d76} /* (13, 14, 5) {real, imag} */,
  {32'hbe14b843, 32'hbd807fd0} /* (13, 14, 4) {real, imag} */,
  {32'h3c3c3e48, 32'h3ce4a0ea} /* (13, 14, 3) {real, imag} */,
  {32'h3f839641, 32'h3e457762} /* (13, 14, 2) {real, imag} */,
  {32'hc051ba7e, 32'hbe813898} /* (13, 14, 1) {real, imag} */,
  {32'hc00f0074, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'hc033aec8, 32'h3e36a98c} /* (13, 13, 31) {real, imag} */,
  {32'h3f7c793e, 32'hbe0f8d31} /* (13, 13, 30) {real, imag} */,
  {32'h3d847450, 32'h3d93e452} /* (13, 13, 29) {real, imag} */,
  {32'hbe03b72c, 32'h3e06f499} /* (13, 13, 28) {real, imag} */,
  {32'h3d968b76, 32'hbdb9e43c} /* (13, 13, 27) {real, imag} */,
  {32'h3cb77b91, 32'hbdcea07e} /* (13, 13, 26) {real, imag} */,
  {32'h3cfaaad5, 32'h3acb99c8} /* (13, 13, 25) {real, imag} */,
  {32'hbd788a0b, 32'hbceddf67} /* (13, 13, 24) {real, imag} */,
  {32'h3d06295f, 32'h3d948eb8} /* (13, 13, 23) {real, imag} */,
  {32'hbcdd8e53, 32'hbd84092d} /* (13, 13, 22) {real, imag} */,
  {32'h3d3c3a04, 32'hbe026bf4} /* (13, 13, 21) {real, imag} */,
  {32'hbcc5e5fc, 32'h3c45a940} /* (13, 13, 20) {real, imag} */,
  {32'hbcf5c558, 32'h3cf21ac0} /* (13, 13, 19) {real, imag} */,
  {32'hbd4355af, 32'h3ca3dbe2} /* (13, 13, 18) {real, imag} */,
  {32'h3cec049a, 32'hbced5135} /* (13, 13, 17) {real, imag} */,
  {32'hbc99b4f2, 32'h00000000} /* (13, 13, 16) {real, imag} */,
  {32'h3cec049a, 32'h3ced5135} /* (13, 13, 15) {real, imag} */,
  {32'hbd4355af, 32'hbca3dbe2} /* (13, 13, 14) {real, imag} */,
  {32'hbcf5c558, 32'hbcf21ac0} /* (13, 13, 13) {real, imag} */,
  {32'hbcc5e5fc, 32'hbc45a940} /* (13, 13, 12) {real, imag} */,
  {32'h3d3c3a04, 32'h3e026bf4} /* (13, 13, 11) {real, imag} */,
  {32'hbcdd8e53, 32'h3d84092d} /* (13, 13, 10) {real, imag} */,
  {32'h3d06295f, 32'hbd948eb8} /* (13, 13, 9) {real, imag} */,
  {32'hbd788a0b, 32'h3ceddf67} /* (13, 13, 8) {real, imag} */,
  {32'h3cfaaad5, 32'hbacb99c8} /* (13, 13, 7) {real, imag} */,
  {32'h3cb77b91, 32'h3dcea07e} /* (13, 13, 6) {real, imag} */,
  {32'h3d968b76, 32'h3db9e43c} /* (13, 13, 5) {real, imag} */,
  {32'hbe03b72c, 32'hbe06f499} /* (13, 13, 4) {real, imag} */,
  {32'h3d847450, 32'hbd93e452} /* (13, 13, 3) {real, imag} */,
  {32'h3f7c793e, 32'h3e0f8d31} /* (13, 13, 2) {real, imag} */,
  {32'hc033aec8, 32'hbe36a98c} /* (13, 13, 1) {real, imag} */,
  {32'hbfe0a9a2, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'hc0112cee, 32'h3d4229b0} /* (13, 12, 31) {real, imag} */,
  {32'h3f4aa16a, 32'h3c1a2190} /* (13, 12, 30) {real, imag} */,
  {32'h3dfbe731, 32'h3d212043} /* (13, 12, 29) {real, imag} */,
  {32'hbe281aae, 32'h3e8e8584} /* (13, 12, 28) {real, imag} */,
  {32'h3e7a9bd6, 32'hbdf5c150} /* (13, 12, 27) {real, imag} */,
  {32'h3de7dbfe, 32'hbddd8428} /* (13, 12, 26) {real, imag} */,
  {32'hbc9a5d58, 32'h3cc4e8da} /* (13, 12, 25) {real, imag} */,
  {32'h3daca27a, 32'hbe660848} /* (13, 12, 24) {real, imag} */,
  {32'hbd6d1090, 32'h3df9917f} /* (13, 12, 23) {real, imag} */,
  {32'hbcd88568, 32'hbc3e289a} /* (13, 12, 22) {real, imag} */,
  {32'h3c444d60, 32'h3cc10fe6} /* (13, 12, 21) {real, imag} */,
  {32'h3caf70f6, 32'h3dbc5cf4} /* (13, 12, 20) {real, imag} */,
  {32'hbd617f84, 32'hbcf5aa52} /* (13, 12, 19) {real, imag} */,
  {32'hbd4199c2, 32'hbc5755de} /* (13, 12, 18) {real, imag} */,
  {32'h3d804114, 32'hbd48552f} /* (13, 12, 17) {real, imag} */,
  {32'h3c6c656a, 32'h00000000} /* (13, 12, 16) {real, imag} */,
  {32'h3d804114, 32'h3d48552f} /* (13, 12, 15) {real, imag} */,
  {32'hbd4199c2, 32'h3c5755de} /* (13, 12, 14) {real, imag} */,
  {32'hbd617f84, 32'h3cf5aa52} /* (13, 12, 13) {real, imag} */,
  {32'h3caf70f6, 32'hbdbc5cf4} /* (13, 12, 12) {real, imag} */,
  {32'h3c444d60, 32'hbcc10fe6} /* (13, 12, 11) {real, imag} */,
  {32'hbcd88568, 32'h3c3e289a} /* (13, 12, 10) {real, imag} */,
  {32'hbd6d1090, 32'hbdf9917f} /* (13, 12, 9) {real, imag} */,
  {32'h3daca27a, 32'h3e660848} /* (13, 12, 8) {real, imag} */,
  {32'hbc9a5d58, 32'hbcc4e8da} /* (13, 12, 7) {real, imag} */,
  {32'h3de7dbfe, 32'h3ddd8428} /* (13, 12, 6) {real, imag} */,
  {32'h3e7a9bd6, 32'h3df5c150} /* (13, 12, 5) {real, imag} */,
  {32'hbe281aae, 32'hbe8e8584} /* (13, 12, 4) {real, imag} */,
  {32'h3dfbe731, 32'hbd212043} /* (13, 12, 3) {real, imag} */,
  {32'h3f4aa16a, 32'hbc1a2190} /* (13, 12, 2) {real, imag} */,
  {32'hc0112cee, 32'hbd4229b0} /* (13, 12, 1) {real, imag} */,
  {32'hbf8607fd, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'hbfa00a02, 32'hbe52bcb4} /* (13, 11, 31) {real, imag} */,
  {32'h3f0e621e, 32'hbcdcac58} /* (13, 11, 30) {real, imag} */,
  {32'h3daead44, 32'h3d93d19c} /* (13, 11, 29) {real, imag} */,
  {32'hbdcb7a57, 32'h3e227f78} /* (13, 11, 28) {real, imag} */,
  {32'h3d48e170, 32'hbe1973ac} /* (13, 11, 27) {real, imag} */,
  {32'h3d5de284, 32'h3d3b5646} /* (13, 11, 26) {real, imag} */,
  {32'hbdba5231, 32'hbe09c449} /* (13, 11, 25) {real, imag} */,
  {32'h3d973328, 32'h3d217d5d} /* (13, 11, 24) {real, imag} */,
  {32'h3cadf052, 32'h3dd71394} /* (13, 11, 23) {real, imag} */,
  {32'hbdb0e89f, 32'h3dac127c} /* (13, 11, 22) {real, imag} */,
  {32'hbd8e315e, 32'hbd9097a4} /* (13, 11, 21) {real, imag} */,
  {32'h3d1c5ecb, 32'hbc5ab03a} /* (13, 11, 20) {real, imag} */,
  {32'h3d93a6dd, 32'hbd843cb8} /* (13, 11, 19) {real, imag} */,
  {32'h3d04b3fa, 32'hbd9be80a} /* (13, 11, 18) {real, imag} */,
  {32'hbd3da60e, 32'h3c71f660} /* (13, 11, 17) {real, imag} */,
  {32'hbdc2ac4b, 32'h00000000} /* (13, 11, 16) {real, imag} */,
  {32'hbd3da60e, 32'hbc71f660} /* (13, 11, 15) {real, imag} */,
  {32'h3d04b3fa, 32'h3d9be80a} /* (13, 11, 14) {real, imag} */,
  {32'h3d93a6dd, 32'h3d843cb8} /* (13, 11, 13) {real, imag} */,
  {32'h3d1c5ecb, 32'h3c5ab03a} /* (13, 11, 12) {real, imag} */,
  {32'hbd8e315e, 32'h3d9097a4} /* (13, 11, 11) {real, imag} */,
  {32'hbdb0e89f, 32'hbdac127c} /* (13, 11, 10) {real, imag} */,
  {32'h3cadf052, 32'hbdd71394} /* (13, 11, 9) {real, imag} */,
  {32'h3d973328, 32'hbd217d5d} /* (13, 11, 8) {real, imag} */,
  {32'hbdba5231, 32'h3e09c449} /* (13, 11, 7) {real, imag} */,
  {32'h3d5de284, 32'hbd3b5646} /* (13, 11, 6) {real, imag} */,
  {32'h3d48e170, 32'h3e1973ac} /* (13, 11, 5) {real, imag} */,
  {32'hbdcb7a57, 32'hbe227f78} /* (13, 11, 4) {real, imag} */,
  {32'h3daead44, 32'hbd93d19c} /* (13, 11, 3) {real, imag} */,
  {32'h3f0e621e, 32'h3cdcac58} /* (13, 11, 2) {real, imag} */,
  {32'hbfa00a02, 32'h3e52bcb4} /* (13, 11, 1) {real, imag} */,
  {32'hbe50bd94, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'h3ef2d436, 32'hbee52bb4} /* (13, 10, 31) {real, imag} */,
  {32'h3d6c8090, 32'hbc1300e0} /* (13, 10, 30) {real, imag} */,
  {32'hbdcd52ae, 32'hbcb92d46} /* (13, 10, 29) {real, imag} */,
  {32'h3cede728, 32'hbd9d4182} /* (13, 10, 28) {real, imag} */,
  {32'hbdcaa302, 32'hbd112e0c} /* (13, 10, 27) {real, imag} */,
  {32'hbdb0893a, 32'h3d6265f0} /* (13, 10, 26) {real, imag} */,
  {32'h3d0fd926, 32'hbdba83a7} /* (13, 10, 25) {real, imag} */,
  {32'hbd0c10a0, 32'h3d7f5894} /* (13, 10, 24) {real, imag} */,
  {32'h3a57bb00, 32'hbe25ee10} /* (13, 10, 23) {real, imag} */,
  {32'h3ca8f99f, 32'h3c8205ab} /* (13, 10, 22) {real, imag} */,
  {32'hbdbe73b3, 32'hbd7bef8f} /* (13, 10, 21) {real, imag} */,
  {32'hbda900aa, 32'h3d3aee4d} /* (13, 10, 20) {real, imag} */,
  {32'h3cbeaef9, 32'hbc8697b2} /* (13, 10, 19) {real, imag} */,
  {32'hbddd5171, 32'h3d7fdcb4} /* (13, 10, 18) {real, imag} */,
  {32'h3d40eaec, 32'h3da1b1df} /* (13, 10, 17) {real, imag} */,
  {32'hbc10f4b6, 32'h00000000} /* (13, 10, 16) {real, imag} */,
  {32'h3d40eaec, 32'hbda1b1df} /* (13, 10, 15) {real, imag} */,
  {32'hbddd5171, 32'hbd7fdcb4} /* (13, 10, 14) {real, imag} */,
  {32'h3cbeaef9, 32'h3c8697b2} /* (13, 10, 13) {real, imag} */,
  {32'hbda900aa, 32'hbd3aee4d} /* (13, 10, 12) {real, imag} */,
  {32'hbdbe73b3, 32'h3d7bef8f} /* (13, 10, 11) {real, imag} */,
  {32'h3ca8f99f, 32'hbc8205ab} /* (13, 10, 10) {real, imag} */,
  {32'h3a57bb00, 32'h3e25ee10} /* (13, 10, 9) {real, imag} */,
  {32'hbd0c10a0, 32'hbd7f5894} /* (13, 10, 8) {real, imag} */,
  {32'h3d0fd926, 32'h3dba83a7} /* (13, 10, 7) {real, imag} */,
  {32'hbdb0893a, 32'hbd6265f0} /* (13, 10, 6) {real, imag} */,
  {32'hbdcaa302, 32'h3d112e0c} /* (13, 10, 5) {real, imag} */,
  {32'h3cede728, 32'h3d9d4182} /* (13, 10, 4) {real, imag} */,
  {32'hbdcd52ae, 32'h3cb92d46} /* (13, 10, 3) {real, imag} */,
  {32'h3d6c8090, 32'h3c1300e0} /* (13, 10, 2) {real, imag} */,
  {32'h3ef2d436, 32'h3ee52bb4} /* (13, 10, 1) {real, imag} */,
  {32'h3f83f277, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h3fc99f1e, 32'hbf2b5b13} /* (13, 9, 31) {real, imag} */,
  {32'hbf311026, 32'h3e8ca72c} /* (13, 9, 30) {real, imag} */,
  {32'hbda50862, 32'h3caefd5c} /* (13, 9, 29) {real, imag} */,
  {32'h3d164af2, 32'h3cc561d8} /* (13, 9, 28) {real, imag} */,
  {32'hbda9b058, 32'h3d43fea8} /* (13, 9, 27) {real, imag} */,
  {32'h3bd47ea8, 32'hbb94a704} /* (13, 9, 26) {real, imag} */,
  {32'h3d9ae296, 32'h3d50a77e} /* (13, 9, 25) {real, imag} */,
  {32'h3d819444, 32'h3cf2a8e8} /* (13, 9, 24) {real, imag} */,
  {32'h3c013244, 32'h3b7f19b0} /* (13, 9, 23) {real, imag} */,
  {32'hbc95868e, 32'hbd620c2b} /* (13, 9, 22) {real, imag} */,
  {32'hbdf772a8, 32'h3dfc0f0e} /* (13, 9, 21) {real, imag} */,
  {32'h3d148d92, 32'hbdc8cca0} /* (13, 9, 20) {real, imag} */,
  {32'h3e103c51, 32'hbcd4a0bc} /* (13, 9, 19) {real, imag} */,
  {32'hbdaa03d1, 32'h3d9ed6db} /* (13, 9, 18) {real, imag} */,
  {32'h3dbd44d0, 32'h3d1a07da} /* (13, 9, 17) {real, imag} */,
  {32'hbdc249b9, 32'h00000000} /* (13, 9, 16) {real, imag} */,
  {32'h3dbd44d0, 32'hbd1a07da} /* (13, 9, 15) {real, imag} */,
  {32'hbdaa03d1, 32'hbd9ed6db} /* (13, 9, 14) {real, imag} */,
  {32'h3e103c51, 32'h3cd4a0bc} /* (13, 9, 13) {real, imag} */,
  {32'h3d148d92, 32'h3dc8cca0} /* (13, 9, 12) {real, imag} */,
  {32'hbdf772a8, 32'hbdfc0f0e} /* (13, 9, 11) {real, imag} */,
  {32'hbc95868e, 32'h3d620c2b} /* (13, 9, 10) {real, imag} */,
  {32'h3c013244, 32'hbb7f19b0} /* (13, 9, 9) {real, imag} */,
  {32'h3d819444, 32'hbcf2a8e8} /* (13, 9, 8) {real, imag} */,
  {32'h3d9ae296, 32'hbd50a77e} /* (13, 9, 7) {real, imag} */,
  {32'h3bd47ea8, 32'h3b94a704} /* (13, 9, 6) {real, imag} */,
  {32'hbda9b058, 32'hbd43fea8} /* (13, 9, 5) {real, imag} */,
  {32'h3d164af2, 32'hbcc561d8} /* (13, 9, 4) {real, imag} */,
  {32'hbda50862, 32'hbcaefd5c} /* (13, 9, 3) {real, imag} */,
  {32'hbf311026, 32'hbe8ca72c} /* (13, 9, 2) {real, imag} */,
  {32'h3fc99f1e, 32'h3f2b5b13} /* (13, 9, 1) {real, imag} */,
  {32'h3ff6d6b0, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'h4009b4e7, 32'hbf52f380} /* (13, 8, 31) {real, imag} */,
  {32'hbf56ed5e, 32'h3ee9d665} /* (13, 8, 30) {real, imag} */,
  {32'hbdb50594, 32'h3d02408e} /* (13, 8, 29) {real, imag} */,
  {32'h3e038ce6, 32'h3c7b9ee4} /* (13, 8, 28) {real, imag} */,
  {32'hbda8c523, 32'h3daf28d2} /* (13, 8, 27) {real, imag} */,
  {32'hbd17ab99, 32'h3d779ea8} /* (13, 8, 26) {real, imag} */,
  {32'h3c4293c4, 32'hbdc8a8c7} /* (13, 8, 25) {real, imag} */,
  {32'hbc916c78, 32'h3d86b3c9} /* (13, 8, 24) {real, imag} */,
  {32'hbda79dda, 32'hbde77c3a} /* (13, 8, 23) {real, imag} */,
  {32'hbdbdcb37, 32'hbcb93d37} /* (13, 8, 22) {real, imag} */,
  {32'hbc5dcd48, 32'h3d69ecb0} /* (13, 8, 21) {real, imag} */,
  {32'hbce9ab98, 32'hbd535447} /* (13, 8, 20) {real, imag} */,
  {32'h3d08ec76, 32'hbc8c137a} /* (13, 8, 19) {real, imag} */,
  {32'h3d21b9e4, 32'hbb5a9988} /* (13, 8, 18) {real, imag} */,
  {32'h3c426c48, 32'h3cd5430b} /* (13, 8, 17) {real, imag} */,
  {32'h3cf13f36, 32'h00000000} /* (13, 8, 16) {real, imag} */,
  {32'h3c426c48, 32'hbcd5430b} /* (13, 8, 15) {real, imag} */,
  {32'h3d21b9e4, 32'h3b5a9988} /* (13, 8, 14) {real, imag} */,
  {32'h3d08ec76, 32'h3c8c137a} /* (13, 8, 13) {real, imag} */,
  {32'hbce9ab98, 32'h3d535447} /* (13, 8, 12) {real, imag} */,
  {32'hbc5dcd48, 32'hbd69ecb0} /* (13, 8, 11) {real, imag} */,
  {32'hbdbdcb37, 32'h3cb93d37} /* (13, 8, 10) {real, imag} */,
  {32'hbda79dda, 32'h3de77c3a} /* (13, 8, 9) {real, imag} */,
  {32'hbc916c78, 32'hbd86b3c9} /* (13, 8, 8) {real, imag} */,
  {32'h3c4293c4, 32'h3dc8a8c7} /* (13, 8, 7) {real, imag} */,
  {32'hbd17ab99, 32'hbd779ea8} /* (13, 8, 6) {real, imag} */,
  {32'hbda8c523, 32'hbdaf28d2} /* (13, 8, 5) {real, imag} */,
  {32'h3e038ce6, 32'hbc7b9ee4} /* (13, 8, 4) {real, imag} */,
  {32'hbdb50594, 32'hbd02408e} /* (13, 8, 3) {real, imag} */,
  {32'hbf56ed5e, 32'hbee9d665} /* (13, 8, 2) {real, imag} */,
  {32'h4009b4e7, 32'h3f52f380} /* (13, 8, 1) {real, imag} */,
  {32'h40216ccc, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'h402068e2, 32'hbf92fb18} /* (13, 7, 31) {real, imag} */,
  {32'hbf672d8c, 32'h3f1fc6a2} /* (13, 7, 30) {real, imag} */,
  {32'hbe1398e4, 32'h3e13a6bc} /* (13, 7, 29) {real, imag} */,
  {32'h3e56d473, 32'hbe1acee6} /* (13, 7, 28) {real, imag} */,
  {32'hbe46aa70, 32'h3de804d0} /* (13, 7, 27) {real, imag} */,
  {32'hbd269f70, 32'h3e198cb0} /* (13, 7, 26) {real, imag} */,
  {32'h3d963921, 32'hbdee5ab5} /* (13, 7, 25) {real, imag} */,
  {32'hbdfad5db, 32'hbc117fcc} /* (13, 7, 24) {real, imag} */,
  {32'hbc210aac, 32'h3b568f10} /* (13, 7, 23) {real, imag} */,
  {32'h3da08e80, 32'h3b837908} /* (13, 7, 22) {real, imag} */,
  {32'hbdf8ba2e, 32'h3e262ab2} /* (13, 7, 21) {real, imag} */,
  {32'hbc5edd4a, 32'hbd753cd7} /* (13, 7, 20) {real, imag} */,
  {32'hbc95a992, 32'hbd9b1eb1} /* (13, 7, 19) {real, imag} */,
  {32'hbb790018, 32'h3d00d682} /* (13, 7, 18) {real, imag} */,
  {32'hbbe8bbf0, 32'h3d953000} /* (13, 7, 17) {real, imag} */,
  {32'h3d11d12a, 32'h00000000} /* (13, 7, 16) {real, imag} */,
  {32'hbbe8bbf0, 32'hbd953000} /* (13, 7, 15) {real, imag} */,
  {32'hbb790018, 32'hbd00d682} /* (13, 7, 14) {real, imag} */,
  {32'hbc95a992, 32'h3d9b1eb1} /* (13, 7, 13) {real, imag} */,
  {32'hbc5edd4a, 32'h3d753cd7} /* (13, 7, 12) {real, imag} */,
  {32'hbdf8ba2e, 32'hbe262ab2} /* (13, 7, 11) {real, imag} */,
  {32'h3da08e80, 32'hbb837908} /* (13, 7, 10) {real, imag} */,
  {32'hbc210aac, 32'hbb568f10} /* (13, 7, 9) {real, imag} */,
  {32'hbdfad5db, 32'h3c117fcc} /* (13, 7, 8) {real, imag} */,
  {32'h3d963921, 32'h3dee5ab5} /* (13, 7, 7) {real, imag} */,
  {32'hbd269f70, 32'hbe198cb0} /* (13, 7, 6) {real, imag} */,
  {32'hbe46aa70, 32'hbde804d0} /* (13, 7, 5) {real, imag} */,
  {32'h3e56d473, 32'h3e1acee6} /* (13, 7, 4) {real, imag} */,
  {32'hbe1398e4, 32'hbe13a6bc} /* (13, 7, 3) {real, imag} */,
  {32'hbf672d8c, 32'hbf1fc6a2} /* (13, 7, 2) {real, imag} */,
  {32'h402068e2, 32'h3f92fb18} /* (13, 7, 1) {real, imag} */,
  {32'h403d0a14, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'h4022b7fa, 32'hbfd1e92e} /* (13, 6, 31) {real, imag} */,
  {32'hbf442454, 32'h3f2d64c8} /* (13, 6, 30) {real, imag} */,
  {32'hbde9a58a, 32'h3dc5702a} /* (13, 6, 29) {real, imag} */,
  {32'h3d8a18d2, 32'hbdfe6a62} /* (13, 6, 28) {real, imag} */,
  {32'hbe2c7636, 32'h3e202db7} /* (13, 6, 27) {real, imag} */,
  {32'h3d990362, 32'h3cee17dd} /* (13, 6, 26) {real, imag} */,
  {32'h3cc614b5, 32'hbcddffaa} /* (13, 6, 25) {real, imag} */,
  {32'hbcb6b30c, 32'h3c08a008} /* (13, 6, 24) {real, imag} */,
  {32'h3dba350a, 32'hbcdeb4c3} /* (13, 6, 23) {real, imag} */,
  {32'hbc660b2c, 32'hbd62c020} /* (13, 6, 22) {real, imag} */,
  {32'hbdb36d8a, 32'h3d2ebc56} /* (13, 6, 21) {real, imag} */,
  {32'hbd1797fc, 32'h3d8cd5dc} /* (13, 6, 20) {real, imag} */,
  {32'hbc81bbd5, 32'hbd01b1f8} /* (13, 6, 19) {real, imag} */,
  {32'h3c8adbed, 32'hbd01e4a4} /* (13, 6, 18) {real, imag} */,
  {32'h3c074ad8, 32'hbd929c61} /* (13, 6, 17) {real, imag} */,
  {32'h3cdcf287, 32'h00000000} /* (13, 6, 16) {real, imag} */,
  {32'h3c074ad8, 32'h3d929c61} /* (13, 6, 15) {real, imag} */,
  {32'h3c8adbed, 32'h3d01e4a4} /* (13, 6, 14) {real, imag} */,
  {32'hbc81bbd5, 32'h3d01b1f8} /* (13, 6, 13) {real, imag} */,
  {32'hbd1797fc, 32'hbd8cd5dc} /* (13, 6, 12) {real, imag} */,
  {32'hbdb36d8a, 32'hbd2ebc56} /* (13, 6, 11) {real, imag} */,
  {32'hbc660b2c, 32'h3d62c020} /* (13, 6, 10) {real, imag} */,
  {32'h3dba350a, 32'h3cdeb4c3} /* (13, 6, 9) {real, imag} */,
  {32'hbcb6b30c, 32'hbc08a008} /* (13, 6, 8) {real, imag} */,
  {32'h3cc614b5, 32'h3cddffaa} /* (13, 6, 7) {real, imag} */,
  {32'h3d990362, 32'hbcee17dd} /* (13, 6, 6) {real, imag} */,
  {32'hbe2c7636, 32'hbe202db7} /* (13, 6, 5) {real, imag} */,
  {32'h3d8a18d2, 32'h3dfe6a62} /* (13, 6, 4) {real, imag} */,
  {32'hbde9a58a, 32'hbdc5702a} /* (13, 6, 3) {real, imag} */,
  {32'hbf442454, 32'hbf2d64c8} /* (13, 6, 2) {real, imag} */,
  {32'h4022b7fa, 32'h3fd1e92e} /* (13, 6, 1) {real, imag} */,
  {32'h40571d72, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'h401b783c, 32'hc013e397} /* (13, 5, 31) {real, imag} */,
  {32'hbe3a40d8, 32'h3f5234ff} /* (13, 5, 30) {real, imag} */,
  {32'hbe0bb87a, 32'h3d53be3a} /* (13, 5, 29) {real, imag} */,
  {32'hbe05fe5d, 32'h3d8f0591} /* (13, 5, 28) {real, imag} */,
  {32'hbe4641ab, 32'hbc8c2a8c} /* (13, 5, 27) {real, imag} */,
  {32'h3e12ee3b, 32'h3c22eb4f} /* (13, 5, 26) {real, imag} */,
  {32'hbd05b59c, 32'hbdcf5146} /* (13, 5, 25) {real, imag} */,
  {32'hbc0ae21c, 32'h3e15cd25} /* (13, 5, 24) {real, imag} */,
  {32'hbd827a76, 32'hbd416b2a} /* (13, 5, 23) {real, imag} */,
  {32'hbcf46296, 32'h3ccdb22a} /* (13, 5, 22) {real, imag} */,
  {32'h3ba7f000, 32'h3cbcc153} /* (13, 5, 21) {real, imag} */,
  {32'h3d5ca67c, 32'h3ce70e5c} /* (13, 5, 20) {real, imag} */,
  {32'h3d0bc30c, 32'hbba8b360} /* (13, 5, 19) {real, imag} */,
  {32'hbd4464f9, 32'h3c72f81d} /* (13, 5, 18) {real, imag} */,
  {32'h3cbaf0db, 32'hbd1106b6} /* (13, 5, 17) {real, imag} */,
  {32'hbe0e8202, 32'h00000000} /* (13, 5, 16) {real, imag} */,
  {32'h3cbaf0db, 32'h3d1106b6} /* (13, 5, 15) {real, imag} */,
  {32'hbd4464f9, 32'hbc72f81d} /* (13, 5, 14) {real, imag} */,
  {32'h3d0bc30c, 32'h3ba8b360} /* (13, 5, 13) {real, imag} */,
  {32'h3d5ca67c, 32'hbce70e5c} /* (13, 5, 12) {real, imag} */,
  {32'h3ba7f000, 32'hbcbcc153} /* (13, 5, 11) {real, imag} */,
  {32'hbcf46296, 32'hbccdb22a} /* (13, 5, 10) {real, imag} */,
  {32'hbd827a76, 32'h3d416b2a} /* (13, 5, 9) {real, imag} */,
  {32'hbc0ae21c, 32'hbe15cd25} /* (13, 5, 8) {real, imag} */,
  {32'hbd05b59c, 32'h3dcf5146} /* (13, 5, 7) {real, imag} */,
  {32'h3e12ee3b, 32'hbc22eb4f} /* (13, 5, 6) {real, imag} */,
  {32'hbe4641ab, 32'h3c8c2a8c} /* (13, 5, 5) {real, imag} */,
  {32'hbe05fe5d, 32'hbd8f0591} /* (13, 5, 4) {real, imag} */,
  {32'hbe0bb87a, 32'hbd53be3a} /* (13, 5, 3) {real, imag} */,
  {32'hbe3a40d8, 32'hbf5234ff} /* (13, 5, 2) {real, imag} */,
  {32'h401b783c, 32'h4013e397} /* (13, 5, 1) {real, imag} */,
  {32'h406c3f1f, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h400e485a, 32'hc03b300e} /* (13, 4, 31) {real, imag} */,
  {32'h3dfe2590, 32'h3f8a3ed4} /* (13, 4, 30) {real, imag} */,
  {32'hbd6820a0, 32'h3dca6ca4} /* (13, 4, 29) {real, imag} */,
  {32'hbe2aed44, 32'h3d669064} /* (13, 4, 28) {real, imag} */,
  {32'hbe8067aa, 32'hbda390a6} /* (13, 4, 27) {real, imag} */,
  {32'h3dd37ca1, 32'h3db7cc38} /* (13, 4, 26) {real, imag} */,
  {32'hbdb8b890, 32'hbdccd902} /* (13, 4, 25) {real, imag} */,
  {32'h3cf5cec9, 32'h3daf3f3b} /* (13, 4, 24) {real, imag} */,
  {32'hbcfd8574, 32'h3c9537b5} /* (13, 4, 23) {real, imag} */,
  {32'hbcb7a222, 32'h3c8d68c4} /* (13, 4, 22) {real, imag} */,
  {32'hbcd68a2f, 32'hbd26e0ad} /* (13, 4, 21) {real, imag} */,
  {32'h3d89e5d8, 32'hbd46b407} /* (13, 4, 20) {real, imag} */,
  {32'hbd456a5f, 32'h3ce335c0} /* (13, 4, 19) {real, imag} */,
  {32'h3d60f924, 32'hbd64e228} /* (13, 4, 18) {real, imag} */,
  {32'hbc9c0b65, 32'h3cf79544} /* (13, 4, 17) {real, imag} */,
  {32'hbd8b682f, 32'h00000000} /* (13, 4, 16) {real, imag} */,
  {32'hbc9c0b65, 32'hbcf79544} /* (13, 4, 15) {real, imag} */,
  {32'h3d60f924, 32'h3d64e228} /* (13, 4, 14) {real, imag} */,
  {32'hbd456a5f, 32'hbce335c0} /* (13, 4, 13) {real, imag} */,
  {32'h3d89e5d8, 32'h3d46b407} /* (13, 4, 12) {real, imag} */,
  {32'hbcd68a2f, 32'h3d26e0ad} /* (13, 4, 11) {real, imag} */,
  {32'hbcb7a222, 32'hbc8d68c4} /* (13, 4, 10) {real, imag} */,
  {32'hbcfd8574, 32'hbc9537b5} /* (13, 4, 9) {real, imag} */,
  {32'h3cf5cec9, 32'hbdaf3f3b} /* (13, 4, 8) {real, imag} */,
  {32'hbdb8b890, 32'h3dccd902} /* (13, 4, 7) {real, imag} */,
  {32'h3dd37ca1, 32'hbdb7cc38} /* (13, 4, 6) {real, imag} */,
  {32'hbe8067aa, 32'h3da390a6} /* (13, 4, 5) {real, imag} */,
  {32'hbe2aed44, 32'hbd669064} /* (13, 4, 4) {real, imag} */,
  {32'hbd6820a0, 32'hbdca6ca4} /* (13, 4, 3) {real, imag} */,
  {32'h3dfe2590, 32'hbf8a3ed4} /* (13, 4, 2) {real, imag} */,
  {32'h400e485a, 32'h403b300e} /* (13, 4, 1) {real, imag} */,
  {32'h40822e7f, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'h4016776d, 32'hc04611c2} /* (13, 3, 31) {real, imag} */,
  {32'h3dafdb30, 32'h3f866c82} /* (13, 3, 30) {real, imag} */,
  {32'hbe76639f, 32'h3e1d58f3} /* (13, 3, 29) {real, imag} */,
  {32'hbd7f020f, 32'h3da90fd7} /* (13, 3, 28) {real, imag} */,
  {32'hbe1b40df, 32'hbd9be44e} /* (13, 3, 27) {real, imag} */,
  {32'h3c9a7710, 32'h3c6f3130} /* (13, 3, 26) {real, imag} */,
  {32'h3d80adb9, 32'hbdba4074} /* (13, 3, 25) {real, imag} */,
  {32'h3deab7b0, 32'h3cadc308} /* (13, 3, 24) {real, imag} */,
  {32'h3d82bb4b, 32'hbdb0459e} /* (13, 3, 23) {real, imag} */,
  {32'hbd3f4619, 32'h3d19e218} /* (13, 3, 22) {real, imag} */,
  {32'hbd15ca34, 32'h3e0327a1} /* (13, 3, 21) {real, imag} */,
  {32'hbd1ba82c, 32'hbd05c600} /* (13, 3, 20) {real, imag} */,
  {32'h3d9a7e5a, 32'hbd292563} /* (13, 3, 19) {real, imag} */,
  {32'hbda41618, 32'h3dae9c3a} /* (13, 3, 18) {real, imag} */,
  {32'h3c937db2, 32'hbd3979d6} /* (13, 3, 17) {real, imag} */,
  {32'h3e1e4310, 32'h00000000} /* (13, 3, 16) {real, imag} */,
  {32'h3c937db2, 32'h3d3979d6} /* (13, 3, 15) {real, imag} */,
  {32'hbda41618, 32'hbdae9c3a} /* (13, 3, 14) {real, imag} */,
  {32'h3d9a7e5a, 32'h3d292563} /* (13, 3, 13) {real, imag} */,
  {32'hbd1ba82c, 32'h3d05c600} /* (13, 3, 12) {real, imag} */,
  {32'hbd15ca34, 32'hbe0327a1} /* (13, 3, 11) {real, imag} */,
  {32'hbd3f4619, 32'hbd19e218} /* (13, 3, 10) {real, imag} */,
  {32'h3d82bb4b, 32'h3db0459e} /* (13, 3, 9) {real, imag} */,
  {32'h3deab7b0, 32'hbcadc308} /* (13, 3, 8) {real, imag} */,
  {32'h3d80adb9, 32'h3dba4074} /* (13, 3, 7) {real, imag} */,
  {32'h3c9a7710, 32'hbc6f3130} /* (13, 3, 6) {real, imag} */,
  {32'hbe1b40df, 32'h3d9be44e} /* (13, 3, 5) {real, imag} */,
  {32'hbd7f020f, 32'hbda90fd7} /* (13, 3, 4) {real, imag} */,
  {32'hbe76639f, 32'hbe1d58f3} /* (13, 3, 3) {real, imag} */,
  {32'h3dafdb30, 32'hbf866c82} /* (13, 3, 2) {real, imag} */,
  {32'h4016776d, 32'h404611c2} /* (13, 3, 1) {real, imag} */,
  {32'h4081e5f3, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h401b704e, 32'hc043605f} /* (13, 2, 31) {real, imag} */,
  {32'h3dd68090, 32'h3f582af8} /* (13, 2, 30) {real, imag} */,
  {32'hbe8de468, 32'h3e130b33} /* (13, 2, 29) {real, imag} */,
  {32'hbe375759, 32'h3e56c2d2} /* (13, 2, 28) {real, imag} */,
  {32'hbe2ae879, 32'hbe148a6a} /* (13, 2, 27) {real, imag} */,
  {32'h3ce991c8, 32'h3c503c58} /* (13, 2, 26) {real, imag} */,
  {32'hbcc8800e, 32'h3d6ac5e0} /* (13, 2, 25) {real, imag} */,
  {32'h3dd9d028, 32'h3dc3ef1a} /* (13, 2, 24) {real, imag} */,
  {32'hbde6fa0e, 32'h3d8c9116} /* (13, 2, 23) {real, imag} */,
  {32'hbbd5b340, 32'hbc0e9d28} /* (13, 2, 22) {real, imag} */,
  {32'hbd5c77ce, 32'h3d34c343} /* (13, 2, 21) {real, imag} */,
  {32'h3dd5fd44, 32'hbe11b75d} /* (13, 2, 20) {real, imag} */,
  {32'hbd170556, 32'hbdd9611b} /* (13, 2, 19) {real, imag} */,
  {32'hbd3a7f2c, 32'hbcf2a282} /* (13, 2, 18) {real, imag} */,
  {32'h3d7c80fc, 32'h3d3a83d0} /* (13, 2, 17) {real, imag} */,
  {32'h3d5a0fde, 32'h00000000} /* (13, 2, 16) {real, imag} */,
  {32'h3d7c80fc, 32'hbd3a83d0} /* (13, 2, 15) {real, imag} */,
  {32'hbd3a7f2c, 32'h3cf2a282} /* (13, 2, 14) {real, imag} */,
  {32'hbd170556, 32'h3dd9611b} /* (13, 2, 13) {real, imag} */,
  {32'h3dd5fd44, 32'h3e11b75d} /* (13, 2, 12) {real, imag} */,
  {32'hbd5c77ce, 32'hbd34c343} /* (13, 2, 11) {real, imag} */,
  {32'hbbd5b340, 32'h3c0e9d28} /* (13, 2, 10) {real, imag} */,
  {32'hbde6fa0e, 32'hbd8c9116} /* (13, 2, 9) {real, imag} */,
  {32'h3dd9d028, 32'hbdc3ef1a} /* (13, 2, 8) {real, imag} */,
  {32'hbcc8800e, 32'hbd6ac5e0} /* (13, 2, 7) {real, imag} */,
  {32'h3ce991c8, 32'hbc503c58} /* (13, 2, 6) {real, imag} */,
  {32'hbe2ae879, 32'h3e148a6a} /* (13, 2, 5) {real, imag} */,
  {32'hbe375759, 32'hbe56c2d2} /* (13, 2, 4) {real, imag} */,
  {32'hbe8de468, 32'hbe130b33} /* (13, 2, 3) {real, imag} */,
  {32'h3dd68090, 32'hbf582af8} /* (13, 2, 2) {real, imag} */,
  {32'h401b704e, 32'h4043605f} /* (13, 2, 1) {real, imag} */,
  {32'h40851f8a, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h40169a59, 32'hc0339fd1} /* (13, 1, 31) {real, imag} */,
  {32'h3e0fb7b0, 32'h3f4647b0} /* (13, 1, 30) {real, imag} */,
  {32'hbe12fb81, 32'h3db25605} /* (13, 1, 29) {real, imag} */,
  {32'hbdeab47b, 32'h3e57b9e9} /* (13, 1, 28) {real, imag} */,
  {32'hbe5459fc, 32'hbd0b68b4} /* (13, 1, 27) {real, imag} */,
  {32'h3d681bd0, 32'hbcc151a8} /* (13, 1, 26) {real, imag} */,
  {32'h3d05fae5, 32'h3d3f6334} /* (13, 1, 25) {real, imag} */,
  {32'h3dd739e4, 32'h3d533740} /* (13, 1, 24) {real, imag} */,
  {32'hbe05df20, 32'h3deb8e86} /* (13, 1, 23) {real, imag} */,
  {32'hbd6fc7c0, 32'h3dd702f6} /* (13, 1, 22) {real, imag} */,
  {32'hbcb801d9, 32'hbe16d1bb} /* (13, 1, 21) {real, imag} */,
  {32'h3d2ca888, 32'hbd41e521} /* (13, 1, 20) {real, imag} */,
  {32'h3cc4d943, 32'hbc14f838} /* (13, 1, 19) {real, imag} */,
  {32'h3d9b4c78, 32'h3d064dea} /* (13, 1, 18) {real, imag} */,
  {32'hbd656904, 32'h3c4e2ad2} /* (13, 1, 17) {real, imag} */,
  {32'hbda61462, 32'h00000000} /* (13, 1, 16) {real, imag} */,
  {32'hbd656904, 32'hbc4e2ad2} /* (13, 1, 15) {real, imag} */,
  {32'h3d9b4c78, 32'hbd064dea} /* (13, 1, 14) {real, imag} */,
  {32'h3cc4d943, 32'h3c14f838} /* (13, 1, 13) {real, imag} */,
  {32'h3d2ca888, 32'h3d41e521} /* (13, 1, 12) {real, imag} */,
  {32'hbcb801d9, 32'h3e16d1bb} /* (13, 1, 11) {real, imag} */,
  {32'hbd6fc7c0, 32'hbdd702f6} /* (13, 1, 10) {real, imag} */,
  {32'hbe05df20, 32'hbdeb8e86} /* (13, 1, 9) {real, imag} */,
  {32'h3dd739e4, 32'hbd533740} /* (13, 1, 8) {real, imag} */,
  {32'h3d05fae5, 32'hbd3f6334} /* (13, 1, 7) {real, imag} */,
  {32'h3d681bd0, 32'h3cc151a8} /* (13, 1, 6) {real, imag} */,
  {32'hbe5459fc, 32'h3d0b68b4} /* (13, 1, 5) {real, imag} */,
  {32'hbdeab47b, 32'hbe57b9e9} /* (13, 1, 4) {real, imag} */,
  {32'hbe12fb81, 32'hbdb25605} /* (13, 1, 3) {real, imag} */,
  {32'h3e0fb7b0, 32'hbf4647b0} /* (13, 1, 2) {real, imag} */,
  {32'h40169a59, 32'h40339fd1} /* (13, 1, 1) {real, imag} */,
  {32'h40789eee, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h401b2866, 32'hc014bc3c} /* (13, 0, 31) {real, imag} */,
  {32'hbe146fa4, 32'h3f225e6a} /* (13, 0, 30) {real, imag} */,
  {32'hbd8c6e1f, 32'h3c76ed4c} /* (13, 0, 29) {real, imag} */,
  {32'hbd7a4123, 32'h3e3f5a24} /* (13, 0, 28) {real, imag} */,
  {32'hbc1f5f00, 32'h3c18b4c4} /* (13, 0, 27) {real, imag} */,
  {32'hbc9e7989, 32'h3cc36d7f} /* (13, 0, 26) {real, imag} */,
  {32'h3d99b581, 32'hbdc60eda} /* (13, 0, 25) {real, imag} */,
  {32'h3dc33b48, 32'h3c6f7e6c} /* (13, 0, 24) {real, imag} */,
  {32'h3c6bfabc, 32'hbc861b3c} /* (13, 0, 23) {real, imag} */,
  {32'hbd298a9b, 32'h3d9081a4} /* (13, 0, 22) {real, imag} */,
  {32'h3dddf547, 32'hbd03b44a} /* (13, 0, 21) {real, imag} */,
  {32'hbc1ea800, 32'h3d43ecf4} /* (13, 0, 20) {real, imag} */,
  {32'h3d19aa53, 32'h3b97ca2c} /* (13, 0, 19) {real, imag} */,
  {32'hbbd90132, 32'h3ce9a982} /* (13, 0, 18) {real, imag} */,
  {32'h3cb0b243, 32'h3d3f83c4} /* (13, 0, 17) {real, imag} */,
  {32'hbcfb8fa0, 32'h00000000} /* (13, 0, 16) {real, imag} */,
  {32'h3cb0b243, 32'hbd3f83c4} /* (13, 0, 15) {real, imag} */,
  {32'hbbd90132, 32'hbce9a982} /* (13, 0, 14) {real, imag} */,
  {32'h3d19aa53, 32'hbb97ca2c} /* (13, 0, 13) {real, imag} */,
  {32'hbc1ea800, 32'hbd43ecf4} /* (13, 0, 12) {real, imag} */,
  {32'h3dddf547, 32'h3d03b44a} /* (13, 0, 11) {real, imag} */,
  {32'hbd298a9b, 32'hbd9081a4} /* (13, 0, 10) {real, imag} */,
  {32'h3c6bfabc, 32'h3c861b3c} /* (13, 0, 9) {real, imag} */,
  {32'h3dc33b48, 32'hbc6f7e6c} /* (13, 0, 8) {real, imag} */,
  {32'h3d99b581, 32'h3dc60eda} /* (13, 0, 7) {real, imag} */,
  {32'hbc9e7989, 32'hbcc36d7f} /* (13, 0, 6) {real, imag} */,
  {32'hbc1f5f00, 32'hbc18b4c4} /* (13, 0, 5) {real, imag} */,
  {32'hbd7a4123, 32'hbe3f5a24} /* (13, 0, 4) {real, imag} */,
  {32'hbd8c6e1f, 32'hbc76ed4c} /* (13, 0, 3) {real, imag} */,
  {32'hbe146fa4, 32'hbf225e6a} /* (13, 0, 2) {real, imag} */,
  {32'h401b2866, 32'h4014bc3c} /* (13, 0, 1) {real, imag} */,
  {32'h406f85db, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h4062dca8, 32'hbffe1114} /* (12, 31, 31) {real, imag} */,
  {32'hbf3e1f30, 32'h3f05257c} /* (12, 31, 30) {real, imag} */,
  {32'hbde214d3, 32'h3d4782a0} /* (12, 31, 29) {real, imag} */,
  {32'h3d8011f0, 32'h3db31132} /* (12, 31, 28) {real, imag} */,
  {32'hbe24e98e, 32'hbc363688} /* (12, 31, 27) {real, imag} */,
  {32'h3d6fd8a4, 32'hbbb4e7a6} /* (12, 31, 26) {real, imag} */,
  {32'hbcc0f072, 32'hbce0f5d0} /* (12, 31, 25) {real, imag} */,
  {32'hbdd6702b, 32'h3c9b1306} /* (12, 31, 24) {real, imag} */,
  {32'hbd5098ac, 32'hbc4d36a4} /* (12, 31, 23) {real, imag} */,
  {32'h3c92b884, 32'hbd20775d} /* (12, 31, 22) {real, imag} */,
  {32'h3c9083be, 32'hbb063130} /* (12, 31, 21) {real, imag} */,
  {32'hbd611bd5, 32'hbd160a7a} /* (12, 31, 20) {real, imag} */,
  {32'hbc1bf298, 32'hbd3fb5d2} /* (12, 31, 19) {real, imag} */,
  {32'hbcca0d17, 32'hbcb12e2b} /* (12, 31, 18) {real, imag} */,
  {32'h3c9fe09c, 32'h3c3887e5} /* (12, 31, 17) {real, imag} */,
  {32'h3d960a7c, 32'h00000000} /* (12, 31, 16) {real, imag} */,
  {32'h3c9fe09c, 32'hbc3887e5} /* (12, 31, 15) {real, imag} */,
  {32'hbcca0d17, 32'h3cb12e2b} /* (12, 31, 14) {real, imag} */,
  {32'hbc1bf298, 32'h3d3fb5d2} /* (12, 31, 13) {real, imag} */,
  {32'hbd611bd5, 32'h3d160a7a} /* (12, 31, 12) {real, imag} */,
  {32'h3c9083be, 32'h3b063130} /* (12, 31, 11) {real, imag} */,
  {32'h3c92b884, 32'h3d20775d} /* (12, 31, 10) {real, imag} */,
  {32'hbd5098ac, 32'h3c4d36a4} /* (12, 31, 9) {real, imag} */,
  {32'hbdd6702b, 32'hbc9b1306} /* (12, 31, 8) {real, imag} */,
  {32'hbcc0f072, 32'h3ce0f5d0} /* (12, 31, 7) {real, imag} */,
  {32'h3d6fd8a4, 32'h3bb4e7a6} /* (12, 31, 6) {real, imag} */,
  {32'hbe24e98e, 32'h3c363688} /* (12, 31, 5) {real, imag} */,
  {32'h3d8011f0, 32'hbdb31132} /* (12, 31, 4) {real, imag} */,
  {32'hbde214d3, 32'hbd4782a0} /* (12, 31, 3) {real, imag} */,
  {32'hbf3e1f30, 32'hbf05257c} /* (12, 31, 2) {real, imag} */,
  {32'h4062dca8, 32'h3ffe1114} /* (12, 31, 1) {real, imag} */,
  {32'h409754de, 32'h00000000} /* (12, 31, 0) {real, imag} */,
  {32'h40802c75, 32'hbfbb559a} /* (12, 30, 31) {real, imag} */,
  {32'hbf9b914c, 32'h3efd5d01} /* (12, 30, 30) {real, imag} */,
  {32'h3cf935f8, 32'h3dba8350} /* (12, 30, 29) {real, imag} */,
  {32'h3d9a323a, 32'hbd5fb1a2} /* (12, 30, 28) {real, imag} */,
  {32'hbe9594e0, 32'hbc6f8608} /* (12, 30, 27) {real, imag} */,
  {32'h3d20048d, 32'hbd6959ca} /* (12, 30, 26) {real, imag} */,
  {32'h3c5bc9b8, 32'hbdcb1dc8} /* (12, 30, 25) {real, imag} */,
  {32'hbe00eef4, 32'h3c2bfd04} /* (12, 30, 24) {real, imag} */,
  {32'hbd3c2130, 32'hbcfdd50d} /* (12, 30, 23) {real, imag} */,
  {32'hbb9bf254, 32'h3d32701e} /* (12, 30, 22) {real, imag} */,
  {32'hbdade723, 32'h3bd48e4e} /* (12, 30, 21) {real, imag} */,
  {32'h3a2faf80, 32'h3cceaf39} /* (12, 30, 20) {real, imag} */,
  {32'h3d85c932, 32'h3ce6eb7c} /* (12, 30, 19) {real, imag} */,
  {32'h3c211920, 32'hbd3541d0} /* (12, 30, 18) {real, imag} */,
  {32'h3c14ccfc, 32'h3c5ac87e} /* (12, 30, 17) {real, imag} */,
  {32'h3dbdb6ce, 32'h00000000} /* (12, 30, 16) {real, imag} */,
  {32'h3c14ccfc, 32'hbc5ac87e} /* (12, 30, 15) {real, imag} */,
  {32'h3c211920, 32'h3d3541d0} /* (12, 30, 14) {real, imag} */,
  {32'h3d85c932, 32'hbce6eb7c} /* (12, 30, 13) {real, imag} */,
  {32'h3a2faf80, 32'hbcceaf39} /* (12, 30, 12) {real, imag} */,
  {32'hbdade723, 32'hbbd48e4e} /* (12, 30, 11) {real, imag} */,
  {32'hbb9bf254, 32'hbd32701e} /* (12, 30, 10) {real, imag} */,
  {32'hbd3c2130, 32'h3cfdd50d} /* (12, 30, 9) {real, imag} */,
  {32'hbe00eef4, 32'hbc2bfd04} /* (12, 30, 8) {real, imag} */,
  {32'h3c5bc9b8, 32'h3dcb1dc8} /* (12, 30, 7) {real, imag} */,
  {32'h3d20048d, 32'h3d6959ca} /* (12, 30, 6) {real, imag} */,
  {32'hbe9594e0, 32'h3c6f8608} /* (12, 30, 5) {real, imag} */,
  {32'h3d9a323a, 32'h3d5fb1a2} /* (12, 30, 4) {real, imag} */,
  {32'h3cf935f8, 32'hbdba8350} /* (12, 30, 3) {real, imag} */,
  {32'hbf9b914c, 32'hbefd5d01} /* (12, 30, 2) {real, imag} */,
  {32'h40802c75, 32'h3fbb559a} /* (12, 30, 1) {real, imag} */,
  {32'h40a10627, 32'h00000000} /* (12, 30, 0) {real, imag} */,
  {32'h408d1089, 32'hbf9f0e13} /* (12, 29, 31) {real, imag} */,
  {32'hbfbca606, 32'h3efa2828} /* (12, 29, 30) {real, imag} */,
  {32'h3c8a14a0, 32'h3db57ea2} /* (12, 29, 29) {real, imag} */,
  {32'h3e03e162, 32'hbe449ba3} /* (12, 29, 28) {real, imag} */,
  {32'hbe687f36, 32'hbcf8ad50} /* (12, 29, 27) {real, imag} */,
  {32'h3cdafbb6, 32'h3d52ddba} /* (12, 29, 26) {real, imag} */,
  {32'hbda166e6, 32'hbd377c3d} /* (12, 29, 25) {real, imag} */,
  {32'hbdef8d02, 32'hbccd0368} /* (12, 29, 24) {real, imag} */,
  {32'h3bc530c2, 32'h3bf92e30} /* (12, 29, 23) {real, imag} */,
  {32'hbceeac34, 32'hbb865d80} /* (12, 29, 22) {real, imag} */,
  {32'h3d770cce, 32'h3ce27409} /* (12, 29, 21) {real, imag} */,
  {32'hbd9be1e4, 32'h3dc50a13} /* (12, 29, 20) {real, imag} */,
  {32'h3d7ac29f, 32'h3db81470} /* (12, 29, 19) {real, imag} */,
  {32'h3d12da61, 32'h3daf1ba8} /* (12, 29, 18) {real, imag} */,
  {32'hbc21fdea, 32'h3b64f560} /* (12, 29, 17) {real, imag} */,
  {32'hbd5abac2, 32'h00000000} /* (12, 29, 16) {real, imag} */,
  {32'hbc21fdea, 32'hbb64f560} /* (12, 29, 15) {real, imag} */,
  {32'h3d12da61, 32'hbdaf1ba8} /* (12, 29, 14) {real, imag} */,
  {32'h3d7ac29f, 32'hbdb81470} /* (12, 29, 13) {real, imag} */,
  {32'hbd9be1e4, 32'hbdc50a13} /* (12, 29, 12) {real, imag} */,
  {32'h3d770cce, 32'hbce27409} /* (12, 29, 11) {real, imag} */,
  {32'hbceeac34, 32'h3b865d80} /* (12, 29, 10) {real, imag} */,
  {32'h3bc530c2, 32'hbbf92e30} /* (12, 29, 9) {real, imag} */,
  {32'hbdef8d02, 32'h3ccd0368} /* (12, 29, 8) {real, imag} */,
  {32'hbda166e6, 32'h3d377c3d} /* (12, 29, 7) {real, imag} */,
  {32'h3cdafbb6, 32'hbd52ddba} /* (12, 29, 6) {real, imag} */,
  {32'hbe687f36, 32'h3cf8ad50} /* (12, 29, 5) {real, imag} */,
  {32'h3e03e162, 32'h3e449ba3} /* (12, 29, 4) {real, imag} */,
  {32'h3c8a14a0, 32'hbdb57ea2} /* (12, 29, 3) {real, imag} */,
  {32'hbfbca606, 32'hbefa2828} /* (12, 29, 2) {real, imag} */,
  {32'h408d1089, 32'h3f9f0e13} /* (12, 29, 1) {real, imag} */,
  {32'h40a09f1d, 32'h00000000} /* (12, 29, 0) {real, imag} */,
  {32'h40977443, 32'hbf8aead2} /* (12, 28, 31) {real, imag} */,
  {32'hbfca5662, 32'h3e92cd8a} /* (12, 28, 30) {real, imag} */,
  {32'hbd590de3, 32'h3d8696a6} /* (12, 28, 29) {real, imag} */,
  {32'h3e07d336, 32'hbe6c589d} /* (12, 28, 28) {real, imag} */,
  {32'hbe51146d, 32'h3d0c5081} /* (12, 28, 27) {real, imag} */,
  {32'hbc2562bd, 32'hbcf7980f} /* (12, 28, 26) {real, imag} */,
  {32'hbb644350, 32'h3d70df96} /* (12, 28, 25) {real, imag} */,
  {32'hbdffd0cd, 32'h3ce1b714} /* (12, 28, 24) {real, imag} */,
  {32'hbb6959d0, 32'h3dff780c} /* (12, 28, 23) {real, imag} */,
  {32'hbc208d60, 32'h3e0ff931} /* (12, 28, 22) {real, imag} */,
  {32'h3d8726db, 32'h3d265d25} /* (12, 28, 21) {real, imag} */,
  {32'hbd1255b9, 32'h3bd1ac1c} /* (12, 28, 20) {real, imag} */,
  {32'hbdfc743a, 32'hbcfa9714} /* (12, 28, 19) {real, imag} */,
  {32'h3d41ec22, 32'hbcaad4ec} /* (12, 28, 18) {real, imag} */,
  {32'h3da261d4, 32'hbd9af4cc} /* (12, 28, 17) {real, imag} */,
  {32'h3ce20aa2, 32'h00000000} /* (12, 28, 16) {real, imag} */,
  {32'h3da261d4, 32'h3d9af4cc} /* (12, 28, 15) {real, imag} */,
  {32'h3d41ec22, 32'h3caad4ec} /* (12, 28, 14) {real, imag} */,
  {32'hbdfc743a, 32'h3cfa9714} /* (12, 28, 13) {real, imag} */,
  {32'hbd1255b9, 32'hbbd1ac1c} /* (12, 28, 12) {real, imag} */,
  {32'h3d8726db, 32'hbd265d25} /* (12, 28, 11) {real, imag} */,
  {32'hbc208d60, 32'hbe0ff931} /* (12, 28, 10) {real, imag} */,
  {32'hbb6959d0, 32'hbdff780c} /* (12, 28, 9) {real, imag} */,
  {32'hbdffd0cd, 32'hbce1b714} /* (12, 28, 8) {real, imag} */,
  {32'hbb644350, 32'hbd70df96} /* (12, 28, 7) {real, imag} */,
  {32'hbc2562bd, 32'h3cf7980f} /* (12, 28, 6) {real, imag} */,
  {32'hbe51146d, 32'hbd0c5081} /* (12, 28, 5) {real, imag} */,
  {32'h3e07d336, 32'h3e6c589d} /* (12, 28, 4) {real, imag} */,
  {32'hbd590de3, 32'hbd8696a6} /* (12, 28, 3) {real, imag} */,
  {32'hbfca5662, 32'hbe92cd8a} /* (12, 28, 2) {real, imag} */,
  {32'h40977443, 32'h3f8aead2} /* (12, 28, 1) {real, imag} */,
  {32'h409baf19, 32'h00000000} /* (12, 28, 0) {real, imag} */,
  {32'h409bd260, 32'hbf6e34e9} /* (12, 27, 31) {real, imag} */,
  {32'hbfd0e6c1, 32'h3e093a12} /* (12, 27, 30) {real, imag} */,
  {32'h3bc05c70, 32'hbd9ec3c2} /* (12, 27, 29) {real, imag} */,
  {32'h3d5e3e3e, 32'hbe8f432e} /* (12, 27, 28) {real, imag} */,
  {32'hbe04b16c, 32'h3db98940} /* (12, 27, 27) {real, imag} */,
  {32'hbc2303e4, 32'h3db8334e} /* (12, 27, 26) {real, imag} */,
  {32'h3c8d02ad, 32'hbc6de920} /* (12, 27, 25) {real, imag} */,
  {32'hbd2239a4, 32'h3e30bb64} /* (12, 27, 24) {real, imag} */,
  {32'hbdcd7672, 32'hbd5d0d67} /* (12, 27, 23) {real, imag} */,
  {32'h3cc774a8, 32'h3da7f2cd} /* (12, 27, 22) {real, imag} */,
  {32'hbc9da452, 32'hbb3f5640} /* (12, 27, 21) {real, imag} */,
  {32'h3e0a649e, 32'h3dc18f96} /* (12, 27, 20) {real, imag} */,
  {32'hbc3c966a, 32'h3de09433} /* (12, 27, 19) {real, imag} */,
  {32'hbca238c9, 32'hbb911f24} /* (12, 27, 18) {real, imag} */,
  {32'h3d6d5bd2, 32'h3c602e90} /* (12, 27, 17) {real, imag} */,
  {32'h3baf9bb4, 32'h00000000} /* (12, 27, 16) {real, imag} */,
  {32'h3d6d5bd2, 32'hbc602e90} /* (12, 27, 15) {real, imag} */,
  {32'hbca238c9, 32'h3b911f24} /* (12, 27, 14) {real, imag} */,
  {32'hbc3c966a, 32'hbde09433} /* (12, 27, 13) {real, imag} */,
  {32'h3e0a649e, 32'hbdc18f96} /* (12, 27, 12) {real, imag} */,
  {32'hbc9da452, 32'h3b3f5640} /* (12, 27, 11) {real, imag} */,
  {32'h3cc774a8, 32'hbda7f2cd} /* (12, 27, 10) {real, imag} */,
  {32'hbdcd7672, 32'h3d5d0d67} /* (12, 27, 9) {real, imag} */,
  {32'hbd2239a4, 32'hbe30bb64} /* (12, 27, 8) {real, imag} */,
  {32'h3c8d02ad, 32'h3c6de920} /* (12, 27, 7) {real, imag} */,
  {32'hbc2303e4, 32'hbdb8334e} /* (12, 27, 6) {real, imag} */,
  {32'hbe04b16c, 32'hbdb98940} /* (12, 27, 5) {real, imag} */,
  {32'h3d5e3e3e, 32'h3e8f432e} /* (12, 27, 4) {real, imag} */,
  {32'h3bc05c70, 32'h3d9ec3c2} /* (12, 27, 3) {real, imag} */,
  {32'hbfd0e6c1, 32'hbe093a12} /* (12, 27, 2) {real, imag} */,
  {32'h409bd260, 32'h3f6e34e9} /* (12, 27, 1) {real, imag} */,
  {32'h409702f1, 32'h00000000} /* (12, 27, 0) {real, imag} */,
  {32'h4093491a, 32'hbf53bc34} /* (12, 26, 31) {real, imag} */,
  {32'hbfda71ea, 32'h3e32b962} /* (12, 26, 30) {real, imag} */,
  {32'h3d89c3d1, 32'hbdad5688} /* (12, 26, 29) {real, imag} */,
  {32'h3e43d45a, 32'hbd00e8e6} /* (12, 26, 28) {real, imag} */,
  {32'hbe0dac78, 32'h3e19b875} /* (12, 26, 27) {real, imag} */,
  {32'hbdcc7d90, 32'h3b6ec970} /* (12, 26, 26) {real, imag} */,
  {32'h3caea0ec, 32'hbe0dac98} /* (12, 26, 25) {real, imag} */,
  {32'h3bce6e9c, 32'h3e24cf60} /* (12, 26, 24) {real, imag} */,
  {32'hbcbbac51, 32'h3d1ea458} /* (12, 26, 23) {real, imag} */,
  {32'h3cebeb2b, 32'hbd793b0a} /* (12, 26, 22) {real, imag} */,
  {32'h3c7c2118, 32'h3d267fe0} /* (12, 26, 21) {real, imag} */,
  {32'hbd139dd1, 32'h3d9db610} /* (12, 26, 20) {real, imag} */,
  {32'h3d1b080c, 32'h3d7ff571} /* (12, 26, 19) {real, imag} */,
  {32'hbcd63aa4, 32'hbcd968a4} /* (12, 26, 18) {real, imag} */,
  {32'hbcb74629, 32'hbcfba346} /* (12, 26, 17) {real, imag} */,
  {32'hbcbf309b, 32'h00000000} /* (12, 26, 16) {real, imag} */,
  {32'hbcb74629, 32'h3cfba346} /* (12, 26, 15) {real, imag} */,
  {32'hbcd63aa4, 32'h3cd968a4} /* (12, 26, 14) {real, imag} */,
  {32'h3d1b080c, 32'hbd7ff571} /* (12, 26, 13) {real, imag} */,
  {32'hbd139dd1, 32'hbd9db610} /* (12, 26, 12) {real, imag} */,
  {32'h3c7c2118, 32'hbd267fe0} /* (12, 26, 11) {real, imag} */,
  {32'h3cebeb2b, 32'h3d793b0a} /* (12, 26, 10) {real, imag} */,
  {32'hbcbbac51, 32'hbd1ea458} /* (12, 26, 9) {real, imag} */,
  {32'h3bce6e9c, 32'hbe24cf60} /* (12, 26, 8) {real, imag} */,
  {32'h3caea0ec, 32'h3e0dac98} /* (12, 26, 7) {real, imag} */,
  {32'hbdcc7d90, 32'hbb6ec970} /* (12, 26, 6) {real, imag} */,
  {32'hbe0dac78, 32'hbe19b875} /* (12, 26, 5) {real, imag} */,
  {32'h3e43d45a, 32'h3d00e8e6} /* (12, 26, 4) {real, imag} */,
  {32'h3d89c3d1, 32'h3dad5688} /* (12, 26, 3) {real, imag} */,
  {32'hbfda71ea, 32'hbe32b962} /* (12, 26, 2) {real, imag} */,
  {32'h4093491a, 32'h3f53bc34} /* (12, 26, 1) {real, imag} */,
  {32'h408f1f7e, 32'h00000000} /* (12, 26, 0) {real, imag} */,
  {32'h408bb832, 32'hbf336552} /* (12, 25, 31) {real, imag} */,
  {32'hbfd37076, 32'h3e0ebfca} /* (12, 25, 30) {real, imag} */,
  {32'h3cd2d36c, 32'h3d15a9f6} /* (12, 25, 29) {real, imag} */,
  {32'h3e39a86e, 32'hbd8bd2a6} /* (12, 25, 28) {real, imag} */,
  {32'hbddcfdaa, 32'h3e63277d} /* (12, 25, 27) {real, imag} */,
  {32'hbe3ebff5, 32'hbd920086} /* (12, 25, 26) {real, imag} */,
  {32'h3d52147c, 32'h3cfcc7c8} /* (12, 25, 25) {real, imag} */,
  {32'hbdb06a92, 32'h3df03f4d} /* (12, 25, 24) {real, imag} */,
  {32'h3d7200d2, 32'h3a770700} /* (12, 25, 23) {real, imag} */,
  {32'hbdc8a890, 32'hbe184f53} /* (12, 25, 22) {real, imag} */,
  {32'hbdac7276, 32'h3d34e23a} /* (12, 25, 21) {real, imag} */,
  {32'hbcefe602, 32'h3dd40928} /* (12, 25, 20) {real, imag} */,
  {32'h3ca31c12, 32'hbd29d1e2} /* (12, 25, 19) {real, imag} */,
  {32'h3b9d0944, 32'h3cad2ea3} /* (12, 25, 18) {real, imag} */,
  {32'h3d172d0d, 32'hbd9f4a68} /* (12, 25, 17) {real, imag} */,
  {32'h3d877a74, 32'h00000000} /* (12, 25, 16) {real, imag} */,
  {32'h3d172d0d, 32'h3d9f4a68} /* (12, 25, 15) {real, imag} */,
  {32'h3b9d0944, 32'hbcad2ea3} /* (12, 25, 14) {real, imag} */,
  {32'h3ca31c12, 32'h3d29d1e2} /* (12, 25, 13) {real, imag} */,
  {32'hbcefe602, 32'hbdd40928} /* (12, 25, 12) {real, imag} */,
  {32'hbdac7276, 32'hbd34e23a} /* (12, 25, 11) {real, imag} */,
  {32'hbdc8a890, 32'h3e184f53} /* (12, 25, 10) {real, imag} */,
  {32'h3d7200d2, 32'hba770700} /* (12, 25, 9) {real, imag} */,
  {32'hbdb06a92, 32'hbdf03f4d} /* (12, 25, 8) {real, imag} */,
  {32'h3d52147c, 32'hbcfcc7c8} /* (12, 25, 7) {real, imag} */,
  {32'hbe3ebff5, 32'h3d920086} /* (12, 25, 6) {real, imag} */,
  {32'hbddcfdaa, 32'hbe63277d} /* (12, 25, 5) {real, imag} */,
  {32'h3e39a86e, 32'h3d8bd2a6} /* (12, 25, 4) {real, imag} */,
  {32'h3cd2d36c, 32'hbd15a9f6} /* (12, 25, 3) {real, imag} */,
  {32'hbfd37076, 32'hbe0ebfca} /* (12, 25, 2) {real, imag} */,
  {32'h408bb832, 32'h3f336552} /* (12, 25, 1) {real, imag} */,
  {32'h407f8be7, 32'h00000000} /* (12, 25, 0) {real, imag} */,
  {32'h407ae782, 32'hbf09ac1e} /* (12, 24, 31) {real, imag} */,
  {32'hbfc1f575, 32'h3e422592} /* (12, 24, 30) {real, imag} */,
  {32'hbdc71e04, 32'hbd30e1b9} /* (12, 24, 29) {real, imag} */,
  {32'h3e5b5ce8, 32'hbd8ca465} /* (12, 24, 28) {real, imag} */,
  {32'hbda79677, 32'h3e489e52} /* (12, 24, 27) {real, imag} */,
  {32'hbe179ed8, 32'hbd7423a0} /* (12, 24, 26) {real, imag} */,
  {32'h3db7459c, 32'hbcf71943} /* (12, 24, 25) {real, imag} */,
  {32'hbd939b62, 32'h3e4679e2} /* (12, 24, 24) {real, imag} */,
  {32'h3db55f1a, 32'h3d6973be} /* (12, 24, 23) {real, imag} */,
  {32'h3cb78d62, 32'hbe1e7976} /* (12, 24, 22) {real, imag} */,
  {32'hbd15b72b, 32'h3dab42c7} /* (12, 24, 21) {real, imag} */,
  {32'h3c7cfa28, 32'hbcf297b4} /* (12, 24, 20) {real, imag} */,
  {32'hbbc7a8a0, 32'hbdabc475} /* (12, 24, 19) {real, imag} */,
  {32'h3cd0f8c3, 32'hbc9b271e} /* (12, 24, 18) {real, imag} */,
  {32'h3bbab9e4, 32'h3d2bf532} /* (12, 24, 17) {real, imag} */,
  {32'h3af5ba20, 32'h00000000} /* (12, 24, 16) {real, imag} */,
  {32'h3bbab9e4, 32'hbd2bf532} /* (12, 24, 15) {real, imag} */,
  {32'h3cd0f8c3, 32'h3c9b271e} /* (12, 24, 14) {real, imag} */,
  {32'hbbc7a8a0, 32'h3dabc475} /* (12, 24, 13) {real, imag} */,
  {32'h3c7cfa28, 32'h3cf297b4} /* (12, 24, 12) {real, imag} */,
  {32'hbd15b72b, 32'hbdab42c7} /* (12, 24, 11) {real, imag} */,
  {32'h3cb78d62, 32'h3e1e7976} /* (12, 24, 10) {real, imag} */,
  {32'h3db55f1a, 32'hbd6973be} /* (12, 24, 9) {real, imag} */,
  {32'hbd939b62, 32'hbe4679e2} /* (12, 24, 8) {real, imag} */,
  {32'h3db7459c, 32'h3cf71943} /* (12, 24, 7) {real, imag} */,
  {32'hbe179ed8, 32'h3d7423a0} /* (12, 24, 6) {real, imag} */,
  {32'hbda79677, 32'hbe489e52} /* (12, 24, 5) {real, imag} */,
  {32'h3e5b5ce8, 32'h3d8ca465} /* (12, 24, 4) {real, imag} */,
  {32'hbdc71e04, 32'h3d30e1b9} /* (12, 24, 3) {real, imag} */,
  {32'hbfc1f575, 32'hbe422592} /* (12, 24, 2) {real, imag} */,
  {32'h407ae782, 32'h3f09ac1e} /* (12, 24, 1) {real, imag} */,
  {32'h40588330, 32'h00000000} /* (12, 24, 0) {real, imag} */,
  {32'h404cdd4d, 32'hbeff7483} /* (12, 23, 31) {real, imag} */,
  {32'hbf973298, 32'h3e2cbfa7} /* (12, 23, 30) {real, imag} */,
  {32'hbdf17597, 32'hbd062a82} /* (12, 23, 29) {real, imag} */,
  {32'h3e25dbd5, 32'hbe33a8cf} /* (12, 23, 28) {real, imag} */,
  {32'hbe681963, 32'h3d877658} /* (12, 23, 27) {real, imag} */,
  {32'hbd4aa5cb, 32'h3c8644a1} /* (12, 23, 26) {real, imag} */,
  {32'hbbd84ca4, 32'hbce49194} /* (12, 23, 25) {real, imag} */,
  {32'hbc02901e, 32'h3d6b23fe} /* (12, 23, 24) {real, imag} */,
  {32'hbd9ea9d4, 32'h3d8acc25} /* (12, 23, 23) {real, imag} */,
  {32'h3d0f9cdf, 32'h3d932a49} /* (12, 23, 22) {real, imag} */,
  {32'h3d77d3e5, 32'h3d62c04a} /* (12, 23, 21) {real, imag} */,
  {32'hbd62c994, 32'h3d098d84} /* (12, 23, 20) {real, imag} */,
  {32'h3d52d5ba, 32'h3bee4440} /* (12, 23, 19) {real, imag} */,
  {32'hbb93d6a0, 32'hbb7b7bb0} /* (12, 23, 18) {real, imag} */,
  {32'h3c6980f2, 32'hbd84cd3e} /* (12, 23, 17) {real, imag} */,
  {32'hbd1c6080, 32'h00000000} /* (12, 23, 16) {real, imag} */,
  {32'h3c6980f2, 32'h3d84cd3e} /* (12, 23, 15) {real, imag} */,
  {32'hbb93d6a0, 32'h3b7b7bb0} /* (12, 23, 14) {real, imag} */,
  {32'h3d52d5ba, 32'hbbee4440} /* (12, 23, 13) {real, imag} */,
  {32'hbd62c994, 32'hbd098d84} /* (12, 23, 12) {real, imag} */,
  {32'h3d77d3e5, 32'hbd62c04a} /* (12, 23, 11) {real, imag} */,
  {32'h3d0f9cdf, 32'hbd932a49} /* (12, 23, 10) {real, imag} */,
  {32'hbd9ea9d4, 32'hbd8acc25} /* (12, 23, 9) {real, imag} */,
  {32'hbc02901e, 32'hbd6b23fe} /* (12, 23, 8) {real, imag} */,
  {32'hbbd84ca4, 32'h3ce49194} /* (12, 23, 7) {real, imag} */,
  {32'hbd4aa5cb, 32'hbc8644a1} /* (12, 23, 6) {real, imag} */,
  {32'hbe681963, 32'hbd877658} /* (12, 23, 5) {real, imag} */,
  {32'h3e25dbd5, 32'h3e33a8cf} /* (12, 23, 4) {real, imag} */,
  {32'hbdf17597, 32'h3d062a82} /* (12, 23, 3) {real, imag} */,
  {32'hbf973298, 32'hbe2cbfa7} /* (12, 23, 2) {real, imag} */,
  {32'h404cdd4d, 32'h3eff7483} /* (12, 23, 1) {real, imag} */,
  {32'h40284369, 32'h00000000} /* (12, 23, 0) {real, imag} */,
  {32'h4015661e, 32'hbe9c888f} /* (12, 22, 31) {real, imag} */,
  {32'hbf4fcd15, 32'h3e54b89e} /* (12, 22, 30) {real, imag} */,
  {32'hbd57e2c2, 32'hbcbebde2} /* (12, 22, 29) {real, imag} */,
  {32'h3eac0825, 32'hbe3c6a4e} /* (12, 22, 28) {real, imag} */,
  {32'hbe8e7d5a, 32'h3e68e7a8} /* (12, 22, 27) {real, imag} */,
  {32'hbe20d61c, 32'hbd736e6d} /* (12, 22, 26) {real, imag} */,
  {32'h3e0e42ea, 32'h3bea7be8} /* (12, 22, 25) {real, imag} */,
  {32'hbe0e6251, 32'hbc19bc2c} /* (12, 22, 24) {real, imag} */,
  {32'hbdc93aaa, 32'h3dc9fedf} /* (12, 22, 23) {real, imag} */,
  {32'h3db3f2d9, 32'h3cab91e9} /* (12, 22, 22) {real, imag} */,
  {32'hbda3ec6a, 32'h3cbd98b4} /* (12, 22, 21) {real, imag} */,
  {32'hbd3dccf2, 32'h3d1c17f5} /* (12, 22, 20) {real, imag} */,
  {32'h3b146460, 32'h3c8d6ebf} /* (12, 22, 19) {real, imag} */,
  {32'h3d0bde1c, 32'hbc28b978} /* (12, 22, 18) {real, imag} */,
  {32'h3db92176, 32'h3d191198} /* (12, 22, 17) {real, imag} */,
  {32'hbdfd70d2, 32'h00000000} /* (12, 22, 16) {real, imag} */,
  {32'h3db92176, 32'hbd191198} /* (12, 22, 15) {real, imag} */,
  {32'h3d0bde1c, 32'h3c28b978} /* (12, 22, 14) {real, imag} */,
  {32'h3b146460, 32'hbc8d6ebf} /* (12, 22, 13) {real, imag} */,
  {32'hbd3dccf2, 32'hbd1c17f5} /* (12, 22, 12) {real, imag} */,
  {32'hbda3ec6a, 32'hbcbd98b4} /* (12, 22, 11) {real, imag} */,
  {32'h3db3f2d9, 32'hbcab91e9} /* (12, 22, 10) {real, imag} */,
  {32'hbdc93aaa, 32'hbdc9fedf} /* (12, 22, 9) {real, imag} */,
  {32'hbe0e6251, 32'h3c19bc2c} /* (12, 22, 8) {real, imag} */,
  {32'h3e0e42ea, 32'hbbea7be8} /* (12, 22, 7) {real, imag} */,
  {32'hbe20d61c, 32'h3d736e6d} /* (12, 22, 6) {real, imag} */,
  {32'hbe8e7d5a, 32'hbe68e7a8} /* (12, 22, 5) {real, imag} */,
  {32'h3eac0825, 32'h3e3c6a4e} /* (12, 22, 4) {real, imag} */,
  {32'hbd57e2c2, 32'h3cbebde2} /* (12, 22, 3) {real, imag} */,
  {32'hbf4fcd15, 32'hbe54b89e} /* (12, 22, 2) {real, imag} */,
  {32'h4015661e, 32'h3e9c888f} /* (12, 22, 1) {real, imag} */,
  {32'h3fe815af, 32'h00000000} /* (12, 22, 0) {real, imag} */,
  {32'h3f3c8e7c, 32'h3bbee100} /* (12, 21, 31) {real, imag} */,
  {32'hbe78b440, 32'h3c4d0a60} /* (12, 21, 30) {real, imag} */,
  {32'hbd3b3ecf, 32'hbc3efeae} /* (12, 21, 29) {real, imag} */,
  {32'h3e3f8de4, 32'hbc7ec510} /* (12, 21, 28) {real, imag} */,
  {32'hbe260b0a, 32'h3de31250} /* (12, 21, 27) {real, imag} */,
  {32'hbdab5b1e, 32'h3c41025e} /* (12, 21, 26) {real, imag} */,
  {32'h3d135774, 32'hbc941bd4} /* (12, 21, 25) {real, imag} */,
  {32'hbdcbf3a8, 32'h3b4ec0bc} /* (12, 21, 24) {real, imag} */,
  {32'h3d72d1a5, 32'h3bc846fa} /* (12, 21, 23) {real, imag} */,
  {32'hbccbfd5a, 32'hbdc2c8df} /* (12, 21, 22) {real, imag} */,
  {32'hbdc699ea, 32'h3caa8fe2} /* (12, 21, 21) {real, imag} */,
  {32'hbd347020, 32'hbd774280} /* (12, 21, 20) {real, imag} */,
  {32'hbcb29244, 32'h3c98b10b} /* (12, 21, 19) {real, imag} */,
  {32'hbbb47ae4, 32'h3cc30518} /* (12, 21, 18) {real, imag} */,
  {32'hbcff46e4, 32'h3c94ad3a} /* (12, 21, 17) {real, imag} */,
  {32'h3e02e420, 32'h00000000} /* (12, 21, 16) {real, imag} */,
  {32'hbcff46e4, 32'hbc94ad3a} /* (12, 21, 15) {real, imag} */,
  {32'hbbb47ae4, 32'hbcc30518} /* (12, 21, 14) {real, imag} */,
  {32'hbcb29244, 32'hbc98b10b} /* (12, 21, 13) {real, imag} */,
  {32'hbd347020, 32'h3d774280} /* (12, 21, 12) {real, imag} */,
  {32'hbdc699ea, 32'hbcaa8fe2} /* (12, 21, 11) {real, imag} */,
  {32'hbccbfd5a, 32'h3dc2c8df} /* (12, 21, 10) {real, imag} */,
  {32'h3d72d1a5, 32'hbbc846fa} /* (12, 21, 9) {real, imag} */,
  {32'hbdcbf3a8, 32'hbb4ec0bc} /* (12, 21, 8) {real, imag} */,
  {32'h3d135774, 32'h3c941bd4} /* (12, 21, 7) {real, imag} */,
  {32'hbdab5b1e, 32'hbc41025e} /* (12, 21, 6) {real, imag} */,
  {32'hbe260b0a, 32'hbde31250} /* (12, 21, 5) {real, imag} */,
  {32'h3e3f8de4, 32'h3c7ec510} /* (12, 21, 4) {real, imag} */,
  {32'hbd3b3ecf, 32'h3c3efeae} /* (12, 21, 3) {real, imag} */,
  {32'hbe78b440, 32'hbc4d0a60} /* (12, 21, 2) {real, imag} */,
  {32'h3f3c8e7c, 32'hbbbee100} /* (12, 21, 1) {real, imag} */,
  {32'h3f2db1ad, 32'h00000000} /* (12, 21, 0) {real, imag} */,
  {32'hbf9515b8, 32'h3e5316a4} /* (12, 20, 31) {real, imag} */,
  {32'h3f1ac181, 32'hbe13305f} /* (12, 20, 30) {real, imag} */,
  {32'hbe00b7b5, 32'h3c91908a} /* (12, 20, 29) {real, imag} */,
  {32'hbd53da1a, 32'h3e3ca5da} /* (12, 20, 28) {real, imag} */,
  {32'h3e53ddca, 32'hbd208e58} /* (12, 20, 27) {real, imag} */,
  {32'h3cfcd5d8, 32'h3c97b207} /* (12, 20, 26) {real, imag} */,
  {32'hbd8ad458, 32'hbc052148} /* (12, 20, 25) {real, imag} */,
  {32'h3dc2d10c, 32'hbcd85544} /* (12, 20, 24) {real, imag} */,
  {32'h3d725482, 32'hbd0b3e0e} /* (12, 20, 23) {real, imag} */,
  {32'hbdcd1afc, 32'h3d73d632} /* (12, 20, 22) {real, imag} */,
  {32'h3dc0dba5, 32'hbc761f44} /* (12, 20, 21) {real, imag} */,
  {32'hbc42fd6c, 32'hbda4b0c2} /* (12, 20, 20) {real, imag} */,
  {32'h3cca90ad, 32'hbd68e476} /* (12, 20, 19) {real, imag} */,
  {32'hbdae779d, 32'h3ca2333a} /* (12, 20, 18) {real, imag} */,
  {32'h3d34cda2, 32'hbdd85af7} /* (12, 20, 17) {real, imag} */,
  {32'hbc980dc2, 32'h00000000} /* (12, 20, 16) {real, imag} */,
  {32'h3d34cda2, 32'h3dd85af7} /* (12, 20, 15) {real, imag} */,
  {32'hbdae779d, 32'hbca2333a} /* (12, 20, 14) {real, imag} */,
  {32'h3cca90ad, 32'h3d68e476} /* (12, 20, 13) {real, imag} */,
  {32'hbc42fd6c, 32'h3da4b0c2} /* (12, 20, 12) {real, imag} */,
  {32'h3dc0dba5, 32'h3c761f44} /* (12, 20, 11) {real, imag} */,
  {32'hbdcd1afc, 32'hbd73d632} /* (12, 20, 10) {real, imag} */,
  {32'h3d725482, 32'h3d0b3e0e} /* (12, 20, 9) {real, imag} */,
  {32'h3dc2d10c, 32'h3cd85544} /* (12, 20, 8) {real, imag} */,
  {32'hbd8ad458, 32'h3c052148} /* (12, 20, 7) {real, imag} */,
  {32'h3cfcd5d8, 32'hbc97b207} /* (12, 20, 6) {real, imag} */,
  {32'h3e53ddca, 32'h3d208e58} /* (12, 20, 5) {real, imag} */,
  {32'hbd53da1a, 32'hbe3ca5da} /* (12, 20, 4) {real, imag} */,
  {32'hbe00b7b5, 32'hbc91908a} /* (12, 20, 3) {real, imag} */,
  {32'h3f1ac181, 32'h3e13305f} /* (12, 20, 2) {real, imag} */,
  {32'hbf9515b8, 32'hbe5316a4} /* (12, 20, 1) {real, imag} */,
  {32'hbf5728fe, 32'h00000000} /* (12, 20, 0) {real, imag} */,
  {32'hc014c6b1, 32'h3e847d78} /* (12, 19, 31) {real, imag} */,
  {32'h3f85a3ec, 32'hbe6a2a15} /* (12, 19, 30) {real, imag} */,
  {32'hbdd16014, 32'h3c340602} /* (12, 19, 29) {real, imag} */,
  {32'hbdcac844, 32'h3d6ade06} /* (12, 19, 28) {real, imag} */,
  {32'h3e33ff7b, 32'h3cc0d4ae} /* (12, 19, 27) {real, imag} */,
  {32'hbd8cda5c, 32'hbd00ce83} /* (12, 19, 26) {real, imag} */,
  {32'hbdbca94e, 32'h3d8424b2} /* (12, 19, 25) {real, imag} */,
  {32'h3ddefd2b, 32'hbe3dc0e7} /* (12, 19, 24) {real, imag} */,
  {32'h3cc70835, 32'hbd1ea360} /* (12, 19, 23) {real, imag} */,
  {32'hbc7d7fd8, 32'hbde02748} /* (12, 19, 22) {real, imag} */,
  {32'h3da67cf8, 32'hbd99350d} /* (12, 19, 21) {real, imag} */,
  {32'h3d8180c0, 32'h3c915414} /* (12, 19, 20) {real, imag} */,
  {32'hbc536a84, 32'h3d0fc56a} /* (12, 19, 19) {real, imag} */,
  {32'hbde3cdeb, 32'hbdd4a0e6} /* (12, 19, 18) {real, imag} */,
  {32'hbd7b285f, 32'hbc49c9c8} /* (12, 19, 17) {real, imag} */,
  {32'hbbe76e0c, 32'h00000000} /* (12, 19, 16) {real, imag} */,
  {32'hbd7b285f, 32'h3c49c9c8} /* (12, 19, 15) {real, imag} */,
  {32'hbde3cdeb, 32'h3dd4a0e6} /* (12, 19, 14) {real, imag} */,
  {32'hbc536a84, 32'hbd0fc56a} /* (12, 19, 13) {real, imag} */,
  {32'h3d8180c0, 32'hbc915414} /* (12, 19, 12) {real, imag} */,
  {32'h3da67cf8, 32'h3d99350d} /* (12, 19, 11) {real, imag} */,
  {32'hbc7d7fd8, 32'h3de02748} /* (12, 19, 10) {real, imag} */,
  {32'h3cc70835, 32'h3d1ea360} /* (12, 19, 9) {real, imag} */,
  {32'h3ddefd2b, 32'h3e3dc0e7} /* (12, 19, 8) {real, imag} */,
  {32'hbdbca94e, 32'hbd8424b2} /* (12, 19, 7) {real, imag} */,
  {32'hbd8cda5c, 32'h3d00ce83} /* (12, 19, 6) {real, imag} */,
  {32'h3e33ff7b, 32'hbcc0d4ae} /* (12, 19, 5) {real, imag} */,
  {32'hbdcac844, 32'hbd6ade06} /* (12, 19, 4) {real, imag} */,
  {32'hbdd16014, 32'hbc340602} /* (12, 19, 3) {real, imag} */,
  {32'h3f85a3ec, 32'h3e6a2a15} /* (12, 19, 2) {real, imag} */,
  {32'hc014c6b1, 32'hbe847d78} /* (12, 19, 1) {real, imag} */,
  {32'hbfdef6e4, 32'h00000000} /* (12, 19, 0) {real, imag} */,
  {32'hc0490edd, 32'h3ee8c616} /* (12, 18, 31) {real, imag} */,
  {32'h3fa4e7e4, 32'hbe8328b1} /* (12, 18, 30) {real, imag} */,
  {32'hbc980178, 32'h3c61b008} /* (12, 18, 29) {real, imag} */,
  {32'hbd93b25c, 32'h3e09b374} /* (12, 18, 28) {real, imag} */,
  {32'h3ea9d41c, 32'hbe197dfc} /* (12, 18, 27) {real, imag} */,
  {32'hbd75d68c, 32'h3cb87a34} /* (12, 18, 26) {real, imag} */,
  {32'h3c8bbbf6, 32'hbceacdc6} /* (12, 18, 25) {real, imag} */,
  {32'h3cd70136, 32'hbdcb5eaa} /* (12, 18, 24) {real, imag} */,
  {32'h3de6aa66, 32'h3d363788} /* (12, 18, 23) {real, imag} */,
  {32'hbda42020, 32'h3d8d8a4d} /* (12, 18, 22) {real, imag} */,
  {32'hbd0fdf4f, 32'hbd9e487e} /* (12, 18, 21) {real, imag} */,
  {32'hbd18580a, 32'h3d855ced} /* (12, 18, 20) {real, imag} */,
  {32'h3c945cee, 32'h3e0a6f55} /* (12, 18, 19) {real, imag} */,
  {32'h3c9e6448, 32'hbdc93f72} /* (12, 18, 18) {real, imag} */,
  {32'hbd2a10cc, 32'h3d507e48} /* (12, 18, 17) {real, imag} */,
  {32'h3d926c80, 32'h00000000} /* (12, 18, 16) {real, imag} */,
  {32'hbd2a10cc, 32'hbd507e48} /* (12, 18, 15) {real, imag} */,
  {32'h3c9e6448, 32'h3dc93f72} /* (12, 18, 14) {real, imag} */,
  {32'h3c945cee, 32'hbe0a6f55} /* (12, 18, 13) {real, imag} */,
  {32'hbd18580a, 32'hbd855ced} /* (12, 18, 12) {real, imag} */,
  {32'hbd0fdf4f, 32'h3d9e487e} /* (12, 18, 11) {real, imag} */,
  {32'hbda42020, 32'hbd8d8a4d} /* (12, 18, 10) {real, imag} */,
  {32'h3de6aa66, 32'hbd363788} /* (12, 18, 9) {real, imag} */,
  {32'h3cd70136, 32'h3dcb5eaa} /* (12, 18, 8) {real, imag} */,
  {32'h3c8bbbf6, 32'h3ceacdc6} /* (12, 18, 7) {real, imag} */,
  {32'hbd75d68c, 32'hbcb87a34} /* (12, 18, 6) {real, imag} */,
  {32'h3ea9d41c, 32'h3e197dfc} /* (12, 18, 5) {real, imag} */,
  {32'hbd93b25c, 32'hbe09b374} /* (12, 18, 4) {real, imag} */,
  {32'hbc980178, 32'hbc61b008} /* (12, 18, 3) {real, imag} */,
  {32'h3fa4e7e4, 32'h3e8328b1} /* (12, 18, 2) {real, imag} */,
  {32'hc0490edd, 32'hbee8c616} /* (12, 18, 1) {real, imag} */,
  {32'hc01fd213, 32'h00000000} /* (12, 18, 0) {real, imag} */,
  {32'hc06c6054, 32'h3efe8a6d} /* (12, 17, 31) {real, imag} */,
  {32'h3fbbf0e9, 32'hbe6fd60a} /* (12, 17, 30) {real, imag} */,
  {32'h3de237ab, 32'h3c3c84c2} /* (12, 17, 29) {real, imag} */,
  {32'h3d1f3cfc, 32'h3da1cdb6} /* (12, 17, 28) {real, imag} */,
  {32'h3eac8af7, 32'hbdcc8709} /* (12, 17, 27) {real, imag} */,
  {32'h3cd007e4, 32'hbdac40b0} /* (12, 17, 26) {real, imag} */,
  {32'hbde7a44d, 32'h3bcf8860} /* (12, 17, 25) {real, imag} */,
  {32'hbac53a00, 32'h3c9feaae} /* (12, 17, 24) {real, imag} */,
  {32'hbdb47806, 32'h3dd75d19} /* (12, 17, 23) {real, imag} */,
  {32'hbd2cc61e, 32'hbcb17276} /* (12, 17, 22) {real, imag} */,
  {32'h3d8a28ce, 32'h3c65559a} /* (12, 17, 21) {real, imag} */,
  {32'hbd4ee68b, 32'hbc5b3ed6} /* (12, 17, 20) {real, imag} */,
  {32'h3d11c668, 32'hbd6d9096} /* (12, 17, 19) {real, imag} */,
  {32'hbd3e7b43, 32'hbda870c7} /* (12, 17, 18) {real, imag} */,
  {32'hbd3656be, 32'h3ce4b494} /* (12, 17, 17) {real, imag} */,
  {32'hbd307148, 32'h00000000} /* (12, 17, 16) {real, imag} */,
  {32'hbd3656be, 32'hbce4b494} /* (12, 17, 15) {real, imag} */,
  {32'hbd3e7b43, 32'h3da870c7} /* (12, 17, 14) {real, imag} */,
  {32'h3d11c668, 32'h3d6d9096} /* (12, 17, 13) {real, imag} */,
  {32'hbd4ee68b, 32'h3c5b3ed6} /* (12, 17, 12) {real, imag} */,
  {32'h3d8a28ce, 32'hbc65559a} /* (12, 17, 11) {real, imag} */,
  {32'hbd2cc61e, 32'h3cb17276} /* (12, 17, 10) {real, imag} */,
  {32'hbdb47806, 32'hbdd75d19} /* (12, 17, 9) {real, imag} */,
  {32'hbac53a00, 32'hbc9feaae} /* (12, 17, 8) {real, imag} */,
  {32'hbde7a44d, 32'hbbcf8860} /* (12, 17, 7) {real, imag} */,
  {32'h3cd007e4, 32'h3dac40b0} /* (12, 17, 6) {real, imag} */,
  {32'h3eac8af7, 32'h3dcc8709} /* (12, 17, 5) {real, imag} */,
  {32'h3d1f3cfc, 32'hbda1cdb6} /* (12, 17, 4) {real, imag} */,
  {32'h3de237ab, 32'hbc3c84c2} /* (12, 17, 3) {real, imag} */,
  {32'h3fbbf0e9, 32'h3e6fd60a} /* (12, 17, 2) {real, imag} */,
  {32'hc06c6054, 32'hbefe8a6d} /* (12, 17, 1) {real, imag} */,
  {32'hc036137e, 32'h00000000} /* (12, 17, 0) {real, imag} */,
  {32'hc07fd375, 32'h3f04760e} /* (12, 16, 31) {real, imag} */,
  {32'h3fc2a904, 32'hbe5c3a96} /* (12, 16, 30) {real, imag} */,
  {32'h3d573853, 32'hbdc91d08} /* (12, 16, 29) {real, imag} */,
  {32'hbe6569f0, 32'h3dcb0b0a} /* (12, 16, 28) {real, imag} */,
  {32'h3e817905, 32'h3d5700b0} /* (12, 16, 27) {real, imag} */,
  {32'hbd90e458, 32'hbc9a5346} /* (12, 16, 26) {real, imag} */,
  {32'hbd857760, 32'hbc5a2ecc} /* (12, 16, 25) {real, imag} */,
  {32'h3dbfb4e1, 32'h3d18e2fc} /* (12, 16, 24) {real, imag} */,
  {32'hbdb810b0, 32'hbd766848} /* (12, 16, 23) {real, imag} */,
  {32'hbd9b5d4c, 32'hbd4db47b} /* (12, 16, 22) {real, imag} */,
  {32'hbd3713b4, 32'hbdc1a592} /* (12, 16, 21) {real, imag} */,
  {32'h3d1a701d, 32'hbd905dbb} /* (12, 16, 20) {real, imag} */,
  {32'hbcf75645, 32'h3b4c8330} /* (12, 16, 19) {real, imag} */,
  {32'h3d6fee55, 32'hbcf96acc} /* (12, 16, 18) {real, imag} */,
  {32'hbcc1a800, 32'hbd5aaa66} /* (12, 16, 17) {real, imag} */,
  {32'h3d90c604, 32'h00000000} /* (12, 16, 16) {real, imag} */,
  {32'hbcc1a800, 32'h3d5aaa66} /* (12, 16, 15) {real, imag} */,
  {32'h3d6fee55, 32'h3cf96acc} /* (12, 16, 14) {real, imag} */,
  {32'hbcf75645, 32'hbb4c8330} /* (12, 16, 13) {real, imag} */,
  {32'h3d1a701d, 32'h3d905dbb} /* (12, 16, 12) {real, imag} */,
  {32'hbd3713b4, 32'h3dc1a592} /* (12, 16, 11) {real, imag} */,
  {32'hbd9b5d4c, 32'h3d4db47b} /* (12, 16, 10) {real, imag} */,
  {32'hbdb810b0, 32'h3d766848} /* (12, 16, 9) {real, imag} */,
  {32'h3dbfb4e1, 32'hbd18e2fc} /* (12, 16, 8) {real, imag} */,
  {32'hbd857760, 32'h3c5a2ecc} /* (12, 16, 7) {real, imag} */,
  {32'hbd90e458, 32'h3c9a5346} /* (12, 16, 6) {real, imag} */,
  {32'h3e817905, 32'hbd5700b0} /* (12, 16, 5) {real, imag} */,
  {32'hbe6569f0, 32'hbdcb0b0a} /* (12, 16, 4) {real, imag} */,
  {32'h3d573853, 32'h3dc91d08} /* (12, 16, 3) {real, imag} */,
  {32'h3fc2a904, 32'h3e5c3a96} /* (12, 16, 2) {real, imag} */,
  {32'hc07fd375, 32'hbf04760e} /* (12, 16, 1) {real, imag} */,
  {32'hc03d5b76, 32'h00000000} /* (12, 16, 0) {real, imag} */,
  {32'hc08030aa, 32'h3ee639d3} /* (12, 15, 31) {real, imag} */,
  {32'h3fb6392b, 32'hbe35350a} /* (12, 15, 30) {real, imag} */,
  {32'h3d767e06, 32'hbd5fbce4} /* (12, 15, 29) {real, imag} */,
  {32'hbe6a1985, 32'h3da2028a} /* (12, 15, 28) {real, imag} */,
  {32'h3dbe9265, 32'hbda35a27} /* (12, 15, 27) {real, imag} */,
  {32'hbd93c2a6, 32'hbd95787a} /* (12, 15, 26) {real, imag} */,
  {32'hbd4b2dfe, 32'hbdc0d77c} /* (12, 15, 25) {real, imag} */,
  {32'hbd2d1730, 32'h3c25f00a} /* (12, 15, 24) {real, imag} */,
  {32'hbdb77566, 32'h3d3d9286} /* (12, 15, 23) {real, imag} */,
  {32'hbd5fe576, 32'h3cfc8c62} /* (12, 15, 22) {real, imag} */,
  {32'h3c859a1a, 32'hbc9f4e99} /* (12, 15, 21) {real, imag} */,
  {32'hbc84d00e, 32'hbd829c26} /* (12, 15, 20) {real, imag} */,
  {32'h3c313ac0, 32'hbd85cb51} /* (12, 15, 19) {real, imag} */,
  {32'h3c0f8ea0, 32'hbcd1c81d} /* (12, 15, 18) {real, imag} */,
  {32'hbd5c7326, 32'hbc234bcf} /* (12, 15, 17) {real, imag} */,
  {32'hbdb7e92a, 32'h00000000} /* (12, 15, 16) {real, imag} */,
  {32'hbd5c7326, 32'h3c234bcf} /* (12, 15, 15) {real, imag} */,
  {32'h3c0f8ea0, 32'h3cd1c81d} /* (12, 15, 14) {real, imag} */,
  {32'h3c313ac0, 32'h3d85cb51} /* (12, 15, 13) {real, imag} */,
  {32'hbc84d00e, 32'h3d829c26} /* (12, 15, 12) {real, imag} */,
  {32'h3c859a1a, 32'h3c9f4e99} /* (12, 15, 11) {real, imag} */,
  {32'hbd5fe576, 32'hbcfc8c62} /* (12, 15, 10) {real, imag} */,
  {32'hbdb77566, 32'hbd3d9286} /* (12, 15, 9) {real, imag} */,
  {32'hbd2d1730, 32'hbc25f00a} /* (12, 15, 8) {real, imag} */,
  {32'hbd4b2dfe, 32'h3dc0d77c} /* (12, 15, 7) {real, imag} */,
  {32'hbd93c2a6, 32'h3d95787a} /* (12, 15, 6) {real, imag} */,
  {32'h3dbe9265, 32'h3da35a27} /* (12, 15, 5) {real, imag} */,
  {32'hbe6a1985, 32'hbda2028a} /* (12, 15, 4) {real, imag} */,
  {32'h3d767e06, 32'h3d5fbce4} /* (12, 15, 3) {real, imag} */,
  {32'h3fb6392b, 32'h3e35350a} /* (12, 15, 2) {real, imag} */,
  {32'hc08030aa, 32'hbee639d3} /* (12, 15, 1) {real, imag} */,
  {32'hc044275e, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'hc076f82f, 32'h3ebf44c2} /* (12, 14, 31) {real, imag} */,
  {32'h3fa846ec, 32'hbe7a9ce6} /* (12, 14, 30) {real, imag} */,
  {32'h3c9b9f08, 32'h3dae4e8a} /* (12, 14, 29) {real, imag} */,
  {32'hbe879cbd, 32'h3e207894} /* (12, 14, 28) {real, imag} */,
  {32'hbdb37a30, 32'hbe33d408} /* (12, 14, 27) {real, imag} */,
  {32'hbd7dc5d6, 32'hbe46b52c} /* (12, 14, 26) {real, imag} */,
  {32'hbd266de1, 32'h3cbc3352} /* (12, 14, 25) {real, imag} */,
  {32'h3cffda32, 32'hbc1c4fe4} /* (12, 14, 24) {real, imag} */,
  {32'hbb9cbc88, 32'h3c07be56} /* (12, 14, 23) {real, imag} */,
  {32'hbd925afc, 32'hbd6ff2be} /* (12, 14, 22) {real, imag} */,
  {32'h3d531925, 32'hbe102bcf} /* (12, 14, 21) {real, imag} */,
  {32'hbc0438be, 32'hbca1723d} /* (12, 14, 20) {real, imag} */,
  {32'h3d826a16, 32'h3cd4ef00} /* (12, 14, 19) {real, imag} */,
  {32'hbd1eac3e, 32'hbd4b4029} /* (12, 14, 18) {real, imag} */,
  {32'hbb014758, 32'h3c835d1c} /* (12, 14, 17) {real, imag} */,
  {32'h3cb737d6, 32'h00000000} /* (12, 14, 16) {real, imag} */,
  {32'hbb014758, 32'hbc835d1c} /* (12, 14, 15) {real, imag} */,
  {32'hbd1eac3e, 32'h3d4b4029} /* (12, 14, 14) {real, imag} */,
  {32'h3d826a16, 32'hbcd4ef00} /* (12, 14, 13) {real, imag} */,
  {32'hbc0438be, 32'h3ca1723d} /* (12, 14, 12) {real, imag} */,
  {32'h3d531925, 32'h3e102bcf} /* (12, 14, 11) {real, imag} */,
  {32'hbd925afc, 32'h3d6ff2be} /* (12, 14, 10) {real, imag} */,
  {32'hbb9cbc88, 32'hbc07be56} /* (12, 14, 9) {real, imag} */,
  {32'h3cffda32, 32'h3c1c4fe4} /* (12, 14, 8) {real, imag} */,
  {32'hbd266de1, 32'hbcbc3352} /* (12, 14, 7) {real, imag} */,
  {32'hbd7dc5d6, 32'h3e46b52c} /* (12, 14, 6) {real, imag} */,
  {32'hbdb37a30, 32'h3e33d408} /* (12, 14, 5) {real, imag} */,
  {32'hbe879cbd, 32'hbe207894} /* (12, 14, 4) {real, imag} */,
  {32'h3c9b9f08, 32'hbdae4e8a} /* (12, 14, 3) {real, imag} */,
  {32'h3fa846ec, 32'h3e7a9ce6} /* (12, 14, 2) {real, imag} */,
  {32'hc076f82f, 32'hbebf44c2} /* (12, 14, 1) {real, imag} */,
  {32'hc035be81, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'hc058e24b, 32'h3e9704c8} /* (12, 13, 31) {real, imag} */,
  {32'h3f8f9cb0, 32'hbe44e0df} /* (12, 13, 30) {real, imag} */,
  {32'hbe01c3a6, 32'h3ceae699} /* (12, 13, 29) {real, imag} */,
  {32'hbe45344a, 32'h3e67fa72} /* (12, 13, 28) {real, imag} */,
  {32'h3e713c95, 32'hbde06428} /* (12, 13, 27) {real, imag} */,
  {32'h3d39dee5, 32'hbdfc5c32} /* (12, 13, 26) {real, imag} */,
  {32'h3c827e4e, 32'hbd07396a} /* (12, 13, 25) {real, imag} */,
  {32'hbc6adc30, 32'hbd5f9244} /* (12, 13, 24) {real, imag} */,
  {32'h3d582a54, 32'hbbecad20} /* (12, 13, 23) {real, imag} */,
  {32'hbd00a19a, 32'h3ad62c00} /* (12, 13, 22) {real, imag} */,
  {32'h3e37cc58, 32'hbe01aa15} /* (12, 13, 21) {real, imag} */,
  {32'h3d268746, 32'hbcd42e60} /* (12, 13, 20) {real, imag} */,
  {32'hbd815c3c, 32'h3d0c3a6a} /* (12, 13, 19) {real, imag} */,
  {32'h3c62c268, 32'hbb928f40} /* (12, 13, 18) {real, imag} */,
  {32'hbd84a976, 32'hbcc4f144} /* (12, 13, 17) {real, imag} */,
  {32'hbc0738fe, 32'h00000000} /* (12, 13, 16) {real, imag} */,
  {32'hbd84a976, 32'h3cc4f144} /* (12, 13, 15) {real, imag} */,
  {32'h3c62c268, 32'h3b928f40} /* (12, 13, 14) {real, imag} */,
  {32'hbd815c3c, 32'hbd0c3a6a} /* (12, 13, 13) {real, imag} */,
  {32'h3d268746, 32'h3cd42e60} /* (12, 13, 12) {real, imag} */,
  {32'h3e37cc58, 32'h3e01aa15} /* (12, 13, 11) {real, imag} */,
  {32'hbd00a19a, 32'hbad62c00} /* (12, 13, 10) {real, imag} */,
  {32'h3d582a54, 32'h3becad20} /* (12, 13, 9) {real, imag} */,
  {32'hbc6adc30, 32'h3d5f9244} /* (12, 13, 8) {real, imag} */,
  {32'h3c827e4e, 32'h3d07396a} /* (12, 13, 7) {real, imag} */,
  {32'h3d39dee5, 32'h3dfc5c32} /* (12, 13, 6) {real, imag} */,
  {32'h3e713c95, 32'h3de06428} /* (12, 13, 5) {real, imag} */,
  {32'hbe45344a, 32'hbe67fa72} /* (12, 13, 4) {real, imag} */,
  {32'hbe01c3a6, 32'hbceae699} /* (12, 13, 3) {real, imag} */,
  {32'h3f8f9cb0, 32'h3e44e0df} /* (12, 13, 2) {real, imag} */,
  {32'hc058e24b, 32'hbe9704c8} /* (12, 13, 1) {real, imag} */,
  {32'hc0143ef8, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'hc02a58cd, 32'hbd617d50} /* (12, 12, 31) {real, imag} */,
  {32'h3f85598e, 32'hbdbebf0a} /* (12, 12, 30) {real, imag} */,
  {32'hbd4c0223, 32'h3d29de97} /* (12, 12, 29) {real, imag} */,
  {32'hbd4c5052, 32'h3e72cc84} /* (12, 12, 28) {real, imag} */,
  {32'h3e15a5de, 32'hbd0e7e88} /* (12, 12, 27) {real, imag} */,
  {32'h3d756748, 32'h3cb6d3b1} /* (12, 12, 26) {real, imag} */,
  {32'hbbfeab08, 32'hbdb89063} /* (12, 12, 25) {real, imag} */,
  {32'h3d7aa519, 32'hbcce50da} /* (12, 12, 24) {real, imag} */,
  {32'h3da574a1, 32'h3e067210} /* (12, 12, 23) {real, imag} */,
  {32'h3d33282c, 32'h3dc01637} /* (12, 12, 22) {real, imag} */,
  {32'hbb4eb9e0, 32'hbd6f9283} /* (12, 12, 21) {real, imag} */,
  {32'h3c7f5746, 32'hbcf0a341} /* (12, 12, 20) {real, imag} */,
  {32'hbc6c1e6a, 32'hbb69cb40} /* (12, 12, 19) {real, imag} */,
  {32'h3d57e6d6, 32'hbd3e93f1} /* (12, 12, 18) {real, imag} */,
  {32'h3cb2eba1, 32'hbcacb0f4} /* (12, 12, 17) {real, imag} */,
  {32'h3d85014a, 32'h00000000} /* (12, 12, 16) {real, imag} */,
  {32'h3cb2eba1, 32'h3cacb0f4} /* (12, 12, 15) {real, imag} */,
  {32'h3d57e6d6, 32'h3d3e93f1} /* (12, 12, 14) {real, imag} */,
  {32'hbc6c1e6a, 32'h3b69cb40} /* (12, 12, 13) {real, imag} */,
  {32'h3c7f5746, 32'h3cf0a341} /* (12, 12, 12) {real, imag} */,
  {32'hbb4eb9e0, 32'h3d6f9283} /* (12, 12, 11) {real, imag} */,
  {32'h3d33282c, 32'hbdc01637} /* (12, 12, 10) {real, imag} */,
  {32'h3da574a1, 32'hbe067210} /* (12, 12, 9) {real, imag} */,
  {32'h3d7aa519, 32'h3cce50da} /* (12, 12, 8) {real, imag} */,
  {32'hbbfeab08, 32'h3db89063} /* (12, 12, 7) {real, imag} */,
  {32'h3d756748, 32'hbcb6d3b1} /* (12, 12, 6) {real, imag} */,
  {32'h3e15a5de, 32'h3d0e7e88} /* (12, 12, 5) {real, imag} */,
  {32'hbd4c5052, 32'hbe72cc84} /* (12, 12, 4) {real, imag} */,
  {32'hbd4c0223, 32'hbd29de97} /* (12, 12, 3) {real, imag} */,
  {32'h3f85598e, 32'h3dbebf0a} /* (12, 12, 2) {real, imag} */,
  {32'hc02a58cd, 32'h3d617d50} /* (12, 12, 1) {real, imag} */,
  {32'hbfc60e37, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'hbfa7e048, 32'hbebef370} /* (12, 11, 31) {real, imag} */,
  {32'h3f27fb40, 32'hbdc6f88c} /* (12, 11, 30) {real, imag} */,
  {32'hbd1c17c3, 32'h3ce38241} /* (12, 11, 29) {real, imag} */,
  {32'hbe416198, 32'h3db93cde} /* (12, 11, 28) {real, imag} */,
  {32'h3e0f6d1a, 32'hbc02b71c} /* (12, 11, 27) {real, imag} */,
  {32'hbd67fd0c, 32'hbc8d37f3} /* (12, 11, 26) {real, imag} */,
  {32'hbde30d0e, 32'hbd47b4b0} /* (12, 11, 25) {real, imag} */,
  {32'hbbd2f280, 32'hbce50464} /* (12, 11, 24) {real, imag} */,
  {32'h3dfef6da, 32'hbb9eb7ca} /* (12, 11, 23) {real, imag} */,
  {32'h3afd4278, 32'h3c093528} /* (12, 11, 22) {real, imag} */,
  {32'hb9274f00, 32'hbe0aed68} /* (12, 11, 21) {real, imag} */,
  {32'h3d624eb4, 32'hbcc81030} /* (12, 11, 20) {real, imag} */,
  {32'h3c83c1c8, 32'h399f3940} /* (12, 11, 19) {real, imag} */,
  {32'hbd2b3280, 32'hbd600ab4} /* (12, 11, 18) {real, imag} */,
  {32'hbd33e1e8, 32'hbc872caa} /* (12, 11, 17) {real, imag} */,
  {32'hbd4ccb0a, 32'h00000000} /* (12, 11, 16) {real, imag} */,
  {32'hbd33e1e8, 32'h3c872caa} /* (12, 11, 15) {real, imag} */,
  {32'hbd2b3280, 32'h3d600ab4} /* (12, 11, 14) {real, imag} */,
  {32'h3c83c1c8, 32'hb99f3940} /* (12, 11, 13) {real, imag} */,
  {32'h3d624eb4, 32'h3cc81030} /* (12, 11, 12) {real, imag} */,
  {32'hb9274f00, 32'h3e0aed68} /* (12, 11, 11) {real, imag} */,
  {32'h3afd4278, 32'hbc093528} /* (12, 11, 10) {real, imag} */,
  {32'h3dfef6da, 32'h3b9eb7ca} /* (12, 11, 9) {real, imag} */,
  {32'hbbd2f280, 32'h3ce50464} /* (12, 11, 8) {real, imag} */,
  {32'hbde30d0e, 32'h3d47b4b0} /* (12, 11, 7) {real, imag} */,
  {32'hbd67fd0c, 32'h3c8d37f3} /* (12, 11, 6) {real, imag} */,
  {32'h3e0f6d1a, 32'h3c02b71c} /* (12, 11, 5) {real, imag} */,
  {32'hbe416198, 32'hbdb93cde} /* (12, 11, 4) {real, imag} */,
  {32'hbd1c17c3, 32'hbce38241} /* (12, 11, 3) {real, imag} */,
  {32'h3f27fb40, 32'h3dc6f88c} /* (12, 11, 2) {real, imag} */,
  {32'hbfa7e048, 32'h3ebef370} /* (12, 11, 1) {real, imag} */,
  {32'hbebd3d1a, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'h3f032b2f, 32'hbf0d2dc0} /* (12, 10, 31) {real, imag} */,
  {32'hbdd05c28, 32'h3d97e4b4} /* (12, 10, 30) {real, imag} */,
  {32'hbe3d5562, 32'h3c2da794} /* (12, 10, 29) {real, imag} */,
  {32'hbd0d48b8, 32'hbcab1dc0} /* (12, 10, 28) {real, imag} */,
  {32'h3d214f78, 32'h3cd74180} /* (12, 10, 27) {real, imag} */,
  {32'h3d298a38, 32'h3d44ac49} /* (12, 10, 26) {real, imag} */,
  {32'h3dc89c1b, 32'h3c54282c} /* (12, 10, 25) {real, imag} */,
  {32'h3d79be70, 32'h3d940c50} /* (12, 10, 24) {real, imag} */,
  {32'hbc543080, 32'h3ce38894} /* (12, 10, 23) {real, imag} */,
  {32'hbdfae425, 32'h3d0d0be0} /* (12, 10, 22) {real, imag} */,
  {32'hbd382064, 32'h3acac050} /* (12, 10, 21) {real, imag} */,
  {32'h3c4ff688, 32'h3d801dec} /* (12, 10, 20) {real, imag} */,
  {32'h3de095ff, 32'hbd5b0884} /* (12, 10, 19) {real, imag} */,
  {32'h3cb5426c, 32'h3dd19595} /* (12, 10, 18) {real, imag} */,
  {32'hbceb2067, 32'hbc6ed289} /* (12, 10, 17) {real, imag} */,
  {32'hbc2df750, 32'h00000000} /* (12, 10, 16) {real, imag} */,
  {32'hbceb2067, 32'h3c6ed289} /* (12, 10, 15) {real, imag} */,
  {32'h3cb5426c, 32'hbdd19595} /* (12, 10, 14) {real, imag} */,
  {32'h3de095ff, 32'h3d5b0884} /* (12, 10, 13) {real, imag} */,
  {32'h3c4ff688, 32'hbd801dec} /* (12, 10, 12) {real, imag} */,
  {32'hbd382064, 32'hbacac050} /* (12, 10, 11) {real, imag} */,
  {32'hbdfae425, 32'hbd0d0be0} /* (12, 10, 10) {real, imag} */,
  {32'hbc543080, 32'hbce38894} /* (12, 10, 9) {real, imag} */,
  {32'h3d79be70, 32'hbd940c50} /* (12, 10, 8) {real, imag} */,
  {32'h3dc89c1b, 32'hbc54282c} /* (12, 10, 7) {real, imag} */,
  {32'h3d298a38, 32'hbd44ac49} /* (12, 10, 6) {real, imag} */,
  {32'h3d214f78, 32'hbcd74180} /* (12, 10, 5) {real, imag} */,
  {32'hbd0d48b8, 32'h3cab1dc0} /* (12, 10, 4) {real, imag} */,
  {32'hbe3d5562, 32'hbc2da794} /* (12, 10, 3) {real, imag} */,
  {32'hbdd05c28, 32'hbd97e4b4} /* (12, 10, 2) {real, imag} */,
  {32'h3f032b2f, 32'h3f0d2dc0} /* (12, 10, 1) {real, imag} */,
  {32'h3f94d5db, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h3fd7d9d2, 32'hbf6ecea6} /* (12, 9, 31) {real, imag} */,
  {32'hbf458c21, 32'h3e7568fd} /* (12, 9, 30) {real, imag} */,
  {32'hbda2aab1, 32'hbd6516f6} /* (12, 9, 29) {real, imag} */,
  {32'h3dd8df02, 32'hbcb0e5d8} /* (12, 9, 28) {real, imag} */,
  {32'hbd51782c, 32'h3dcf0d18} /* (12, 9, 27) {real, imag} */,
  {32'h3c6ff214, 32'h3c13ddfe} /* (12, 9, 26) {real, imag} */,
  {32'h3d2856c4, 32'h3cab57e4} /* (12, 9, 25) {real, imag} */,
  {32'h3cfab33d, 32'h3d413d86} /* (12, 9, 24) {real, imag} */,
  {32'hbbfe01c8, 32'h389a3400} /* (12, 9, 23) {real, imag} */,
  {32'hbda85936, 32'hbd64d036} /* (12, 9, 22) {real, imag} */,
  {32'hbc0f6e9c, 32'h3bdca45c} /* (12, 9, 21) {real, imag} */,
  {32'hbd0c97ac, 32'h3ae08340} /* (12, 9, 20) {real, imag} */,
  {32'hbcb43345, 32'h3d638dea} /* (12, 9, 19) {real, imag} */,
  {32'hbd9b33aa, 32'h3d888ca6} /* (12, 9, 18) {real, imag} */,
  {32'hbce7efa3, 32'h3c766c7a} /* (12, 9, 17) {real, imag} */,
  {32'hbc3a550b, 32'h00000000} /* (12, 9, 16) {real, imag} */,
  {32'hbce7efa3, 32'hbc766c7a} /* (12, 9, 15) {real, imag} */,
  {32'hbd9b33aa, 32'hbd888ca6} /* (12, 9, 14) {real, imag} */,
  {32'hbcb43345, 32'hbd638dea} /* (12, 9, 13) {real, imag} */,
  {32'hbd0c97ac, 32'hbae08340} /* (12, 9, 12) {real, imag} */,
  {32'hbc0f6e9c, 32'hbbdca45c} /* (12, 9, 11) {real, imag} */,
  {32'hbda85936, 32'h3d64d036} /* (12, 9, 10) {real, imag} */,
  {32'hbbfe01c8, 32'hb89a3400} /* (12, 9, 9) {real, imag} */,
  {32'h3cfab33d, 32'hbd413d86} /* (12, 9, 8) {real, imag} */,
  {32'h3d2856c4, 32'hbcab57e4} /* (12, 9, 7) {real, imag} */,
  {32'h3c6ff214, 32'hbc13ddfe} /* (12, 9, 6) {real, imag} */,
  {32'hbd51782c, 32'hbdcf0d18} /* (12, 9, 5) {real, imag} */,
  {32'h3dd8df02, 32'h3cb0e5d8} /* (12, 9, 4) {real, imag} */,
  {32'hbda2aab1, 32'h3d6516f6} /* (12, 9, 3) {real, imag} */,
  {32'hbf458c21, 32'hbe7568fd} /* (12, 9, 2) {real, imag} */,
  {32'h3fd7d9d2, 32'h3f6ecea6} /* (12, 9, 1) {real, imag} */,
  {32'h400f6fc7, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'h4018b00e, 32'hbfa86951} /* (12, 8, 31) {real, imag} */,
  {32'hbf8d1383, 32'h3eb8aa0d} /* (12, 8, 30) {real, imag} */,
  {32'hbc18c42c, 32'h3b0d02b0} /* (12, 8, 29) {real, imag} */,
  {32'h3d921f54, 32'hbc803d20} /* (12, 8, 28) {real, imag} */,
  {32'hbd8ca2ed, 32'hbc5604d0} /* (12, 8, 27) {real, imag} */,
  {32'hbd088ffa, 32'h3d995f14} /* (12, 8, 26) {real, imag} */,
  {32'h3dba8aa0, 32'hbc6ef97a} /* (12, 8, 25) {real, imag} */,
  {32'h3d851e5c, 32'h3d6bb588} /* (12, 8, 24) {real, imag} */,
  {32'h3c4b591c, 32'hbdda00a7} /* (12, 8, 23) {real, imag} */,
  {32'hbcb171f8, 32'h3d52e765} /* (12, 8, 22) {real, imag} */,
  {32'hbd1eaa25, 32'h3dc227f7} /* (12, 8, 21) {real, imag} */,
  {32'h3dab1ff1, 32'hbdb99c77} /* (12, 8, 20) {real, imag} */,
  {32'hbe0df228, 32'hbd82181b} /* (12, 8, 19) {real, imag} */,
  {32'hbd35d4e2, 32'h3e006396} /* (12, 8, 18) {real, imag} */,
  {32'h3ce2c23d, 32'h3d31466a} /* (12, 8, 17) {real, imag} */,
  {32'h3d258655, 32'h00000000} /* (12, 8, 16) {real, imag} */,
  {32'h3ce2c23d, 32'hbd31466a} /* (12, 8, 15) {real, imag} */,
  {32'hbd35d4e2, 32'hbe006396} /* (12, 8, 14) {real, imag} */,
  {32'hbe0df228, 32'h3d82181b} /* (12, 8, 13) {real, imag} */,
  {32'h3dab1ff1, 32'h3db99c77} /* (12, 8, 12) {real, imag} */,
  {32'hbd1eaa25, 32'hbdc227f7} /* (12, 8, 11) {real, imag} */,
  {32'hbcb171f8, 32'hbd52e765} /* (12, 8, 10) {real, imag} */,
  {32'h3c4b591c, 32'h3dda00a7} /* (12, 8, 9) {real, imag} */,
  {32'h3d851e5c, 32'hbd6bb588} /* (12, 8, 8) {real, imag} */,
  {32'h3dba8aa0, 32'h3c6ef97a} /* (12, 8, 7) {real, imag} */,
  {32'hbd088ffa, 32'hbd995f14} /* (12, 8, 6) {real, imag} */,
  {32'hbd8ca2ed, 32'h3c5604d0} /* (12, 8, 5) {real, imag} */,
  {32'h3d921f54, 32'h3c803d20} /* (12, 8, 4) {real, imag} */,
  {32'hbc18c42c, 32'hbb0d02b0} /* (12, 8, 3) {real, imag} */,
  {32'hbf8d1383, 32'hbeb8aa0d} /* (12, 8, 2) {real, imag} */,
  {32'h4018b00e, 32'h3fa86951} /* (12, 8, 1) {real, imag} */,
  {32'h40459d50, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'h403e2617, 32'hbfc2854b} /* (12, 7, 31) {real, imag} */,
  {32'hbf80ffb2, 32'h3f2e5b4e} /* (12, 7, 30) {real, imag} */,
  {32'hbd66e1be, 32'h3c99dce3} /* (12, 7, 29) {real, imag} */,
  {32'h3d25e830, 32'hbccb8c36} /* (12, 7, 28) {real, imag} */,
  {32'hbe4efa0d, 32'h3de42cd6} /* (12, 7, 27) {real, imag} */,
  {32'hbc379c70, 32'hbbd60020} /* (12, 7, 26) {real, imag} */,
  {32'h3d79df14, 32'hbe18d811} /* (12, 7, 25) {real, imag} */,
  {32'hbc4ba194, 32'h3df23279} /* (12, 7, 24) {real, imag} */,
  {32'h3d712840, 32'hbd846928} /* (12, 7, 23) {real, imag} */,
  {32'hbd1e3680, 32'h3e38246d} /* (12, 7, 22) {real, imag} */,
  {32'hbdfa98d2, 32'h3d3cd110} /* (12, 7, 21) {real, imag} */,
  {32'h3d098933, 32'h3b26bc60} /* (12, 7, 20) {real, imag} */,
  {32'hbd33649f, 32'h3cc61e58} /* (12, 7, 19) {real, imag} */,
  {32'hbd27531e, 32'hbcea7c4b} /* (12, 7, 18) {real, imag} */,
  {32'h3cb3dd4c, 32'hbdbfcdec} /* (12, 7, 17) {real, imag} */,
  {32'h3d9d9584, 32'h00000000} /* (12, 7, 16) {real, imag} */,
  {32'h3cb3dd4c, 32'h3dbfcdec} /* (12, 7, 15) {real, imag} */,
  {32'hbd27531e, 32'h3cea7c4b} /* (12, 7, 14) {real, imag} */,
  {32'hbd33649f, 32'hbcc61e58} /* (12, 7, 13) {real, imag} */,
  {32'h3d098933, 32'hbb26bc60} /* (12, 7, 12) {real, imag} */,
  {32'hbdfa98d2, 32'hbd3cd110} /* (12, 7, 11) {real, imag} */,
  {32'hbd1e3680, 32'hbe38246d} /* (12, 7, 10) {real, imag} */,
  {32'h3d712840, 32'h3d846928} /* (12, 7, 9) {real, imag} */,
  {32'hbc4ba194, 32'hbdf23279} /* (12, 7, 8) {real, imag} */,
  {32'h3d79df14, 32'h3e18d811} /* (12, 7, 7) {real, imag} */,
  {32'hbc379c70, 32'h3bd60020} /* (12, 7, 6) {real, imag} */,
  {32'hbe4efa0d, 32'hbde42cd6} /* (12, 7, 5) {real, imag} */,
  {32'h3d25e830, 32'h3ccb8c36} /* (12, 7, 4) {real, imag} */,
  {32'hbd66e1be, 32'hbc99dce3} /* (12, 7, 3) {real, imag} */,
  {32'hbf80ffb2, 32'hbf2e5b4e} /* (12, 7, 2) {real, imag} */,
  {32'h403e2617, 32'h3fc2854b} /* (12, 7, 1) {real, imag} */,
  {32'h406419cd, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'h404822df, 32'hc003120f} /* (12, 6, 31) {real, imag} */,
  {32'hbf56e734, 32'h3f6156a6} /* (12, 6, 30) {real, imag} */,
  {32'hbd527f4a, 32'h3d911164} /* (12, 6, 29) {real, imag} */,
  {32'h3cf5dc50, 32'h3d3a2e6c} /* (12, 6, 28) {real, imag} */,
  {32'hbdbfccbc, 32'h3e5d57c3} /* (12, 6, 27) {real, imag} */,
  {32'hbd06d749, 32'h3cce791a} /* (12, 6, 26) {real, imag} */,
  {32'hbd8471e3, 32'hbd9a7386} /* (12, 6, 25) {real, imag} */,
  {32'hbc9687c1, 32'h3cbc665c} /* (12, 6, 24) {real, imag} */,
  {32'h3d1d540c, 32'h3db189b4} /* (12, 6, 23) {real, imag} */,
  {32'hbdaf6567, 32'hbd8edd93} /* (12, 6, 22) {real, imag} */,
  {32'h3ca4ecc6, 32'hbc04cc90} /* (12, 6, 21) {real, imag} */,
  {32'hbd2fcd4f, 32'hbd41136e} /* (12, 6, 20) {real, imag} */,
  {32'h3d80840c, 32'h3cde3afe} /* (12, 6, 19) {real, imag} */,
  {32'hbdbdab36, 32'h3c76e524} /* (12, 6, 18) {real, imag} */,
  {32'h3d815cce, 32'hbb83f24a} /* (12, 6, 17) {real, imag} */,
  {32'hbdab2299, 32'h00000000} /* (12, 6, 16) {real, imag} */,
  {32'h3d815cce, 32'h3b83f24a} /* (12, 6, 15) {real, imag} */,
  {32'hbdbdab36, 32'hbc76e524} /* (12, 6, 14) {real, imag} */,
  {32'h3d80840c, 32'hbcde3afe} /* (12, 6, 13) {real, imag} */,
  {32'hbd2fcd4f, 32'h3d41136e} /* (12, 6, 12) {real, imag} */,
  {32'h3ca4ecc6, 32'h3c04cc90} /* (12, 6, 11) {real, imag} */,
  {32'hbdaf6567, 32'h3d8edd93} /* (12, 6, 10) {real, imag} */,
  {32'h3d1d540c, 32'hbdb189b4} /* (12, 6, 9) {real, imag} */,
  {32'hbc9687c1, 32'hbcbc665c} /* (12, 6, 8) {real, imag} */,
  {32'hbd8471e3, 32'h3d9a7386} /* (12, 6, 7) {real, imag} */,
  {32'hbd06d749, 32'hbcce791a} /* (12, 6, 6) {real, imag} */,
  {32'hbdbfccbc, 32'hbe5d57c3} /* (12, 6, 5) {real, imag} */,
  {32'h3cf5dc50, 32'hbd3a2e6c} /* (12, 6, 4) {real, imag} */,
  {32'hbd527f4a, 32'hbd911164} /* (12, 6, 3) {real, imag} */,
  {32'hbf56e734, 32'hbf6156a6} /* (12, 6, 2) {real, imag} */,
  {32'h404822df, 32'h4003120f} /* (12, 6, 1) {real, imag} */,
  {32'h4081e0b4, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'h403cc780, 32'hc0344f84} /* (12, 5, 31) {real, imag} */,
  {32'hbe98da8c, 32'h3f768e20} /* (12, 5, 30) {real, imag} */,
  {32'hbe1bc4dc, 32'h3c9560a9} /* (12, 5, 29) {real, imag} */,
  {32'hbd32d10e, 32'h3e307685} /* (12, 5, 28) {real, imag} */,
  {32'hbe344a30, 32'h3d267845} /* (12, 5, 27) {real, imag} */,
  {32'hbdb6fd54, 32'h3de42a66} /* (12, 5, 26) {real, imag} */,
  {32'h3d46b376, 32'hbd58d756} /* (12, 5, 25) {real, imag} */,
  {32'h3b2da780, 32'h3dc4dcf5} /* (12, 5, 24) {real, imag} */,
  {32'hbce36bea, 32'hbdaa9f78} /* (12, 5, 23) {real, imag} */,
  {32'h3bd8fad6, 32'h3d691ae2} /* (12, 5, 22) {real, imag} */,
  {32'h3d6da40d, 32'hbd214106} /* (12, 5, 21) {real, imag} */,
  {32'hbc347390, 32'hbd39b718} /* (12, 5, 20) {real, imag} */,
  {32'hbb7be420, 32'h3d4ad4f2} /* (12, 5, 19) {real, imag} */,
  {32'h3c0d7542, 32'h3d3cb2d8} /* (12, 5, 18) {real, imag} */,
  {32'hbd057f76, 32'hbd67ecd4} /* (12, 5, 17) {real, imag} */,
  {32'hbc02c3a6, 32'h00000000} /* (12, 5, 16) {real, imag} */,
  {32'hbd057f76, 32'h3d67ecd4} /* (12, 5, 15) {real, imag} */,
  {32'h3c0d7542, 32'hbd3cb2d8} /* (12, 5, 14) {real, imag} */,
  {32'hbb7be420, 32'hbd4ad4f2} /* (12, 5, 13) {real, imag} */,
  {32'hbc347390, 32'h3d39b718} /* (12, 5, 12) {real, imag} */,
  {32'h3d6da40d, 32'h3d214106} /* (12, 5, 11) {real, imag} */,
  {32'h3bd8fad6, 32'hbd691ae2} /* (12, 5, 10) {real, imag} */,
  {32'hbce36bea, 32'h3daa9f78} /* (12, 5, 9) {real, imag} */,
  {32'h3b2da780, 32'hbdc4dcf5} /* (12, 5, 8) {real, imag} */,
  {32'h3d46b376, 32'h3d58d756} /* (12, 5, 7) {real, imag} */,
  {32'hbdb6fd54, 32'hbde42a66} /* (12, 5, 6) {real, imag} */,
  {32'hbe344a30, 32'hbd267845} /* (12, 5, 5) {real, imag} */,
  {32'hbd32d10e, 32'hbe307685} /* (12, 5, 4) {real, imag} */,
  {32'hbe1bc4dc, 32'hbc9560a9} /* (12, 5, 3) {real, imag} */,
  {32'hbe98da8c, 32'hbf768e20} /* (12, 5, 2) {real, imag} */,
  {32'h403cc780, 32'h40344f84} /* (12, 5, 1) {real, imag} */,
  {32'h409475cf, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'h40329f66, 32'hc05a9417} /* (12, 4, 31) {real, imag} */,
  {32'h3dc0d148, 32'h3f8d91c8} /* (12, 4, 30) {real, imag} */,
  {32'hbddec352, 32'hbd5a6067} /* (12, 4, 29) {real, imag} */,
  {32'hbe19733e, 32'h3e5dbe73} /* (12, 4, 28) {real, imag} */,
  {32'hbe21f723, 32'hbb95957a} /* (12, 4, 27) {real, imag} */,
  {32'hbb4b2ecc, 32'h3d50de60} /* (12, 4, 26) {real, imag} */,
  {32'hbd7c11d5, 32'hbe115aac} /* (12, 4, 25) {real, imag} */,
  {32'hbd2dc94e, 32'h3d84047f} /* (12, 4, 24) {real, imag} */,
  {32'hbd118c63, 32'h3d297ae8} /* (12, 4, 23) {real, imag} */,
  {32'hbd98e930, 32'h3dbc38be} /* (12, 4, 22) {real, imag} */,
  {32'h3ca33f13, 32'h3d8a50e2} /* (12, 4, 21) {real, imag} */,
  {32'hbc63042d, 32'hbb3e72d8} /* (12, 4, 20) {real, imag} */,
  {32'hbce2a060, 32'h3d302edc} /* (12, 4, 19) {real, imag} */,
  {32'h3da34903, 32'hbd7f3678} /* (12, 4, 18) {real, imag} */,
  {32'hbbe91748, 32'hbd2888fc} /* (12, 4, 17) {real, imag} */,
  {32'hbc61e553, 32'h00000000} /* (12, 4, 16) {real, imag} */,
  {32'hbbe91748, 32'h3d2888fc} /* (12, 4, 15) {real, imag} */,
  {32'h3da34903, 32'h3d7f3678} /* (12, 4, 14) {real, imag} */,
  {32'hbce2a060, 32'hbd302edc} /* (12, 4, 13) {real, imag} */,
  {32'hbc63042d, 32'h3b3e72d8} /* (12, 4, 12) {real, imag} */,
  {32'h3ca33f13, 32'hbd8a50e2} /* (12, 4, 11) {real, imag} */,
  {32'hbd98e930, 32'hbdbc38be} /* (12, 4, 10) {real, imag} */,
  {32'hbd118c63, 32'hbd297ae8} /* (12, 4, 9) {real, imag} */,
  {32'hbd2dc94e, 32'hbd84047f} /* (12, 4, 8) {real, imag} */,
  {32'hbd7c11d5, 32'h3e115aac} /* (12, 4, 7) {real, imag} */,
  {32'hbb4b2ecc, 32'hbd50de60} /* (12, 4, 6) {real, imag} */,
  {32'hbe21f723, 32'h3b95957a} /* (12, 4, 5) {real, imag} */,
  {32'hbe19733e, 32'hbe5dbe73} /* (12, 4, 4) {real, imag} */,
  {32'hbddec352, 32'h3d5a6067} /* (12, 4, 3) {real, imag} */,
  {32'h3dc0d148, 32'hbf8d91c8} /* (12, 4, 2) {real, imag} */,
  {32'h40329f66, 32'h405a9417} /* (12, 4, 1) {real, imag} */,
  {32'h409d5885, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'h402f6746, 32'hc066e0d6} /* (12, 3, 31) {real, imag} */,
  {32'h3e584dd8, 32'h3f8a072c} /* (12, 3, 30) {real, imag} */,
  {32'hbd439e5e, 32'h3d86a304} /* (12, 3, 29) {real, imag} */,
  {32'hbe50dcae, 32'h3dd2ac4a} /* (12, 3, 28) {real, imag} */,
  {32'hbe8caebd, 32'hbe3b0c58} /* (12, 3, 27) {real, imag} */,
  {32'hbd9efbe4, 32'h3d19fb18} /* (12, 3, 26) {real, imag} */,
  {32'h3c50414c, 32'hbdc540d6} /* (12, 3, 25) {real, imag} */,
  {32'h3d36975d, 32'h3e1fdb4d} /* (12, 3, 24) {real, imag} */,
  {32'hbcd7fd9a, 32'h3df32f41} /* (12, 3, 23) {real, imag} */,
  {32'hbbd84ef0, 32'h3db2fc14} /* (12, 3, 22) {real, imag} */,
  {32'hbe0f8c18, 32'hbce4a8bd} /* (12, 3, 21) {real, imag} */,
  {32'hbb30c850, 32'hbd8ebb6d} /* (12, 3, 20) {real, imag} */,
  {32'h3d490af7, 32'hbd86a1a0} /* (12, 3, 19) {real, imag} */,
  {32'h3d5c1843, 32'hbd980de6} /* (12, 3, 18) {real, imag} */,
  {32'hbcb1ec21, 32'h3d1d3450} /* (12, 3, 17) {real, imag} */,
  {32'hbd36538e, 32'h00000000} /* (12, 3, 16) {real, imag} */,
  {32'hbcb1ec21, 32'hbd1d3450} /* (12, 3, 15) {real, imag} */,
  {32'h3d5c1843, 32'h3d980de6} /* (12, 3, 14) {real, imag} */,
  {32'h3d490af7, 32'h3d86a1a0} /* (12, 3, 13) {real, imag} */,
  {32'hbb30c850, 32'h3d8ebb6d} /* (12, 3, 12) {real, imag} */,
  {32'hbe0f8c18, 32'h3ce4a8bd} /* (12, 3, 11) {real, imag} */,
  {32'hbbd84ef0, 32'hbdb2fc14} /* (12, 3, 10) {real, imag} */,
  {32'hbcd7fd9a, 32'hbdf32f41} /* (12, 3, 9) {real, imag} */,
  {32'h3d36975d, 32'hbe1fdb4d} /* (12, 3, 8) {real, imag} */,
  {32'h3c50414c, 32'h3dc540d6} /* (12, 3, 7) {real, imag} */,
  {32'hbd9efbe4, 32'hbd19fb18} /* (12, 3, 6) {real, imag} */,
  {32'hbe8caebd, 32'h3e3b0c58} /* (12, 3, 5) {real, imag} */,
  {32'hbe50dcae, 32'hbdd2ac4a} /* (12, 3, 4) {real, imag} */,
  {32'hbd439e5e, 32'hbd86a304} /* (12, 3, 3) {real, imag} */,
  {32'h3e584dd8, 32'hbf8a072c} /* (12, 3, 2) {real, imag} */,
  {32'h402f6746, 32'h4066e0d6} /* (12, 3, 1) {real, imag} */,
  {32'h409ee0f3, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'h403760de, 32'hc06741bf} /* (12, 2, 31) {real, imag} */,
  {32'h3e4fef2c, 32'h3f84beb1} /* (12, 2, 30) {real, imag} */,
  {32'hbe379a89, 32'h3e0e763e} /* (12, 2, 29) {real, imag} */,
  {32'hbd0d36ed, 32'h3e8c8b66} /* (12, 2, 28) {real, imag} */,
  {32'hbe6113e8, 32'hbe5815d4} /* (12, 2, 27) {real, imag} */,
  {32'hbdbd77de, 32'hbdd44e3b} /* (12, 2, 26) {real, imag} */,
  {32'h3d8b27a3, 32'h3e010385} /* (12, 2, 25) {real, imag} */,
  {32'h3dc90ff5, 32'hbcdcc79a} /* (12, 2, 24) {real, imag} */,
  {32'h3b271e28, 32'h3d7bc4a0} /* (12, 2, 23) {real, imag} */,
  {32'hbcb0fd5b, 32'h3d70cbb2} /* (12, 2, 22) {real, imag} */,
  {32'hbdd1abe5, 32'hbb6fe4fc} /* (12, 2, 21) {real, imag} */,
  {32'hbe0ccea4, 32'h3d1e61ae} /* (12, 2, 20) {real, imag} */,
  {32'hbcf1303d, 32'h3cb5f6ca} /* (12, 2, 19) {real, imag} */,
  {32'h3dcba75d, 32'hbdbde6c2} /* (12, 2, 18) {real, imag} */,
  {32'hbd69e379, 32'h3c39cea8} /* (12, 2, 17) {real, imag} */,
  {32'h3d32a3a9, 32'h00000000} /* (12, 2, 16) {real, imag} */,
  {32'hbd69e379, 32'hbc39cea8} /* (12, 2, 15) {real, imag} */,
  {32'h3dcba75d, 32'h3dbde6c2} /* (12, 2, 14) {real, imag} */,
  {32'hbcf1303d, 32'hbcb5f6ca} /* (12, 2, 13) {real, imag} */,
  {32'hbe0ccea4, 32'hbd1e61ae} /* (12, 2, 12) {real, imag} */,
  {32'hbdd1abe5, 32'h3b6fe4fc} /* (12, 2, 11) {real, imag} */,
  {32'hbcb0fd5b, 32'hbd70cbb2} /* (12, 2, 10) {real, imag} */,
  {32'h3b271e28, 32'hbd7bc4a0} /* (12, 2, 9) {real, imag} */,
  {32'h3dc90ff5, 32'h3cdcc79a} /* (12, 2, 8) {real, imag} */,
  {32'h3d8b27a3, 32'hbe010385} /* (12, 2, 7) {real, imag} */,
  {32'hbdbd77de, 32'h3dd44e3b} /* (12, 2, 6) {real, imag} */,
  {32'hbe6113e8, 32'h3e5815d4} /* (12, 2, 5) {real, imag} */,
  {32'hbd0d36ed, 32'hbe8c8b66} /* (12, 2, 4) {real, imag} */,
  {32'hbe379a89, 32'hbe0e763e} /* (12, 2, 3) {real, imag} */,
  {32'h3e4fef2c, 32'hbf84beb1} /* (12, 2, 2) {real, imag} */,
  {32'h403760de, 32'h406741bf} /* (12, 2, 1) {real, imag} */,
  {32'h40a3092f, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'h403d4878, 32'hc057b7e6} /* (12, 1, 31) {real, imag} */,
  {32'h3de6732c, 32'h3f75a3bc} /* (12, 1, 30) {real, imag} */,
  {32'hbc3b2f38, 32'h3d18c204} /* (12, 1, 29) {real, imag} */,
  {32'hbd476dc5, 32'h3ec6b49a} /* (12, 1, 28) {real, imag} */,
  {32'hbe0f828a, 32'hbe7f90f6} /* (12, 1, 27) {real, imag} */,
  {32'h3d37e3ba, 32'hbcd1d58e} /* (12, 1, 26) {real, imag} */,
  {32'hbbb1f5c8, 32'h3aab81e8} /* (12, 1, 25) {real, imag} */,
  {32'h3df7f591, 32'hbc08c313} /* (12, 1, 24) {real, imag} */,
  {32'hbd5469b2, 32'hbbe49f48} /* (12, 1, 23) {real, imag} */,
  {32'hbd75e322, 32'h3da79224} /* (12, 1, 22) {real, imag} */,
  {32'h3baf02a8, 32'h3dbfee74} /* (12, 1, 21) {real, imag} */,
  {32'hbc56c224, 32'hbaf747b0} /* (12, 1, 20) {real, imag} */,
  {32'hbd9c3c93, 32'h3d8c57bb} /* (12, 1, 19) {real, imag} */,
  {32'h3d4923a0, 32'hbda0767f} /* (12, 1, 18) {real, imag} */,
  {32'hbd028754, 32'h3ca865fa} /* (12, 1, 17) {real, imag} */,
  {32'hbc8133cf, 32'h00000000} /* (12, 1, 16) {real, imag} */,
  {32'hbd028754, 32'hbca865fa} /* (12, 1, 15) {real, imag} */,
  {32'h3d4923a0, 32'h3da0767f} /* (12, 1, 14) {real, imag} */,
  {32'hbd9c3c93, 32'hbd8c57bb} /* (12, 1, 13) {real, imag} */,
  {32'hbc56c224, 32'h3af747b0} /* (12, 1, 12) {real, imag} */,
  {32'h3baf02a8, 32'hbdbfee74} /* (12, 1, 11) {real, imag} */,
  {32'hbd75e322, 32'hbda79224} /* (12, 1, 10) {real, imag} */,
  {32'hbd5469b2, 32'h3be49f48} /* (12, 1, 9) {real, imag} */,
  {32'h3df7f591, 32'h3c08c313} /* (12, 1, 8) {real, imag} */,
  {32'hbbb1f5c8, 32'hbaab81e8} /* (12, 1, 7) {real, imag} */,
  {32'h3d37e3ba, 32'h3cd1d58e} /* (12, 1, 6) {real, imag} */,
  {32'hbe0f828a, 32'h3e7f90f6} /* (12, 1, 5) {real, imag} */,
  {32'hbd476dc5, 32'hbec6b49a} /* (12, 1, 4) {real, imag} */,
  {32'hbc3b2f38, 32'hbd18c204} /* (12, 1, 3) {real, imag} */,
  {32'h3de6732c, 32'hbf75a3bc} /* (12, 1, 2) {real, imag} */,
  {32'h403d4878, 32'h4057b7e6} /* (12, 1, 1) {real, imag} */,
  {32'h409d5512, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'h4044c76b, 32'hc02e1f7a} /* (12, 0, 31) {real, imag} */,
  {32'hbea5ab4a, 32'h3f4609da} /* (12, 0, 30) {real, imag} */,
  {32'hbd03fe81, 32'h3ca4037a} /* (12, 0, 29) {real, imag} */,
  {32'hbd9fe4ec, 32'h3e1d9537} /* (12, 0, 28) {real, imag} */,
  {32'hbe09acfd, 32'hbe04e283} /* (12, 0, 27) {real, imag} */,
  {32'hbc58c004, 32'h3c281081} /* (12, 0, 26) {real, imag} */,
  {32'h3c916512, 32'hbda1d93e} /* (12, 0, 25) {real, imag} */,
  {32'h3d8fa6ad, 32'hbcae1f61} /* (12, 0, 24) {real, imag} */,
  {32'hbd6d54e8, 32'h3c2d4df6} /* (12, 0, 23) {real, imag} */,
  {32'h3d36a2e5, 32'h3ccf0dda} /* (12, 0, 22) {real, imag} */,
  {32'h3cbcdddd, 32'h3bc86938} /* (12, 0, 21) {real, imag} */,
  {32'h3cf72efe, 32'hbcde3644} /* (12, 0, 20) {real, imag} */,
  {32'hbc29f64a, 32'h3d874d10} /* (12, 0, 19) {real, imag} */,
  {32'h3ca75f9e, 32'h3d0ba462} /* (12, 0, 18) {real, imag} */,
  {32'h3d2c2264, 32'h3cbc1e9f} /* (12, 0, 17) {real, imag} */,
  {32'hbd43449d, 32'h00000000} /* (12, 0, 16) {real, imag} */,
  {32'h3d2c2264, 32'hbcbc1e9f} /* (12, 0, 15) {real, imag} */,
  {32'h3ca75f9e, 32'hbd0ba462} /* (12, 0, 14) {real, imag} */,
  {32'hbc29f64a, 32'hbd874d10} /* (12, 0, 13) {real, imag} */,
  {32'h3cf72efe, 32'h3cde3644} /* (12, 0, 12) {real, imag} */,
  {32'h3cbcdddd, 32'hbbc86938} /* (12, 0, 11) {real, imag} */,
  {32'h3d36a2e5, 32'hbccf0dda} /* (12, 0, 10) {real, imag} */,
  {32'hbd6d54e8, 32'hbc2d4df6} /* (12, 0, 9) {real, imag} */,
  {32'h3d8fa6ad, 32'h3cae1f61} /* (12, 0, 8) {real, imag} */,
  {32'h3c916512, 32'h3da1d93e} /* (12, 0, 7) {real, imag} */,
  {32'hbc58c004, 32'hbc281081} /* (12, 0, 6) {real, imag} */,
  {32'hbe09acfd, 32'h3e04e283} /* (12, 0, 5) {real, imag} */,
  {32'hbd9fe4ec, 32'hbe1d9537} /* (12, 0, 4) {real, imag} */,
  {32'hbd03fe81, 32'hbca4037a} /* (12, 0, 3) {real, imag} */,
  {32'hbea5ab4a, 32'hbf4609da} /* (12, 0, 2) {real, imag} */,
  {32'h4044c76b, 32'h402e1f7a} /* (12, 0, 1) {real, imag} */,
  {32'h40984ff7, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h4080b08d, 32'hc01085c2} /* (11, 31, 31) {real, imag} */,
  {32'hbf56c99d, 32'h3f379a39} /* (11, 31, 30) {real, imag} */,
  {32'hbd304cb4, 32'h3d1dedc0} /* (11, 31, 29) {real, imag} */,
  {32'h3d957d51, 32'h3da3c13a} /* (11, 31, 28) {real, imag} */,
  {32'hbe0bf696, 32'h3ce7b6b0} /* (11, 31, 27) {real, imag} */,
  {32'hbc9aee78, 32'hbcdabf22} /* (11, 31, 26) {real, imag} */,
  {32'h3dccc25e, 32'hbd5f191c} /* (11, 31, 25) {real, imag} */,
  {32'hbdd4801f, 32'h3d67c1e0} /* (11, 31, 24) {real, imag} */,
  {32'h3ae4da80, 32'hbd07e114} /* (11, 31, 23) {real, imag} */,
  {32'h3d054503, 32'h3c3e8d5c} /* (11, 31, 22) {real, imag} */,
  {32'h3d2054be, 32'h3c999196} /* (11, 31, 21) {real, imag} */,
  {32'h3cded65b, 32'hbd4c16ea} /* (11, 31, 20) {real, imag} */,
  {32'h3dd2a29c, 32'hbd887d0f} /* (11, 31, 19) {real, imag} */,
  {32'h3d232323, 32'h3d5aea96} /* (11, 31, 18) {real, imag} */,
  {32'h3cb9c876, 32'hbdb0934e} /* (11, 31, 17) {real, imag} */,
  {32'h3e09728f, 32'h00000000} /* (11, 31, 16) {real, imag} */,
  {32'h3cb9c876, 32'h3db0934e} /* (11, 31, 15) {real, imag} */,
  {32'h3d232323, 32'hbd5aea96} /* (11, 31, 14) {real, imag} */,
  {32'h3dd2a29c, 32'h3d887d0f} /* (11, 31, 13) {real, imag} */,
  {32'h3cded65b, 32'h3d4c16ea} /* (11, 31, 12) {real, imag} */,
  {32'h3d2054be, 32'hbc999196} /* (11, 31, 11) {real, imag} */,
  {32'h3d054503, 32'hbc3e8d5c} /* (11, 31, 10) {real, imag} */,
  {32'h3ae4da80, 32'h3d07e114} /* (11, 31, 9) {real, imag} */,
  {32'hbdd4801f, 32'hbd67c1e0} /* (11, 31, 8) {real, imag} */,
  {32'h3dccc25e, 32'h3d5f191c} /* (11, 31, 7) {real, imag} */,
  {32'hbc9aee78, 32'h3cdabf22} /* (11, 31, 6) {real, imag} */,
  {32'hbe0bf696, 32'hbce7b6b0} /* (11, 31, 5) {real, imag} */,
  {32'h3d957d51, 32'hbda3c13a} /* (11, 31, 4) {real, imag} */,
  {32'hbd304cb4, 32'hbd1dedc0} /* (11, 31, 3) {real, imag} */,
  {32'hbf56c99d, 32'hbf379a39} /* (11, 31, 2) {real, imag} */,
  {32'h4080b08d, 32'h401085c2} /* (11, 31, 1) {real, imag} */,
  {32'h40a9f1cd, 32'h00000000} /* (11, 31, 0) {real, imag} */,
  {32'h408feef9, 32'hbfd98c4c} /* (11, 30, 31) {real, imag} */,
  {32'hbfad3eae, 32'h3f310ca8} /* (11, 30, 30) {real, imag} */,
  {32'hbcf26293, 32'h3dad15b2} /* (11, 30, 29) {real, imag} */,
  {32'h3d97e14b, 32'h3da9ce3a} /* (11, 30, 28) {real, imag} */,
  {32'hbe1f48e0, 32'hbdab3c99} /* (11, 30, 27) {real, imag} */,
  {32'h3cb0d48c, 32'hbe1b1c58} /* (11, 30, 26) {real, imag} */,
  {32'h3d608967, 32'h3d4c865b} /* (11, 30, 25) {real, imag} */,
  {32'hbca9e22c, 32'hbaeca420} /* (11, 30, 24) {real, imag} */,
  {32'hbd21224d, 32'hbdb9a630} /* (11, 30, 23) {real, imag} */,
  {32'h3d13b73d, 32'hbca4a33c} /* (11, 30, 22) {real, imag} */,
  {32'hbdb819de, 32'h3d82f6e6} /* (11, 30, 21) {real, imag} */,
  {32'hbcd5efe8, 32'hbe035f9e} /* (11, 30, 20) {real, imag} */,
  {32'hbc7847d0, 32'hbd1a932f} /* (11, 30, 19) {real, imag} */,
  {32'h3c8a477a, 32'hbba6c69a} /* (11, 30, 18) {real, imag} */,
  {32'h3c9144ad, 32'hbc826e21} /* (11, 30, 17) {real, imag} */,
  {32'h3d5edeb6, 32'h00000000} /* (11, 30, 16) {real, imag} */,
  {32'h3c9144ad, 32'h3c826e21} /* (11, 30, 15) {real, imag} */,
  {32'h3c8a477a, 32'h3ba6c69a} /* (11, 30, 14) {real, imag} */,
  {32'hbc7847d0, 32'h3d1a932f} /* (11, 30, 13) {real, imag} */,
  {32'hbcd5efe8, 32'h3e035f9e} /* (11, 30, 12) {real, imag} */,
  {32'hbdb819de, 32'hbd82f6e6} /* (11, 30, 11) {real, imag} */,
  {32'h3d13b73d, 32'h3ca4a33c} /* (11, 30, 10) {real, imag} */,
  {32'hbd21224d, 32'h3db9a630} /* (11, 30, 9) {real, imag} */,
  {32'hbca9e22c, 32'h3aeca420} /* (11, 30, 8) {real, imag} */,
  {32'h3d608967, 32'hbd4c865b} /* (11, 30, 7) {real, imag} */,
  {32'h3cb0d48c, 32'h3e1b1c58} /* (11, 30, 6) {real, imag} */,
  {32'hbe1f48e0, 32'h3dab3c99} /* (11, 30, 5) {real, imag} */,
  {32'h3d97e14b, 32'hbda9ce3a} /* (11, 30, 4) {real, imag} */,
  {32'hbcf26293, 32'hbdad15b2} /* (11, 30, 3) {real, imag} */,
  {32'hbfad3eae, 32'hbf310ca8} /* (11, 30, 2) {real, imag} */,
  {32'h408feef9, 32'h3fd98c4c} /* (11, 30, 1) {real, imag} */,
  {32'h40b00b9b, 32'h00000000} /* (11, 30, 0) {real, imag} */,
  {32'h409892e6, 32'hbfb245c2} /* (11, 29, 31) {real, imag} */,
  {32'hbfb8fc2c, 32'h3f08e4b9} /* (11, 29, 30) {real, imag} */,
  {32'h3d33475d, 32'h3aab3c50} /* (11, 29, 29) {real, imag} */,
  {32'h3e373972, 32'hbd9b6327} /* (11, 29, 28) {real, imag} */,
  {32'hbe784552, 32'hbce64ce9} /* (11, 29, 27) {real, imag} */,
  {32'h3c8a0b14, 32'hbd4bacec} /* (11, 29, 26) {real, imag} */,
  {32'hbc58b272, 32'h3d7a85f4} /* (11, 29, 25) {real, imag} */,
  {32'hbcffffce, 32'h3cdd7e6c} /* (11, 29, 24) {real, imag} */,
  {32'hbcd7de8c, 32'hbc7b9dc4} /* (11, 29, 23) {real, imag} */,
  {32'h3d465da2, 32'h3cedbe04} /* (11, 29, 22) {real, imag} */,
  {32'hbd06a812, 32'hbc95ad96} /* (11, 29, 21) {real, imag} */,
  {32'hbc25b563, 32'h3caa4e6a} /* (11, 29, 20) {real, imag} */,
  {32'hbd7d4eae, 32'h3d31b2c2} /* (11, 29, 19) {real, imag} */,
  {32'hbd20c1c1, 32'h3ade2240} /* (11, 29, 18) {real, imag} */,
  {32'h3c892ce4, 32'h3c10533c} /* (11, 29, 17) {real, imag} */,
  {32'h3d179d6e, 32'h00000000} /* (11, 29, 16) {real, imag} */,
  {32'h3c892ce4, 32'hbc10533c} /* (11, 29, 15) {real, imag} */,
  {32'hbd20c1c1, 32'hbade2240} /* (11, 29, 14) {real, imag} */,
  {32'hbd7d4eae, 32'hbd31b2c2} /* (11, 29, 13) {real, imag} */,
  {32'hbc25b563, 32'hbcaa4e6a} /* (11, 29, 12) {real, imag} */,
  {32'hbd06a812, 32'h3c95ad96} /* (11, 29, 11) {real, imag} */,
  {32'h3d465da2, 32'hbcedbe04} /* (11, 29, 10) {real, imag} */,
  {32'hbcd7de8c, 32'h3c7b9dc4} /* (11, 29, 9) {real, imag} */,
  {32'hbcffffce, 32'hbcdd7e6c} /* (11, 29, 8) {real, imag} */,
  {32'hbc58b272, 32'hbd7a85f4} /* (11, 29, 7) {real, imag} */,
  {32'h3c8a0b14, 32'h3d4bacec} /* (11, 29, 6) {real, imag} */,
  {32'hbe784552, 32'h3ce64ce9} /* (11, 29, 5) {real, imag} */,
  {32'h3e373972, 32'h3d9b6327} /* (11, 29, 4) {real, imag} */,
  {32'h3d33475d, 32'hbaab3c50} /* (11, 29, 3) {real, imag} */,
  {32'hbfb8fc2c, 32'hbf08e4b9} /* (11, 29, 2) {real, imag} */,
  {32'h409892e6, 32'h3fb245c2} /* (11, 29, 1) {real, imag} */,
  {32'h40b01a21, 32'h00000000} /* (11, 29, 0) {real, imag} */,
  {32'h40a4369e, 32'hbf985aed} /* (11, 28, 31) {real, imag} */,
  {32'hbfd36833, 32'h3ec6d004} /* (11, 28, 30) {real, imag} */,
  {32'h3d7e63ee, 32'h3df51838} /* (11, 28, 29) {real, imag} */,
  {32'h3dafe1a6, 32'hbdea9b94} /* (11, 28, 28) {real, imag} */,
  {32'hbe492f4c, 32'h3d9541fa} /* (11, 28, 27) {real, imag} */,
  {32'h3bd17a5e, 32'h3d55db24} /* (11, 28, 26) {real, imag} */,
  {32'h3ca57227, 32'hbd99eb31} /* (11, 28, 25) {real, imag} */,
  {32'hbe1012c3, 32'h3d362322} /* (11, 28, 24) {real, imag} */,
  {32'hbcf6e1dc, 32'h3ddf66c4} /* (11, 28, 23) {real, imag} */,
  {32'hbcc97f6e, 32'hbca26a82} /* (11, 28, 22) {real, imag} */,
  {32'hbc0ece18, 32'hbc87efbd} /* (11, 28, 21) {real, imag} */,
  {32'h3d96a614, 32'h3d55c302} /* (11, 28, 20) {real, imag} */,
  {32'hbd9b1e8e, 32'hbc1cdf34} /* (11, 28, 19) {real, imag} */,
  {32'h3cf0732e, 32'hbbe7a68c} /* (11, 28, 18) {real, imag} */,
  {32'h3cab9ca8, 32'hbda7b7f0} /* (11, 28, 17) {real, imag} */,
  {32'hbd18f0ca, 32'h00000000} /* (11, 28, 16) {real, imag} */,
  {32'h3cab9ca8, 32'h3da7b7f0} /* (11, 28, 15) {real, imag} */,
  {32'h3cf0732e, 32'h3be7a68c} /* (11, 28, 14) {real, imag} */,
  {32'hbd9b1e8e, 32'h3c1cdf34} /* (11, 28, 13) {real, imag} */,
  {32'h3d96a614, 32'hbd55c302} /* (11, 28, 12) {real, imag} */,
  {32'hbc0ece18, 32'h3c87efbd} /* (11, 28, 11) {real, imag} */,
  {32'hbcc97f6e, 32'h3ca26a82} /* (11, 28, 10) {real, imag} */,
  {32'hbcf6e1dc, 32'hbddf66c4} /* (11, 28, 9) {real, imag} */,
  {32'hbe1012c3, 32'hbd362322} /* (11, 28, 8) {real, imag} */,
  {32'h3ca57227, 32'h3d99eb31} /* (11, 28, 7) {real, imag} */,
  {32'h3bd17a5e, 32'hbd55db24} /* (11, 28, 6) {real, imag} */,
  {32'hbe492f4c, 32'hbd9541fa} /* (11, 28, 5) {real, imag} */,
  {32'h3dafe1a6, 32'h3dea9b94} /* (11, 28, 4) {real, imag} */,
  {32'h3d7e63ee, 32'hbdf51838} /* (11, 28, 3) {real, imag} */,
  {32'hbfd36833, 32'hbec6d004} /* (11, 28, 2) {real, imag} */,
  {32'h40a4369e, 32'h3f985aed} /* (11, 28, 1) {real, imag} */,
  {32'h40acf012, 32'h00000000} /* (11, 28, 0) {real, imag} */,
  {32'h40a8072f, 32'hbf80ab34} /* (11, 27, 31) {real, imag} */,
  {32'hbfe9f8aa, 32'h3e94683e} /* (11, 27, 30) {real, imag} */,
  {32'hbcd11656, 32'h3def62ea} /* (11, 27, 29) {real, imag} */,
  {32'h3e1ed6a8, 32'hbe808ee0} /* (11, 27, 28) {real, imag} */,
  {32'hbe17835e, 32'h3c9788bc} /* (11, 27, 27) {real, imag} */,
  {32'hbd31ec7b, 32'h3d928ee0} /* (11, 27, 26) {real, imag} */,
  {32'hbc008b68, 32'hbe06941a} /* (11, 27, 25) {real, imag} */,
  {32'hbd75da3e, 32'h3d4d9bc7} /* (11, 27, 24) {real, imag} */,
  {32'h3b8092d8, 32'h3dc3ed70} /* (11, 27, 23) {real, imag} */,
  {32'h3e2d46a5, 32'h3d837b2b} /* (11, 27, 22) {real, imag} */,
  {32'h3d13e9ce, 32'hbba09510} /* (11, 27, 21) {real, imag} */,
  {32'hbe17fe92, 32'hbd7e9b8e} /* (11, 27, 20) {real, imag} */,
  {32'hbd71a93a, 32'h3cba16a8} /* (11, 27, 19) {real, imag} */,
  {32'hbd67eaa2, 32'hbd38b1cf} /* (11, 27, 18) {real, imag} */,
  {32'h3d3c8b57, 32'hbd83584b} /* (11, 27, 17) {real, imag} */,
  {32'h3c28104c, 32'h00000000} /* (11, 27, 16) {real, imag} */,
  {32'h3d3c8b57, 32'h3d83584b} /* (11, 27, 15) {real, imag} */,
  {32'hbd67eaa2, 32'h3d38b1cf} /* (11, 27, 14) {real, imag} */,
  {32'hbd71a93a, 32'hbcba16a8} /* (11, 27, 13) {real, imag} */,
  {32'hbe17fe92, 32'h3d7e9b8e} /* (11, 27, 12) {real, imag} */,
  {32'h3d13e9ce, 32'h3ba09510} /* (11, 27, 11) {real, imag} */,
  {32'h3e2d46a5, 32'hbd837b2b} /* (11, 27, 10) {real, imag} */,
  {32'h3b8092d8, 32'hbdc3ed70} /* (11, 27, 9) {real, imag} */,
  {32'hbd75da3e, 32'hbd4d9bc7} /* (11, 27, 8) {real, imag} */,
  {32'hbc008b68, 32'h3e06941a} /* (11, 27, 7) {real, imag} */,
  {32'hbd31ec7b, 32'hbd928ee0} /* (11, 27, 6) {real, imag} */,
  {32'hbe17835e, 32'hbc9788bc} /* (11, 27, 5) {real, imag} */,
  {32'h3e1ed6a8, 32'h3e808ee0} /* (11, 27, 4) {real, imag} */,
  {32'hbcd11656, 32'hbdef62ea} /* (11, 27, 3) {real, imag} */,
  {32'hbfe9f8aa, 32'hbe94683e} /* (11, 27, 2) {real, imag} */,
  {32'h40a8072f, 32'h3f80ab34} /* (11, 27, 1) {real, imag} */,
  {32'h40a9eb1e, 32'h00000000} /* (11, 27, 0) {real, imag} */,
  {32'h40a3bb95, 32'hbf59615c} /* (11, 26, 31) {real, imag} */,
  {32'hbfe4ee89, 32'h3e594b68} /* (11, 26, 30) {real, imag} */,
  {32'h3d1918da, 32'hbd39dc5a} /* (11, 26, 29) {real, imag} */,
  {32'h3e12cb89, 32'hbdba22ac} /* (11, 26, 28) {real, imag} */,
  {32'hbe0b3f12, 32'h3bf53e80} /* (11, 26, 27) {real, imag} */,
  {32'hbdcbde0e, 32'h3d84d911} /* (11, 26, 26) {real, imag} */,
  {32'h3ce96ad0, 32'hbd5f22ef} /* (11, 26, 25) {real, imag} */,
  {32'h3c8bc2cf, 32'h3d890ba5} /* (11, 26, 24) {real, imag} */,
  {32'hbae21570, 32'h3d327a35} /* (11, 26, 23) {real, imag} */,
  {32'h3c0da4d4, 32'h3d747bfe} /* (11, 26, 22) {real, imag} */,
  {32'h3cc35e6c, 32'h3d858859} /* (11, 26, 21) {real, imag} */,
  {32'h3d0a7c1a, 32'h3c457661} /* (11, 26, 20) {real, imag} */,
  {32'h3d99b736, 32'h3c9fdce0} /* (11, 26, 19) {real, imag} */,
  {32'h3d2d628e, 32'h3bfe51f8} /* (11, 26, 18) {real, imag} */,
  {32'hbac6fe00, 32'h3b686520} /* (11, 26, 17) {real, imag} */,
  {32'h3c054b01, 32'h00000000} /* (11, 26, 16) {real, imag} */,
  {32'hbac6fe00, 32'hbb686520} /* (11, 26, 15) {real, imag} */,
  {32'h3d2d628e, 32'hbbfe51f8} /* (11, 26, 14) {real, imag} */,
  {32'h3d99b736, 32'hbc9fdce0} /* (11, 26, 13) {real, imag} */,
  {32'h3d0a7c1a, 32'hbc457661} /* (11, 26, 12) {real, imag} */,
  {32'h3cc35e6c, 32'hbd858859} /* (11, 26, 11) {real, imag} */,
  {32'h3c0da4d4, 32'hbd747bfe} /* (11, 26, 10) {real, imag} */,
  {32'hbae21570, 32'hbd327a35} /* (11, 26, 9) {real, imag} */,
  {32'h3c8bc2cf, 32'hbd890ba5} /* (11, 26, 8) {real, imag} */,
  {32'h3ce96ad0, 32'h3d5f22ef} /* (11, 26, 7) {real, imag} */,
  {32'hbdcbde0e, 32'hbd84d911} /* (11, 26, 6) {real, imag} */,
  {32'hbe0b3f12, 32'hbbf53e80} /* (11, 26, 5) {real, imag} */,
  {32'h3e12cb89, 32'h3dba22ac} /* (11, 26, 4) {real, imag} */,
  {32'h3d1918da, 32'h3d39dc5a} /* (11, 26, 3) {real, imag} */,
  {32'hbfe4ee89, 32'hbe594b68} /* (11, 26, 2) {real, imag} */,
  {32'h40a3bb95, 32'h3f59615c} /* (11, 26, 1) {real, imag} */,
  {32'h40a0d45a, 32'h00000000} /* (11, 26, 0) {real, imag} */,
  {32'h40992ebd, 32'hbf0c8d9f} /* (11, 25, 31) {real, imag} */,
  {32'hbfe9af5e, 32'h3e6ffb28} /* (11, 25, 30) {real, imag} */,
  {32'hbdafa8e6, 32'h3d89dbce} /* (11, 25, 29) {real, imag} */,
  {32'h3da6f63a, 32'hbe025fba} /* (11, 25, 28) {real, imag} */,
  {32'hbdf00b29, 32'h3e615f36} /* (11, 25, 27) {real, imag} */,
  {32'hbe6c8b17, 32'hbe207fbc} /* (11, 25, 26) {real, imag} */,
  {32'h3dc97c9d, 32'h3d50e0db} /* (11, 25, 25) {real, imag} */,
  {32'hbc933eaa, 32'h3d84038f} /* (11, 25, 24) {real, imag} */,
  {32'h3dd64bca, 32'h3d6b00aa} /* (11, 25, 23) {real, imag} */,
  {32'hbcd959ea, 32'hbd72fff0} /* (11, 25, 22) {real, imag} */,
  {32'hbdaf23d8, 32'hbcdbbca0} /* (11, 25, 21) {real, imag} */,
  {32'hbcc2a7ee, 32'h3c382c03} /* (11, 25, 20) {real, imag} */,
  {32'h3d658973, 32'h3cd21afb} /* (11, 25, 19) {real, imag} */,
  {32'h3d072c40, 32'hbd7978e3} /* (11, 25, 18) {real, imag} */,
  {32'h3cf9c750, 32'h3cec00a7} /* (11, 25, 17) {real, imag} */,
  {32'hbd4897d8, 32'h00000000} /* (11, 25, 16) {real, imag} */,
  {32'h3cf9c750, 32'hbcec00a7} /* (11, 25, 15) {real, imag} */,
  {32'h3d072c40, 32'h3d7978e3} /* (11, 25, 14) {real, imag} */,
  {32'h3d658973, 32'hbcd21afb} /* (11, 25, 13) {real, imag} */,
  {32'hbcc2a7ee, 32'hbc382c03} /* (11, 25, 12) {real, imag} */,
  {32'hbdaf23d8, 32'h3cdbbca0} /* (11, 25, 11) {real, imag} */,
  {32'hbcd959ea, 32'h3d72fff0} /* (11, 25, 10) {real, imag} */,
  {32'h3dd64bca, 32'hbd6b00aa} /* (11, 25, 9) {real, imag} */,
  {32'hbc933eaa, 32'hbd84038f} /* (11, 25, 8) {real, imag} */,
  {32'h3dc97c9d, 32'hbd50e0db} /* (11, 25, 7) {real, imag} */,
  {32'hbe6c8b17, 32'h3e207fbc} /* (11, 25, 6) {real, imag} */,
  {32'hbdf00b29, 32'hbe615f36} /* (11, 25, 5) {real, imag} */,
  {32'h3da6f63a, 32'h3e025fba} /* (11, 25, 4) {real, imag} */,
  {32'hbdafa8e6, 32'hbd89dbce} /* (11, 25, 3) {real, imag} */,
  {32'hbfe9af5e, 32'hbe6ffb28} /* (11, 25, 2) {real, imag} */,
  {32'h40992ebd, 32'h3f0c8d9f} /* (11, 25, 1) {real, imag} */,
  {32'h40921d2f, 32'h00000000} /* (11, 25, 0) {real, imag} */,
  {32'h40886e20, 32'hbe3b7598} /* (11, 24, 31) {real, imag} */,
  {32'hbfd9014c, 32'h3da605b4} /* (11, 24, 30) {real, imag} */,
  {32'hbe196de2, 32'h3deee5f2} /* (11, 24, 29) {real, imag} */,
  {32'h3e2abec4, 32'hbdec349c} /* (11, 24, 28) {real, imag} */,
  {32'hbe85be13, 32'h3e5733ca} /* (11, 24, 27) {real, imag} */,
  {32'hbddfb9e2, 32'hbdbb6a0a} /* (11, 24, 26) {real, imag} */,
  {32'h3c2b0804, 32'h3d183ff6} /* (11, 24, 25) {real, imag} */,
  {32'hbd8c2594, 32'hbda710c4} /* (11, 24, 24) {real, imag} */,
  {32'h3cb5ee20, 32'hbd60b637} /* (11, 24, 23) {real, imag} */,
  {32'h3c2f4644, 32'hbda5d554} /* (11, 24, 22) {real, imag} */,
  {32'hbdba27a4, 32'h3d6d4d72} /* (11, 24, 21) {real, imag} */,
  {32'h3d93b79e, 32'h3dda0844} /* (11, 24, 20) {real, imag} */,
  {32'hbd737652, 32'hbcb53674} /* (11, 24, 19) {real, imag} */,
  {32'h3db087b6, 32'hbc13bba8} /* (11, 24, 18) {real, imag} */,
  {32'hbd52ee2a, 32'h3ce003d2} /* (11, 24, 17) {real, imag} */,
  {32'hbd2371bc, 32'h00000000} /* (11, 24, 16) {real, imag} */,
  {32'hbd52ee2a, 32'hbce003d2} /* (11, 24, 15) {real, imag} */,
  {32'h3db087b6, 32'h3c13bba8} /* (11, 24, 14) {real, imag} */,
  {32'hbd737652, 32'h3cb53674} /* (11, 24, 13) {real, imag} */,
  {32'h3d93b79e, 32'hbdda0844} /* (11, 24, 12) {real, imag} */,
  {32'hbdba27a4, 32'hbd6d4d72} /* (11, 24, 11) {real, imag} */,
  {32'h3c2f4644, 32'h3da5d554} /* (11, 24, 10) {real, imag} */,
  {32'h3cb5ee20, 32'h3d60b637} /* (11, 24, 9) {real, imag} */,
  {32'hbd8c2594, 32'h3da710c4} /* (11, 24, 8) {real, imag} */,
  {32'h3c2b0804, 32'hbd183ff6} /* (11, 24, 7) {real, imag} */,
  {32'hbddfb9e2, 32'h3dbb6a0a} /* (11, 24, 6) {real, imag} */,
  {32'hbe85be13, 32'hbe5733ca} /* (11, 24, 5) {real, imag} */,
  {32'h3e2abec4, 32'h3dec349c} /* (11, 24, 4) {real, imag} */,
  {32'hbe196de2, 32'hbdeee5f2} /* (11, 24, 3) {real, imag} */,
  {32'hbfd9014c, 32'hbda605b4} /* (11, 24, 2) {real, imag} */,
  {32'h40886e20, 32'h3e3b7598} /* (11, 24, 1) {real, imag} */,
  {32'h407c5762, 32'h00000000} /* (11, 24, 0) {real, imag} */,
  {32'h4060f4ae, 32'hbdfc9778} /* (11, 23, 31) {real, imag} */,
  {32'hbfa1f1e1, 32'h3d6691e4} /* (11, 23, 30) {real, imag} */,
  {32'hbdb58568, 32'h3d8dcccd} /* (11, 23, 29) {real, imag} */,
  {32'h3e4bd4b8, 32'hbe086ec6} /* (11, 23, 28) {real, imag} */,
  {32'hbe58ecee, 32'h3e2c3746} /* (11, 23, 27) {real, imag} */,
  {32'hbc62a1e4, 32'hbd519c4b} /* (11, 23, 26) {real, imag} */,
  {32'h3cf0f60c, 32'hbd5d5cad} /* (11, 23, 25) {real, imag} */,
  {32'hbd0a3671, 32'h3d2e763a} /* (11, 23, 24) {real, imag} */,
  {32'hbc8ee8f2, 32'hbbbda1be} /* (11, 23, 23) {real, imag} */,
  {32'hbb7eb010, 32'hbbe89370} /* (11, 23, 22) {real, imag} */,
  {32'h3d1d70ac, 32'h3df117da} /* (11, 23, 21) {real, imag} */,
  {32'hb9a10500, 32'h3c008c00} /* (11, 23, 20) {real, imag} */,
  {32'hbd842f6a, 32'h3b309a20} /* (11, 23, 19) {real, imag} */,
  {32'h3cb85313, 32'h3ced3d1e} /* (11, 23, 18) {real, imag} */,
  {32'hbc487a93, 32'h3d1254b2} /* (11, 23, 17) {real, imag} */,
  {32'hbd0e7ff8, 32'h00000000} /* (11, 23, 16) {real, imag} */,
  {32'hbc487a93, 32'hbd1254b2} /* (11, 23, 15) {real, imag} */,
  {32'h3cb85313, 32'hbced3d1e} /* (11, 23, 14) {real, imag} */,
  {32'hbd842f6a, 32'hbb309a20} /* (11, 23, 13) {real, imag} */,
  {32'hb9a10500, 32'hbc008c00} /* (11, 23, 12) {real, imag} */,
  {32'h3d1d70ac, 32'hbdf117da} /* (11, 23, 11) {real, imag} */,
  {32'hbb7eb010, 32'h3be89370} /* (11, 23, 10) {real, imag} */,
  {32'hbc8ee8f2, 32'h3bbda1be} /* (11, 23, 9) {real, imag} */,
  {32'hbd0a3671, 32'hbd2e763a} /* (11, 23, 8) {real, imag} */,
  {32'h3cf0f60c, 32'h3d5d5cad} /* (11, 23, 7) {real, imag} */,
  {32'hbc62a1e4, 32'h3d519c4b} /* (11, 23, 6) {real, imag} */,
  {32'hbe58ecee, 32'hbe2c3746} /* (11, 23, 5) {real, imag} */,
  {32'h3e4bd4b8, 32'h3e086ec6} /* (11, 23, 4) {real, imag} */,
  {32'hbdb58568, 32'hbd8dcccd} /* (11, 23, 3) {real, imag} */,
  {32'hbfa1f1e1, 32'hbd6691e4} /* (11, 23, 2) {real, imag} */,
  {32'h4060f4ae, 32'h3dfc9778} /* (11, 23, 1) {real, imag} */,
  {32'h4045cda9, 32'h00000000} /* (11, 23, 0) {real, imag} */,
  {32'h4019e123, 32'hbe359606} /* (11, 22, 31) {real, imag} */,
  {32'hbf52d5e6, 32'h3d3bb2f4} /* (11, 22, 30) {real, imag} */,
  {32'hbb0295b8, 32'h3c54a4ee} /* (11, 22, 29) {real, imag} */,
  {32'h3e98e5f4, 32'hbe2131b9} /* (11, 22, 28) {real, imag} */,
  {32'hbe47fbba, 32'h3e5c6774} /* (11, 22, 27) {real, imag} */,
  {32'hbd67d6ef, 32'h3dbdd8f0} /* (11, 22, 26) {real, imag} */,
  {32'h3dd31df9, 32'hbcff5538} /* (11, 22, 25) {real, imag} */,
  {32'hbdbf5ac4, 32'h3e1f56c7} /* (11, 22, 24) {real, imag} */,
  {32'h3c6c8953, 32'h3cfed07c} /* (11, 22, 23) {real, imag} */,
  {32'hbc920760, 32'h3d39cbe2} /* (11, 22, 22) {real, imag} */,
  {32'h3d961812, 32'h3dacb5a3} /* (11, 22, 21) {real, imag} */,
  {32'hbd5ae8f6, 32'h3c352ae4} /* (11, 22, 20) {real, imag} */,
  {32'h3cb1c95a, 32'h3d503266} /* (11, 22, 19) {real, imag} */,
  {32'hbd2a0da0, 32'h3ccc554b} /* (11, 22, 18) {real, imag} */,
  {32'h3d037e89, 32'hbd2c4c2b} /* (11, 22, 17) {real, imag} */,
  {32'h3cde6b42, 32'h00000000} /* (11, 22, 16) {real, imag} */,
  {32'h3d037e89, 32'h3d2c4c2b} /* (11, 22, 15) {real, imag} */,
  {32'hbd2a0da0, 32'hbccc554b} /* (11, 22, 14) {real, imag} */,
  {32'h3cb1c95a, 32'hbd503266} /* (11, 22, 13) {real, imag} */,
  {32'hbd5ae8f6, 32'hbc352ae4} /* (11, 22, 12) {real, imag} */,
  {32'h3d961812, 32'hbdacb5a3} /* (11, 22, 11) {real, imag} */,
  {32'hbc920760, 32'hbd39cbe2} /* (11, 22, 10) {real, imag} */,
  {32'h3c6c8953, 32'hbcfed07c} /* (11, 22, 9) {real, imag} */,
  {32'hbdbf5ac4, 32'hbe1f56c7} /* (11, 22, 8) {real, imag} */,
  {32'h3dd31df9, 32'h3cff5538} /* (11, 22, 7) {real, imag} */,
  {32'hbd67d6ef, 32'hbdbdd8f0} /* (11, 22, 6) {real, imag} */,
  {32'hbe47fbba, 32'hbe5c6774} /* (11, 22, 5) {real, imag} */,
  {32'h3e98e5f4, 32'h3e2131b9} /* (11, 22, 4) {real, imag} */,
  {32'hbb0295b8, 32'hbc54a4ee} /* (11, 22, 3) {real, imag} */,
  {32'hbf52d5e6, 32'hbd3bb2f4} /* (11, 22, 2) {real, imag} */,
  {32'h4019e123, 32'h3e359606} /* (11, 22, 1) {real, imag} */,
  {32'h40019cb3, 32'h00000000} /* (11, 22, 0) {real, imag} */,
  {32'h3f5b784e, 32'hbd750a60} /* (11, 21, 31) {real, imag} */,
  {32'hbe21b0e4, 32'hbd8d0462} /* (11, 21, 30) {real, imag} */,
  {32'hbdd02d80, 32'h3d4092de} /* (11, 21, 29) {real, imag} */,
  {32'hbcb90fe6, 32'hbcc93eac} /* (11, 21, 28) {real, imag} */,
  {32'hbdf27622, 32'h3d8debb9} /* (11, 21, 27) {real, imag} */,
  {32'h3d2f0588, 32'h3ced9024} /* (11, 21, 26) {real, imag} */,
  {32'hbd3292e0, 32'h3e006249} /* (11, 21, 25) {real, imag} */,
  {32'h3db39ebb, 32'h3d8b8f8e} /* (11, 21, 24) {real, imag} */,
  {32'h3d68daaa, 32'hbcd7d8d6} /* (11, 21, 23) {real, imag} */,
  {32'hbd3c2add, 32'hbdab4bf4} /* (11, 21, 22) {real, imag} */,
  {32'h3a269680, 32'h3d635284} /* (11, 21, 21) {real, imag} */,
  {32'hbd31d8e2, 32'h3d4ffa2b} /* (11, 21, 20) {real, imag} */,
  {32'hbd1ed1fd, 32'hbc5513fb} /* (11, 21, 19) {real, imag} */,
  {32'hbd934198, 32'h3d82a30e} /* (11, 21, 18) {real, imag} */,
  {32'hbbf6d1c6, 32'hbb0e03a8} /* (11, 21, 17) {real, imag} */,
  {32'hbc5f0d54, 32'h00000000} /* (11, 21, 16) {real, imag} */,
  {32'hbbf6d1c6, 32'h3b0e03a8} /* (11, 21, 15) {real, imag} */,
  {32'hbd934198, 32'hbd82a30e} /* (11, 21, 14) {real, imag} */,
  {32'hbd1ed1fd, 32'h3c5513fb} /* (11, 21, 13) {real, imag} */,
  {32'hbd31d8e2, 32'hbd4ffa2b} /* (11, 21, 12) {real, imag} */,
  {32'h3a269680, 32'hbd635284} /* (11, 21, 11) {real, imag} */,
  {32'hbd3c2add, 32'h3dab4bf4} /* (11, 21, 10) {real, imag} */,
  {32'h3d68daaa, 32'h3cd7d8d6} /* (11, 21, 9) {real, imag} */,
  {32'h3db39ebb, 32'hbd8b8f8e} /* (11, 21, 8) {real, imag} */,
  {32'hbd3292e0, 32'hbe006249} /* (11, 21, 7) {real, imag} */,
  {32'h3d2f0588, 32'hbced9024} /* (11, 21, 6) {real, imag} */,
  {32'hbdf27622, 32'hbd8debb9} /* (11, 21, 5) {real, imag} */,
  {32'hbcb90fe6, 32'h3cc93eac} /* (11, 21, 4) {real, imag} */,
  {32'hbdd02d80, 32'hbd4092de} /* (11, 21, 3) {real, imag} */,
  {32'hbe21b0e4, 32'h3d8d0462} /* (11, 21, 2) {real, imag} */,
  {32'h3f5b784e, 32'h3d750a60} /* (11, 21, 1) {real, imag} */,
  {32'h3f515a39, 32'h00000000} /* (11, 21, 0) {real, imag} */,
  {32'hbf97f486, 32'h3df16e30} /* (11, 20, 31) {real, imag} */,
  {32'h3f1ce1a6, 32'hbe806376} /* (11, 20, 30) {real, imag} */,
  {32'hbe3c2661, 32'h3d225d5e} /* (11, 20, 29) {real, imag} */,
  {32'hbd6a418c, 32'h3dce53a8} /* (11, 20, 28) {real, imag} */,
  {32'h3d939b2b, 32'hbc605b9a} /* (11, 20, 27) {real, imag} */,
  {32'h3d819af3, 32'h3cf3ef22} /* (11, 20, 26) {real, imag} */,
  {32'hbc9aace8, 32'hbde6e443} /* (11, 20, 25) {real, imag} */,
  {32'h3ddc91b0, 32'hbe3552dc} /* (11, 20, 24) {real, imag} */,
  {32'h3cbe155b, 32'h3d1cb7df} /* (11, 20, 23) {real, imag} */,
  {32'h3d6a132b, 32'hbd20c164} /* (11, 20, 22) {real, imag} */,
  {32'h3deae760, 32'hbccd4016} /* (11, 20, 21) {real, imag} */,
  {32'hbc181001, 32'hbcf282ad} /* (11, 20, 20) {real, imag} */,
  {32'hbdb653d9, 32'h3b9283a4} /* (11, 20, 19) {real, imag} */,
  {32'h3d436582, 32'hbc2b6ba1} /* (11, 20, 18) {real, imag} */,
  {32'h3bc31c60, 32'h3a353e60} /* (11, 20, 17) {real, imag} */,
  {32'hbc46ff1c, 32'h00000000} /* (11, 20, 16) {real, imag} */,
  {32'h3bc31c60, 32'hba353e60} /* (11, 20, 15) {real, imag} */,
  {32'h3d436582, 32'h3c2b6ba1} /* (11, 20, 14) {real, imag} */,
  {32'hbdb653d9, 32'hbb9283a4} /* (11, 20, 13) {real, imag} */,
  {32'hbc181001, 32'h3cf282ad} /* (11, 20, 12) {real, imag} */,
  {32'h3deae760, 32'h3ccd4016} /* (11, 20, 11) {real, imag} */,
  {32'h3d6a132b, 32'h3d20c164} /* (11, 20, 10) {real, imag} */,
  {32'h3cbe155b, 32'hbd1cb7df} /* (11, 20, 9) {real, imag} */,
  {32'h3ddc91b0, 32'h3e3552dc} /* (11, 20, 8) {real, imag} */,
  {32'hbc9aace8, 32'h3de6e443} /* (11, 20, 7) {real, imag} */,
  {32'h3d819af3, 32'hbcf3ef22} /* (11, 20, 6) {real, imag} */,
  {32'h3d939b2b, 32'h3c605b9a} /* (11, 20, 5) {real, imag} */,
  {32'hbd6a418c, 32'hbdce53a8} /* (11, 20, 4) {real, imag} */,
  {32'hbe3c2661, 32'hbd225d5e} /* (11, 20, 3) {real, imag} */,
  {32'h3f1ce1a6, 32'h3e806376} /* (11, 20, 2) {real, imag} */,
  {32'hbf97f486, 32'hbdf16e30} /* (11, 20, 1) {real, imag} */,
  {32'hbf2306cc, 32'h00000000} /* (11, 20, 0) {real, imag} */,
  {32'hc023dafd, 32'h3e9e8b70} /* (11, 19, 31) {real, imag} */,
  {32'h3f8ae62f, 32'hbe791277} /* (11, 19, 30) {real, imag} */,
  {32'hbdbe5a37, 32'h3d54ec4b} /* (11, 19, 29) {real, imag} */,
  {32'hbc0f39a8, 32'hbcbf4b44} /* (11, 19, 28) {real, imag} */,
  {32'h3e1efa18, 32'h3db78bac} /* (11, 19, 27) {real, imag} */,
  {32'h3ded55c8, 32'h3d06ae5e} /* (11, 19, 26) {real, imag} */,
  {32'hbc87b0e9, 32'h3ce8b5a1} /* (11, 19, 25) {real, imag} */,
  {32'h3dd6c262, 32'hbe2329c0} /* (11, 19, 24) {real, imag} */,
  {32'hbdc216a0, 32'h3c857b8a} /* (11, 19, 23) {real, imag} */,
  {32'hbd5dcc3a, 32'hbcc6c538} /* (11, 19, 22) {real, imag} */,
  {32'h3d19aa6e, 32'hbd9ab084} /* (11, 19, 21) {real, imag} */,
  {32'hbdd52d88, 32'hbd025308} /* (11, 19, 20) {real, imag} */,
  {32'h3d100922, 32'h3de34a3e} /* (11, 19, 19) {real, imag} */,
  {32'hbc73f230, 32'hbd5847d5} /* (11, 19, 18) {real, imag} */,
  {32'h3bbaf51b, 32'hbc0e333c} /* (11, 19, 17) {real, imag} */,
  {32'hbd7f22a4, 32'h00000000} /* (11, 19, 16) {real, imag} */,
  {32'h3bbaf51b, 32'h3c0e333c} /* (11, 19, 15) {real, imag} */,
  {32'hbc73f230, 32'h3d5847d5} /* (11, 19, 14) {real, imag} */,
  {32'h3d100922, 32'hbde34a3e} /* (11, 19, 13) {real, imag} */,
  {32'hbdd52d88, 32'h3d025308} /* (11, 19, 12) {real, imag} */,
  {32'h3d19aa6e, 32'h3d9ab084} /* (11, 19, 11) {real, imag} */,
  {32'hbd5dcc3a, 32'h3cc6c538} /* (11, 19, 10) {real, imag} */,
  {32'hbdc216a0, 32'hbc857b8a} /* (11, 19, 9) {real, imag} */,
  {32'h3dd6c262, 32'h3e2329c0} /* (11, 19, 8) {real, imag} */,
  {32'hbc87b0e9, 32'hbce8b5a1} /* (11, 19, 7) {real, imag} */,
  {32'h3ded55c8, 32'hbd06ae5e} /* (11, 19, 6) {real, imag} */,
  {32'h3e1efa18, 32'hbdb78bac} /* (11, 19, 5) {real, imag} */,
  {32'hbc0f39a8, 32'h3cbf4b44} /* (11, 19, 4) {real, imag} */,
  {32'hbdbe5a37, 32'hbd54ec4b} /* (11, 19, 3) {real, imag} */,
  {32'h3f8ae62f, 32'h3e791277} /* (11, 19, 2) {real, imag} */,
  {32'hc023dafd, 32'hbe9e8b70} /* (11, 19, 1) {real, imag} */,
  {32'hbfe2e5e6, 32'h00000000} /* (11, 19, 0) {real, imag} */,
  {32'hc058d576, 32'h3ed063c0} /* (11, 18, 31) {real, imag} */,
  {32'h3fa8962e, 32'hbe5292f3} /* (11, 18, 30) {real, imag} */,
  {32'h3d8582f5, 32'h3da98f3b} /* (11, 18, 29) {real, imag} */,
  {32'hbdc3e468, 32'h3e18c550} /* (11, 18, 28) {real, imag} */,
  {32'h3e40b5c6, 32'h3bfcd790} /* (11, 18, 27) {real, imag} */,
  {32'hbc9b3285, 32'hbe0407cf} /* (11, 18, 26) {real, imag} */,
  {32'h3d224324, 32'h3c813c08} /* (11, 18, 25) {real, imag} */,
  {32'h3e199f30, 32'hbce41bdc} /* (11, 18, 24) {real, imag} */,
  {32'hbd628eda, 32'h3b69c338} /* (11, 18, 23) {real, imag} */,
  {32'h3cd4c5b2, 32'hbd621f2e} /* (11, 18, 22) {real, imag} */,
  {32'h3d86874e, 32'h3d12f798} /* (11, 18, 21) {real, imag} */,
  {32'h3d957c14, 32'h3cc2d669} /* (11, 18, 20) {real, imag} */,
  {32'h3b8891c8, 32'h3d0f95a3} /* (11, 18, 19) {real, imag} */,
  {32'hbdc0189f, 32'hbcc22a18} /* (11, 18, 18) {real, imag} */,
  {32'h3d843177, 32'hbc9f242d} /* (11, 18, 17) {real, imag} */,
  {32'hbd819754, 32'h00000000} /* (11, 18, 16) {real, imag} */,
  {32'h3d843177, 32'h3c9f242d} /* (11, 18, 15) {real, imag} */,
  {32'hbdc0189f, 32'h3cc22a18} /* (11, 18, 14) {real, imag} */,
  {32'h3b8891c8, 32'hbd0f95a3} /* (11, 18, 13) {real, imag} */,
  {32'h3d957c14, 32'hbcc2d669} /* (11, 18, 12) {real, imag} */,
  {32'h3d86874e, 32'hbd12f798} /* (11, 18, 11) {real, imag} */,
  {32'h3cd4c5b2, 32'h3d621f2e} /* (11, 18, 10) {real, imag} */,
  {32'hbd628eda, 32'hbb69c338} /* (11, 18, 9) {real, imag} */,
  {32'h3e199f30, 32'h3ce41bdc} /* (11, 18, 8) {real, imag} */,
  {32'h3d224324, 32'hbc813c08} /* (11, 18, 7) {real, imag} */,
  {32'hbc9b3285, 32'h3e0407cf} /* (11, 18, 6) {real, imag} */,
  {32'h3e40b5c6, 32'hbbfcd790} /* (11, 18, 5) {real, imag} */,
  {32'hbdc3e468, 32'hbe18c550} /* (11, 18, 4) {real, imag} */,
  {32'h3d8582f5, 32'hbda98f3b} /* (11, 18, 3) {real, imag} */,
  {32'h3fa8962e, 32'h3e5292f3} /* (11, 18, 2) {real, imag} */,
  {32'hc058d576, 32'hbed063c0} /* (11, 18, 1) {real, imag} */,
  {32'hc02e3a92, 32'h00000000} /* (11, 18, 0) {real, imag} */,
  {32'hc08204aa, 32'h3eae0266} /* (11, 17, 31) {real, imag} */,
  {32'h3fc712cf, 32'hbedfce92} /* (11, 17, 30) {real, imag} */,
  {32'h3de0e99f, 32'hbe0d9df8} /* (11, 17, 29) {real, imag} */,
  {32'hbd6177b8, 32'h3dbe2b0d} /* (11, 17, 28) {real, imag} */,
  {32'h3eb05931, 32'hbda88e10} /* (11, 17, 27) {real, imag} */,
  {32'hbd910758, 32'hbdb3dc54} /* (11, 17, 26) {real, imag} */,
  {32'h3dc7d0b4, 32'h3ac0f700} /* (11, 17, 25) {real, imag} */,
  {32'h3d1b2752, 32'h3d7de0e1} /* (11, 17, 24) {real, imag} */,
  {32'h3c8012fc, 32'h3dcbe230} /* (11, 17, 23) {real, imag} */,
  {32'hbdec5230, 32'hbcdc4962} /* (11, 17, 22) {real, imag} */,
  {32'hbd569445, 32'hbc284dbb} /* (11, 17, 21) {real, imag} */,
  {32'h3a389120, 32'hbbc31a4c} /* (11, 17, 20) {real, imag} */,
  {32'h3cf40b75, 32'hbd7c3ef5} /* (11, 17, 19) {real, imag} */,
  {32'h3c94e3e4, 32'hbd02040a} /* (11, 17, 18) {real, imag} */,
  {32'hbd39a7f8, 32'h3d88922d} /* (11, 17, 17) {real, imag} */,
  {32'h3d20c96f, 32'h00000000} /* (11, 17, 16) {real, imag} */,
  {32'hbd39a7f8, 32'hbd88922d} /* (11, 17, 15) {real, imag} */,
  {32'h3c94e3e4, 32'h3d02040a} /* (11, 17, 14) {real, imag} */,
  {32'h3cf40b75, 32'h3d7c3ef5} /* (11, 17, 13) {real, imag} */,
  {32'h3a389120, 32'h3bc31a4c} /* (11, 17, 12) {real, imag} */,
  {32'hbd569445, 32'h3c284dbb} /* (11, 17, 11) {real, imag} */,
  {32'hbdec5230, 32'h3cdc4962} /* (11, 17, 10) {real, imag} */,
  {32'h3c8012fc, 32'hbdcbe230} /* (11, 17, 9) {real, imag} */,
  {32'h3d1b2752, 32'hbd7de0e1} /* (11, 17, 8) {real, imag} */,
  {32'h3dc7d0b4, 32'hbac0f700} /* (11, 17, 7) {real, imag} */,
  {32'hbd910758, 32'h3db3dc54} /* (11, 17, 6) {real, imag} */,
  {32'h3eb05931, 32'h3da88e10} /* (11, 17, 5) {real, imag} */,
  {32'hbd6177b8, 32'hbdbe2b0d} /* (11, 17, 4) {real, imag} */,
  {32'h3de0e99f, 32'h3e0d9df8} /* (11, 17, 3) {real, imag} */,
  {32'h3fc712cf, 32'h3edfce92} /* (11, 17, 2) {real, imag} */,
  {32'hc08204aa, 32'hbeae0266} /* (11, 17, 1) {real, imag} */,
  {32'hc0471511, 32'h00000000} /* (11, 17, 0) {real, imag} */,
  {32'hc08bcc0c, 32'h3eab2150} /* (11, 16, 31) {real, imag} */,
  {32'h3fcdffc1, 32'hbe99da60} /* (11, 16, 30) {real, imag} */,
  {32'h3c9eb15c, 32'h3b7b0360} /* (11, 16, 29) {real, imag} */,
  {32'hbe2bb718, 32'hbd965800} /* (11, 16, 28) {real, imag} */,
  {32'h3ea01792, 32'hbe0f6c24} /* (11, 16, 27) {real, imag} */,
  {32'h3d9df442, 32'h3d24a6e0} /* (11, 16, 26) {real, imag} */,
  {32'hbba61d78, 32'h3d2e0100} /* (11, 16, 25) {real, imag} */,
  {32'h3b9b4eac, 32'h3d1e2b0a} /* (11, 16, 24) {real, imag} */,
  {32'hbccd9e07, 32'h3dc1cc32} /* (11, 16, 23) {real, imag} */,
  {32'h3d9a08bf, 32'h3cae4f03} /* (11, 16, 22) {real, imag} */,
  {32'hbbff64d8, 32'hbd46e4d8} /* (11, 16, 21) {real, imag} */,
  {32'hbc740d08, 32'h3d2723a6} /* (11, 16, 20) {real, imag} */,
  {32'hbd07d0ee, 32'hbd618b5c} /* (11, 16, 19) {real, imag} */,
  {32'hbb9fb48e, 32'hbdf58fc6} /* (11, 16, 18) {real, imag} */,
  {32'hbb2afae8, 32'hbccc7937} /* (11, 16, 17) {real, imag} */,
  {32'h3d159ddd, 32'h00000000} /* (11, 16, 16) {real, imag} */,
  {32'hbb2afae8, 32'h3ccc7937} /* (11, 16, 15) {real, imag} */,
  {32'hbb9fb48e, 32'h3df58fc6} /* (11, 16, 14) {real, imag} */,
  {32'hbd07d0ee, 32'h3d618b5c} /* (11, 16, 13) {real, imag} */,
  {32'hbc740d08, 32'hbd2723a6} /* (11, 16, 12) {real, imag} */,
  {32'hbbff64d8, 32'h3d46e4d8} /* (11, 16, 11) {real, imag} */,
  {32'h3d9a08bf, 32'hbcae4f03} /* (11, 16, 10) {real, imag} */,
  {32'hbccd9e07, 32'hbdc1cc32} /* (11, 16, 9) {real, imag} */,
  {32'h3b9b4eac, 32'hbd1e2b0a} /* (11, 16, 8) {real, imag} */,
  {32'hbba61d78, 32'hbd2e0100} /* (11, 16, 7) {real, imag} */,
  {32'h3d9df442, 32'hbd24a6e0} /* (11, 16, 6) {real, imag} */,
  {32'h3ea01792, 32'h3e0f6c24} /* (11, 16, 5) {real, imag} */,
  {32'hbe2bb718, 32'h3d965800} /* (11, 16, 4) {real, imag} */,
  {32'h3c9eb15c, 32'hbb7b0360} /* (11, 16, 3) {real, imag} */,
  {32'h3fcdffc1, 32'h3e99da60} /* (11, 16, 2) {real, imag} */,
  {32'hc08bcc0c, 32'hbeab2150} /* (11, 16, 1) {real, imag} */,
  {32'hc058eb8f, 32'h00000000} /* (11, 16, 0) {real, imag} */,
  {32'hc08cce12, 32'h3e62aa54} /* (11, 15, 31) {real, imag} */,
  {32'h3fc6299f, 32'hbe2c3f94} /* (11, 15, 30) {real, imag} */,
  {32'h3dc5ac13, 32'h3d92cc54} /* (11, 15, 29) {real, imag} */,
  {32'hbe752226, 32'hbd11542e} /* (11, 15, 28) {real, imag} */,
  {32'h3e17c066, 32'hbd0d39c0} /* (11, 15, 27) {real, imag} */,
  {32'h3e3add4e, 32'hbd2eb4dc} /* (11, 15, 26) {real, imag} */,
  {32'hbda54b72, 32'h3b99c940} /* (11, 15, 25) {real, imag} */,
  {32'h3d70b9a6, 32'hbb3eb9f0} /* (11, 15, 24) {real, imag} */,
  {32'h3d512e5c, 32'hbd513c71} /* (11, 15, 23) {real, imag} */,
  {32'hbdb2b3fa, 32'hbdb91586} /* (11, 15, 22) {real, imag} */,
  {32'hbba13068, 32'hbc09d823} /* (11, 15, 21) {real, imag} */,
  {32'h3d15dd8a, 32'hbd213774} /* (11, 15, 20) {real, imag} */,
  {32'hbd4fae2a, 32'h3d14daa3} /* (11, 15, 19) {real, imag} */,
  {32'hbd283d32, 32'hbce03aa5} /* (11, 15, 18) {real, imag} */,
  {32'h3c4408a2, 32'hbcbfeddf} /* (11, 15, 17) {real, imag} */,
  {32'hbd7aa283, 32'h00000000} /* (11, 15, 16) {real, imag} */,
  {32'h3c4408a2, 32'h3cbfeddf} /* (11, 15, 15) {real, imag} */,
  {32'hbd283d32, 32'h3ce03aa5} /* (11, 15, 14) {real, imag} */,
  {32'hbd4fae2a, 32'hbd14daa3} /* (11, 15, 13) {real, imag} */,
  {32'h3d15dd8a, 32'h3d213774} /* (11, 15, 12) {real, imag} */,
  {32'hbba13068, 32'h3c09d823} /* (11, 15, 11) {real, imag} */,
  {32'hbdb2b3fa, 32'h3db91586} /* (11, 15, 10) {real, imag} */,
  {32'h3d512e5c, 32'h3d513c71} /* (11, 15, 9) {real, imag} */,
  {32'h3d70b9a6, 32'h3b3eb9f0} /* (11, 15, 8) {real, imag} */,
  {32'hbda54b72, 32'hbb99c940} /* (11, 15, 7) {real, imag} */,
  {32'h3e3add4e, 32'h3d2eb4dc} /* (11, 15, 6) {real, imag} */,
  {32'h3e17c066, 32'h3d0d39c0} /* (11, 15, 5) {real, imag} */,
  {32'hbe752226, 32'h3d11542e} /* (11, 15, 4) {real, imag} */,
  {32'h3dc5ac13, 32'hbd92cc54} /* (11, 15, 3) {real, imag} */,
  {32'h3fc6299f, 32'h3e2c3f94} /* (11, 15, 2) {real, imag} */,
  {32'hc08cce12, 32'hbe62aa54} /* (11, 15, 1) {real, imag} */,
  {32'hc059130b, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'hc086113b, 32'h3ebe95d0} /* (11, 14, 31) {real, imag} */,
  {32'h3fb04dfa, 32'hbe953202} /* (11, 14, 30) {real, imag} */,
  {32'hbc19e8d8, 32'h3dd59d15} /* (11, 14, 29) {real, imag} */,
  {32'hbe879ff8, 32'h3e05d612} /* (11, 14, 28) {real, imag} */,
  {32'h3e780562, 32'hbe112d46} /* (11, 14, 27) {real, imag} */,
  {32'h3d0e1a22, 32'hbcb992f0} /* (11, 14, 26) {real, imag} */,
  {32'h3dad7235, 32'h3d3cf52c} /* (11, 14, 25) {real, imag} */,
  {32'h3db4adea, 32'hbdd13757} /* (11, 14, 24) {real, imag} */,
  {32'hbcc39b8c, 32'hbc8a6fd7} /* (11, 14, 23) {real, imag} */,
  {32'hbd722825, 32'hbdf40817} /* (11, 14, 22) {real, imag} */,
  {32'h3aacaae0, 32'hbdbf76ee} /* (11, 14, 21) {real, imag} */,
  {32'hbdeef614, 32'h3cc38f9b} /* (11, 14, 20) {real, imag} */,
  {32'h3dafa92e, 32'hbc400494} /* (11, 14, 19) {real, imag} */,
  {32'hbc9c6054, 32'h3abd82d8} /* (11, 14, 18) {real, imag} */,
  {32'hbdaf5eff, 32'hbb85accc} /* (11, 14, 17) {real, imag} */,
  {32'h3d51758a, 32'h00000000} /* (11, 14, 16) {real, imag} */,
  {32'hbdaf5eff, 32'h3b85accc} /* (11, 14, 15) {real, imag} */,
  {32'hbc9c6054, 32'hbabd82d8} /* (11, 14, 14) {real, imag} */,
  {32'h3dafa92e, 32'h3c400494} /* (11, 14, 13) {real, imag} */,
  {32'hbdeef614, 32'hbcc38f9b} /* (11, 14, 12) {real, imag} */,
  {32'h3aacaae0, 32'h3dbf76ee} /* (11, 14, 11) {real, imag} */,
  {32'hbd722825, 32'h3df40817} /* (11, 14, 10) {real, imag} */,
  {32'hbcc39b8c, 32'h3c8a6fd7} /* (11, 14, 9) {real, imag} */,
  {32'h3db4adea, 32'h3dd13757} /* (11, 14, 8) {real, imag} */,
  {32'h3dad7235, 32'hbd3cf52c} /* (11, 14, 7) {real, imag} */,
  {32'h3d0e1a22, 32'h3cb992f0} /* (11, 14, 6) {real, imag} */,
  {32'h3e780562, 32'h3e112d46} /* (11, 14, 5) {real, imag} */,
  {32'hbe879ff8, 32'hbe05d612} /* (11, 14, 4) {real, imag} */,
  {32'hbc19e8d8, 32'hbdd59d15} /* (11, 14, 3) {real, imag} */,
  {32'h3fb04dfa, 32'h3e953202} /* (11, 14, 2) {real, imag} */,
  {32'hc086113b, 32'hbebe95d0} /* (11, 14, 1) {real, imag} */,
  {32'hc0448036, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'hc0650067, 32'h3e8ebf40} /* (11, 13, 31) {real, imag} */,
  {32'h3fa62355, 32'hbdef1812} /* (11, 13, 30) {real, imag} */,
  {32'hbdcffc1d, 32'h3d432759} /* (11, 13, 29) {real, imag} */,
  {32'hbe3d9ae6, 32'h3e829d53} /* (11, 13, 28) {real, imag} */,
  {32'h3dd7b830, 32'hbd63f1af} /* (11, 13, 27) {real, imag} */,
  {32'hbb9b2cb0, 32'h3d08bab0} /* (11, 13, 26) {real, imag} */,
  {32'h3d34b468, 32'h3cc568fb} /* (11, 13, 25) {real, imag} */,
  {32'h3df58d76, 32'hbdd365eb} /* (11, 13, 24) {real, imag} */,
  {32'h3be52318, 32'h3db76640} /* (11, 13, 23) {real, imag} */,
  {32'h3be02ae4, 32'h3d514d54} /* (11, 13, 22) {real, imag} */,
  {32'h3c4c5058, 32'hbc1a8e2c} /* (11, 13, 21) {real, imag} */,
  {32'h3d2e9f78, 32'hbdcd8f38} /* (11, 13, 20) {real, imag} */,
  {32'h3d48fa28, 32'hbe27c4f5} /* (11, 13, 19) {real, imag} */,
  {32'hbcf43954, 32'hbd5e4397} /* (11, 13, 18) {real, imag} */,
  {32'hbc820dfe, 32'h3d5f04b3} /* (11, 13, 17) {real, imag} */,
  {32'hbdb12b56, 32'h00000000} /* (11, 13, 16) {real, imag} */,
  {32'hbc820dfe, 32'hbd5f04b3} /* (11, 13, 15) {real, imag} */,
  {32'hbcf43954, 32'h3d5e4397} /* (11, 13, 14) {real, imag} */,
  {32'h3d48fa28, 32'h3e27c4f5} /* (11, 13, 13) {real, imag} */,
  {32'h3d2e9f78, 32'h3dcd8f38} /* (11, 13, 12) {real, imag} */,
  {32'h3c4c5058, 32'h3c1a8e2c} /* (11, 13, 11) {real, imag} */,
  {32'h3be02ae4, 32'hbd514d54} /* (11, 13, 10) {real, imag} */,
  {32'h3be52318, 32'hbdb76640} /* (11, 13, 9) {real, imag} */,
  {32'h3df58d76, 32'h3dd365eb} /* (11, 13, 8) {real, imag} */,
  {32'h3d34b468, 32'hbcc568fb} /* (11, 13, 7) {real, imag} */,
  {32'hbb9b2cb0, 32'hbd08bab0} /* (11, 13, 6) {real, imag} */,
  {32'h3dd7b830, 32'h3d63f1af} /* (11, 13, 5) {real, imag} */,
  {32'hbe3d9ae6, 32'hbe829d53} /* (11, 13, 4) {real, imag} */,
  {32'hbdcffc1d, 32'hbd432759} /* (11, 13, 3) {real, imag} */,
  {32'h3fa62355, 32'h3def1812} /* (11, 13, 2) {real, imag} */,
  {32'hc0650067, 32'hbe8ebf40} /* (11, 13, 1) {real, imag} */,
  {32'hc01b06ad, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'hc028de1d, 32'hbd72cbe0} /* (11, 12, 31) {real, imag} */,
  {32'h3f8e2ead, 32'hbe1a29cc} /* (11, 12, 30) {real, imag} */,
  {32'hbe3e367f, 32'hbcd2fc24} /* (11, 12, 29) {real, imag} */,
  {32'hbd7412f4, 32'h3e298bec} /* (11, 12, 28) {real, imag} */,
  {32'h3e1f79fc, 32'hbca0ea65} /* (11, 12, 27) {real, imag} */,
  {32'hbd21888e, 32'hbbc1d890} /* (11, 12, 26) {real, imag} */,
  {32'hbd059e29, 32'hbda1627d} /* (11, 12, 25) {real, imag} */,
  {32'h3ce027be, 32'hbcc37eb4} /* (11, 12, 24) {real, imag} */,
  {32'h3cbb8a55, 32'h3c9b7c8a} /* (11, 12, 23) {real, imag} */,
  {32'h3d023d5f, 32'hbcc813a9} /* (11, 12, 22) {real, imag} */,
  {32'h3d2480c0, 32'hbb05b5cc} /* (11, 12, 21) {real, imag} */,
  {32'h3b1cff4c, 32'h3ca0dab5} /* (11, 12, 20) {real, imag} */,
  {32'h3d54e6fe, 32'hbc565a68} /* (11, 12, 19) {real, imag} */,
  {32'h3d5ff536, 32'hbbdd226e} /* (11, 12, 18) {real, imag} */,
  {32'hbd1efff8, 32'h3d3ec45a} /* (11, 12, 17) {real, imag} */,
  {32'h3d000db9, 32'h00000000} /* (11, 12, 16) {real, imag} */,
  {32'hbd1efff8, 32'hbd3ec45a} /* (11, 12, 15) {real, imag} */,
  {32'h3d5ff536, 32'h3bdd226e} /* (11, 12, 14) {real, imag} */,
  {32'h3d54e6fe, 32'h3c565a68} /* (11, 12, 13) {real, imag} */,
  {32'h3b1cff4c, 32'hbca0dab5} /* (11, 12, 12) {real, imag} */,
  {32'h3d2480c0, 32'h3b05b5cc} /* (11, 12, 11) {real, imag} */,
  {32'h3d023d5f, 32'h3cc813a9} /* (11, 12, 10) {real, imag} */,
  {32'h3cbb8a55, 32'hbc9b7c8a} /* (11, 12, 9) {real, imag} */,
  {32'h3ce027be, 32'h3cc37eb4} /* (11, 12, 8) {real, imag} */,
  {32'hbd059e29, 32'h3da1627d} /* (11, 12, 7) {real, imag} */,
  {32'hbd21888e, 32'h3bc1d890} /* (11, 12, 6) {real, imag} */,
  {32'h3e1f79fc, 32'h3ca0ea65} /* (11, 12, 5) {real, imag} */,
  {32'hbd7412f4, 32'hbe298bec} /* (11, 12, 4) {real, imag} */,
  {32'hbe3e367f, 32'h3cd2fc24} /* (11, 12, 3) {real, imag} */,
  {32'h3f8e2ead, 32'h3e1a29cc} /* (11, 12, 2) {real, imag} */,
  {32'hc028de1d, 32'h3d72cbe0} /* (11, 12, 1) {real, imag} */,
  {32'hbfbd667a, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'hbfbb034f, 32'hbe76b2b8} /* (11, 11, 31) {real, imag} */,
  {32'h3f2dace9, 32'hbdf1bb16} /* (11, 11, 30) {real, imag} */,
  {32'hbdacd6ca, 32'hbd7b9c92} /* (11, 11, 29) {real, imag} */,
  {32'hbdf5c60e, 32'h3d8c6571} /* (11, 11, 28) {real, imag} */,
  {32'h3dc8ecd2, 32'h3d238392} /* (11, 11, 27) {real, imag} */,
  {32'h3e38356c, 32'h3d1c427c} /* (11, 11, 26) {real, imag} */,
  {32'h3b471f78, 32'h3c7c4254} /* (11, 11, 25) {real, imag} */,
  {32'h3d74a7de, 32'h3d8a6a5a} /* (11, 11, 24) {real, imag} */,
  {32'hbe0ff10e, 32'h3d88d07c} /* (11, 11, 23) {real, imag} */,
  {32'h3df43b52, 32'hbd89fc02} /* (11, 11, 22) {real, imag} */,
  {32'hbd32be95, 32'hbd58e664} /* (11, 11, 21) {real, imag} */,
  {32'h3c85da85, 32'hbcd9d3b2} /* (11, 11, 20) {real, imag} */,
  {32'hbcd6bebe, 32'hbca7ac50} /* (11, 11, 19) {real, imag} */,
  {32'h3daba90c, 32'h3d1a7c1a} /* (11, 11, 18) {real, imag} */,
  {32'hbcabadf2, 32'hbca5cc99} /* (11, 11, 17) {real, imag} */,
  {32'h3d88e08a, 32'h00000000} /* (11, 11, 16) {real, imag} */,
  {32'hbcabadf2, 32'h3ca5cc99} /* (11, 11, 15) {real, imag} */,
  {32'h3daba90c, 32'hbd1a7c1a} /* (11, 11, 14) {real, imag} */,
  {32'hbcd6bebe, 32'h3ca7ac50} /* (11, 11, 13) {real, imag} */,
  {32'h3c85da85, 32'h3cd9d3b2} /* (11, 11, 12) {real, imag} */,
  {32'hbd32be95, 32'h3d58e664} /* (11, 11, 11) {real, imag} */,
  {32'h3df43b52, 32'h3d89fc02} /* (11, 11, 10) {real, imag} */,
  {32'hbe0ff10e, 32'hbd88d07c} /* (11, 11, 9) {real, imag} */,
  {32'h3d74a7de, 32'hbd8a6a5a} /* (11, 11, 8) {real, imag} */,
  {32'h3b471f78, 32'hbc7c4254} /* (11, 11, 7) {real, imag} */,
  {32'h3e38356c, 32'hbd1c427c} /* (11, 11, 6) {real, imag} */,
  {32'h3dc8ecd2, 32'hbd238392} /* (11, 11, 5) {real, imag} */,
  {32'hbdf5c60e, 32'hbd8c6571} /* (11, 11, 4) {real, imag} */,
  {32'hbdacd6ca, 32'h3d7b9c92} /* (11, 11, 3) {real, imag} */,
  {32'h3f2dace9, 32'h3df1bb16} /* (11, 11, 2) {real, imag} */,
  {32'hbfbb034f, 32'h3e76b2b8} /* (11, 11, 1) {real, imag} */,
  {32'hbe9dfa72, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'h3ed6abf8, 32'hbf2c8c28} /* (11, 10, 31) {real, imag} */,
  {32'hbe960b07, 32'h3e2e397d} /* (11, 10, 30) {real, imag} */,
  {32'h3c8bf029, 32'hbd802946} /* (11, 10, 29) {real, imag} */,
  {32'hbd1beabc, 32'hbe7e30d7} /* (11, 10, 28) {real, imag} */,
  {32'hbcdd0204, 32'h3e281fb8} /* (11, 10, 27) {real, imag} */,
  {32'h3e1bee4f, 32'hbc5e4ad4} /* (11, 10, 26) {real, imag} */,
  {32'hbc164078, 32'h3ccdbc5c} /* (11, 10, 25) {real, imag} */,
  {32'h3c5b0d94, 32'h3d8a219e} /* (11, 10, 24) {real, imag} */,
  {32'h3d10760a, 32'h3c3ddd5b} /* (11, 10, 23) {real, imag} */,
  {32'hbbec0c10, 32'h3b568700} /* (11, 10, 22) {real, imag} */,
  {32'hbd83cb38, 32'h3dda94f5} /* (11, 10, 21) {real, imag} */,
  {32'hbd5852fa, 32'h3da1f98a} /* (11, 10, 20) {real, imag} */,
  {32'hbd2f2f87, 32'hbc790da8} /* (11, 10, 19) {real, imag} */,
  {32'h3d982a38, 32'hbcca535b} /* (11, 10, 18) {real, imag} */,
  {32'hbc37abb4, 32'h3ca45dfe} /* (11, 10, 17) {real, imag} */,
  {32'hbd829e62, 32'h00000000} /* (11, 10, 16) {real, imag} */,
  {32'hbc37abb4, 32'hbca45dfe} /* (11, 10, 15) {real, imag} */,
  {32'h3d982a38, 32'h3cca535b} /* (11, 10, 14) {real, imag} */,
  {32'hbd2f2f87, 32'h3c790da8} /* (11, 10, 13) {real, imag} */,
  {32'hbd5852fa, 32'hbda1f98a} /* (11, 10, 12) {real, imag} */,
  {32'hbd83cb38, 32'hbdda94f5} /* (11, 10, 11) {real, imag} */,
  {32'hbbec0c10, 32'hbb568700} /* (11, 10, 10) {real, imag} */,
  {32'h3d10760a, 32'hbc3ddd5b} /* (11, 10, 9) {real, imag} */,
  {32'h3c5b0d94, 32'hbd8a219e} /* (11, 10, 8) {real, imag} */,
  {32'hbc164078, 32'hbccdbc5c} /* (11, 10, 7) {real, imag} */,
  {32'h3e1bee4f, 32'h3c5e4ad4} /* (11, 10, 6) {real, imag} */,
  {32'hbcdd0204, 32'hbe281fb8} /* (11, 10, 5) {real, imag} */,
  {32'hbd1beabc, 32'h3e7e30d7} /* (11, 10, 4) {real, imag} */,
  {32'h3c8bf029, 32'h3d802946} /* (11, 10, 3) {real, imag} */,
  {32'hbe960b07, 32'hbe2e397d} /* (11, 10, 2) {real, imag} */,
  {32'h3ed6abf8, 32'h3f2c8c28} /* (11, 10, 1) {real, imag} */,
  {32'h3fb08b26, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h3fe5fbec, 32'hbf856cca} /* (11, 9, 31) {real, imag} */,
  {32'hbf4e1142, 32'h3e9a51d4} /* (11, 9, 30) {real, imag} */,
  {32'hbda89b66, 32'hbe34ee74} /* (11, 9, 29) {real, imag} */,
  {32'h3cc023e4, 32'hbdd756eb} /* (11, 9, 28) {real, imag} */,
  {32'hbdcb68b0, 32'h3e2ee31e} /* (11, 9, 27) {real, imag} */,
  {32'hbd7fedb1, 32'h3daa8596} /* (11, 9, 26) {real, imag} */,
  {32'h3d27a76c, 32'hbcb9c792} /* (11, 9, 25) {real, imag} */,
  {32'hbd4db223, 32'hba3d5ba0} /* (11, 9, 24) {real, imag} */,
  {32'h3dbcbf9e, 32'hbcc90fa4} /* (11, 9, 23) {real, imag} */,
  {32'h3d9e5754, 32'h3da54814} /* (11, 9, 22) {real, imag} */,
  {32'h3d46375a, 32'h3cd90570} /* (11, 9, 21) {real, imag} */,
  {32'hbd779c3c, 32'hbc6ec1be} /* (11, 9, 20) {real, imag} */,
  {32'hb89ce600, 32'hba9f9ea0} /* (11, 9, 19) {real, imag} */,
  {32'h3d3ed226, 32'h3c3243e5} /* (11, 9, 18) {real, imag} */,
  {32'h3b9b86d6, 32'hbd388b2e} /* (11, 9, 17) {real, imag} */,
  {32'hbd0ddcc4, 32'h00000000} /* (11, 9, 16) {real, imag} */,
  {32'h3b9b86d6, 32'h3d388b2e} /* (11, 9, 15) {real, imag} */,
  {32'h3d3ed226, 32'hbc3243e5} /* (11, 9, 14) {real, imag} */,
  {32'hb89ce600, 32'h3a9f9ea0} /* (11, 9, 13) {real, imag} */,
  {32'hbd779c3c, 32'h3c6ec1be} /* (11, 9, 12) {real, imag} */,
  {32'h3d46375a, 32'hbcd90570} /* (11, 9, 11) {real, imag} */,
  {32'h3d9e5754, 32'hbda54814} /* (11, 9, 10) {real, imag} */,
  {32'h3dbcbf9e, 32'h3cc90fa4} /* (11, 9, 9) {real, imag} */,
  {32'hbd4db223, 32'h3a3d5ba0} /* (11, 9, 8) {real, imag} */,
  {32'h3d27a76c, 32'h3cb9c792} /* (11, 9, 7) {real, imag} */,
  {32'hbd7fedb1, 32'hbdaa8596} /* (11, 9, 6) {real, imag} */,
  {32'hbdcb68b0, 32'hbe2ee31e} /* (11, 9, 5) {real, imag} */,
  {32'h3cc023e4, 32'h3dd756eb} /* (11, 9, 4) {real, imag} */,
  {32'hbda89b66, 32'h3e34ee74} /* (11, 9, 3) {real, imag} */,
  {32'hbf4e1142, 32'hbe9a51d4} /* (11, 9, 2) {real, imag} */,
  {32'h3fe5fbec, 32'h3f856cca} /* (11, 9, 1) {real, imag} */,
  {32'h40270ea7, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h40288c0e, 32'hbfb82421} /* (11, 8, 31) {real, imag} */,
  {32'hbf81fbe8, 32'h3ec81375} /* (11, 8, 30) {real, imag} */,
  {32'hbd9348f1, 32'hbaad8b20} /* (11, 8, 29) {real, imag} */,
  {32'hbd2504ee, 32'h3b8ea248} /* (11, 8, 28) {real, imag} */,
  {32'hbcf1a7d0, 32'h3e3289a6} /* (11, 8, 27) {real, imag} */,
  {32'hbc156e08, 32'h3db3c908} /* (11, 8, 26) {real, imag} */,
  {32'h3dddfec6, 32'hbcfda4dc} /* (11, 8, 25) {real, imag} */,
  {32'hbc753754, 32'h3d3f8ab7} /* (11, 8, 24) {real, imag} */,
  {32'hbdbde8cc, 32'h3dbcd9f2} /* (11, 8, 23) {real, imag} */,
  {32'h3ce8a05a, 32'h3db5d450} /* (11, 8, 22) {real, imag} */,
  {32'hbd335a38, 32'hbdaae65b} /* (11, 8, 21) {real, imag} */,
  {32'h3dc52680, 32'h3b126a30} /* (11, 8, 20) {real, imag} */,
  {32'h3cc06ded, 32'h3de1c5a5} /* (11, 8, 19) {real, imag} */,
  {32'hbc727b64, 32'h3d28170c} /* (11, 8, 18) {real, imag} */,
  {32'hbc8100ec, 32'hbcf39bee} /* (11, 8, 17) {real, imag} */,
  {32'h3d80a0dc, 32'h00000000} /* (11, 8, 16) {real, imag} */,
  {32'hbc8100ec, 32'h3cf39bee} /* (11, 8, 15) {real, imag} */,
  {32'hbc727b64, 32'hbd28170c} /* (11, 8, 14) {real, imag} */,
  {32'h3cc06ded, 32'hbde1c5a5} /* (11, 8, 13) {real, imag} */,
  {32'h3dc52680, 32'hbb126a30} /* (11, 8, 12) {real, imag} */,
  {32'hbd335a38, 32'h3daae65b} /* (11, 8, 11) {real, imag} */,
  {32'h3ce8a05a, 32'hbdb5d450} /* (11, 8, 10) {real, imag} */,
  {32'hbdbde8cc, 32'hbdbcd9f2} /* (11, 8, 9) {real, imag} */,
  {32'hbc753754, 32'hbd3f8ab7} /* (11, 8, 8) {real, imag} */,
  {32'h3dddfec6, 32'h3cfda4dc} /* (11, 8, 7) {real, imag} */,
  {32'hbc156e08, 32'hbdb3c908} /* (11, 8, 6) {real, imag} */,
  {32'hbcf1a7d0, 32'hbe3289a6} /* (11, 8, 5) {real, imag} */,
  {32'hbd2504ee, 32'hbb8ea248} /* (11, 8, 4) {real, imag} */,
  {32'hbd9348f1, 32'h3aad8b20} /* (11, 8, 3) {real, imag} */,
  {32'hbf81fbe8, 32'hbec81375} /* (11, 8, 2) {real, imag} */,
  {32'h40288c0e, 32'h3fb82421} /* (11, 8, 1) {real, imag} */,
  {32'h405dfc1c, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h404bb402, 32'hbfe0965c} /* (11, 7, 31) {real, imag} */,
  {32'hbf8f0cc0, 32'h3f442982} /* (11, 7, 30) {real, imag} */,
  {32'hbe089056, 32'h3c886258} /* (11, 7, 29) {real, imag} */,
  {32'hbc81219e, 32'hbd82199f} /* (11, 7, 28) {real, imag} */,
  {32'hbd93228b, 32'h3e38830e} /* (11, 7, 27) {real, imag} */,
  {32'h3ce9c7e8, 32'hbcdd3980} /* (11, 7, 26) {real, imag} */,
  {32'hbda2fb27, 32'hbdda1eda} /* (11, 7, 25) {real, imag} */,
  {32'hbda2a13c, 32'hbc686ff8} /* (11, 7, 24) {real, imag} */,
  {32'hbc093a14, 32'hbdf07473} /* (11, 7, 23) {real, imag} */,
  {32'hbc27e314, 32'hbcf0d704} /* (11, 7, 22) {real, imag} */,
  {32'h3c5b521c, 32'h3c80b948} /* (11, 7, 21) {real, imag} */,
  {32'h3c8f2242, 32'hbcaa66c6} /* (11, 7, 20) {real, imag} */,
  {32'h3d1a30e5, 32'hbda27291} /* (11, 7, 19) {real, imag} */,
  {32'hb9c44f40, 32'hbc9c5e66} /* (11, 7, 18) {real, imag} */,
  {32'h3c6174c3, 32'h3d0ad10c} /* (11, 7, 17) {real, imag} */,
  {32'hbddf2c3c, 32'h00000000} /* (11, 7, 16) {real, imag} */,
  {32'h3c6174c3, 32'hbd0ad10c} /* (11, 7, 15) {real, imag} */,
  {32'hb9c44f40, 32'h3c9c5e66} /* (11, 7, 14) {real, imag} */,
  {32'h3d1a30e5, 32'h3da27291} /* (11, 7, 13) {real, imag} */,
  {32'h3c8f2242, 32'h3caa66c6} /* (11, 7, 12) {real, imag} */,
  {32'h3c5b521c, 32'hbc80b948} /* (11, 7, 11) {real, imag} */,
  {32'hbc27e314, 32'h3cf0d704} /* (11, 7, 10) {real, imag} */,
  {32'hbc093a14, 32'h3df07473} /* (11, 7, 9) {real, imag} */,
  {32'hbda2a13c, 32'h3c686ff8} /* (11, 7, 8) {real, imag} */,
  {32'hbda2fb27, 32'h3dda1eda} /* (11, 7, 7) {real, imag} */,
  {32'h3ce9c7e8, 32'h3cdd3980} /* (11, 7, 6) {real, imag} */,
  {32'hbd93228b, 32'hbe38830e} /* (11, 7, 5) {real, imag} */,
  {32'hbc81219e, 32'h3d82199f} /* (11, 7, 4) {real, imag} */,
  {32'hbe089056, 32'hbc886258} /* (11, 7, 3) {real, imag} */,
  {32'hbf8f0cc0, 32'hbf442982} /* (11, 7, 2) {real, imag} */,
  {32'h404bb402, 32'h3fe0965c} /* (11, 7, 1) {real, imag} */,
  {32'h4087d105, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'h4063f9fe, 32'hc00ded8b} /* (11, 6, 31) {real, imag} */,
  {32'hbf71d296, 32'h3f626d2c} /* (11, 6, 30) {real, imag} */,
  {32'hbe01cf78, 32'hbd7634d6} /* (11, 6, 29) {real, imag} */,
  {32'h3e04d311, 32'hbcd17fca} /* (11, 6, 28) {real, imag} */,
  {32'hbc7bb5f8, 32'h3eac66ac} /* (11, 6, 27) {real, imag} */,
  {32'hbc212dfc, 32'hbd300c18} /* (11, 6, 26) {real, imag} */,
  {32'hbd3286b8, 32'hbd67c09d} /* (11, 6, 25) {real, imag} */,
  {32'h3d61b9ae, 32'hbd1a1fcc} /* (11, 6, 24) {real, imag} */,
  {32'h3d082afc, 32'h3c90fc78} /* (11, 6, 23) {real, imag} */,
  {32'hbc76413c, 32'h3de79725} /* (11, 6, 22) {real, imag} */,
  {32'hbd96f14f, 32'h3d1040b0} /* (11, 6, 21) {real, imag} */,
  {32'h3d0c0a8a, 32'hbb2200f4} /* (11, 6, 20) {real, imag} */,
  {32'hbdb48d0e, 32'hbca2d488} /* (11, 6, 19) {real, imag} */,
  {32'hbdc9a4f1, 32'h3dab30b0} /* (11, 6, 18) {real, imag} */,
  {32'h3e00da10, 32'hbd778d34} /* (11, 6, 17) {real, imag} */,
  {32'hbc2db9c7, 32'h00000000} /* (11, 6, 16) {real, imag} */,
  {32'h3e00da10, 32'h3d778d34} /* (11, 6, 15) {real, imag} */,
  {32'hbdc9a4f1, 32'hbdab30b0} /* (11, 6, 14) {real, imag} */,
  {32'hbdb48d0e, 32'h3ca2d488} /* (11, 6, 13) {real, imag} */,
  {32'h3d0c0a8a, 32'h3b2200f4} /* (11, 6, 12) {real, imag} */,
  {32'hbd96f14f, 32'hbd1040b0} /* (11, 6, 11) {real, imag} */,
  {32'hbc76413c, 32'hbde79725} /* (11, 6, 10) {real, imag} */,
  {32'h3d082afc, 32'hbc90fc78} /* (11, 6, 9) {real, imag} */,
  {32'h3d61b9ae, 32'h3d1a1fcc} /* (11, 6, 8) {real, imag} */,
  {32'hbd3286b8, 32'h3d67c09d} /* (11, 6, 7) {real, imag} */,
  {32'hbc212dfc, 32'h3d300c18} /* (11, 6, 6) {real, imag} */,
  {32'hbc7bb5f8, 32'hbeac66ac} /* (11, 6, 5) {real, imag} */,
  {32'h3e04d311, 32'h3cd17fca} /* (11, 6, 4) {real, imag} */,
  {32'hbe01cf78, 32'h3d7634d6} /* (11, 6, 3) {real, imag} */,
  {32'hbf71d296, 32'hbf626d2c} /* (11, 6, 2) {real, imag} */,
  {32'h4063f9fe, 32'h400ded8b} /* (11, 6, 1) {real, imag} */,
  {32'h40939a96, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'h4058882e, 32'hc044569a} /* (11, 5, 31) {real, imag} */,
  {32'hbebdb656, 32'h3f8370ea} /* (11, 5, 30) {real, imag} */,
  {32'hbd8d4df4, 32'hbb98c720} /* (11, 5, 29) {real, imag} */,
  {32'hbc88a920, 32'h3e931310} /* (11, 5, 28) {real, imag} */,
  {32'hbe000df8, 32'h3e2f33e2} /* (11, 5, 27) {real, imag} */,
  {32'hbdff891e, 32'h3de2a8c0} /* (11, 5, 26) {real, imag} */,
  {32'h3dbbbcff, 32'hbe0ca2c0} /* (11, 5, 25) {real, imag} */,
  {32'hbd196676, 32'hbd322e75} /* (11, 5, 24) {real, imag} */,
  {32'hbddc2b7c, 32'h3e00d962} /* (11, 5, 23) {real, imag} */,
  {32'h3d364b54, 32'h3cb4198c} /* (11, 5, 22) {real, imag} */,
  {32'hbd441eba, 32'h3e01c14e} /* (11, 5, 21) {real, imag} */,
  {32'h3d272bd8, 32'hbd92a601} /* (11, 5, 20) {real, imag} */,
  {32'h3da46517, 32'h3d3da068} /* (11, 5, 19) {real, imag} */,
  {32'hbd941577, 32'hbc0ae22c} /* (11, 5, 18) {real, imag} */,
  {32'hbd48d605, 32'hbcfbb98c} /* (11, 5, 17) {real, imag} */,
  {32'hbd8c5ca6, 32'h00000000} /* (11, 5, 16) {real, imag} */,
  {32'hbd48d605, 32'h3cfbb98c} /* (11, 5, 15) {real, imag} */,
  {32'hbd941577, 32'h3c0ae22c} /* (11, 5, 14) {real, imag} */,
  {32'h3da46517, 32'hbd3da068} /* (11, 5, 13) {real, imag} */,
  {32'h3d272bd8, 32'h3d92a601} /* (11, 5, 12) {real, imag} */,
  {32'hbd441eba, 32'hbe01c14e} /* (11, 5, 11) {real, imag} */,
  {32'h3d364b54, 32'hbcb4198c} /* (11, 5, 10) {real, imag} */,
  {32'hbddc2b7c, 32'hbe00d962} /* (11, 5, 9) {real, imag} */,
  {32'hbd196676, 32'h3d322e75} /* (11, 5, 8) {real, imag} */,
  {32'h3dbbbcff, 32'h3e0ca2c0} /* (11, 5, 7) {real, imag} */,
  {32'hbdff891e, 32'hbde2a8c0} /* (11, 5, 6) {real, imag} */,
  {32'hbe000df8, 32'hbe2f33e2} /* (11, 5, 5) {real, imag} */,
  {32'hbc88a920, 32'hbe931310} /* (11, 5, 4) {real, imag} */,
  {32'hbd8d4df4, 32'h3b98c720} /* (11, 5, 3) {real, imag} */,
  {32'hbebdb656, 32'hbf8370ea} /* (11, 5, 2) {real, imag} */,
  {32'h4058882e, 32'h4044569a} /* (11, 5, 1) {real, imag} */,
  {32'h40a29b4a, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h403ce750, 32'hc06c6448} /* (11, 4, 31) {real, imag} */,
  {32'h3e0e30b8, 32'h3fa68d34} /* (11, 4, 30) {real, imag} */,
  {32'hbda20c4d, 32'h3cfb2cf8} /* (11, 4, 29) {real, imag} */,
  {32'hbe13fca8, 32'h3e5b073a} /* (11, 4, 28) {real, imag} */,
  {32'hbe610d2a, 32'hbdd60b20} /* (11, 4, 27) {real, imag} */,
  {32'h3c861a18, 32'h3d5b9080} /* (11, 4, 26) {real, imag} */,
  {32'hbd8e103a, 32'hbd64546d} /* (11, 4, 25) {real, imag} */,
  {32'hbd41b4f5, 32'h3e1f7878} /* (11, 4, 24) {real, imag} */,
  {32'hbd2200b6, 32'hbd6f0550} /* (11, 4, 23) {real, imag} */,
  {32'h3e16f171, 32'h3ca2049c} /* (11, 4, 22) {real, imag} */,
  {32'hbd64442c, 32'hbc93aa9d} /* (11, 4, 21) {real, imag} */,
  {32'hbd473ce8, 32'h3d8f3e81} /* (11, 4, 20) {real, imag} */,
  {32'h3d7f1afb, 32'h3c3374aa} /* (11, 4, 19) {real, imag} */,
  {32'h3d93dfe6, 32'h3d413840} /* (11, 4, 18) {real, imag} */,
  {32'hbd957354, 32'hbceec611} /* (11, 4, 17) {real, imag} */,
  {32'hbb5b7140, 32'h00000000} /* (11, 4, 16) {real, imag} */,
  {32'hbd957354, 32'h3ceec611} /* (11, 4, 15) {real, imag} */,
  {32'h3d93dfe6, 32'hbd413840} /* (11, 4, 14) {real, imag} */,
  {32'h3d7f1afb, 32'hbc3374aa} /* (11, 4, 13) {real, imag} */,
  {32'hbd473ce8, 32'hbd8f3e81} /* (11, 4, 12) {real, imag} */,
  {32'hbd64442c, 32'h3c93aa9d} /* (11, 4, 11) {real, imag} */,
  {32'h3e16f171, 32'hbca2049c} /* (11, 4, 10) {real, imag} */,
  {32'hbd2200b6, 32'h3d6f0550} /* (11, 4, 9) {real, imag} */,
  {32'hbd41b4f5, 32'hbe1f7878} /* (11, 4, 8) {real, imag} */,
  {32'hbd8e103a, 32'h3d64546d} /* (11, 4, 7) {real, imag} */,
  {32'h3c861a18, 32'hbd5b9080} /* (11, 4, 6) {real, imag} */,
  {32'hbe610d2a, 32'h3dd60b20} /* (11, 4, 5) {real, imag} */,
  {32'hbe13fca8, 32'hbe5b073a} /* (11, 4, 4) {real, imag} */,
  {32'hbda20c4d, 32'hbcfb2cf8} /* (11, 4, 3) {real, imag} */,
  {32'h3e0e30b8, 32'hbfa68d34} /* (11, 4, 2) {real, imag} */,
  {32'h403ce750, 32'h406c6448} /* (11, 4, 1) {real, imag} */,
  {32'h40b0555a, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h4046af41, 32'hc07ec301} /* (11, 3, 31) {real, imag} */,
  {32'h3e7a0814, 32'h3f8ef4be} /* (11, 3, 30) {real, imag} */,
  {32'hbdc23cc6, 32'hbd34ddca} /* (11, 3, 29) {real, imag} */,
  {32'hbe2a6e72, 32'h3e6ab9fe} /* (11, 3, 28) {real, imag} */,
  {32'hbe758d2e, 32'hbdb5d2ff} /* (11, 3, 27) {real, imag} */,
  {32'hbd66ed88, 32'h3d852599} /* (11, 3, 26) {real, imag} */,
  {32'hbd0d0264, 32'h3c3dcce8} /* (11, 3, 25) {real, imag} */,
  {32'h3cfca5ee, 32'h3dcf4001} /* (11, 3, 24) {real, imag} */,
  {32'h3d2798e4, 32'h3d8a4f96} /* (11, 3, 23) {real, imag} */,
  {32'h3d18feb8, 32'h3d3f900e} /* (11, 3, 22) {real, imag} */,
  {32'hbda1cfcf, 32'hbd15df2a} /* (11, 3, 21) {real, imag} */,
  {32'hbc1fb56b, 32'h3cd6c49e} /* (11, 3, 20) {real, imag} */,
  {32'hbd22c0f8, 32'hbe152d12} /* (11, 3, 19) {real, imag} */,
  {32'h3db5dff0, 32'hbcc002f4} /* (11, 3, 18) {real, imag} */,
  {32'hbd2edfb6, 32'h3c00c9e2} /* (11, 3, 17) {real, imag} */,
  {32'hbbce491c, 32'h00000000} /* (11, 3, 16) {real, imag} */,
  {32'hbd2edfb6, 32'hbc00c9e2} /* (11, 3, 15) {real, imag} */,
  {32'h3db5dff0, 32'h3cc002f4} /* (11, 3, 14) {real, imag} */,
  {32'hbd22c0f8, 32'h3e152d12} /* (11, 3, 13) {real, imag} */,
  {32'hbc1fb56b, 32'hbcd6c49e} /* (11, 3, 12) {real, imag} */,
  {32'hbda1cfcf, 32'h3d15df2a} /* (11, 3, 11) {real, imag} */,
  {32'h3d18feb8, 32'hbd3f900e} /* (11, 3, 10) {real, imag} */,
  {32'h3d2798e4, 32'hbd8a4f96} /* (11, 3, 9) {real, imag} */,
  {32'h3cfca5ee, 32'hbdcf4001} /* (11, 3, 8) {real, imag} */,
  {32'hbd0d0264, 32'hbc3dcce8} /* (11, 3, 7) {real, imag} */,
  {32'hbd66ed88, 32'hbd852599} /* (11, 3, 6) {real, imag} */,
  {32'hbe758d2e, 32'h3db5d2ff} /* (11, 3, 5) {real, imag} */,
  {32'hbe2a6e72, 32'hbe6ab9fe} /* (11, 3, 4) {real, imag} */,
  {32'hbdc23cc6, 32'h3d34ddca} /* (11, 3, 3) {real, imag} */,
  {32'h3e7a0814, 32'hbf8ef4be} /* (11, 3, 2) {real, imag} */,
  {32'h4046af41, 32'h407ec301} /* (11, 3, 1) {real, imag} */,
  {32'h40ae2263, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'h404e644a, 32'hc07ce094} /* (11, 2, 31) {real, imag} */,
  {32'h3e81981a, 32'h3f8e95dd} /* (11, 2, 30) {real, imag} */,
  {32'hbd331baa, 32'hbbd80c58} /* (11, 2, 29) {real, imag} */,
  {32'hbe4f1ba4, 32'h3eac5bdc} /* (11, 2, 28) {real, imag} */,
  {32'hbe80a36c, 32'hbd890c33} /* (11, 2, 27) {real, imag} */,
  {32'hbe1113c6, 32'h3c828d68} /* (11, 2, 26) {real, imag} */,
  {32'h3c5ea0dc, 32'hbbeaa828} /* (11, 2, 25) {real, imag} */,
  {32'h3e11dd34, 32'h3c5a57e8} /* (11, 2, 24) {real, imag} */,
  {32'hba960e60, 32'hbbb24c88} /* (11, 2, 23) {real, imag} */,
  {32'hbd8d2aa8, 32'h3dacfc09} /* (11, 2, 22) {real, imag} */,
  {32'hbcf9f58a, 32'hbd560cd0} /* (11, 2, 21) {real, imag} */,
  {32'hbde8b59a, 32'hbd33280a} /* (11, 2, 20) {real, imag} */,
  {32'hbd5fb0fa, 32'hbd62e5a7} /* (11, 2, 19) {real, imag} */,
  {32'h3d566bcb, 32'h3cf04e52} /* (11, 2, 18) {real, imag} */,
  {32'h3cea59b5, 32'hbcb1732b} /* (11, 2, 17) {real, imag} */,
  {32'hbd017f78, 32'h00000000} /* (11, 2, 16) {real, imag} */,
  {32'h3cea59b5, 32'h3cb1732b} /* (11, 2, 15) {real, imag} */,
  {32'h3d566bcb, 32'hbcf04e52} /* (11, 2, 14) {real, imag} */,
  {32'hbd5fb0fa, 32'h3d62e5a7} /* (11, 2, 13) {real, imag} */,
  {32'hbde8b59a, 32'h3d33280a} /* (11, 2, 12) {real, imag} */,
  {32'hbcf9f58a, 32'h3d560cd0} /* (11, 2, 11) {real, imag} */,
  {32'hbd8d2aa8, 32'hbdacfc09} /* (11, 2, 10) {real, imag} */,
  {32'hba960e60, 32'h3bb24c88} /* (11, 2, 9) {real, imag} */,
  {32'h3e11dd34, 32'hbc5a57e8} /* (11, 2, 8) {real, imag} */,
  {32'h3c5ea0dc, 32'h3beaa828} /* (11, 2, 7) {real, imag} */,
  {32'hbe1113c6, 32'hbc828d68} /* (11, 2, 6) {real, imag} */,
  {32'hbe80a36c, 32'h3d890c33} /* (11, 2, 5) {real, imag} */,
  {32'hbe4f1ba4, 32'hbeac5bdc} /* (11, 2, 4) {real, imag} */,
  {32'hbd331baa, 32'h3bd80c58} /* (11, 2, 3) {real, imag} */,
  {32'h3e81981a, 32'hbf8e95dd} /* (11, 2, 2) {real, imag} */,
  {32'h404e644a, 32'h407ce094} /* (11, 2, 1) {real, imag} */,
  {32'h40acc3c1, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'h4056c645, 32'hc06b2684} /* (11, 1, 31) {real, imag} */,
  {32'h3cf975a0, 32'h3f658441} /* (11, 1, 30) {real, imag} */,
  {32'hbde87718, 32'hbd7aec52} /* (11, 1, 29) {real, imag} */,
  {32'hbe26201c, 32'h3e889cd6} /* (11, 1, 28) {real, imag} */,
  {32'hbe28681a, 32'hbda44c48} /* (11, 1, 27) {real, imag} */,
  {32'hbd39430e, 32'hbaca2b60} /* (11, 1, 26) {real, imag} */,
  {32'h3dfb4a52, 32'h3d8a2af4} /* (11, 1, 25) {real, imag} */,
  {32'h3da6922b, 32'h3d13e642} /* (11, 1, 24) {real, imag} */,
  {32'hbd7e5b56, 32'h3ba1bbe4} /* (11, 1, 23) {real, imag} */,
  {32'hbd4b4343, 32'h3dc1ce9e} /* (11, 1, 22) {real, imag} */,
  {32'h3ce414f8, 32'h3c9af38e} /* (11, 1, 21) {real, imag} */,
  {32'h3d86ac02, 32'hbbaa04ec} /* (11, 1, 20) {real, imag} */,
  {32'hbd82c902, 32'h3d8e390d} /* (11, 1, 19) {real, imag} */,
  {32'h3d296b4d, 32'hbcd53664} /* (11, 1, 18) {real, imag} */,
  {32'hbd15fa2d, 32'h3cce4715} /* (11, 1, 17) {real, imag} */,
  {32'h3ceb74fa, 32'h00000000} /* (11, 1, 16) {real, imag} */,
  {32'hbd15fa2d, 32'hbcce4715} /* (11, 1, 15) {real, imag} */,
  {32'h3d296b4d, 32'h3cd53664} /* (11, 1, 14) {real, imag} */,
  {32'hbd82c902, 32'hbd8e390d} /* (11, 1, 13) {real, imag} */,
  {32'h3d86ac02, 32'h3baa04ec} /* (11, 1, 12) {real, imag} */,
  {32'h3ce414f8, 32'hbc9af38e} /* (11, 1, 11) {real, imag} */,
  {32'hbd4b4343, 32'hbdc1ce9e} /* (11, 1, 10) {real, imag} */,
  {32'hbd7e5b56, 32'hbba1bbe4} /* (11, 1, 9) {real, imag} */,
  {32'h3da6922b, 32'hbd13e642} /* (11, 1, 8) {real, imag} */,
  {32'h3dfb4a52, 32'hbd8a2af4} /* (11, 1, 7) {real, imag} */,
  {32'hbd39430e, 32'h3aca2b60} /* (11, 1, 6) {real, imag} */,
  {32'hbe28681a, 32'h3da44c48} /* (11, 1, 5) {real, imag} */,
  {32'hbe26201c, 32'hbe889cd6} /* (11, 1, 4) {real, imag} */,
  {32'hbde87718, 32'h3d7aec52} /* (11, 1, 3) {real, imag} */,
  {32'h3cf975a0, 32'hbf658441} /* (11, 1, 2) {real, imag} */,
  {32'h4056c645, 32'h406b2684} /* (11, 1, 1) {real, imag} */,
  {32'h40aff029, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h405f585d, 32'hc03ec240} /* (11, 0, 31) {real, imag} */,
  {32'hbe7ae2c8, 32'h3f357374} /* (11, 0, 30) {real, imag} */,
  {32'hbdc71d06, 32'h3beb32a8} /* (11, 0, 29) {real, imag} */,
  {32'hbd408f62, 32'h3e844a58} /* (11, 0, 28) {real, imag} */,
  {32'hbe0fc678, 32'hbd714990} /* (11, 0, 27) {real, imag} */,
  {32'h3c2faa1c, 32'h3d92fc0b} /* (11, 0, 26) {real, imag} */,
  {32'h3dae3f6c, 32'h3d269cec} /* (11, 0, 25) {real, imag} */,
  {32'h3c9b300b, 32'h3b441fc0} /* (11, 0, 24) {real, imag} */,
  {32'hbd847834, 32'h3c76d9cc} /* (11, 0, 23) {real, imag} */,
  {32'h3b20a3c0, 32'hbd176552} /* (11, 0, 22) {real, imag} */,
  {32'hbd3a1a22, 32'h3d14e170} /* (11, 0, 21) {real, imag} */,
  {32'h3d45405e, 32'h3ccf4230} /* (11, 0, 20) {real, imag} */,
  {32'hbc31e72c, 32'h3b745b00} /* (11, 0, 19) {real, imag} */,
  {32'h3c987108, 32'hbb6b7910} /* (11, 0, 18) {real, imag} */,
  {32'hbb141d48, 32'h3bb4d244} /* (11, 0, 17) {real, imag} */,
  {32'hbda3a182, 32'h00000000} /* (11, 0, 16) {real, imag} */,
  {32'hbb141d48, 32'hbbb4d244} /* (11, 0, 15) {real, imag} */,
  {32'h3c987108, 32'h3b6b7910} /* (11, 0, 14) {real, imag} */,
  {32'hbc31e72c, 32'hbb745b00} /* (11, 0, 13) {real, imag} */,
  {32'h3d45405e, 32'hbccf4230} /* (11, 0, 12) {real, imag} */,
  {32'hbd3a1a22, 32'hbd14e170} /* (11, 0, 11) {real, imag} */,
  {32'h3b20a3c0, 32'h3d176552} /* (11, 0, 10) {real, imag} */,
  {32'hbd847834, 32'hbc76d9cc} /* (11, 0, 9) {real, imag} */,
  {32'h3c9b300b, 32'hbb441fc0} /* (11, 0, 8) {real, imag} */,
  {32'h3dae3f6c, 32'hbd269cec} /* (11, 0, 7) {real, imag} */,
  {32'h3c2faa1c, 32'hbd92fc0b} /* (11, 0, 6) {real, imag} */,
  {32'hbe0fc678, 32'h3d714990} /* (11, 0, 5) {real, imag} */,
  {32'hbd408f62, 32'hbe844a58} /* (11, 0, 4) {real, imag} */,
  {32'hbdc71d06, 32'hbbeb32a8} /* (11, 0, 3) {real, imag} */,
  {32'hbe7ae2c8, 32'hbf357374} /* (11, 0, 2) {real, imag} */,
  {32'h405f585d, 32'h403ec240} /* (11, 0, 1) {real, imag} */,
  {32'h40ac3538, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h4080f03b, 32'hc018cf90} /* (10, 31, 31) {real, imag} */,
  {32'hbf54b627, 32'h3f469b0e} /* (10, 31, 30) {real, imag} */,
  {32'hbb346ea0, 32'hbd2e20ef} /* (10, 31, 29) {real, imag} */,
  {32'h3e10d49a, 32'h3d0c2e20} /* (10, 31, 28) {real, imag} */,
  {32'hbe01bdfc, 32'hbcb267ac} /* (10, 31, 27) {real, imag} */,
  {32'h3cef7eeb, 32'h3e055efe} /* (10, 31, 26) {real, imag} */,
  {32'h3d4ee255, 32'h3c36b9e8} /* (10, 31, 25) {real, imag} */,
  {32'hbd2713be, 32'h3d7fe6a7} /* (10, 31, 24) {real, imag} */,
  {32'h3d9c96bc, 32'hbc0f7858} /* (10, 31, 23) {real, imag} */,
  {32'hbc934bfc, 32'h3ca8e942} /* (10, 31, 22) {real, imag} */,
  {32'h3c9df37e, 32'h3ce166aa} /* (10, 31, 21) {real, imag} */,
  {32'h3c194538, 32'h3e1091d6} /* (10, 31, 20) {real, imag} */,
  {32'hbcbd73f3, 32'hbbeb0974} /* (10, 31, 19) {real, imag} */,
  {32'hbc38286c, 32'hbafa8a60} /* (10, 31, 18) {real, imag} */,
  {32'hbb588d80, 32'hbd33fb30} /* (10, 31, 17) {real, imag} */,
  {32'hbc30c1d8, 32'h00000000} /* (10, 31, 16) {real, imag} */,
  {32'hbb588d80, 32'h3d33fb30} /* (10, 31, 15) {real, imag} */,
  {32'hbc38286c, 32'h3afa8a60} /* (10, 31, 14) {real, imag} */,
  {32'hbcbd73f3, 32'h3beb0974} /* (10, 31, 13) {real, imag} */,
  {32'h3c194538, 32'hbe1091d6} /* (10, 31, 12) {real, imag} */,
  {32'h3c9df37e, 32'hbce166aa} /* (10, 31, 11) {real, imag} */,
  {32'hbc934bfc, 32'hbca8e942} /* (10, 31, 10) {real, imag} */,
  {32'h3d9c96bc, 32'h3c0f7858} /* (10, 31, 9) {real, imag} */,
  {32'hbd2713be, 32'hbd7fe6a7} /* (10, 31, 8) {real, imag} */,
  {32'h3d4ee255, 32'hbc36b9e8} /* (10, 31, 7) {real, imag} */,
  {32'h3cef7eeb, 32'hbe055efe} /* (10, 31, 6) {real, imag} */,
  {32'hbe01bdfc, 32'h3cb267ac} /* (10, 31, 5) {real, imag} */,
  {32'h3e10d49a, 32'hbd0c2e20} /* (10, 31, 4) {real, imag} */,
  {32'hbb346ea0, 32'h3d2e20ef} /* (10, 31, 3) {real, imag} */,
  {32'hbf54b627, 32'hbf469b0e} /* (10, 31, 2) {real, imag} */,
  {32'h4080f03b, 32'h4018cf90} /* (10, 31, 1) {real, imag} */,
  {32'h40b1c50f, 32'h00000000} /* (10, 31, 0) {real, imag} */,
  {32'h4093f067, 32'hbfec31ca} /* (10, 30, 31) {real, imag} */,
  {32'hbf9828da, 32'h3f2d9d26} /* (10, 30, 30) {real, imag} */,
  {32'hbb0abc20, 32'hbe0dc6d4} /* (10, 30, 29) {real, imag} */,
  {32'h3e463534, 32'h3bd79560} /* (10, 30, 28) {real, imag} */,
  {32'hbe699034, 32'h3d3f2b7d} /* (10, 30, 27) {real, imag} */,
  {32'hbd585fb7, 32'h3cb5fb28} /* (10, 30, 26) {real, imag} */,
  {32'h3c439e72, 32'hbc402a00} /* (10, 30, 25) {real, imag} */,
  {32'hbbeb7748, 32'h3d45833d} /* (10, 30, 24) {real, imag} */,
  {32'h3d1ce365, 32'h3d23800f} /* (10, 30, 23) {real, imag} */,
  {32'hbe115f7e, 32'h3c918efc} /* (10, 30, 22) {real, imag} */,
  {32'hbda027e9, 32'hbd796a84} /* (10, 30, 21) {real, imag} */,
  {32'hbcf0e658, 32'h3d8162d9} /* (10, 30, 20) {real, imag} */,
  {32'hbbbf6746, 32'h3cfda1ac} /* (10, 30, 19) {real, imag} */,
  {32'hbd95d5b4, 32'h3cb60816} /* (10, 30, 18) {real, imag} */,
  {32'h3d6b0f87, 32'h3c45dcc9} /* (10, 30, 17) {real, imag} */,
  {32'h3c7ca7e4, 32'h00000000} /* (10, 30, 16) {real, imag} */,
  {32'h3d6b0f87, 32'hbc45dcc9} /* (10, 30, 15) {real, imag} */,
  {32'hbd95d5b4, 32'hbcb60816} /* (10, 30, 14) {real, imag} */,
  {32'hbbbf6746, 32'hbcfda1ac} /* (10, 30, 13) {real, imag} */,
  {32'hbcf0e658, 32'hbd8162d9} /* (10, 30, 12) {real, imag} */,
  {32'hbda027e9, 32'h3d796a84} /* (10, 30, 11) {real, imag} */,
  {32'hbe115f7e, 32'hbc918efc} /* (10, 30, 10) {real, imag} */,
  {32'h3d1ce365, 32'hbd23800f} /* (10, 30, 9) {real, imag} */,
  {32'hbbeb7748, 32'hbd45833d} /* (10, 30, 8) {real, imag} */,
  {32'h3c439e72, 32'h3c402a00} /* (10, 30, 7) {real, imag} */,
  {32'hbd585fb7, 32'hbcb5fb28} /* (10, 30, 6) {real, imag} */,
  {32'hbe699034, 32'hbd3f2b7d} /* (10, 30, 5) {real, imag} */,
  {32'h3e463534, 32'hbbd79560} /* (10, 30, 4) {real, imag} */,
  {32'hbb0abc20, 32'h3e0dc6d4} /* (10, 30, 3) {real, imag} */,
  {32'hbf9828da, 32'hbf2d9d26} /* (10, 30, 2) {real, imag} */,
  {32'h4093f067, 32'h3fec31ca} /* (10, 30, 1) {real, imag} */,
  {32'h40b7c5f9, 32'h00000000} /* (10, 30, 0) {real, imag} */,
  {32'h409dd546, 32'hbfb316ef} /* (10, 29, 31) {real, imag} */,
  {32'hbfafa18c, 32'h3efe0bc5} /* (10, 29, 30) {real, imag} */,
  {32'hbc543ef8, 32'hbc456024} /* (10, 29, 29) {real, imag} */,
  {32'h3e4737f2, 32'hbd146870} /* (10, 29, 28) {real, imag} */,
  {32'hbe265b1e, 32'h3d978710} /* (10, 29, 27) {real, imag} */,
  {32'hbbd8bb88, 32'hbd89dd90} /* (10, 29, 26) {real, imag} */,
  {32'hbb514c84, 32'hbe0a94c4} /* (10, 29, 25) {real, imag} */,
  {32'hbd36b42c, 32'h3d1856bc} /* (10, 29, 24) {real, imag} */,
  {32'hbb7afc9c, 32'hbca1d2f8} /* (10, 29, 23) {real, imag} */,
  {32'h3d6f0a6b, 32'h3dd0241e} /* (10, 29, 22) {real, imag} */,
  {32'hbd5b2780, 32'h3d4721c4} /* (10, 29, 21) {real, imag} */,
  {32'h3ce7ee84, 32'hbcc0411a} /* (10, 29, 20) {real, imag} */,
  {32'hbba08860, 32'hbc477738} /* (10, 29, 19) {real, imag} */,
  {32'hbc401d2c, 32'h3ddde944} /* (10, 29, 18) {real, imag} */,
  {32'hbca63c70, 32'hbcc9f0da} /* (10, 29, 17) {real, imag} */,
  {32'h3ca93b74, 32'h00000000} /* (10, 29, 16) {real, imag} */,
  {32'hbca63c70, 32'h3cc9f0da} /* (10, 29, 15) {real, imag} */,
  {32'hbc401d2c, 32'hbddde944} /* (10, 29, 14) {real, imag} */,
  {32'hbba08860, 32'h3c477738} /* (10, 29, 13) {real, imag} */,
  {32'h3ce7ee84, 32'h3cc0411a} /* (10, 29, 12) {real, imag} */,
  {32'hbd5b2780, 32'hbd4721c4} /* (10, 29, 11) {real, imag} */,
  {32'h3d6f0a6b, 32'hbdd0241e} /* (10, 29, 10) {real, imag} */,
  {32'hbb7afc9c, 32'h3ca1d2f8} /* (10, 29, 9) {real, imag} */,
  {32'hbd36b42c, 32'hbd1856bc} /* (10, 29, 8) {real, imag} */,
  {32'hbb514c84, 32'h3e0a94c4} /* (10, 29, 7) {real, imag} */,
  {32'hbbd8bb88, 32'h3d89dd90} /* (10, 29, 6) {real, imag} */,
  {32'hbe265b1e, 32'hbd978710} /* (10, 29, 5) {real, imag} */,
  {32'h3e4737f2, 32'h3d146870} /* (10, 29, 4) {real, imag} */,
  {32'hbc543ef8, 32'h3c456024} /* (10, 29, 3) {real, imag} */,
  {32'hbfafa18c, 32'hbefe0bc5} /* (10, 29, 2) {real, imag} */,
  {32'h409dd546, 32'h3fb316ef} /* (10, 29, 1) {real, imag} */,
  {32'h40b8a1ca, 32'h00000000} /* (10, 29, 0) {real, imag} */,
  {32'h40a6b1b6, 32'hbf96c8a2} /* (10, 28, 31) {real, imag} */,
  {32'hbfcf4642, 32'h3f027b76} /* (10, 28, 30) {real, imag} */,
  {32'hbbd9e120, 32'h3df028e1} /* (10, 28, 29) {real, imag} */,
  {32'h3e20701d, 32'hbd923742} /* (10, 28, 28) {real, imag} */,
  {32'hbe0686a2, 32'hbd212966} /* (10, 28, 27) {real, imag} */,
  {32'h3d310954, 32'h3c87c5c2} /* (10, 28, 26) {real, imag} */,
  {32'h3daca3a8, 32'hbcd387f8} /* (10, 28, 25) {real, imag} */,
  {32'hbca6013b, 32'h3d547f80} /* (10, 28, 24) {real, imag} */,
  {32'h3ba22588, 32'hbd94bae0} /* (10, 28, 23) {real, imag} */,
  {32'h3cc8781a, 32'h3e0204d1} /* (10, 28, 22) {real, imag} */,
  {32'hbd525054, 32'h3d8e14bc} /* (10, 28, 21) {real, imag} */,
  {32'hbcf95b86, 32'h3daa6660} /* (10, 28, 20) {real, imag} */,
  {32'hbd7f819e, 32'hbd30204e} /* (10, 28, 19) {real, imag} */,
  {32'hbd4e1f12, 32'hbcd2cb7d} /* (10, 28, 18) {real, imag} */,
  {32'h3c129772, 32'h3da56e0a} /* (10, 28, 17) {real, imag} */,
  {32'hba860e8c, 32'h00000000} /* (10, 28, 16) {real, imag} */,
  {32'h3c129772, 32'hbda56e0a} /* (10, 28, 15) {real, imag} */,
  {32'hbd4e1f12, 32'h3cd2cb7d} /* (10, 28, 14) {real, imag} */,
  {32'hbd7f819e, 32'h3d30204e} /* (10, 28, 13) {real, imag} */,
  {32'hbcf95b86, 32'hbdaa6660} /* (10, 28, 12) {real, imag} */,
  {32'hbd525054, 32'hbd8e14bc} /* (10, 28, 11) {real, imag} */,
  {32'h3cc8781a, 32'hbe0204d1} /* (10, 28, 10) {real, imag} */,
  {32'h3ba22588, 32'h3d94bae0} /* (10, 28, 9) {real, imag} */,
  {32'hbca6013b, 32'hbd547f80} /* (10, 28, 8) {real, imag} */,
  {32'h3daca3a8, 32'h3cd387f8} /* (10, 28, 7) {real, imag} */,
  {32'h3d310954, 32'hbc87c5c2} /* (10, 28, 6) {real, imag} */,
  {32'hbe0686a2, 32'h3d212966} /* (10, 28, 5) {real, imag} */,
  {32'h3e20701d, 32'h3d923742} /* (10, 28, 4) {real, imag} */,
  {32'hbbd9e120, 32'hbdf028e1} /* (10, 28, 3) {real, imag} */,
  {32'hbfcf4642, 32'hbf027b76} /* (10, 28, 2) {real, imag} */,
  {32'h40a6b1b6, 32'h3f96c8a2} /* (10, 28, 1) {real, imag} */,
  {32'h40b628e2, 32'h00000000} /* (10, 28, 0) {real, imag} */,
  {32'h40aef8f8, 32'hbf8aca0f} /* (10, 27, 31) {real, imag} */,
  {32'hbfec8f80, 32'h3e9e8ed7} /* (10, 27, 30) {real, imag} */,
  {32'hbd1e0849, 32'h3e19e569} /* (10, 27, 29) {real, imag} */,
  {32'h3dc3923a, 32'hbdd8ce28} /* (10, 27, 28) {real, imag} */,
  {32'hbe165064, 32'hbc90605c} /* (10, 27, 27) {real, imag} */,
  {32'h3bafeb08, 32'h3c81215d} /* (10, 27, 26) {real, imag} */,
  {32'h3e34948d, 32'hbda244dd} /* (10, 27, 25) {real, imag} */,
  {32'hbc55a0d0, 32'h3d825c40} /* (10, 27, 24) {real, imag} */,
  {32'hbd9cb432, 32'h3debbdfe} /* (10, 27, 23) {real, imag} */,
  {32'h3cc44317, 32'h3d3ab8b9} /* (10, 27, 22) {real, imag} */,
  {32'h3da2a73e, 32'h3deed5b0} /* (10, 27, 21) {real, imag} */,
  {32'h3c2e6489, 32'hbd82bd20} /* (10, 27, 20) {real, imag} */,
  {32'h3d6f91b5, 32'hbdedab30} /* (10, 27, 19) {real, imag} */,
  {32'h3bc646e0, 32'hbd98eb06} /* (10, 27, 18) {real, imag} */,
  {32'hbd250540, 32'h3ceaa78a} /* (10, 27, 17) {real, imag} */,
  {32'h3bc392f4, 32'h00000000} /* (10, 27, 16) {real, imag} */,
  {32'hbd250540, 32'hbceaa78a} /* (10, 27, 15) {real, imag} */,
  {32'h3bc646e0, 32'h3d98eb06} /* (10, 27, 14) {real, imag} */,
  {32'h3d6f91b5, 32'h3dedab30} /* (10, 27, 13) {real, imag} */,
  {32'h3c2e6489, 32'h3d82bd20} /* (10, 27, 12) {real, imag} */,
  {32'h3da2a73e, 32'hbdeed5b0} /* (10, 27, 11) {real, imag} */,
  {32'h3cc44317, 32'hbd3ab8b9} /* (10, 27, 10) {real, imag} */,
  {32'hbd9cb432, 32'hbdebbdfe} /* (10, 27, 9) {real, imag} */,
  {32'hbc55a0d0, 32'hbd825c40} /* (10, 27, 8) {real, imag} */,
  {32'h3e34948d, 32'h3da244dd} /* (10, 27, 7) {real, imag} */,
  {32'h3bafeb08, 32'hbc81215d} /* (10, 27, 6) {real, imag} */,
  {32'hbe165064, 32'h3c90605c} /* (10, 27, 5) {real, imag} */,
  {32'h3dc3923a, 32'h3dd8ce28} /* (10, 27, 4) {real, imag} */,
  {32'hbd1e0849, 32'hbe19e569} /* (10, 27, 3) {real, imag} */,
  {32'hbfec8f80, 32'hbe9e8ed7} /* (10, 27, 2) {real, imag} */,
  {32'h40aef8f8, 32'h3f8aca0f} /* (10, 27, 1) {real, imag} */,
  {32'h40b32c28, 32'h00000000} /* (10, 27, 0) {real, imag} */,
  {32'h40a79d8d, 32'hbf2e7222} /* (10, 26, 31) {real, imag} */,
  {32'hbfee9508, 32'h3e5d0ac0} /* (10, 26, 30) {real, imag} */,
  {32'hbc501076, 32'h3d967686} /* (10, 26, 29) {real, imag} */,
  {32'h3e63ce5d, 32'hbd82ccf4} /* (10, 26, 28) {real, imag} */,
  {32'hbe0b4066, 32'h3e081f1f} /* (10, 26, 27) {real, imag} */,
  {32'hbe30252b, 32'hbd78af61} /* (10, 26, 26) {real, imag} */,
  {32'h3c3947d4, 32'h3d375f27} /* (10, 26, 25) {real, imag} */,
  {32'hbe00488f, 32'h3ddc4bbf} /* (10, 26, 24) {real, imag} */,
  {32'h3ddde07c, 32'h3d5ab044} /* (10, 26, 23) {real, imag} */,
  {32'hbd0b4f65, 32'hbd90e732} /* (10, 26, 22) {real, imag} */,
  {32'h3c21c2cc, 32'h3caea934} /* (10, 26, 21) {real, imag} */,
  {32'h3d8b5b5f, 32'h3c450dc0} /* (10, 26, 20) {real, imag} */,
  {32'h3dd65b86, 32'hbe03cc95} /* (10, 26, 19) {real, imag} */,
  {32'h3d80628e, 32'hbdd2881f} /* (10, 26, 18) {real, imag} */,
  {32'hbcd67ac8, 32'h3d216e96} /* (10, 26, 17) {real, imag} */,
  {32'hbd8b3b5c, 32'h00000000} /* (10, 26, 16) {real, imag} */,
  {32'hbcd67ac8, 32'hbd216e96} /* (10, 26, 15) {real, imag} */,
  {32'h3d80628e, 32'h3dd2881f} /* (10, 26, 14) {real, imag} */,
  {32'h3dd65b86, 32'h3e03cc95} /* (10, 26, 13) {real, imag} */,
  {32'h3d8b5b5f, 32'hbc450dc0} /* (10, 26, 12) {real, imag} */,
  {32'h3c21c2cc, 32'hbcaea934} /* (10, 26, 11) {real, imag} */,
  {32'hbd0b4f65, 32'h3d90e732} /* (10, 26, 10) {real, imag} */,
  {32'h3ddde07c, 32'hbd5ab044} /* (10, 26, 9) {real, imag} */,
  {32'hbe00488f, 32'hbddc4bbf} /* (10, 26, 8) {real, imag} */,
  {32'h3c3947d4, 32'hbd375f27} /* (10, 26, 7) {real, imag} */,
  {32'hbe30252b, 32'h3d78af61} /* (10, 26, 6) {real, imag} */,
  {32'hbe0b4066, 32'hbe081f1f} /* (10, 26, 5) {real, imag} */,
  {32'h3e63ce5d, 32'h3d82ccf4} /* (10, 26, 4) {real, imag} */,
  {32'hbc501076, 32'hbd967686} /* (10, 26, 3) {real, imag} */,
  {32'hbfee9508, 32'hbe5d0ac0} /* (10, 26, 2) {real, imag} */,
  {32'h40a79d8d, 32'h3f2e7222} /* (10, 26, 1) {real, imag} */,
  {32'h40a8b93b, 32'h00000000} /* (10, 26, 0) {real, imag} */,
  {32'h4099a6c9, 32'hbec91c94} /* (10, 25, 31) {real, imag} */,
  {32'hbfe887b2, 32'h3e96e2dc} /* (10, 25, 30) {real, imag} */,
  {32'hbd129858, 32'h3c84f95e} /* (10, 25, 29) {real, imag} */,
  {32'h3deb3ff6, 32'hbde1978c} /* (10, 25, 28) {real, imag} */,
  {32'hbdbe79c8, 32'h3da45232} /* (10, 25, 27) {real, imag} */,
  {32'hbd6c63bd, 32'hbdb1df4d} /* (10, 25, 26) {real, imag} */,
  {32'h3b3b9738, 32'h3d8f136e} /* (10, 25, 25) {real, imag} */,
  {32'h3c90ffd9, 32'h3dcbde30} /* (10, 25, 24) {real, imag} */,
  {32'h3d924226, 32'h3d415bef} /* (10, 25, 23) {real, imag} */,
  {32'hbcca6bac, 32'hbdca50ec} /* (10, 25, 22) {real, imag} */,
  {32'hbd64e0aa, 32'hbca03d7f} /* (10, 25, 21) {real, imag} */,
  {32'hbd246f26, 32'hbd2fa6b8} /* (10, 25, 20) {real, imag} */,
  {32'hbc500a6d, 32'h3d3811b4} /* (10, 25, 19) {real, imag} */,
  {32'hbcdcae1c, 32'hbd999d88} /* (10, 25, 18) {real, imag} */,
  {32'hbd4498c7, 32'h3c3add78} /* (10, 25, 17) {real, imag} */,
  {32'hbc5710a8, 32'h00000000} /* (10, 25, 16) {real, imag} */,
  {32'hbd4498c7, 32'hbc3add78} /* (10, 25, 15) {real, imag} */,
  {32'hbcdcae1c, 32'h3d999d88} /* (10, 25, 14) {real, imag} */,
  {32'hbc500a6d, 32'hbd3811b4} /* (10, 25, 13) {real, imag} */,
  {32'hbd246f26, 32'h3d2fa6b8} /* (10, 25, 12) {real, imag} */,
  {32'hbd64e0aa, 32'h3ca03d7f} /* (10, 25, 11) {real, imag} */,
  {32'hbcca6bac, 32'h3dca50ec} /* (10, 25, 10) {real, imag} */,
  {32'h3d924226, 32'hbd415bef} /* (10, 25, 9) {real, imag} */,
  {32'h3c90ffd9, 32'hbdcbde30} /* (10, 25, 8) {real, imag} */,
  {32'h3b3b9738, 32'hbd8f136e} /* (10, 25, 7) {real, imag} */,
  {32'hbd6c63bd, 32'h3db1df4d} /* (10, 25, 6) {real, imag} */,
  {32'hbdbe79c8, 32'hbda45232} /* (10, 25, 5) {real, imag} */,
  {32'h3deb3ff6, 32'h3de1978c} /* (10, 25, 4) {real, imag} */,
  {32'hbd129858, 32'hbc84f95e} /* (10, 25, 3) {real, imag} */,
  {32'hbfe887b2, 32'hbe96e2dc} /* (10, 25, 2) {real, imag} */,
  {32'h4099a6c9, 32'h3ec91c94} /* (10, 25, 1) {real, imag} */,
  {32'h40994bc2, 32'h00000000} /* (10, 25, 0) {real, imag} */,
  {32'h40895a36, 32'hbe6b3350} /* (10, 24, 31) {real, imag} */,
  {32'hbfc23e0f, 32'h3e4da510} /* (10, 24, 30) {real, imag} */,
  {32'hbe408e56, 32'h39bcdf80} /* (10, 24, 29) {real, imag} */,
  {32'h3e81845a, 32'hbce7a988} /* (10, 24, 28) {real, imag} */,
  {32'hbe3d0116, 32'h3e694a81} /* (10, 24, 27) {real, imag} */,
  {32'hbda90ecc, 32'h3dadb81a} /* (10, 24, 26) {real, imag} */,
  {32'h3d8c68a6, 32'hbaf9d600} /* (10, 24, 25) {real, imag} */,
  {32'hbdf28647, 32'h3d260cfa} /* (10, 24, 24) {real, imag} */,
  {32'h3d4072b3, 32'hbd678f7a} /* (10, 24, 23) {real, imag} */,
  {32'h3d81791a, 32'hbd806e7d} /* (10, 24, 22) {real, imag} */,
  {32'hbd955b6d, 32'h3d5dcbff} /* (10, 24, 21) {real, imag} */,
  {32'h3d91c43f, 32'hbdc4efb3} /* (10, 24, 20) {real, imag} */,
  {32'h3d51654a, 32'hbcab9638} /* (10, 24, 19) {real, imag} */,
  {32'h3d98a3f8, 32'hbc16e584} /* (10, 24, 18) {real, imag} */,
  {32'h3d9f6c5e, 32'hbd8790a5} /* (10, 24, 17) {real, imag} */,
  {32'h3d40a552, 32'h00000000} /* (10, 24, 16) {real, imag} */,
  {32'h3d9f6c5e, 32'h3d8790a5} /* (10, 24, 15) {real, imag} */,
  {32'h3d98a3f8, 32'h3c16e584} /* (10, 24, 14) {real, imag} */,
  {32'h3d51654a, 32'h3cab9638} /* (10, 24, 13) {real, imag} */,
  {32'h3d91c43f, 32'h3dc4efb3} /* (10, 24, 12) {real, imag} */,
  {32'hbd955b6d, 32'hbd5dcbff} /* (10, 24, 11) {real, imag} */,
  {32'h3d81791a, 32'h3d806e7d} /* (10, 24, 10) {real, imag} */,
  {32'h3d4072b3, 32'h3d678f7a} /* (10, 24, 9) {real, imag} */,
  {32'hbdf28647, 32'hbd260cfa} /* (10, 24, 8) {real, imag} */,
  {32'h3d8c68a6, 32'h3af9d600} /* (10, 24, 7) {real, imag} */,
  {32'hbda90ecc, 32'hbdadb81a} /* (10, 24, 6) {real, imag} */,
  {32'hbe3d0116, 32'hbe694a81} /* (10, 24, 5) {real, imag} */,
  {32'h3e81845a, 32'h3ce7a988} /* (10, 24, 4) {real, imag} */,
  {32'hbe408e56, 32'hb9bcdf80} /* (10, 24, 3) {real, imag} */,
  {32'hbfc23e0f, 32'hbe4da510} /* (10, 24, 2) {real, imag} */,
  {32'h40895a36, 32'h3e6b3350} /* (10, 24, 1) {real, imag} */,
  {32'h40851561, 32'h00000000} /* (10, 24, 0) {real, imag} */,
  {32'h405dafa0, 32'hbd101ee0} /* (10, 23, 31) {real, imag} */,
  {32'hbfa45294, 32'h3e055d0a} /* (10, 23, 30) {real, imag} */,
  {32'hbe643eb2, 32'h3df1491d} /* (10, 23, 29) {real, imag} */,
  {32'h3ea2a212, 32'hbe0fccd7} /* (10, 23, 28) {real, imag} */,
  {32'hbe5bb39b, 32'h3e9c1384} /* (10, 23, 27) {real, imag} */,
  {32'hbc7a2eec, 32'hbcc89022} /* (10, 23, 26) {real, imag} */,
  {32'h3be1f5d0, 32'hbb526a60} /* (10, 23, 25) {real, imag} */,
  {32'hbda9c799, 32'h3e092064} /* (10, 23, 24) {real, imag} */,
  {32'h3d8b313e, 32'hbd168ac4} /* (10, 23, 23) {real, imag} */,
  {32'h3db271db, 32'hbd9a0eca} /* (10, 23, 22) {real, imag} */,
  {32'hbc94509d, 32'h3e1f4596} /* (10, 23, 21) {real, imag} */,
  {32'h3d317465, 32'h3d640eb8} /* (10, 23, 20) {real, imag} */,
  {32'hbd98e2bf, 32'hbd8ac306} /* (10, 23, 19) {real, imag} */,
  {32'hbd06dc6f, 32'h3d13096f} /* (10, 23, 18) {real, imag} */,
  {32'hbb241628, 32'h3c87fd3c} /* (10, 23, 17) {real, imag} */,
  {32'hb80e3400, 32'h00000000} /* (10, 23, 16) {real, imag} */,
  {32'hbb241628, 32'hbc87fd3c} /* (10, 23, 15) {real, imag} */,
  {32'hbd06dc6f, 32'hbd13096f} /* (10, 23, 14) {real, imag} */,
  {32'hbd98e2bf, 32'h3d8ac306} /* (10, 23, 13) {real, imag} */,
  {32'h3d317465, 32'hbd640eb8} /* (10, 23, 12) {real, imag} */,
  {32'hbc94509d, 32'hbe1f4596} /* (10, 23, 11) {real, imag} */,
  {32'h3db271db, 32'h3d9a0eca} /* (10, 23, 10) {real, imag} */,
  {32'h3d8b313e, 32'h3d168ac4} /* (10, 23, 9) {real, imag} */,
  {32'hbda9c799, 32'hbe092064} /* (10, 23, 8) {real, imag} */,
  {32'h3be1f5d0, 32'h3b526a60} /* (10, 23, 7) {real, imag} */,
  {32'hbc7a2eec, 32'h3cc89022} /* (10, 23, 6) {real, imag} */,
  {32'hbe5bb39b, 32'hbe9c1384} /* (10, 23, 5) {real, imag} */,
  {32'h3ea2a212, 32'h3e0fccd7} /* (10, 23, 4) {real, imag} */,
  {32'hbe643eb2, 32'hbdf1491d} /* (10, 23, 3) {real, imag} */,
  {32'hbfa45294, 32'hbe055d0a} /* (10, 23, 2) {real, imag} */,
  {32'h405dafa0, 32'h3d101ee0} /* (10, 23, 1) {real, imag} */,
  {32'h40513cf4, 32'h00000000} /* (10, 23, 0) {real, imag} */,
  {32'h401b0e92, 32'hbde9904c} /* (10, 22, 31) {real, imag} */,
  {32'hbf5220f2, 32'h3dec1e2a} /* (10, 22, 30) {real, imag} */,
  {32'hbe0230c2, 32'h3e156bd6} /* (10, 22, 29) {real, imag} */,
  {32'h3e3bbb67, 32'hbca4e6dc} /* (10, 22, 28) {real, imag} */,
  {32'hbe51dee8, 32'h3d8a42ca} /* (10, 22, 27) {real, imag} */,
  {32'h3dc44452, 32'h3d65f7f0} /* (10, 22, 26) {real, imag} */,
  {32'hbe361fde, 32'hbcbfdf74} /* (10, 22, 25) {real, imag} */,
  {32'hbd8c0b40, 32'h3d51a38e} /* (10, 22, 24) {real, imag} */,
  {32'hbbaca9dc, 32'hba950aa0} /* (10, 22, 23) {real, imag} */,
  {32'hbd015257, 32'hbddd64e8} /* (10, 22, 22) {real, imag} */,
  {32'h3cc22396, 32'h3c745ec9} /* (10, 22, 21) {real, imag} */,
  {32'hbd63b494, 32'hbd74ca72} /* (10, 22, 20) {real, imag} */,
  {32'h3d08746d, 32'h3c43b09c} /* (10, 22, 19) {real, imag} */,
  {32'h3d677ef1, 32'h3d8a8378} /* (10, 22, 18) {real, imag} */,
  {32'h3d2d3d70, 32'hbb95ad94} /* (10, 22, 17) {real, imag} */,
  {32'h3daf7758, 32'h00000000} /* (10, 22, 16) {real, imag} */,
  {32'h3d2d3d70, 32'h3b95ad94} /* (10, 22, 15) {real, imag} */,
  {32'h3d677ef1, 32'hbd8a8378} /* (10, 22, 14) {real, imag} */,
  {32'h3d08746d, 32'hbc43b09c} /* (10, 22, 13) {real, imag} */,
  {32'hbd63b494, 32'h3d74ca72} /* (10, 22, 12) {real, imag} */,
  {32'h3cc22396, 32'hbc745ec9} /* (10, 22, 11) {real, imag} */,
  {32'hbd015257, 32'h3ddd64e8} /* (10, 22, 10) {real, imag} */,
  {32'hbbaca9dc, 32'h3a950aa0} /* (10, 22, 9) {real, imag} */,
  {32'hbd8c0b40, 32'hbd51a38e} /* (10, 22, 8) {real, imag} */,
  {32'hbe361fde, 32'h3cbfdf74} /* (10, 22, 7) {real, imag} */,
  {32'h3dc44452, 32'hbd65f7f0} /* (10, 22, 6) {real, imag} */,
  {32'hbe51dee8, 32'hbd8a42ca} /* (10, 22, 5) {real, imag} */,
  {32'h3e3bbb67, 32'h3ca4e6dc} /* (10, 22, 4) {real, imag} */,
  {32'hbe0230c2, 32'hbe156bd6} /* (10, 22, 3) {real, imag} */,
  {32'hbf5220f2, 32'hbdec1e2a} /* (10, 22, 2) {real, imag} */,
  {32'h401b0e92, 32'h3de9904c} /* (10, 22, 1) {real, imag} */,
  {32'h400afd88, 32'h00000000} /* (10, 22, 0) {real, imag} */,
  {32'h3f2f3040, 32'hbdb83a24} /* (10, 21, 31) {real, imag} */,
  {32'hbe3bd36e, 32'hbb3b7980} /* (10, 21, 30) {real, imag} */,
  {32'hbcc4880e, 32'h3d98e9de} /* (10, 21, 29) {real, imag} */,
  {32'h3db75536, 32'hbd8a7289} /* (10, 21, 28) {real, imag} */,
  {32'hbe3c9fc6, 32'h3d1fadc2} /* (10, 21, 27) {real, imag} */,
  {32'h3de8524c, 32'h3c930bf7} /* (10, 21, 26) {real, imag} */,
  {32'hbce72246, 32'hbd8c6292} /* (10, 21, 25) {real, imag} */,
  {32'hbd836b6a, 32'h3d615fc0} /* (10, 21, 24) {real, imag} */,
  {32'hbd5a140c, 32'h3d91def4} /* (10, 21, 23) {real, imag} */,
  {32'hbd3049aa, 32'hbd0585cf} /* (10, 21, 22) {real, imag} */,
  {32'h3d151d41, 32'h3da6bc14} /* (10, 21, 21) {real, imag} */,
  {32'h3d9b72e7, 32'hbd2ff6dd} /* (10, 21, 20) {real, imag} */,
  {32'h3d1735af, 32'h3d2d2411} /* (10, 21, 19) {real, imag} */,
  {32'h3d3b73ee, 32'hbbf01afa} /* (10, 21, 18) {real, imag} */,
  {32'h3d6da5be, 32'h3cd4e52e} /* (10, 21, 17) {real, imag} */,
  {32'hbc29c02a, 32'h00000000} /* (10, 21, 16) {real, imag} */,
  {32'h3d6da5be, 32'hbcd4e52e} /* (10, 21, 15) {real, imag} */,
  {32'h3d3b73ee, 32'h3bf01afa} /* (10, 21, 14) {real, imag} */,
  {32'h3d1735af, 32'hbd2d2411} /* (10, 21, 13) {real, imag} */,
  {32'h3d9b72e7, 32'h3d2ff6dd} /* (10, 21, 12) {real, imag} */,
  {32'h3d151d41, 32'hbda6bc14} /* (10, 21, 11) {real, imag} */,
  {32'hbd3049aa, 32'h3d0585cf} /* (10, 21, 10) {real, imag} */,
  {32'hbd5a140c, 32'hbd91def4} /* (10, 21, 9) {real, imag} */,
  {32'hbd836b6a, 32'hbd615fc0} /* (10, 21, 8) {real, imag} */,
  {32'hbce72246, 32'h3d8c6292} /* (10, 21, 7) {real, imag} */,
  {32'h3de8524c, 32'hbc930bf7} /* (10, 21, 6) {real, imag} */,
  {32'hbe3c9fc6, 32'hbd1fadc2} /* (10, 21, 5) {real, imag} */,
  {32'h3db75536, 32'h3d8a7289} /* (10, 21, 4) {real, imag} */,
  {32'hbcc4880e, 32'hbd98e9de} /* (10, 21, 3) {real, imag} */,
  {32'hbe3bd36e, 32'h3b3b7980} /* (10, 21, 2) {real, imag} */,
  {32'h3f2f3040, 32'h3db83a24} /* (10, 21, 1) {real, imag} */,
  {32'h3f6f4988, 32'h00000000} /* (10, 21, 0) {real, imag} */,
  {32'hbfa872a6, 32'h3de724b8} /* (10, 20, 31) {real, imag} */,
  {32'h3f1e1a40, 32'hbe924854} /* (10, 20, 30) {real, imag} */,
  {32'hbd8f0d60, 32'h3bf924c0} /* (10, 20, 29) {real, imag} */,
  {32'hbe4558de, 32'hbd04a954} /* (10, 20, 28) {real, imag} */,
  {32'h3d78acc8, 32'h3da43bbf} /* (10, 20, 27) {real, imag} */,
  {32'h3d694556, 32'hbe0b6ff9} /* (10, 20, 26) {real, imag} */,
  {32'h3b8b8f48, 32'h3d0e41b6} /* (10, 20, 25) {real, imag} */,
  {32'h3d546e18, 32'hbd0947df} /* (10, 20, 24) {real, imag} */,
  {32'hbd99c178, 32'h3c888b51} /* (10, 20, 23) {real, imag} */,
  {32'h3ca61f23, 32'hbd101020} /* (10, 20, 22) {real, imag} */,
  {32'hbc6034fa, 32'hbd1cef4e} /* (10, 20, 21) {real, imag} */,
  {32'hbba90a48, 32'hbc719544} /* (10, 20, 20) {real, imag} */,
  {32'hbdd5566c, 32'hbdb24178} /* (10, 20, 19) {real, imag} */,
  {32'h3d21e2b0, 32'hbdab0552} /* (10, 20, 18) {real, imag} */,
  {32'h3d367b08, 32'hbcb7d40f} /* (10, 20, 17) {real, imag} */,
  {32'hbc6c4d3e, 32'h00000000} /* (10, 20, 16) {real, imag} */,
  {32'h3d367b08, 32'h3cb7d40f} /* (10, 20, 15) {real, imag} */,
  {32'h3d21e2b0, 32'h3dab0552} /* (10, 20, 14) {real, imag} */,
  {32'hbdd5566c, 32'h3db24178} /* (10, 20, 13) {real, imag} */,
  {32'hbba90a48, 32'h3c719544} /* (10, 20, 12) {real, imag} */,
  {32'hbc6034fa, 32'h3d1cef4e} /* (10, 20, 11) {real, imag} */,
  {32'h3ca61f23, 32'h3d101020} /* (10, 20, 10) {real, imag} */,
  {32'hbd99c178, 32'hbc888b51} /* (10, 20, 9) {real, imag} */,
  {32'h3d546e18, 32'h3d0947df} /* (10, 20, 8) {real, imag} */,
  {32'h3b8b8f48, 32'hbd0e41b6} /* (10, 20, 7) {real, imag} */,
  {32'h3d694556, 32'h3e0b6ff9} /* (10, 20, 6) {real, imag} */,
  {32'h3d78acc8, 32'hbda43bbf} /* (10, 20, 5) {real, imag} */,
  {32'hbe4558de, 32'h3d04a954} /* (10, 20, 4) {real, imag} */,
  {32'hbd8f0d60, 32'hbbf924c0} /* (10, 20, 3) {real, imag} */,
  {32'h3f1e1a40, 32'h3e924854} /* (10, 20, 2) {real, imag} */,
  {32'hbfa872a6, 32'hbde724b8} /* (10, 20, 1) {real, imag} */,
  {32'hbf10e206, 32'h00000000} /* (10, 20, 0) {real, imag} */,
  {32'hc02b8027, 32'h3ebe2790} /* (10, 19, 31) {real, imag} */,
  {32'h3f80ce54, 32'hbeab1fcd} /* (10, 19, 30) {real, imag} */,
  {32'hbe0b7e36, 32'h3da0547c} /* (10, 19, 29) {real, imag} */,
  {32'hbdabc276, 32'h3dc1e131} /* (10, 19, 28) {real, imag} */,
  {32'h3de3f0d0, 32'h3cb1e204} /* (10, 19, 27) {real, imag} */,
  {32'h3d21af82, 32'hbd7c98fa} /* (10, 19, 26) {real, imag} */,
  {32'hbd570d99, 32'h3baa0f50} /* (10, 19, 25) {real, imag} */,
  {32'h3d8d2829, 32'hbd7e8e72} /* (10, 19, 24) {real, imag} */,
  {32'hbc18e873, 32'hbda89234} /* (10, 19, 23) {real, imag} */,
  {32'h3d1b403e, 32'hbcdca57c} /* (10, 19, 22) {real, imag} */,
  {32'h3d945c52, 32'hbc8aa892} /* (10, 19, 21) {real, imag} */,
  {32'h3c956078, 32'h3d10ed90} /* (10, 19, 20) {real, imag} */,
  {32'hbce31c94, 32'h3a7195a0} /* (10, 19, 19) {real, imag} */,
  {32'hbc5f1693, 32'h3d7de251} /* (10, 19, 18) {real, imag} */,
  {32'hbd0d2002, 32'hbd889e5c} /* (10, 19, 17) {real, imag} */,
  {32'hb9ad69c0, 32'h00000000} /* (10, 19, 16) {real, imag} */,
  {32'hbd0d2002, 32'h3d889e5c} /* (10, 19, 15) {real, imag} */,
  {32'hbc5f1693, 32'hbd7de251} /* (10, 19, 14) {real, imag} */,
  {32'hbce31c94, 32'hba7195a0} /* (10, 19, 13) {real, imag} */,
  {32'h3c956078, 32'hbd10ed90} /* (10, 19, 12) {real, imag} */,
  {32'h3d945c52, 32'h3c8aa892} /* (10, 19, 11) {real, imag} */,
  {32'h3d1b403e, 32'h3cdca57c} /* (10, 19, 10) {real, imag} */,
  {32'hbc18e873, 32'h3da89234} /* (10, 19, 9) {real, imag} */,
  {32'h3d8d2829, 32'h3d7e8e72} /* (10, 19, 8) {real, imag} */,
  {32'hbd570d99, 32'hbbaa0f50} /* (10, 19, 7) {real, imag} */,
  {32'h3d21af82, 32'h3d7c98fa} /* (10, 19, 6) {real, imag} */,
  {32'h3de3f0d0, 32'hbcb1e204} /* (10, 19, 5) {real, imag} */,
  {32'hbdabc276, 32'hbdc1e131} /* (10, 19, 4) {real, imag} */,
  {32'hbe0b7e36, 32'hbda0547c} /* (10, 19, 3) {real, imag} */,
  {32'h3f80ce54, 32'h3eab1fcd} /* (10, 19, 2) {real, imag} */,
  {32'hc02b8027, 32'hbebe2790} /* (10, 19, 1) {real, imag} */,
  {32'hbfe9e0f7, 32'h00000000} /* (10, 19, 0) {real, imag} */,
  {32'hc067cf78, 32'h3ea3eca6} /* (10, 18, 31) {real, imag} */,
  {32'h3faffd84, 32'hbed3d923} /* (10, 18, 30) {real, imag} */,
  {32'h3dab600f, 32'h3e5c23f8} /* (10, 18, 29) {real, imag} */,
  {32'hbe1e1ab6, 32'h3d35363c} /* (10, 18, 28) {real, imag} */,
  {32'h3e0a0924, 32'hbda9e1da} /* (10, 18, 27) {real, imag} */,
  {32'h3dc90e8e, 32'hbd31d8fe} /* (10, 18, 26) {real, imag} */,
  {32'hbd8385fc, 32'h3d42131a} /* (10, 18, 25) {real, imag} */,
  {32'h3d0a51cc, 32'h3bef9440} /* (10, 18, 24) {real, imag} */,
  {32'hbd876c10, 32'h3dda33f0} /* (10, 18, 23) {real, imag} */,
  {32'h3d844687, 32'hbd965f77} /* (10, 18, 22) {real, imag} */,
  {32'h3e0037e0, 32'hbd8ebfdf} /* (10, 18, 21) {real, imag} */,
  {32'hbd850334, 32'hbcef88b5} /* (10, 18, 20) {real, imag} */,
  {32'hbcc7499c, 32'hbd42b1a6} /* (10, 18, 19) {real, imag} */,
  {32'hbc3808d8, 32'hbe17a3a6} /* (10, 18, 18) {real, imag} */,
  {32'hbd009f84, 32'hbd16b921} /* (10, 18, 17) {real, imag} */,
  {32'hbdc4f10e, 32'h00000000} /* (10, 18, 16) {real, imag} */,
  {32'hbd009f84, 32'h3d16b921} /* (10, 18, 15) {real, imag} */,
  {32'hbc3808d8, 32'h3e17a3a6} /* (10, 18, 14) {real, imag} */,
  {32'hbcc7499c, 32'h3d42b1a6} /* (10, 18, 13) {real, imag} */,
  {32'hbd850334, 32'h3cef88b5} /* (10, 18, 12) {real, imag} */,
  {32'h3e0037e0, 32'h3d8ebfdf} /* (10, 18, 11) {real, imag} */,
  {32'h3d844687, 32'h3d965f77} /* (10, 18, 10) {real, imag} */,
  {32'hbd876c10, 32'hbdda33f0} /* (10, 18, 9) {real, imag} */,
  {32'h3d0a51cc, 32'hbbef9440} /* (10, 18, 8) {real, imag} */,
  {32'hbd8385fc, 32'hbd42131a} /* (10, 18, 7) {real, imag} */,
  {32'h3dc90e8e, 32'h3d31d8fe} /* (10, 18, 6) {real, imag} */,
  {32'h3e0a0924, 32'h3da9e1da} /* (10, 18, 5) {real, imag} */,
  {32'hbe1e1ab6, 32'hbd35363c} /* (10, 18, 4) {real, imag} */,
  {32'h3dab600f, 32'hbe5c23f8} /* (10, 18, 3) {real, imag} */,
  {32'h3faffd84, 32'h3ed3d923} /* (10, 18, 2) {real, imag} */,
  {32'hc067cf78, 32'hbea3eca6} /* (10, 18, 1) {real, imag} */,
  {32'hc0324c5a, 32'h00000000} /* (10, 18, 0) {real, imag} */,
  {32'hc085e513, 32'h3eb310d8} /* (10, 17, 31) {real, imag} */,
  {32'h3fd83e41, 32'hbec57f21} /* (10, 17, 30) {real, imag} */,
  {32'h3c29c31c, 32'h3d5887cb} /* (10, 17, 29) {real, imag} */,
  {32'hbe5d90ec, 32'h3b008ba0} /* (10, 17, 28) {real, imag} */,
  {32'h3e74a34a, 32'hbe5b98f5} /* (10, 17, 27) {real, imag} */,
  {32'hbd345198, 32'hbc848e70} /* (10, 17, 26) {real, imag} */,
  {32'h3d535d40, 32'hbd12243e} /* (10, 17, 25) {real, imag} */,
  {32'h3dcc9a53, 32'hbda051be} /* (10, 17, 24) {real, imag} */,
  {32'h3d0627c6, 32'h3df22bef} /* (10, 17, 23) {real, imag} */,
  {32'hbdafe2dd, 32'h3d4db0b9} /* (10, 17, 22) {real, imag} */,
  {32'h3d24ac32, 32'hbd930a32} /* (10, 17, 21) {real, imag} */,
  {32'hbdc26d6a, 32'h398e1600} /* (10, 17, 20) {real, imag} */,
  {32'hbc97c075, 32'h3cfed3e0} /* (10, 17, 19) {real, imag} */,
  {32'h3d88a794, 32'h3ba254dc} /* (10, 17, 18) {real, imag} */,
  {32'hbd3dde0a, 32'h3d747035} /* (10, 17, 17) {real, imag} */,
  {32'hbcd127c7, 32'h00000000} /* (10, 17, 16) {real, imag} */,
  {32'hbd3dde0a, 32'hbd747035} /* (10, 17, 15) {real, imag} */,
  {32'h3d88a794, 32'hbba254dc} /* (10, 17, 14) {real, imag} */,
  {32'hbc97c075, 32'hbcfed3e0} /* (10, 17, 13) {real, imag} */,
  {32'hbdc26d6a, 32'hb98e1600} /* (10, 17, 12) {real, imag} */,
  {32'h3d24ac32, 32'h3d930a32} /* (10, 17, 11) {real, imag} */,
  {32'hbdafe2dd, 32'hbd4db0b9} /* (10, 17, 10) {real, imag} */,
  {32'h3d0627c6, 32'hbdf22bef} /* (10, 17, 9) {real, imag} */,
  {32'h3dcc9a53, 32'h3da051be} /* (10, 17, 8) {real, imag} */,
  {32'h3d535d40, 32'h3d12243e} /* (10, 17, 7) {real, imag} */,
  {32'hbd345198, 32'h3c848e70} /* (10, 17, 6) {real, imag} */,
  {32'h3e74a34a, 32'h3e5b98f5} /* (10, 17, 5) {real, imag} */,
  {32'hbe5d90ec, 32'hbb008ba0} /* (10, 17, 4) {real, imag} */,
  {32'h3c29c31c, 32'hbd5887cb} /* (10, 17, 3) {real, imag} */,
  {32'h3fd83e41, 32'h3ec57f21} /* (10, 17, 2) {real, imag} */,
  {32'hc085e513, 32'hbeb310d8} /* (10, 17, 1) {real, imag} */,
  {32'hc0569797, 32'h00000000} /* (10, 17, 0) {real, imag} */,
  {32'hc08e7ff8, 32'h3ec4e814} /* (10, 16, 31) {real, imag} */,
  {32'h3fd476f2, 32'hbe3b7824} /* (10, 16, 30) {real, imag} */,
  {32'hbc382708, 32'h3c8c3b1a} /* (10, 16, 29) {real, imag} */,
  {32'hbe4652b7, 32'hbd9149f0} /* (10, 16, 28) {real, imag} */,
  {32'h3e8e2f00, 32'hbe2e465b} /* (10, 16, 27) {real, imag} */,
  {32'h3c8355ec, 32'hbd9ab080} /* (10, 16, 26) {real, imag} */,
  {32'h3cd7a34c, 32'hbd117aa3} /* (10, 16, 25) {real, imag} */,
  {32'h3d9bbe3c, 32'h3cfa03fa} /* (10, 16, 24) {real, imag} */,
  {32'h3da37cd0, 32'h3c59fdc6} /* (10, 16, 23) {real, imag} */,
  {32'h3d4c177b, 32'h3cb04017} /* (10, 16, 22) {real, imag} */,
  {32'hbc9a9b20, 32'hbd3e82d9} /* (10, 16, 21) {real, imag} */,
  {32'h3da261e1, 32'hbca60eb6} /* (10, 16, 20) {real, imag} */,
  {32'hbdcba40f, 32'h3c20a0f1} /* (10, 16, 19) {real, imag} */,
  {32'h3cb635c0, 32'h3d38d194} /* (10, 16, 18) {real, imag} */,
  {32'hbc60937b, 32'h3d829e9c} /* (10, 16, 17) {real, imag} */,
  {32'hbd612b11, 32'h00000000} /* (10, 16, 16) {real, imag} */,
  {32'hbc60937b, 32'hbd829e9c} /* (10, 16, 15) {real, imag} */,
  {32'h3cb635c0, 32'hbd38d194} /* (10, 16, 14) {real, imag} */,
  {32'hbdcba40f, 32'hbc20a0f1} /* (10, 16, 13) {real, imag} */,
  {32'h3da261e1, 32'h3ca60eb6} /* (10, 16, 12) {real, imag} */,
  {32'hbc9a9b20, 32'h3d3e82d9} /* (10, 16, 11) {real, imag} */,
  {32'h3d4c177b, 32'hbcb04017} /* (10, 16, 10) {real, imag} */,
  {32'h3da37cd0, 32'hbc59fdc6} /* (10, 16, 9) {real, imag} */,
  {32'h3d9bbe3c, 32'hbcfa03fa} /* (10, 16, 8) {real, imag} */,
  {32'h3cd7a34c, 32'h3d117aa3} /* (10, 16, 7) {real, imag} */,
  {32'h3c8355ec, 32'h3d9ab080} /* (10, 16, 6) {real, imag} */,
  {32'h3e8e2f00, 32'h3e2e465b} /* (10, 16, 5) {real, imag} */,
  {32'hbe4652b7, 32'h3d9149f0} /* (10, 16, 4) {real, imag} */,
  {32'hbc382708, 32'hbc8c3b1a} /* (10, 16, 3) {real, imag} */,
  {32'h3fd476f2, 32'h3e3b7824} /* (10, 16, 2) {real, imag} */,
  {32'hc08e7ff8, 32'hbec4e814} /* (10, 16, 1) {real, imag} */,
  {32'hc05776ad, 32'h00000000} /* (10, 16, 0) {real, imag} */,
  {32'hc08faf05, 32'h3e5c04a0} /* (10, 15, 31) {real, imag} */,
  {32'h3fc84831, 32'hbe246806} /* (10, 15, 30) {real, imag} */,
  {32'h3d6a336b, 32'h3b110b90} /* (10, 15, 29) {real, imag} */,
  {32'hbe98a5fe, 32'hbd1654f6} /* (10, 15, 28) {real, imag} */,
  {32'h3e58a0da, 32'hbdfc59de} /* (10, 15, 27) {real, imag} */,
  {32'h3e16f426, 32'hba359c00} /* (10, 15, 26) {real, imag} */,
  {32'hbd5d965e, 32'h3c9207c0} /* (10, 15, 25) {real, imag} */,
  {32'h3d21b5d2, 32'h3cdde882} /* (10, 15, 24) {real, imag} */,
  {32'h3d2cc6f2, 32'hbdb5202b} /* (10, 15, 23) {real, imag} */,
  {32'hb783d000, 32'hbda39a30} /* (10, 15, 22) {real, imag} */,
  {32'h3db09791, 32'h3c44b97c} /* (10, 15, 21) {real, imag} */,
  {32'h3a762bc0, 32'hbc519680} /* (10, 15, 20) {real, imag} */,
  {32'h3cf07015, 32'h3d1b4a38} /* (10, 15, 19) {real, imag} */,
  {32'h3d99020c, 32'hbcf88ccb} /* (10, 15, 18) {real, imag} */,
  {32'hbd703bcc, 32'hbc2d478c} /* (10, 15, 17) {real, imag} */,
  {32'hbc12a8aa, 32'h00000000} /* (10, 15, 16) {real, imag} */,
  {32'hbd703bcc, 32'h3c2d478c} /* (10, 15, 15) {real, imag} */,
  {32'h3d99020c, 32'h3cf88ccb} /* (10, 15, 14) {real, imag} */,
  {32'h3cf07015, 32'hbd1b4a38} /* (10, 15, 13) {real, imag} */,
  {32'h3a762bc0, 32'h3c519680} /* (10, 15, 12) {real, imag} */,
  {32'h3db09791, 32'hbc44b97c} /* (10, 15, 11) {real, imag} */,
  {32'hb783d000, 32'h3da39a30} /* (10, 15, 10) {real, imag} */,
  {32'h3d2cc6f2, 32'h3db5202b} /* (10, 15, 9) {real, imag} */,
  {32'h3d21b5d2, 32'hbcdde882} /* (10, 15, 8) {real, imag} */,
  {32'hbd5d965e, 32'hbc9207c0} /* (10, 15, 7) {real, imag} */,
  {32'h3e16f426, 32'h3a359c00} /* (10, 15, 6) {real, imag} */,
  {32'h3e58a0da, 32'h3dfc59de} /* (10, 15, 5) {real, imag} */,
  {32'hbe98a5fe, 32'h3d1654f6} /* (10, 15, 4) {real, imag} */,
  {32'h3d6a336b, 32'hbb110b90} /* (10, 15, 3) {real, imag} */,
  {32'h3fc84831, 32'h3e246806} /* (10, 15, 2) {real, imag} */,
  {32'hc08faf05, 32'hbe5c04a0} /* (10, 15, 1) {real, imag} */,
  {32'hc059e171, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'hc0845abe, 32'h3e450a04} /* (10, 14, 31) {real, imag} */,
  {32'h3fb32544, 32'hbe56de32} /* (10, 14, 30) {real, imag} */,
  {32'h3cdb16ed, 32'h3caba214} /* (10, 14, 29) {real, imag} */,
  {32'hbe6b6f32, 32'h3d31e854} /* (10, 14, 28) {real, imag} */,
  {32'h3d8dabd1, 32'hbdde5ef2} /* (10, 14, 27) {real, imag} */,
  {32'h3b854518, 32'h3d7cfd16} /* (10, 14, 26) {real, imag} */,
  {32'hbd680894, 32'hbd330f0e} /* (10, 14, 25) {real, imag} */,
  {32'hbdae1248, 32'hbe1ddc52} /* (10, 14, 24) {real, imag} */,
  {32'hbc38c4d4, 32'hbd377c71} /* (10, 14, 23) {real, imag} */,
  {32'hbd10eee4, 32'h3d943ca7} /* (10, 14, 22) {real, imag} */,
  {32'hbd40192a, 32'hbdbb1529} /* (10, 14, 21) {real, imag} */,
  {32'h3d187d55, 32'hbcc322cf} /* (10, 14, 20) {real, imag} */,
  {32'h3b235774, 32'hbd61fe04} /* (10, 14, 19) {real, imag} */,
  {32'hbcf302c8, 32'hbd85d9d0} /* (10, 14, 18) {real, imag} */,
  {32'hbc5eb6da, 32'h3c03eb25} /* (10, 14, 17) {real, imag} */,
  {32'hbc862f8a, 32'h00000000} /* (10, 14, 16) {real, imag} */,
  {32'hbc5eb6da, 32'hbc03eb25} /* (10, 14, 15) {real, imag} */,
  {32'hbcf302c8, 32'h3d85d9d0} /* (10, 14, 14) {real, imag} */,
  {32'h3b235774, 32'h3d61fe04} /* (10, 14, 13) {real, imag} */,
  {32'h3d187d55, 32'h3cc322cf} /* (10, 14, 12) {real, imag} */,
  {32'hbd40192a, 32'h3dbb1529} /* (10, 14, 11) {real, imag} */,
  {32'hbd10eee4, 32'hbd943ca7} /* (10, 14, 10) {real, imag} */,
  {32'hbc38c4d4, 32'h3d377c71} /* (10, 14, 9) {real, imag} */,
  {32'hbdae1248, 32'h3e1ddc52} /* (10, 14, 8) {real, imag} */,
  {32'hbd680894, 32'h3d330f0e} /* (10, 14, 7) {real, imag} */,
  {32'h3b854518, 32'hbd7cfd16} /* (10, 14, 6) {real, imag} */,
  {32'h3d8dabd1, 32'h3dde5ef2} /* (10, 14, 5) {real, imag} */,
  {32'hbe6b6f32, 32'hbd31e854} /* (10, 14, 4) {real, imag} */,
  {32'h3cdb16ed, 32'hbcaba214} /* (10, 14, 3) {real, imag} */,
  {32'h3fb32544, 32'h3e56de32} /* (10, 14, 2) {real, imag} */,
  {32'hc0845abe, 32'hbe450a04} /* (10, 14, 1) {real, imag} */,
  {32'hc043bc7e, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'hc05f9a51, 32'h3dce24a0} /* (10, 13, 31) {real, imag} */,
  {32'h3fa261c0, 32'hbe4b4b2e} /* (10, 13, 30) {real, imag} */,
  {32'h3dd92580, 32'hb8af6a00} /* (10, 13, 29) {real, imag} */,
  {32'hbe88563a, 32'h3dd46a81} /* (10, 13, 28) {real, imag} */,
  {32'h3da33492, 32'hbe1d2e9e} /* (10, 13, 27) {real, imag} */,
  {32'h3c74885e, 32'hbd1fac96} /* (10, 13, 26) {real, imag} */,
  {32'hbd82c01c, 32'h3b260d40} /* (10, 13, 25) {real, imag} */,
  {32'hbcae7a48, 32'hbd4d1e5e} /* (10, 13, 24) {real, imag} */,
  {32'hbbab697a, 32'h3d1354ef} /* (10, 13, 23) {real, imag} */,
  {32'hbd5f8b44, 32'hbcef8224} /* (10, 13, 22) {real, imag} */,
  {32'hbc67293c, 32'hbc7fad6b} /* (10, 13, 21) {real, imag} */,
  {32'hbbbdf000, 32'hbdd08dca} /* (10, 13, 20) {real, imag} */,
  {32'hbd75d7f0, 32'hbc91e5dd} /* (10, 13, 19) {real, imag} */,
  {32'h3cdaddbe, 32'hbd161cd3} /* (10, 13, 18) {real, imag} */,
  {32'h3d923537, 32'hbcf5765e} /* (10, 13, 17) {real, imag} */,
  {32'h3cd293ff, 32'h00000000} /* (10, 13, 16) {real, imag} */,
  {32'h3d923537, 32'h3cf5765e} /* (10, 13, 15) {real, imag} */,
  {32'h3cdaddbe, 32'h3d161cd3} /* (10, 13, 14) {real, imag} */,
  {32'hbd75d7f0, 32'h3c91e5dd} /* (10, 13, 13) {real, imag} */,
  {32'hbbbdf000, 32'h3dd08dca} /* (10, 13, 12) {real, imag} */,
  {32'hbc67293c, 32'h3c7fad6b} /* (10, 13, 11) {real, imag} */,
  {32'hbd5f8b44, 32'h3cef8224} /* (10, 13, 10) {real, imag} */,
  {32'hbbab697a, 32'hbd1354ef} /* (10, 13, 9) {real, imag} */,
  {32'hbcae7a48, 32'h3d4d1e5e} /* (10, 13, 8) {real, imag} */,
  {32'hbd82c01c, 32'hbb260d40} /* (10, 13, 7) {real, imag} */,
  {32'h3c74885e, 32'h3d1fac96} /* (10, 13, 6) {real, imag} */,
  {32'h3da33492, 32'h3e1d2e9e} /* (10, 13, 5) {real, imag} */,
  {32'hbe88563a, 32'hbdd46a81} /* (10, 13, 4) {real, imag} */,
  {32'h3dd92580, 32'h38af6a00} /* (10, 13, 3) {real, imag} */,
  {32'h3fa261c0, 32'h3e4b4b2e} /* (10, 13, 2) {real, imag} */,
  {32'hc05f9a51, 32'hbdce24a0} /* (10, 13, 1) {real, imag} */,
  {32'hc01f8d68, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'hc0256d05, 32'hbdbfc158} /* (10, 12, 31) {real, imag} */,
  {32'h3f8d5cdb, 32'hbdae932e} /* (10, 12, 30) {real, imag} */,
  {32'hbd5cf89f, 32'h3b0ef940} /* (10, 12, 29) {real, imag} */,
  {32'hbe5e849e, 32'h3e31ee4f} /* (10, 12, 28) {real, imag} */,
  {32'h3dda4aea, 32'h3c88a16c} /* (10, 12, 27) {real, imag} */,
  {32'h3cf8608d, 32'h3c5dfac4} /* (10, 12, 26) {real, imag} */,
  {32'hbd6eeacd, 32'h3bac8754} /* (10, 12, 25) {real, imag} */,
  {32'h3dac03e2, 32'hbd096e61} /* (10, 12, 24) {real, imag} */,
  {32'hbd28b8fc, 32'hbd09795e} /* (10, 12, 23) {real, imag} */,
  {32'h3d839d7e, 32'hbdae3f7a} /* (10, 12, 22) {real, imag} */,
  {32'hbd87331f, 32'hbde1844d} /* (10, 12, 21) {real, imag} */,
  {32'h3c0520f6, 32'h3da63b44} /* (10, 12, 20) {real, imag} */,
  {32'h3cadf23a, 32'hbc1a4b8c} /* (10, 12, 19) {real, imag} */,
  {32'hbbd87cd0, 32'hbcfbb70a} /* (10, 12, 18) {real, imag} */,
  {32'hbc06c782, 32'hbd5c3f7e} /* (10, 12, 17) {real, imag} */,
  {32'hbceedd5d, 32'h00000000} /* (10, 12, 16) {real, imag} */,
  {32'hbc06c782, 32'h3d5c3f7e} /* (10, 12, 15) {real, imag} */,
  {32'hbbd87cd0, 32'h3cfbb70a} /* (10, 12, 14) {real, imag} */,
  {32'h3cadf23a, 32'h3c1a4b8c} /* (10, 12, 13) {real, imag} */,
  {32'h3c0520f6, 32'hbda63b44} /* (10, 12, 12) {real, imag} */,
  {32'hbd87331f, 32'h3de1844d} /* (10, 12, 11) {real, imag} */,
  {32'h3d839d7e, 32'h3dae3f7a} /* (10, 12, 10) {real, imag} */,
  {32'hbd28b8fc, 32'h3d09795e} /* (10, 12, 9) {real, imag} */,
  {32'h3dac03e2, 32'h3d096e61} /* (10, 12, 8) {real, imag} */,
  {32'hbd6eeacd, 32'hbbac8754} /* (10, 12, 7) {real, imag} */,
  {32'h3cf8608d, 32'hbc5dfac4} /* (10, 12, 6) {real, imag} */,
  {32'h3dda4aea, 32'hbc88a16c} /* (10, 12, 5) {real, imag} */,
  {32'hbe5e849e, 32'hbe31ee4f} /* (10, 12, 4) {real, imag} */,
  {32'hbd5cf89f, 32'hbb0ef940} /* (10, 12, 3) {real, imag} */,
  {32'h3f8d5cdb, 32'h3dae932e} /* (10, 12, 2) {real, imag} */,
  {32'hc0256d05, 32'h3dbfc158} /* (10, 12, 1) {real, imag} */,
  {32'hbfd85a0d, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hbfb4c768, 32'hbe8be97f} /* (10, 11, 31) {real, imag} */,
  {32'h3f1ce07a, 32'hbc397220} /* (10, 11, 30) {real, imag} */,
  {32'hbd65e3e9, 32'hbd84fa76} /* (10, 11, 29) {real, imag} */,
  {32'hbd09f2d3, 32'hbcfd806c} /* (10, 11, 28) {real, imag} */,
  {32'h3d52398e, 32'hbdbc2ac7} /* (10, 11, 27) {real, imag} */,
  {32'hbd0eabab, 32'hbd24f818} /* (10, 11, 26) {real, imag} */,
  {32'h3c23791c, 32'h3d5a1184} /* (10, 11, 25) {real, imag} */,
  {32'h3d2e737c, 32'hbd753eb6} /* (10, 11, 24) {real, imag} */,
  {32'h3c1ebfb0, 32'h3e0c30e2} /* (10, 11, 23) {real, imag} */,
  {32'hbc8d1975, 32'hbc18e063} /* (10, 11, 22) {real, imag} */,
  {32'h3929b100, 32'h3d02c0ed} /* (10, 11, 21) {real, imag} */,
  {32'h3d9445b5, 32'h3cec415a} /* (10, 11, 20) {real, imag} */,
  {32'h3b4acc10, 32'h3cd5d1b2} /* (10, 11, 19) {real, imag} */,
  {32'h3d4364d8, 32'hbc97fe9e} /* (10, 11, 18) {real, imag} */,
  {32'hbcbf1eb5, 32'h3d57a0b7} /* (10, 11, 17) {real, imag} */,
  {32'hbd332e84, 32'h00000000} /* (10, 11, 16) {real, imag} */,
  {32'hbcbf1eb5, 32'hbd57a0b7} /* (10, 11, 15) {real, imag} */,
  {32'h3d4364d8, 32'h3c97fe9e} /* (10, 11, 14) {real, imag} */,
  {32'h3b4acc10, 32'hbcd5d1b2} /* (10, 11, 13) {real, imag} */,
  {32'h3d9445b5, 32'hbcec415a} /* (10, 11, 12) {real, imag} */,
  {32'h3929b100, 32'hbd02c0ed} /* (10, 11, 11) {real, imag} */,
  {32'hbc8d1975, 32'h3c18e063} /* (10, 11, 10) {real, imag} */,
  {32'h3c1ebfb0, 32'hbe0c30e2} /* (10, 11, 9) {real, imag} */,
  {32'h3d2e737c, 32'h3d753eb6} /* (10, 11, 8) {real, imag} */,
  {32'h3c23791c, 32'hbd5a1184} /* (10, 11, 7) {real, imag} */,
  {32'hbd0eabab, 32'h3d24f818} /* (10, 11, 6) {real, imag} */,
  {32'h3d52398e, 32'h3dbc2ac7} /* (10, 11, 5) {real, imag} */,
  {32'hbd09f2d3, 32'h3cfd806c} /* (10, 11, 4) {real, imag} */,
  {32'hbd65e3e9, 32'h3d84fa76} /* (10, 11, 3) {real, imag} */,
  {32'h3f1ce07a, 32'h3c397220} /* (10, 11, 2) {real, imag} */,
  {32'hbfb4c768, 32'h3e8be97f} /* (10, 11, 1) {real, imag} */,
  {32'hbe22a4a0, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h3f061147, 32'hbf24e7ae} /* (10, 10, 31) {real, imag} */,
  {32'hbe9454a3, 32'h3e951d3a} /* (10, 10, 30) {real, imag} */,
  {32'hbe17cf4e, 32'hbdc3ab78} /* (10, 10, 29) {real, imag} */,
  {32'h3accbd80, 32'hbe83277e} /* (10, 10, 28) {real, imag} */,
  {32'hbcc828b0, 32'hbd20d0bc} /* (10, 10, 27) {real, imag} */,
  {32'h3ccf39c8, 32'hbc22eec0} /* (10, 10, 26) {real, imag} */,
  {32'hbd1416e2, 32'h3c6307d7} /* (10, 10, 25) {real, imag} */,
  {32'hbd06d488, 32'h3e066298} /* (10, 10, 24) {real, imag} */,
  {32'h3d7fd6d4, 32'h3cdf2f5a} /* (10, 10, 23) {real, imag} */,
  {32'h3c4ed701, 32'h3e1fac9c} /* (10, 10, 22) {real, imag} */,
  {32'h3dbd648a, 32'h3cd7fd28} /* (10, 10, 21) {real, imag} */,
  {32'hbd509e0c, 32'hbdc4da3b} /* (10, 10, 20) {real, imag} */,
  {32'hbd016c9b, 32'hbcd2531c} /* (10, 10, 19) {real, imag} */,
  {32'h3c5df984, 32'hbd077a34} /* (10, 10, 18) {real, imag} */,
  {32'h3cc75bd9, 32'h3c35b2f0} /* (10, 10, 17) {real, imag} */,
  {32'hbce0b60a, 32'h00000000} /* (10, 10, 16) {real, imag} */,
  {32'h3cc75bd9, 32'hbc35b2f0} /* (10, 10, 15) {real, imag} */,
  {32'h3c5df984, 32'h3d077a34} /* (10, 10, 14) {real, imag} */,
  {32'hbd016c9b, 32'h3cd2531c} /* (10, 10, 13) {real, imag} */,
  {32'hbd509e0c, 32'h3dc4da3b} /* (10, 10, 12) {real, imag} */,
  {32'h3dbd648a, 32'hbcd7fd28} /* (10, 10, 11) {real, imag} */,
  {32'h3c4ed701, 32'hbe1fac9c} /* (10, 10, 10) {real, imag} */,
  {32'h3d7fd6d4, 32'hbcdf2f5a} /* (10, 10, 9) {real, imag} */,
  {32'hbd06d488, 32'hbe066298} /* (10, 10, 8) {real, imag} */,
  {32'hbd1416e2, 32'hbc6307d7} /* (10, 10, 7) {real, imag} */,
  {32'h3ccf39c8, 32'h3c22eec0} /* (10, 10, 6) {real, imag} */,
  {32'hbcc828b0, 32'h3d20d0bc} /* (10, 10, 5) {real, imag} */,
  {32'h3accbd80, 32'h3e83277e} /* (10, 10, 4) {real, imag} */,
  {32'hbe17cf4e, 32'h3dc3ab78} /* (10, 10, 3) {real, imag} */,
  {32'hbe9454a3, 32'hbe951d3a} /* (10, 10, 2) {real, imag} */,
  {32'h3f061147, 32'h3f24e7ae} /* (10, 10, 1) {real, imag} */,
  {32'h3fb4a774, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h3ffe3130, 32'hbf85581f} /* (10, 9, 31) {real, imag} */,
  {32'hbf62e471, 32'h3ea7fb88} /* (10, 9, 30) {real, imag} */,
  {32'hbdc04645, 32'hbd793c36} /* (10, 9, 29) {real, imag} */,
  {32'hbd0311b8, 32'hbe329541} /* (10, 9, 28) {real, imag} */,
  {32'hbdf62e7a, 32'h3e3d2cc1} /* (10, 9, 27) {real, imag} */,
  {32'hbdbbc70a, 32'h3d402047} /* (10, 9, 26) {real, imag} */,
  {32'h3db196c3, 32'hbdd1e515} /* (10, 9, 25) {real, imag} */,
  {32'h3d463d7a, 32'h3d91b4aa} /* (10, 9, 24) {real, imag} */,
  {32'h3d97365e, 32'hbe28969b} /* (10, 9, 23) {real, imag} */,
  {32'h3ce5c993, 32'hbc69aecc} /* (10, 9, 22) {real, imag} */,
  {32'h3c783d5a, 32'hbd16e31a} /* (10, 9, 21) {real, imag} */,
  {32'hbda78064, 32'h3d454298} /* (10, 9, 20) {real, imag} */,
  {32'h3d148a02, 32'h3d0df79a} /* (10, 9, 19) {real, imag} */,
  {32'hbdb2be5a, 32'h3d0506c9} /* (10, 9, 18) {real, imag} */,
  {32'hbd27ea22, 32'h3db40e0c} /* (10, 9, 17) {real, imag} */,
  {32'hbc7f2fe8, 32'h00000000} /* (10, 9, 16) {real, imag} */,
  {32'hbd27ea22, 32'hbdb40e0c} /* (10, 9, 15) {real, imag} */,
  {32'hbdb2be5a, 32'hbd0506c9} /* (10, 9, 14) {real, imag} */,
  {32'h3d148a02, 32'hbd0df79a} /* (10, 9, 13) {real, imag} */,
  {32'hbda78064, 32'hbd454298} /* (10, 9, 12) {real, imag} */,
  {32'h3c783d5a, 32'h3d16e31a} /* (10, 9, 11) {real, imag} */,
  {32'h3ce5c993, 32'h3c69aecc} /* (10, 9, 10) {real, imag} */,
  {32'h3d97365e, 32'h3e28969b} /* (10, 9, 9) {real, imag} */,
  {32'h3d463d7a, 32'hbd91b4aa} /* (10, 9, 8) {real, imag} */,
  {32'h3db196c3, 32'h3dd1e515} /* (10, 9, 7) {real, imag} */,
  {32'hbdbbc70a, 32'hbd402047} /* (10, 9, 6) {real, imag} */,
  {32'hbdf62e7a, 32'hbe3d2cc1} /* (10, 9, 5) {real, imag} */,
  {32'hbd0311b8, 32'h3e329541} /* (10, 9, 4) {real, imag} */,
  {32'hbdc04645, 32'h3d793c36} /* (10, 9, 3) {real, imag} */,
  {32'hbf62e471, 32'hbea7fb88} /* (10, 9, 2) {real, imag} */,
  {32'h3ffe3130, 32'h3f85581f} /* (10, 9, 1) {real, imag} */,
  {32'h4029b276, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'h4036dd56, 32'hbfb1cb86} /* (10, 8, 31) {real, imag} */,
  {32'hbf8c4af5, 32'h3f15bcd2} /* (10, 8, 30) {real, imag} */,
  {32'hbe290e9c, 32'hbd390db5} /* (10, 8, 29) {real, imag} */,
  {32'h3dcc379a, 32'hbd80377a} /* (10, 8, 28) {real, imag} */,
  {32'hbdbc857c, 32'h3e98080c} /* (10, 8, 27) {real, imag} */,
  {32'hbd193eeb, 32'h3d43c8a8} /* (10, 8, 26) {real, imag} */,
  {32'h3d6ac400, 32'hbd35ca8c} /* (10, 8, 25) {real, imag} */,
  {32'hbc1fbbb8, 32'h3d34e6ea} /* (10, 8, 24) {real, imag} */,
  {32'hbdb92752, 32'h3c811b65} /* (10, 8, 23) {real, imag} */,
  {32'h3dad48fc, 32'h3cd59ecf} /* (10, 8, 22) {real, imag} */,
  {32'h3d672e87, 32'h3de3966e} /* (10, 8, 21) {real, imag} */,
  {32'hbd3dab82, 32'hbabe80c0} /* (10, 8, 20) {real, imag} */,
  {32'h3d691df2, 32'hbdc15522} /* (10, 8, 19) {real, imag} */,
  {32'h3d865188, 32'hbd6525cb} /* (10, 8, 18) {real, imag} */,
  {32'hbb3caff0, 32'hbcff548c} /* (10, 8, 17) {real, imag} */,
  {32'hbd32ea2a, 32'h00000000} /* (10, 8, 16) {real, imag} */,
  {32'hbb3caff0, 32'h3cff548c} /* (10, 8, 15) {real, imag} */,
  {32'h3d865188, 32'h3d6525cb} /* (10, 8, 14) {real, imag} */,
  {32'h3d691df2, 32'h3dc15522} /* (10, 8, 13) {real, imag} */,
  {32'hbd3dab82, 32'h3abe80c0} /* (10, 8, 12) {real, imag} */,
  {32'h3d672e87, 32'hbde3966e} /* (10, 8, 11) {real, imag} */,
  {32'h3dad48fc, 32'hbcd59ecf} /* (10, 8, 10) {real, imag} */,
  {32'hbdb92752, 32'hbc811b65} /* (10, 8, 9) {real, imag} */,
  {32'hbc1fbbb8, 32'hbd34e6ea} /* (10, 8, 8) {real, imag} */,
  {32'h3d6ac400, 32'h3d35ca8c} /* (10, 8, 7) {real, imag} */,
  {32'hbd193eeb, 32'hbd43c8a8} /* (10, 8, 6) {real, imag} */,
  {32'hbdbc857c, 32'hbe98080c} /* (10, 8, 5) {real, imag} */,
  {32'h3dcc379a, 32'h3d80377a} /* (10, 8, 4) {real, imag} */,
  {32'hbe290e9c, 32'h3d390db5} /* (10, 8, 3) {real, imag} */,
  {32'hbf8c4af5, 32'hbf15bcd2} /* (10, 8, 2) {real, imag} */,
  {32'h4036dd56, 32'h3fb1cb86} /* (10, 8, 1) {real, imag} */,
  {32'h40673684, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h405c8472, 32'hbfece771} /* (10, 7, 31) {real, imag} */,
  {32'hbf8a94ce, 32'h3f53c128} /* (10, 7, 30) {real, imag} */,
  {32'hbdffcb12, 32'hbda966fe} /* (10, 7, 29) {real, imag} */,
  {32'h3d15c80c, 32'hbe0d24b1} /* (10, 7, 28) {real, imag} */,
  {32'hbddac2a0, 32'h3e541cef} /* (10, 7, 27) {real, imag} */,
  {32'hbdced70e, 32'h3db7423d} /* (10, 7, 26) {real, imag} */,
  {32'hbbb63acc, 32'hbd153db0} /* (10, 7, 25) {real, imag} */,
  {32'hbcdbd001, 32'hbc49ed94} /* (10, 7, 24) {real, imag} */,
  {32'h3d52c1ab, 32'h3ca6fa82} /* (10, 7, 23) {real, imag} */,
  {32'h3e085b3e, 32'h3de2db70} /* (10, 7, 22) {real, imag} */,
  {32'hbce0fefd, 32'h3d4c70b2} /* (10, 7, 21) {real, imag} */,
  {32'h3cc3ccbc, 32'h3c0227a6} /* (10, 7, 20) {real, imag} */,
  {32'h3b384a1c, 32'hbd35efc6} /* (10, 7, 19) {real, imag} */,
  {32'hbe0c1a1c, 32'h3a96c6a0} /* (10, 7, 18) {real, imag} */,
  {32'hbd768931, 32'hbc9c0be8} /* (10, 7, 17) {real, imag} */,
  {32'hbdc5834b, 32'h00000000} /* (10, 7, 16) {real, imag} */,
  {32'hbd768931, 32'h3c9c0be8} /* (10, 7, 15) {real, imag} */,
  {32'hbe0c1a1c, 32'hba96c6a0} /* (10, 7, 14) {real, imag} */,
  {32'h3b384a1c, 32'h3d35efc6} /* (10, 7, 13) {real, imag} */,
  {32'h3cc3ccbc, 32'hbc0227a6} /* (10, 7, 12) {real, imag} */,
  {32'hbce0fefd, 32'hbd4c70b2} /* (10, 7, 11) {real, imag} */,
  {32'h3e085b3e, 32'hbde2db70} /* (10, 7, 10) {real, imag} */,
  {32'h3d52c1ab, 32'hbca6fa82} /* (10, 7, 9) {real, imag} */,
  {32'hbcdbd001, 32'h3c49ed94} /* (10, 7, 8) {real, imag} */,
  {32'hbbb63acc, 32'h3d153db0} /* (10, 7, 7) {real, imag} */,
  {32'hbdced70e, 32'hbdb7423d} /* (10, 7, 6) {real, imag} */,
  {32'hbddac2a0, 32'hbe541cef} /* (10, 7, 5) {real, imag} */,
  {32'h3d15c80c, 32'h3e0d24b1} /* (10, 7, 4) {real, imag} */,
  {32'hbdffcb12, 32'h3da966fe} /* (10, 7, 3) {real, imag} */,
  {32'hbf8a94ce, 32'hbf53c128} /* (10, 7, 2) {real, imag} */,
  {32'h405c8472, 32'h3fece771} /* (10, 7, 1) {real, imag} */,
  {32'h408d9ada, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h4067af3a, 32'hc01b0e78} /* (10, 6, 31) {real, imag} */,
  {32'hbf5349f4, 32'h3f813d6b} /* (10, 6, 30) {real, imag} */,
  {32'hbcdbe2e5, 32'h3d12284d} /* (10, 6, 29) {real, imag} */,
  {32'hbc9b5938, 32'h3d0cf8c4} /* (10, 6, 28) {real, imag} */,
  {32'hbdd0c6c1, 32'h3ddb88be} /* (10, 6, 27) {real, imag} */,
  {32'h3d5478e4, 32'hbb9e8d98} /* (10, 6, 26) {real, imag} */,
  {32'h3d3d75ff, 32'hbba67198} /* (10, 6, 25) {real, imag} */,
  {32'hbc1c7490, 32'hbb85c8d0} /* (10, 6, 24) {real, imag} */,
  {32'h3d875360, 32'hbdab8772} /* (10, 6, 23) {real, imag} */,
  {32'h3d06aabf, 32'h3ad6f9c0} /* (10, 6, 22) {real, imag} */,
  {32'hbcbb0426, 32'h3d94449c} /* (10, 6, 21) {real, imag} */,
  {32'hbb9acab0, 32'hbd12c77a} /* (10, 6, 20) {real, imag} */,
  {32'hbb50a8f0, 32'h3bef1fa0} /* (10, 6, 19) {real, imag} */,
  {32'hbdac0f00, 32'h3d8d2c27} /* (10, 6, 18) {real, imag} */,
  {32'h3c92b702, 32'h3c6e799f} /* (10, 6, 17) {real, imag} */,
  {32'hbd699bc0, 32'h00000000} /* (10, 6, 16) {real, imag} */,
  {32'h3c92b702, 32'hbc6e799f} /* (10, 6, 15) {real, imag} */,
  {32'hbdac0f00, 32'hbd8d2c27} /* (10, 6, 14) {real, imag} */,
  {32'hbb50a8f0, 32'hbbef1fa0} /* (10, 6, 13) {real, imag} */,
  {32'hbb9acab0, 32'h3d12c77a} /* (10, 6, 12) {real, imag} */,
  {32'hbcbb0426, 32'hbd94449c} /* (10, 6, 11) {real, imag} */,
  {32'h3d06aabf, 32'hbad6f9c0} /* (10, 6, 10) {real, imag} */,
  {32'h3d875360, 32'h3dab8772} /* (10, 6, 9) {real, imag} */,
  {32'hbc1c7490, 32'h3b85c8d0} /* (10, 6, 8) {real, imag} */,
  {32'h3d3d75ff, 32'h3ba67198} /* (10, 6, 7) {real, imag} */,
  {32'h3d5478e4, 32'h3b9e8d98} /* (10, 6, 6) {real, imag} */,
  {32'hbdd0c6c1, 32'hbddb88be} /* (10, 6, 5) {real, imag} */,
  {32'hbc9b5938, 32'hbd0cf8c4} /* (10, 6, 4) {real, imag} */,
  {32'hbcdbe2e5, 32'hbd12284d} /* (10, 6, 3) {real, imag} */,
  {32'hbf5349f4, 32'hbf813d6b} /* (10, 6, 2) {real, imag} */,
  {32'h4067af3a, 32'h401b0e78} /* (10, 6, 1) {real, imag} */,
  {32'h40a09f19, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'h40599ed3, 32'hc04b7a08} /* (10, 5, 31) {real, imag} */,
  {32'hbeded632, 32'h3f94388f} /* (10, 5, 30) {real, imag} */,
  {32'hbdfc3d0c, 32'hbc85c088} /* (10, 5, 29) {real, imag} */,
  {32'hbabd8aa0, 32'h3e5883b0} /* (10, 5, 28) {real, imag} */,
  {32'hbdf663c9, 32'h3e5fa416} /* (10, 5, 27) {real, imag} */,
  {32'h3d4ae169, 32'hbcd601c7} /* (10, 5, 26) {real, imag} */,
  {32'h3ca16208, 32'hbce17894} /* (10, 5, 25) {real, imag} */,
  {32'hbda21ae4, 32'h3e178d3a} /* (10, 5, 24) {real, imag} */,
  {32'hbdcc7c32, 32'hbcfb253a} /* (10, 5, 23) {real, imag} */,
  {32'h3c81c9e9, 32'h3db23cb6} /* (10, 5, 22) {real, imag} */,
  {32'hbdbb0962, 32'hbc5cfefc} /* (10, 5, 21) {real, imag} */,
  {32'hbc833020, 32'hbd00c51d} /* (10, 5, 20) {real, imag} */,
  {32'h3d29200f, 32'h3c928c12} /* (10, 5, 19) {real, imag} */,
  {32'h3d31e00e, 32'h3c62b9c4} /* (10, 5, 18) {real, imag} */,
  {32'hbc31e263, 32'hbda52c1c} /* (10, 5, 17) {real, imag} */,
  {32'hbd76b446, 32'h00000000} /* (10, 5, 16) {real, imag} */,
  {32'hbc31e263, 32'h3da52c1c} /* (10, 5, 15) {real, imag} */,
  {32'h3d31e00e, 32'hbc62b9c4} /* (10, 5, 14) {real, imag} */,
  {32'h3d29200f, 32'hbc928c12} /* (10, 5, 13) {real, imag} */,
  {32'hbc833020, 32'h3d00c51d} /* (10, 5, 12) {real, imag} */,
  {32'hbdbb0962, 32'h3c5cfefc} /* (10, 5, 11) {real, imag} */,
  {32'h3c81c9e9, 32'hbdb23cb6} /* (10, 5, 10) {real, imag} */,
  {32'hbdcc7c32, 32'h3cfb253a} /* (10, 5, 9) {real, imag} */,
  {32'hbda21ae4, 32'hbe178d3a} /* (10, 5, 8) {real, imag} */,
  {32'h3ca16208, 32'h3ce17894} /* (10, 5, 7) {real, imag} */,
  {32'h3d4ae169, 32'h3cd601c7} /* (10, 5, 6) {real, imag} */,
  {32'hbdf663c9, 32'hbe5fa416} /* (10, 5, 5) {real, imag} */,
  {32'hbabd8aa0, 32'hbe5883b0} /* (10, 5, 4) {real, imag} */,
  {32'hbdfc3d0c, 32'h3c85c088} /* (10, 5, 3) {real, imag} */,
  {32'hbeded632, 32'hbf94388f} /* (10, 5, 2) {real, imag} */,
  {32'h40599ed3, 32'h404b7a08} /* (10, 5, 1) {real, imag} */,
  {32'h40adf68c, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h40533099, 32'hc06a8f63} /* (10, 4, 31) {real, imag} */,
  {32'hbc004e80, 32'h3f938523} /* (10, 4, 30) {real, imag} */,
  {32'hbdd5bd80, 32'h3b884890} /* (10, 4, 29) {real, imag} */,
  {32'hbda4cf24, 32'h3e7ab093} /* (10, 4, 28) {real, imag} */,
  {32'hbde5032a, 32'h3dc61b3d} /* (10, 4, 27) {real, imag} */,
  {32'h3d6a5648, 32'h3d59dfd9} /* (10, 4, 26) {real, imag} */,
  {32'h3d4aca35, 32'hbdb64626} /* (10, 4, 25) {real, imag} */,
  {32'hbda7c35f, 32'h3e4902c2} /* (10, 4, 24) {real, imag} */,
  {32'hbc7cf468, 32'hbda8346c} /* (10, 4, 23) {real, imag} */,
  {32'h39c10420, 32'h3dc715f7} /* (10, 4, 22) {real, imag} */,
  {32'hbcea7031, 32'hbd34f119} /* (10, 4, 21) {real, imag} */,
  {32'hbc869b3e, 32'h3d9ad18a} /* (10, 4, 20) {real, imag} */,
  {32'hb99b9040, 32'hbd0cfd50} /* (10, 4, 19) {real, imag} */,
  {32'h3ce7ef98, 32'h3d2c3576} /* (10, 4, 18) {real, imag} */,
  {32'hbd3302ae, 32'h3be504a8} /* (10, 4, 17) {real, imag} */,
  {32'h3c4eaec4, 32'h00000000} /* (10, 4, 16) {real, imag} */,
  {32'hbd3302ae, 32'hbbe504a8} /* (10, 4, 15) {real, imag} */,
  {32'h3ce7ef98, 32'hbd2c3576} /* (10, 4, 14) {real, imag} */,
  {32'hb99b9040, 32'h3d0cfd50} /* (10, 4, 13) {real, imag} */,
  {32'hbc869b3e, 32'hbd9ad18a} /* (10, 4, 12) {real, imag} */,
  {32'hbcea7031, 32'h3d34f119} /* (10, 4, 11) {real, imag} */,
  {32'h39c10420, 32'hbdc715f7} /* (10, 4, 10) {real, imag} */,
  {32'hbc7cf468, 32'h3da8346c} /* (10, 4, 9) {real, imag} */,
  {32'hbda7c35f, 32'hbe4902c2} /* (10, 4, 8) {real, imag} */,
  {32'h3d4aca35, 32'h3db64626} /* (10, 4, 7) {real, imag} */,
  {32'h3d6a5648, 32'hbd59dfd9} /* (10, 4, 6) {real, imag} */,
  {32'hbde5032a, 32'hbdc61b3d} /* (10, 4, 5) {real, imag} */,
  {32'hbda4cf24, 32'hbe7ab093} /* (10, 4, 4) {real, imag} */,
  {32'hbdd5bd80, 32'hbb884890} /* (10, 4, 3) {real, imag} */,
  {32'hbc004e80, 32'hbf938523} /* (10, 4, 2) {real, imag} */,
  {32'h40533099, 32'h406a8f63} /* (10, 4, 1) {real, imag} */,
  {32'h40b6f506, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'h4052a8e4, 32'hc07ff964} /* (10, 3, 31) {real, imag} */,
  {32'h3e6e834c, 32'h3f9cea44} /* (10, 3, 30) {real, imag} */,
  {32'hbc6135b0, 32'h3e02421e} /* (10, 3, 29) {real, imag} */,
  {32'hbe2e6d5c, 32'h3e92d0dc} /* (10, 3, 28) {real, imag} */,
  {32'hbe3d53f2, 32'hbd853614} /* (10, 3, 27) {real, imag} */,
  {32'hbd84b8f0, 32'h3d59c730} /* (10, 3, 26) {real, imag} */,
  {32'h3c0ff9f9, 32'h3d2f6c11} /* (10, 3, 25) {real, imag} */,
  {32'h3df0ffc6, 32'h3e14dfe1} /* (10, 3, 24) {real, imag} */,
  {32'hbcb68718, 32'hbe0773f5} /* (10, 3, 23) {real, imag} */,
  {32'hbd11807f, 32'hbbc6fbe0} /* (10, 3, 22) {real, imag} */,
  {32'hbb6dda58, 32'h3da95434} /* (10, 3, 21) {real, imag} */,
  {32'hbd574df8, 32'h3a401df0} /* (10, 3, 20) {real, imag} */,
  {32'hbd2f3fde, 32'hbdaf7991} /* (10, 3, 19) {real, imag} */,
  {32'hbc7d2a86, 32'h3da1a2e0} /* (10, 3, 18) {real, imag} */,
  {32'h3db4e5bc, 32'h3c66073c} /* (10, 3, 17) {real, imag} */,
  {32'h3e13a2dc, 32'h00000000} /* (10, 3, 16) {real, imag} */,
  {32'h3db4e5bc, 32'hbc66073c} /* (10, 3, 15) {real, imag} */,
  {32'hbc7d2a86, 32'hbda1a2e0} /* (10, 3, 14) {real, imag} */,
  {32'hbd2f3fde, 32'h3daf7991} /* (10, 3, 13) {real, imag} */,
  {32'hbd574df8, 32'hba401df0} /* (10, 3, 12) {real, imag} */,
  {32'hbb6dda58, 32'hbda95434} /* (10, 3, 11) {real, imag} */,
  {32'hbd11807f, 32'h3bc6fbe0} /* (10, 3, 10) {real, imag} */,
  {32'hbcb68718, 32'h3e0773f5} /* (10, 3, 9) {real, imag} */,
  {32'h3df0ffc6, 32'hbe14dfe1} /* (10, 3, 8) {real, imag} */,
  {32'h3c0ff9f9, 32'hbd2f6c11} /* (10, 3, 7) {real, imag} */,
  {32'hbd84b8f0, 32'hbd59c730} /* (10, 3, 6) {real, imag} */,
  {32'hbe3d53f2, 32'h3d853614} /* (10, 3, 5) {real, imag} */,
  {32'hbe2e6d5c, 32'hbe92d0dc} /* (10, 3, 4) {real, imag} */,
  {32'hbc6135b0, 32'hbe02421e} /* (10, 3, 3) {real, imag} */,
  {32'h3e6e834c, 32'hbf9cea44} /* (10, 3, 2) {real, imag} */,
  {32'h4052a8e4, 32'h407ff964} /* (10, 3, 1) {real, imag} */,
  {32'h40b7e3a4, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'h405171fe, 32'hc0814cc4} /* (10, 2, 31) {real, imag} */,
  {32'h3e8c4717, 32'h3f995146} /* (10, 2, 30) {real, imag} */,
  {32'hbdf60ed9, 32'h3b8cffd0} /* (10, 2, 29) {real, imag} */,
  {32'hbe273098, 32'h3eb4af38} /* (10, 2, 28) {real, imag} */,
  {32'hbe1053bc, 32'hbe088da5} /* (10, 2, 27) {real, imag} */,
  {32'hbd760a03, 32'h3db50860} /* (10, 2, 26) {real, imag} */,
  {32'h3cea5f7d, 32'h3bde5ba8} /* (10, 2, 25) {real, imag} */,
  {32'h3d543e7b, 32'h3dac5d5a} /* (10, 2, 24) {real, imag} */,
  {32'hbdb038e8, 32'hbd14c231} /* (10, 2, 23) {real, imag} */,
  {32'h3df871fb, 32'hbd12a883} /* (10, 2, 22) {real, imag} */,
  {32'hbc8813b4, 32'h3cc7d628} /* (10, 2, 21) {real, imag} */,
  {32'h3c8a20c8, 32'h3c8db71f} /* (10, 2, 20) {real, imag} */,
  {32'h3c70fd0f, 32'h3d4489ec} /* (10, 2, 19) {real, imag} */,
  {32'h3c7d2be8, 32'hbca3b33e} /* (10, 2, 18) {real, imag} */,
  {32'h3d51fff7, 32'hbce48b18} /* (10, 2, 17) {real, imag} */,
  {32'hbdc8eb42, 32'h00000000} /* (10, 2, 16) {real, imag} */,
  {32'h3d51fff7, 32'h3ce48b18} /* (10, 2, 15) {real, imag} */,
  {32'h3c7d2be8, 32'h3ca3b33e} /* (10, 2, 14) {real, imag} */,
  {32'h3c70fd0f, 32'hbd4489ec} /* (10, 2, 13) {real, imag} */,
  {32'h3c8a20c8, 32'hbc8db71f} /* (10, 2, 12) {real, imag} */,
  {32'hbc8813b4, 32'hbcc7d628} /* (10, 2, 11) {real, imag} */,
  {32'h3df871fb, 32'h3d12a883} /* (10, 2, 10) {real, imag} */,
  {32'hbdb038e8, 32'h3d14c231} /* (10, 2, 9) {real, imag} */,
  {32'h3d543e7b, 32'hbdac5d5a} /* (10, 2, 8) {real, imag} */,
  {32'h3cea5f7d, 32'hbbde5ba8} /* (10, 2, 7) {real, imag} */,
  {32'hbd760a03, 32'hbdb50860} /* (10, 2, 6) {real, imag} */,
  {32'hbe1053bc, 32'h3e088da5} /* (10, 2, 5) {real, imag} */,
  {32'hbe273098, 32'hbeb4af38} /* (10, 2, 4) {real, imag} */,
  {32'hbdf60ed9, 32'hbb8cffd0} /* (10, 2, 3) {real, imag} */,
  {32'h3e8c4717, 32'hbf995146} /* (10, 2, 2) {real, imag} */,
  {32'h405171fe, 32'h40814cc4} /* (10, 2, 1) {real, imag} */,
  {32'h40b1a273, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'h405cce8c, 32'hc0700414} /* (10, 1, 31) {real, imag} */,
  {32'h3d58e1b0, 32'h3f840658} /* (10, 1, 30) {real, imag} */,
  {32'hbe64d818, 32'hbe15a417} /* (10, 1, 29) {real, imag} */,
  {32'hbda1dc1b, 32'h3ebd4f8c} /* (10, 1, 28) {real, imag} */,
  {32'hbe452764, 32'hbd7d14a6} /* (10, 1, 27) {real, imag} */,
  {32'hbd957245, 32'h3d661a22} /* (10, 1, 26) {real, imag} */,
  {32'h3d00e6a7, 32'h3c1f12f8} /* (10, 1, 25) {real, imag} */,
  {32'h3d896a7f, 32'h3c8d7caa} /* (10, 1, 24) {real, imag} */,
  {32'h3c94fc92, 32'h3d403ac6} /* (10, 1, 23) {real, imag} */,
  {32'hbd96106b, 32'hbbfe4d47} /* (10, 1, 22) {real, imag} */,
  {32'h3d43964d, 32'hbcad895a} /* (10, 1, 21) {real, imag} */,
  {32'h3bf33b10, 32'h3d4cf6f5} /* (10, 1, 20) {real, imag} */,
  {32'hbd801d03, 32'hbd378c60} /* (10, 1, 19) {real, imag} */,
  {32'h3c6f8404, 32'h3c20e584} /* (10, 1, 18) {real, imag} */,
  {32'hbd14a176, 32'h3cb40798} /* (10, 1, 17) {real, imag} */,
  {32'hbbcd6ab7, 32'h00000000} /* (10, 1, 16) {real, imag} */,
  {32'hbd14a176, 32'hbcb40798} /* (10, 1, 15) {real, imag} */,
  {32'h3c6f8404, 32'hbc20e584} /* (10, 1, 14) {real, imag} */,
  {32'hbd801d03, 32'h3d378c60} /* (10, 1, 13) {real, imag} */,
  {32'h3bf33b10, 32'hbd4cf6f5} /* (10, 1, 12) {real, imag} */,
  {32'h3d43964d, 32'h3cad895a} /* (10, 1, 11) {real, imag} */,
  {32'hbd96106b, 32'h3bfe4d47} /* (10, 1, 10) {real, imag} */,
  {32'h3c94fc92, 32'hbd403ac6} /* (10, 1, 9) {real, imag} */,
  {32'h3d896a7f, 32'hbc8d7caa} /* (10, 1, 8) {real, imag} */,
  {32'h3d00e6a7, 32'hbc1f12f8} /* (10, 1, 7) {real, imag} */,
  {32'hbd957245, 32'hbd661a22} /* (10, 1, 6) {real, imag} */,
  {32'hbe452764, 32'h3d7d14a6} /* (10, 1, 5) {real, imag} */,
  {32'hbda1dc1b, 32'hbebd4f8c} /* (10, 1, 4) {real, imag} */,
  {32'hbe64d818, 32'h3e15a417} /* (10, 1, 3) {real, imag} */,
  {32'h3d58e1b0, 32'hbf840658} /* (10, 1, 2) {real, imag} */,
  {32'h405cce8c, 32'h40700414} /* (10, 1, 1) {real, imag} */,
  {32'h40b13a39, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h406692e7, 32'hc0409ce6} /* (10, 0, 31) {real, imag} */,
  {32'hbe6298f4, 32'h3f3ae223} /* (10, 0, 30) {real, imag} */,
  {32'hbe25de0a, 32'hbd4480a1} /* (10, 0, 29) {real, imag} */,
  {32'hbd5855e4, 32'h3e764c32} /* (10, 0, 28) {real, imag} */,
  {32'hbe42ec62, 32'hbcaa8060} /* (10, 0, 27) {real, imag} */,
  {32'h39855a00, 32'h3c4067d0} /* (10, 0, 26) {real, imag} */,
  {32'h3d62f2d6, 32'hbc5cc855} /* (10, 0, 25) {real, imag} */,
  {32'h3b8fe5a0, 32'hbcb21fcc} /* (10, 0, 24) {real, imag} */,
  {32'h3c873a0a, 32'hbacb3510} /* (10, 0, 23) {real, imag} */,
  {32'hbd84730e, 32'hbc39438a} /* (10, 0, 22) {real, imag} */,
  {32'h3cccd6f4, 32'h3d2358e5} /* (10, 0, 21) {real, imag} */,
  {32'hbc0c10e8, 32'hbc98a098} /* (10, 0, 20) {real, imag} */,
  {32'h3d3cc8c2, 32'hbc0df9ed} /* (10, 0, 19) {real, imag} */,
  {32'hbbef85b0, 32'h3cd3c590} /* (10, 0, 18) {real, imag} */,
  {32'hbd19ab63, 32'h3a560c00} /* (10, 0, 17) {real, imag} */,
  {32'h3c62e64c, 32'h00000000} /* (10, 0, 16) {real, imag} */,
  {32'hbd19ab63, 32'hba560c00} /* (10, 0, 15) {real, imag} */,
  {32'hbbef85b0, 32'hbcd3c590} /* (10, 0, 14) {real, imag} */,
  {32'h3d3cc8c2, 32'h3c0df9ed} /* (10, 0, 13) {real, imag} */,
  {32'hbc0c10e8, 32'h3c98a098} /* (10, 0, 12) {real, imag} */,
  {32'h3cccd6f4, 32'hbd2358e5} /* (10, 0, 11) {real, imag} */,
  {32'hbd84730e, 32'h3c39438a} /* (10, 0, 10) {real, imag} */,
  {32'h3c873a0a, 32'h3acb3510} /* (10, 0, 9) {real, imag} */,
  {32'h3b8fe5a0, 32'h3cb21fcc} /* (10, 0, 8) {real, imag} */,
  {32'h3d62f2d6, 32'h3c5cc855} /* (10, 0, 7) {real, imag} */,
  {32'h39855a00, 32'hbc4067d0} /* (10, 0, 6) {real, imag} */,
  {32'hbe42ec62, 32'h3caa8060} /* (10, 0, 5) {real, imag} */,
  {32'hbd5855e4, 32'hbe764c32} /* (10, 0, 4) {real, imag} */,
  {32'hbe25de0a, 32'h3d4480a1} /* (10, 0, 3) {real, imag} */,
  {32'hbe6298f4, 32'hbf3ae223} /* (10, 0, 2) {real, imag} */,
  {32'h406692e7, 32'h40409ce6} /* (10, 0, 1) {real, imag} */,
  {32'h40b1008c, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h407763e7, 32'hc0116a1f} /* (9, 31, 31) {real, imag} */,
  {32'hbf55096a, 32'h3f36d006} /* (9, 31, 30) {real, imag} */,
  {32'hbd366328, 32'hbdc3517e} /* (9, 31, 29) {real, imag} */,
  {32'h3dff1a90, 32'h3dcc7c04} /* (9, 31, 28) {real, imag} */,
  {32'hbe2f353b, 32'hbc02c3c8} /* (9, 31, 27) {real, imag} */,
  {32'h3d0c2070, 32'h3d077a6c} /* (9, 31, 26) {real, imag} */,
  {32'hbd086744, 32'h3c78b916} /* (9, 31, 25) {real, imag} */,
  {32'hbd25c60c, 32'hbad358c0} /* (9, 31, 24) {real, imag} */,
  {32'h3d8b0064, 32'h3cae2c48} /* (9, 31, 23) {real, imag} */,
  {32'hbc6e2b1c, 32'h3b8e2ab6} /* (9, 31, 22) {real, imag} */,
  {32'h3ce1e30a, 32'hbc9bc81e} /* (9, 31, 21) {real, imag} */,
  {32'h3d74afa6, 32'hbd34cbe5} /* (9, 31, 20) {real, imag} */,
  {32'h3c3faac0, 32'hbcb9bc2e} /* (9, 31, 19) {real, imag} */,
  {32'hbd4dac79, 32'hbc4e3608} /* (9, 31, 18) {real, imag} */,
  {32'h3abb02d4, 32'h3bbd23f0} /* (9, 31, 17) {real, imag} */,
  {32'hbbc1b1bc, 32'h00000000} /* (9, 31, 16) {real, imag} */,
  {32'h3abb02d4, 32'hbbbd23f0} /* (9, 31, 15) {real, imag} */,
  {32'hbd4dac79, 32'h3c4e3608} /* (9, 31, 14) {real, imag} */,
  {32'h3c3faac0, 32'h3cb9bc2e} /* (9, 31, 13) {real, imag} */,
  {32'h3d74afa6, 32'h3d34cbe5} /* (9, 31, 12) {real, imag} */,
  {32'h3ce1e30a, 32'h3c9bc81e} /* (9, 31, 11) {real, imag} */,
  {32'hbc6e2b1c, 32'hbb8e2ab6} /* (9, 31, 10) {real, imag} */,
  {32'h3d8b0064, 32'hbcae2c48} /* (9, 31, 9) {real, imag} */,
  {32'hbd25c60c, 32'h3ad358c0} /* (9, 31, 8) {real, imag} */,
  {32'hbd086744, 32'hbc78b916} /* (9, 31, 7) {real, imag} */,
  {32'h3d0c2070, 32'hbd077a6c} /* (9, 31, 6) {real, imag} */,
  {32'hbe2f353b, 32'h3c02c3c8} /* (9, 31, 5) {real, imag} */,
  {32'h3dff1a90, 32'hbdcc7c04} /* (9, 31, 4) {real, imag} */,
  {32'hbd366328, 32'h3dc3517e} /* (9, 31, 3) {real, imag} */,
  {32'hbf55096a, 32'hbf36d006} /* (9, 31, 2) {real, imag} */,
  {32'h407763e7, 32'h40116a1f} /* (9, 31, 1) {real, imag} */,
  {32'h40af322b, 32'h00000000} /* (9, 31, 0) {real, imag} */,
  {32'h408ee383, 32'hbfe757d4} /* (9, 30, 31) {real, imag} */,
  {32'hbf95d64e, 32'h3f1d7709} /* (9, 30, 30) {real, imag} */,
  {32'hbd05e090, 32'hbdb42c85} /* (9, 30, 29) {real, imag} */,
  {32'h3e19839a, 32'h3d1a30d0} /* (9, 30, 28) {real, imag} */,
  {32'hbe697fbd, 32'h3c6e3358} /* (9, 30, 27) {real, imag} */,
  {32'h3d19a3cd, 32'hbccc8213} /* (9, 30, 26) {real, imag} */,
  {32'h3d4a027e, 32'h3d7d5495} /* (9, 30, 25) {real, imag} */,
  {32'hbd2b06f6, 32'hbba3e1a0} /* (9, 30, 24) {real, imag} */,
  {32'h3de9e25b, 32'h3c11f938} /* (9, 30, 23) {real, imag} */,
  {32'h3cd2cf8c, 32'h3e018678} /* (9, 30, 22) {real, imag} */,
  {32'hbb85d998, 32'h3dc1d71a} /* (9, 30, 21) {real, imag} */,
  {32'h3e0017da, 32'hbd10619a} /* (9, 30, 20) {real, imag} */,
  {32'h3dbdac41, 32'hbdf833d2} /* (9, 30, 19) {real, imag} */,
  {32'h3c2e4dec, 32'h3cfd1200} /* (9, 30, 18) {real, imag} */,
  {32'hbca47567, 32'hbb86d428} /* (9, 30, 17) {real, imag} */,
  {32'hbc9eca90, 32'h00000000} /* (9, 30, 16) {real, imag} */,
  {32'hbca47567, 32'h3b86d428} /* (9, 30, 15) {real, imag} */,
  {32'h3c2e4dec, 32'hbcfd1200} /* (9, 30, 14) {real, imag} */,
  {32'h3dbdac41, 32'h3df833d2} /* (9, 30, 13) {real, imag} */,
  {32'h3e0017da, 32'h3d10619a} /* (9, 30, 12) {real, imag} */,
  {32'hbb85d998, 32'hbdc1d71a} /* (9, 30, 11) {real, imag} */,
  {32'h3cd2cf8c, 32'hbe018678} /* (9, 30, 10) {real, imag} */,
  {32'h3de9e25b, 32'hbc11f938} /* (9, 30, 9) {real, imag} */,
  {32'hbd2b06f6, 32'h3ba3e1a0} /* (9, 30, 8) {real, imag} */,
  {32'h3d4a027e, 32'hbd7d5495} /* (9, 30, 7) {real, imag} */,
  {32'h3d19a3cd, 32'h3ccc8213} /* (9, 30, 6) {real, imag} */,
  {32'hbe697fbd, 32'hbc6e3358} /* (9, 30, 5) {real, imag} */,
  {32'h3e19839a, 32'hbd1a30d0} /* (9, 30, 4) {real, imag} */,
  {32'hbd05e090, 32'h3db42c85} /* (9, 30, 3) {real, imag} */,
  {32'hbf95d64e, 32'hbf1d7709} /* (9, 30, 2) {real, imag} */,
  {32'h408ee383, 32'h3fe757d4} /* (9, 30, 1) {real, imag} */,
  {32'h40b45a47, 32'h00000000} /* (9, 30, 0) {real, imag} */,
  {32'h409968cd, 32'hbfc09a44} /* (9, 29, 31) {real, imag} */,
  {32'hbfadfaf9, 32'h3f1d52bc} /* (9, 29, 30) {real, imag} */,
  {32'h3d18c36a, 32'hbd88ac1f} /* (9, 29, 29) {real, imag} */,
  {32'h3d5933d7, 32'h3c0119d0} /* (9, 29, 28) {real, imag} */,
  {32'hbe4012a4, 32'hbd8ee97f} /* (9, 29, 27) {real, imag} */,
  {32'hbda88e80, 32'hbb0ac0f0} /* (9, 29, 26) {real, imag} */,
  {32'hbd7975ee, 32'hbe12c82e} /* (9, 29, 25) {real, imag} */,
  {32'hbcf2e1ea, 32'h3d102df0} /* (9, 29, 24) {real, imag} */,
  {32'h3d314df1, 32'hbd8972ca} /* (9, 29, 23) {real, imag} */,
  {32'hbd08806a, 32'h3d7c3bfc} /* (9, 29, 22) {real, imag} */,
  {32'hbd932c0e, 32'h3a861d10} /* (9, 29, 21) {real, imag} */,
  {32'hbbaf3f74, 32'h3dd91383} /* (9, 29, 20) {real, imag} */,
  {32'hbdaf8d86, 32'h3c1bedd8} /* (9, 29, 19) {real, imag} */,
  {32'hbcc43059, 32'h3cebe415} /* (9, 29, 18) {real, imag} */,
  {32'hbbc663a0, 32'hbc556086} /* (9, 29, 17) {real, imag} */,
  {32'hbc839f50, 32'h00000000} /* (9, 29, 16) {real, imag} */,
  {32'hbbc663a0, 32'h3c556086} /* (9, 29, 15) {real, imag} */,
  {32'hbcc43059, 32'hbcebe415} /* (9, 29, 14) {real, imag} */,
  {32'hbdaf8d86, 32'hbc1bedd8} /* (9, 29, 13) {real, imag} */,
  {32'hbbaf3f74, 32'hbdd91383} /* (9, 29, 12) {real, imag} */,
  {32'hbd932c0e, 32'hba861d10} /* (9, 29, 11) {real, imag} */,
  {32'hbd08806a, 32'hbd7c3bfc} /* (9, 29, 10) {real, imag} */,
  {32'h3d314df1, 32'h3d8972ca} /* (9, 29, 9) {real, imag} */,
  {32'hbcf2e1ea, 32'hbd102df0} /* (9, 29, 8) {real, imag} */,
  {32'hbd7975ee, 32'h3e12c82e} /* (9, 29, 7) {real, imag} */,
  {32'hbda88e80, 32'h3b0ac0f0} /* (9, 29, 6) {real, imag} */,
  {32'hbe4012a4, 32'h3d8ee97f} /* (9, 29, 5) {real, imag} */,
  {32'h3d5933d7, 32'hbc0119d0} /* (9, 29, 4) {real, imag} */,
  {32'h3d18c36a, 32'h3d88ac1f} /* (9, 29, 3) {real, imag} */,
  {32'hbfadfaf9, 32'hbf1d52bc} /* (9, 29, 2) {real, imag} */,
  {32'h409968cd, 32'h3fc09a44} /* (9, 29, 1) {real, imag} */,
  {32'h40b1f1cf, 32'h00000000} /* (9, 29, 0) {real, imag} */,
  {32'h40a1369f, 32'hbf8fbcb2} /* (9, 28, 31) {real, imag} */,
  {32'hbfcd74c0, 32'h3f10dcb1} /* (9, 28, 30) {real, imag} */,
  {32'h3e1f7faa, 32'h3c53508c} /* (9, 28, 29) {real, imag} */,
  {32'h3e4366e6, 32'hbda5470c} /* (9, 28, 28) {real, imag} */,
  {32'hbe81f52b, 32'hbd93200f} /* (9, 28, 27) {real, imag} */,
  {32'hbdd6e7a6, 32'hbd334e60} /* (9, 28, 26) {real, imag} */,
  {32'h3ddbbdf6, 32'hbe1c555c} /* (9, 28, 25) {real, imag} */,
  {32'hbcaee018, 32'h3cb42caa} /* (9, 28, 24) {real, imag} */,
  {32'hbdacad8a, 32'hbdd76151} /* (9, 28, 23) {real, imag} */,
  {32'h3a4d73f0, 32'h3c92bc0e} /* (9, 28, 22) {real, imag} */,
  {32'hbdacda0e, 32'h3d87ddc2} /* (9, 28, 21) {real, imag} */,
  {32'h3cb4b1d4, 32'h3d22e449} /* (9, 28, 20) {real, imag} */,
  {32'h3d92801a, 32'h3cfafbb8} /* (9, 28, 19) {real, imag} */,
  {32'hbd85bc66, 32'h3d4739f4} /* (9, 28, 18) {real, imag} */,
  {32'hbe07991f, 32'h3d444e21} /* (9, 28, 17) {real, imag} */,
  {32'h3dabfa5d, 32'h00000000} /* (9, 28, 16) {real, imag} */,
  {32'hbe07991f, 32'hbd444e21} /* (9, 28, 15) {real, imag} */,
  {32'hbd85bc66, 32'hbd4739f4} /* (9, 28, 14) {real, imag} */,
  {32'h3d92801a, 32'hbcfafbb8} /* (9, 28, 13) {real, imag} */,
  {32'h3cb4b1d4, 32'hbd22e449} /* (9, 28, 12) {real, imag} */,
  {32'hbdacda0e, 32'hbd87ddc2} /* (9, 28, 11) {real, imag} */,
  {32'h3a4d73f0, 32'hbc92bc0e} /* (9, 28, 10) {real, imag} */,
  {32'hbdacad8a, 32'h3dd76151} /* (9, 28, 9) {real, imag} */,
  {32'hbcaee018, 32'hbcb42caa} /* (9, 28, 8) {real, imag} */,
  {32'h3ddbbdf6, 32'h3e1c555c} /* (9, 28, 7) {real, imag} */,
  {32'hbdd6e7a6, 32'h3d334e60} /* (9, 28, 6) {real, imag} */,
  {32'hbe81f52b, 32'h3d93200f} /* (9, 28, 5) {real, imag} */,
  {32'h3e4366e6, 32'h3da5470c} /* (9, 28, 4) {real, imag} */,
  {32'h3e1f7faa, 32'hbc53508c} /* (9, 28, 3) {real, imag} */,
  {32'hbfcd74c0, 32'hbf10dcb1} /* (9, 28, 2) {real, imag} */,
  {32'h40a1369f, 32'h3f8fbcb2} /* (9, 28, 1) {real, imag} */,
  {32'h40b10cf8, 32'h00000000} /* (9, 28, 0) {real, imag} */,
  {32'h40a41d81, 32'hbf57b88e} /* (9, 27, 31) {real, imag} */,
  {32'hbfe03bd8, 32'h3ee6f0a2} /* (9, 27, 30) {real, imag} */,
  {32'hbe025fbf, 32'h3dc37b06} /* (9, 27, 29) {real, imag} */,
  {32'h3e9b2bf3, 32'hbd5268b0} /* (9, 27, 28) {real, imag} */,
  {32'hbd829226, 32'hbd309c5c} /* (9, 27, 27) {real, imag} */,
  {32'hbdf755c0, 32'hbbb0d660} /* (9, 27, 26) {real, imag} */,
  {32'h3d71d62b, 32'hbcb1ee84} /* (9, 27, 25) {real, imag} */,
  {32'hbdab39ea, 32'h3dbb994a} /* (9, 27, 24) {real, imag} */,
  {32'h3d9d6f93, 32'h3d2113e3} /* (9, 27, 23) {real, imag} */,
  {32'h3cbe71c6, 32'hba296020} /* (9, 27, 22) {real, imag} */,
  {32'hbd9a33bd, 32'h3c5a8c14} /* (9, 27, 21) {real, imag} */,
  {32'hbd169538, 32'h3d452436} /* (9, 27, 20) {real, imag} */,
  {32'h3dd27e9e, 32'hbce594a0} /* (9, 27, 19) {real, imag} */,
  {32'h3d7145f8, 32'h3d7d0457} /* (9, 27, 18) {real, imag} */,
  {32'hbd65baa3, 32'hbd952f57} /* (9, 27, 17) {real, imag} */,
  {32'hbdcbec3a, 32'h00000000} /* (9, 27, 16) {real, imag} */,
  {32'hbd65baa3, 32'h3d952f57} /* (9, 27, 15) {real, imag} */,
  {32'h3d7145f8, 32'hbd7d0457} /* (9, 27, 14) {real, imag} */,
  {32'h3dd27e9e, 32'h3ce594a0} /* (9, 27, 13) {real, imag} */,
  {32'hbd169538, 32'hbd452436} /* (9, 27, 12) {real, imag} */,
  {32'hbd9a33bd, 32'hbc5a8c14} /* (9, 27, 11) {real, imag} */,
  {32'h3cbe71c6, 32'h3a296020} /* (9, 27, 10) {real, imag} */,
  {32'h3d9d6f93, 32'hbd2113e3} /* (9, 27, 9) {real, imag} */,
  {32'hbdab39ea, 32'hbdbb994a} /* (9, 27, 8) {real, imag} */,
  {32'h3d71d62b, 32'h3cb1ee84} /* (9, 27, 7) {real, imag} */,
  {32'hbdf755c0, 32'h3bb0d660} /* (9, 27, 6) {real, imag} */,
  {32'hbd829226, 32'h3d309c5c} /* (9, 27, 5) {real, imag} */,
  {32'h3e9b2bf3, 32'h3d5268b0} /* (9, 27, 4) {real, imag} */,
  {32'hbe025fbf, 32'hbdc37b06} /* (9, 27, 3) {real, imag} */,
  {32'hbfe03bd8, 32'hbee6f0a2} /* (9, 27, 2) {real, imag} */,
  {32'h40a41d81, 32'h3f57b88e} /* (9, 27, 1) {real, imag} */,
  {32'h40adc4a0, 32'h00000000} /* (9, 27, 0) {real, imag} */,
  {32'h409f97e5, 32'hbf241b26} /* (9, 26, 31) {real, imag} */,
  {32'hbfdde798, 32'h3e84580c} /* (9, 26, 30) {real, imag} */,
  {32'hbd13bf30, 32'h3d950740} /* (9, 26, 29) {real, imag} */,
  {32'h3e4a411a, 32'hbd93511e} /* (9, 26, 28) {real, imag} */,
  {32'hbe2882d4, 32'h3ce880cf} /* (9, 26, 27) {real, imag} */,
  {32'hbd80cde0, 32'h3c533bf8} /* (9, 26, 26) {real, imag} */,
  {32'hbd2672aa, 32'h3bcbcde0} /* (9, 26, 25) {real, imag} */,
  {32'hbc88d24c, 32'h3e482412} /* (9, 26, 24) {real, imag} */,
  {32'h3df35db3, 32'h3b12eb84} /* (9, 26, 23) {real, imag} */,
  {32'hbd6689ba, 32'hbd3bc230} /* (9, 26, 22) {real, imag} */,
  {32'h3d826c1d, 32'h3cf7fcca} /* (9, 26, 21) {real, imag} */,
  {32'h3c18b95f, 32'hbb4f6988} /* (9, 26, 20) {real, imag} */,
  {32'hbdb3296c, 32'hbd022b14} /* (9, 26, 19) {real, imag} */,
  {32'hbd2481e2, 32'hbba5c2b0} /* (9, 26, 18) {real, imag} */,
  {32'h3cc5f9ba, 32'h3cd0e777} /* (9, 26, 17) {real, imag} */,
  {32'h3cc97b48, 32'h00000000} /* (9, 26, 16) {real, imag} */,
  {32'h3cc5f9ba, 32'hbcd0e777} /* (9, 26, 15) {real, imag} */,
  {32'hbd2481e2, 32'h3ba5c2b0} /* (9, 26, 14) {real, imag} */,
  {32'hbdb3296c, 32'h3d022b14} /* (9, 26, 13) {real, imag} */,
  {32'h3c18b95f, 32'h3b4f6988} /* (9, 26, 12) {real, imag} */,
  {32'h3d826c1d, 32'hbcf7fcca} /* (9, 26, 11) {real, imag} */,
  {32'hbd6689ba, 32'h3d3bc230} /* (9, 26, 10) {real, imag} */,
  {32'h3df35db3, 32'hbb12eb84} /* (9, 26, 9) {real, imag} */,
  {32'hbc88d24c, 32'hbe482412} /* (9, 26, 8) {real, imag} */,
  {32'hbd2672aa, 32'hbbcbcde0} /* (9, 26, 7) {real, imag} */,
  {32'hbd80cde0, 32'hbc533bf8} /* (9, 26, 6) {real, imag} */,
  {32'hbe2882d4, 32'hbce880cf} /* (9, 26, 5) {real, imag} */,
  {32'h3e4a411a, 32'h3d93511e} /* (9, 26, 4) {real, imag} */,
  {32'hbd13bf30, 32'hbd950740} /* (9, 26, 3) {real, imag} */,
  {32'hbfdde798, 32'hbe84580c} /* (9, 26, 2) {real, imag} */,
  {32'h409f97e5, 32'h3f241b26} /* (9, 26, 1) {real, imag} */,
  {32'h40a84759, 32'h00000000} /* (9, 26, 0) {real, imag} */,
  {32'h40972706, 32'hbebaa238} /* (9, 25, 31) {real, imag} */,
  {32'hbfcd72f3, 32'h3e873dee} /* (9, 25, 30) {real, imag} */,
  {32'hbdab52b6, 32'h3b8612f0} /* (9, 25, 29) {real, imag} */,
  {32'h3db33a65, 32'hbdd9be1e} /* (9, 25, 28) {real, imag} */,
  {32'hbe505bf4, 32'h3d83abfd} /* (9, 25, 27) {real, imag} */,
  {32'hbd208c60, 32'hbd278e86} /* (9, 25, 26) {real, imag} */,
  {32'h3d82e64c, 32'h3dd8c89c} /* (9, 25, 25) {real, imag} */,
  {32'h3d711a3e, 32'h3e0ad227} /* (9, 25, 24) {real, imag} */,
  {32'h3a449660, 32'hbc6fb2ee} /* (9, 25, 23) {real, imag} */,
  {32'h3d63798f, 32'hbe252f08} /* (9, 25, 22) {real, imag} */,
  {32'h3cff5294, 32'h3d750308} /* (9, 25, 21) {real, imag} */,
  {32'hbd933757, 32'h3cc8e554} /* (9, 25, 20) {real, imag} */,
  {32'hbda3e279, 32'hbc2626ad} /* (9, 25, 19) {real, imag} */,
  {32'h3cc00fe2, 32'h3e0214ae} /* (9, 25, 18) {real, imag} */,
  {32'h3b8f286a, 32'h3c57f966} /* (9, 25, 17) {real, imag} */,
  {32'h3ca56edd, 32'h00000000} /* (9, 25, 16) {real, imag} */,
  {32'h3b8f286a, 32'hbc57f966} /* (9, 25, 15) {real, imag} */,
  {32'h3cc00fe2, 32'hbe0214ae} /* (9, 25, 14) {real, imag} */,
  {32'hbda3e279, 32'h3c2626ad} /* (9, 25, 13) {real, imag} */,
  {32'hbd933757, 32'hbcc8e554} /* (9, 25, 12) {real, imag} */,
  {32'h3cff5294, 32'hbd750308} /* (9, 25, 11) {real, imag} */,
  {32'h3d63798f, 32'h3e252f08} /* (9, 25, 10) {real, imag} */,
  {32'h3a449660, 32'h3c6fb2ee} /* (9, 25, 9) {real, imag} */,
  {32'h3d711a3e, 32'hbe0ad227} /* (9, 25, 8) {real, imag} */,
  {32'h3d82e64c, 32'hbdd8c89c} /* (9, 25, 7) {real, imag} */,
  {32'hbd208c60, 32'h3d278e86} /* (9, 25, 6) {real, imag} */,
  {32'hbe505bf4, 32'hbd83abfd} /* (9, 25, 5) {real, imag} */,
  {32'h3db33a65, 32'h3dd9be1e} /* (9, 25, 4) {real, imag} */,
  {32'hbdab52b6, 32'hbb8612f0} /* (9, 25, 3) {real, imag} */,
  {32'hbfcd72f3, 32'hbe873dee} /* (9, 25, 2) {real, imag} */,
  {32'h40972706, 32'h3ebaa238} /* (9, 25, 1) {real, imag} */,
  {32'h409c3cd4, 32'h00000000} /* (9, 25, 0) {real, imag} */,
  {32'h40818981, 32'hbe1f48e8} /* (9, 24, 31) {real, imag} */,
  {32'hbfb22063, 32'h3e9adee7} /* (9, 24, 30) {real, imag} */,
  {32'hbe43110e, 32'hbe06fed8} /* (9, 24, 29) {real, imag} */,
  {32'h3e967d17, 32'h3c2806e0} /* (9, 24, 28) {real, imag} */,
  {32'hbe637fe7, 32'hbcb27bfd} /* (9, 24, 27) {real, imag} */,
  {32'hbda72041, 32'hbdb0c35b} /* (9, 24, 26) {real, imag} */,
  {32'h3d5f916a, 32'hbdb0f486} /* (9, 24, 25) {real, imag} */,
  {32'hbe4d5843, 32'h3e26df2b} /* (9, 24, 24) {real, imag} */,
  {32'hbd09d3fe, 32'hbe096206} /* (9, 24, 23) {real, imag} */,
  {32'h3a493da0, 32'h3de47727} /* (9, 24, 22) {real, imag} */,
  {32'hbdae5ce6, 32'h3d426866} /* (9, 24, 21) {real, imag} */,
  {32'h3c5f1028, 32'hbca9b786} /* (9, 24, 20) {real, imag} */,
  {32'h3d48fb5a, 32'h3cb60c2d} /* (9, 24, 19) {real, imag} */,
  {32'h3d174c28, 32'h3dd7949b} /* (9, 24, 18) {real, imag} */,
  {32'h3ceff92e, 32'hbcd1c60c} /* (9, 24, 17) {real, imag} */,
  {32'h3d0a79ac, 32'h00000000} /* (9, 24, 16) {real, imag} */,
  {32'h3ceff92e, 32'h3cd1c60c} /* (9, 24, 15) {real, imag} */,
  {32'h3d174c28, 32'hbdd7949b} /* (9, 24, 14) {real, imag} */,
  {32'h3d48fb5a, 32'hbcb60c2d} /* (9, 24, 13) {real, imag} */,
  {32'h3c5f1028, 32'h3ca9b786} /* (9, 24, 12) {real, imag} */,
  {32'hbdae5ce6, 32'hbd426866} /* (9, 24, 11) {real, imag} */,
  {32'h3a493da0, 32'hbde47727} /* (9, 24, 10) {real, imag} */,
  {32'hbd09d3fe, 32'h3e096206} /* (9, 24, 9) {real, imag} */,
  {32'hbe4d5843, 32'hbe26df2b} /* (9, 24, 8) {real, imag} */,
  {32'h3d5f916a, 32'h3db0f486} /* (9, 24, 7) {real, imag} */,
  {32'hbda72041, 32'h3db0c35b} /* (9, 24, 6) {real, imag} */,
  {32'hbe637fe7, 32'h3cb27bfd} /* (9, 24, 5) {real, imag} */,
  {32'h3e967d17, 32'hbc2806e0} /* (9, 24, 4) {real, imag} */,
  {32'hbe43110e, 32'h3e06fed8} /* (9, 24, 3) {real, imag} */,
  {32'hbfb22063, 32'hbe9adee7} /* (9, 24, 2) {real, imag} */,
  {32'h40818981, 32'h3e1f48e8} /* (9, 24, 1) {real, imag} */,
  {32'h4084cf5a, 32'h00000000} /* (9, 24, 0) {real, imag} */,
  {32'h404e33da, 32'hbe33120c} /* (9, 23, 31) {real, imag} */,
  {32'hbf9b486b, 32'h3e72c863} /* (9, 23, 30) {real, imag} */,
  {32'hbdf17542, 32'hbcc5f0eb} /* (9, 23, 29) {real, imag} */,
  {32'h3e804937, 32'hbdd63244} /* (9, 23, 28) {real, imag} */,
  {32'hbe750eaa, 32'h3dffd0be} /* (9, 23, 27) {real, imag} */,
  {32'hbd2606a8, 32'h3d648624} /* (9, 23, 26) {real, imag} */,
  {32'h3da153b9, 32'hbd420dd8} /* (9, 23, 25) {real, imag} */,
  {32'h39d11bc0, 32'h3bb342a8} /* (9, 23, 24) {real, imag} */,
  {32'hbd67e4d5, 32'hbd077cf7} /* (9, 23, 23) {real, imag} */,
  {32'h3c39f7db, 32'h3d9d0b4d} /* (9, 23, 22) {real, imag} */,
  {32'h3c3cc99c, 32'h3d87759c} /* (9, 23, 21) {real, imag} */,
  {32'hbd492794, 32'hbd88176e} /* (9, 23, 20) {real, imag} */,
  {32'hbbd95d72, 32'h3d4de485} /* (9, 23, 19) {real, imag} */,
  {32'hbd15b147, 32'h3d022e40} /* (9, 23, 18) {real, imag} */,
  {32'hbd23988b, 32'hbdbc1242} /* (9, 23, 17) {real, imag} */,
  {32'h3d6ac61e, 32'h00000000} /* (9, 23, 16) {real, imag} */,
  {32'hbd23988b, 32'h3dbc1242} /* (9, 23, 15) {real, imag} */,
  {32'hbd15b147, 32'hbd022e40} /* (9, 23, 14) {real, imag} */,
  {32'hbbd95d72, 32'hbd4de485} /* (9, 23, 13) {real, imag} */,
  {32'hbd492794, 32'h3d88176e} /* (9, 23, 12) {real, imag} */,
  {32'h3c3cc99c, 32'hbd87759c} /* (9, 23, 11) {real, imag} */,
  {32'h3c39f7db, 32'hbd9d0b4d} /* (9, 23, 10) {real, imag} */,
  {32'hbd67e4d5, 32'h3d077cf7} /* (9, 23, 9) {real, imag} */,
  {32'h39d11bc0, 32'hbbb342a8} /* (9, 23, 8) {real, imag} */,
  {32'h3da153b9, 32'h3d420dd8} /* (9, 23, 7) {real, imag} */,
  {32'hbd2606a8, 32'hbd648624} /* (9, 23, 6) {real, imag} */,
  {32'hbe750eaa, 32'hbdffd0be} /* (9, 23, 5) {real, imag} */,
  {32'h3e804937, 32'h3dd63244} /* (9, 23, 4) {real, imag} */,
  {32'hbdf17542, 32'h3cc5f0eb} /* (9, 23, 3) {real, imag} */,
  {32'hbf9b486b, 32'hbe72c863} /* (9, 23, 2) {real, imag} */,
  {32'h404e33da, 32'h3e33120c} /* (9, 23, 1) {real, imag} */,
  {32'h405373fe, 32'h00000000} /* (9, 23, 0) {real, imag} */,
  {32'h400f0cd4, 32'hbe46abc6} /* (9, 22, 31) {real, imag} */,
  {32'hbf55ae5c, 32'h3d996730} /* (9, 22, 30) {real, imag} */,
  {32'hbd72bedc, 32'h3e0928ae} /* (9, 22, 29) {real, imag} */,
  {32'h3d775afe, 32'hbdc0e412} /* (9, 22, 28) {real, imag} */,
  {32'hbea2912c, 32'h3d66bce4} /* (9, 22, 27) {real, imag} */,
  {32'hbd1e9fd0, 32'h3c932362} /* (9, 22, 26) {real, imag} */,
  {32'hbdafa2fb, 32'h3daaacea} /* (9, 22, 25) {real, imag} */,
  {32'hbcb306dc, 32'h3ceff042} /* (9, 22, 24) {real, imag} */,
  {32'hbd6a7d4a, 32'h3d2e5e20} /* (9, 22, 23) {real, imag} */,
  {32'h3d8df493, 32'hbcf3be1d} /* (9, 22, 22) {real, imag} */,
  {32'h3c13c540, 32'hbd81c8ce} /* (9, 22, 21) {real, imag} */,
  {32'h3c6d16c7, 32'hbca6af21} /* (9, 22, 20) {real, imag} */,
  {32'hbd0d7c51, 32'h3aab7b80} /* (9, 22, 19) {real, imag} */,
  {32'h3b85e844, 32'h3d795df4} /* (9, 22, 18) {real, imag} */,
  {32'h3d9afd2f, 32'hbd242ef2} /* (9, 22, 17) {real, imag} */,
  {32'hbdb6cb15, 32'h00000000} /* (9, 22, 16) {real, imag} */,
  {32'h3d9afd2f, 32'h3d242ef2} /* (9, 22, 15) {real, imag} */,
  {32'h3b85e844, 32'hbd795df4} /* (9, 22, 14) {real, imag} */,
  {32'hbd0d7c51, 32'hbaab7b80} /* (9, 22, 13) {real, imag} */,
  {32'h3c6d16c7, 32'h3ca6af21} /* (9, 22, 12) {real, imag} */,
  {32'h3c13c540, 32'h3d81c8ce} /* (9, 22, 11) {real, imag} */,
  {32'h3d8df493, 32'h3cf3be1d} /* (9, 22, 10) {real, imag} */,
  {32'hbd6a7d4a, 32'hbd2e5e20} /* (9, 22, 9) {real, imag} */,
  {32'hbcb306dc, 32'hbceff042} /* (9, 22, 8) {real, imag} */,
  {32'hbdafa2fb, 32'hbdaaacea} /* (9, 22, 7) {real, imag} */,
  {32'hbd1e9fd0, 32'hbc932362} /* (9, 22, 6) {real, imag} */,
  {32'hbea2912c, 32'hbd66bce4} /* (9, 22, 5) {real, imag} */,
  {32'h3d775afe, 32'h3dc0e412} /* (9, 22, 4) {real, imag} */,
  {32'hbd72bedc, 32'hbe0928ae} /* (9, 22, 3) {real, imag} */,
  {32'hbf55ae5c, 32'hbd996730} /* (9, 22, 2) {real, imag} */,
  {32'h400f0cd4, 32'h3e46abc6} /* (9, 22, 1) {real, imag} */,
  {32'h401baa7e, 32'h00000000} /* (9, 22, 0) {real, imag} */,
  {32'h3f2276b1, 32'hbd5207d8} /* (9, 21, 31) {real, imag} */,
  {32'hbe6c9442, 32'hbd03ed84} /* (9, 21, 30) {real, imag} */,
  {32'hbce738eb, 32'h3e443598} /* (9, 21, 29) {real, imag} */,
  {32'h3db56ee3, 32'hbc84ccc4} /* (9, 21, 28) {real, imag} */,
  {32'hbe14cbab, 32'h3d3139ed} /* (9, 21, 27) {real, imag} */,
  {32'h3d3ab74d, 32'hbc088f30} /* (9, 21, 26) {real, imag} */,
  {32'hbdd18561, 32'hbdac569e} /* (9, 21, 25) {real, imag} */,
  {32'hbdbcaa7d, 32'h3e1cb806} /* (9, 21, 24) {real, imag} */,
  {32'hbba7d1f0, 32'hbd36f7b8} /* (9, 21, 23) {real, imag} */,
  {32'hbd328cf8, 32'hbd9bc405} /* (9, 21, 22) {real, imag} */,
  {32'hbdbca0cf, 32'h3d2d4b51} /* (9, 21, 21) {real, imag} */,
  {32'h3d4849da, 32'hbe10aac2} /* (9, 21, 20) {real, imag} */,
  {32'hbd830655, 32'hbd991186} /* (9, 21, 19) {real, imag} */,
  {32'h3dcad2ca, 32'h3d920a09} /* (9, 21, 18) {real, imag} */,
  {32'h3afcb5f8, 32'hbda1270e} /* (9, 21, 17) {real, imag} */,
  {32'h3d6c2087, 32'h00000000} /* (9, 21, 16) {real, imag} */,
  {32'h3afcb5f8, 32'h3da1270e} /* (9, 21, 15) {real, imag} */,
  {32'h3dcad2ca, 32'hbd920a09} /* (9, 21, 14) {real, imag} */,
  {32'hbd830655, 32'h3d991186} /* (9, 21, 13) {real, imag} */,
  {32'h3d4849da, 32'h3e10aac2} /* (9, 21, 12) {real, imag} */,
  {32'hbdbca0cf, 32'hbd2d4b51} /* (9, 21, 11) {real, imag} */,
  {32'hbd328cf8, 32'h3d9bc405} /* (9, 21, 10) {real, imag} */,
  {32'hbba7d1f0, 32'h3d36f7b8} /* (9, 21, 9) {real, imag} */,
  {32'hbdbcaa7d, 32'hbe1cb806} /* (9, 21, 8) {real, imag} */,
  {32'hbdd18561, 32'h3dac569e} /* (9, 21, 7) {real, imag} */,
  {32'h3d3ab74d, 32'h3c088f30} /* (9, 21, 6) {real, imag} */,
  {32'hbe14cbab, 32'hbd3139ed} /* (9, 21, 5) {real, imag} */,
  {32'h3db56ee3, 32'h3c84ccc4} /* (9, 21, 4) {real, imag} */,
  {32'hbce738eb, 32'hbe443598} /* (9, 21, 3) {real, imag} */,
  {32'hbe6c9442, 32'h3d03ed84} /* (9, 21, 2) {real, imag} */,
  {32'h3f2276b1, 32'h3d5207d8} /* (9, 21, 1) {real, imag} */,
  {32'h3f8b0775, 32'h00000000} /* (9, 21, 0) {real, imag} */,
  {32'hbfa37382, 32'h3de5c240} /* (9, 20, 31) {real, imag} */,
  {32'h3efa8a88, 32'hbe772e4f} /* (9, 20, 30) {real, imag} */,
  {32'h3c862aa4, 32'h3e16a083} /* (9, 20, 29) {real, imag} */,
  {32'hbe316a45, 32'hbd4c269c} /* (9, 20, 28) {real, imag} */,
  {32'h3d9fae32, 32'hbd019336} /* (9, 20, 27) {real, imag} */,
  {32'h3df8b1cc, 32'hbc89f9e3} /* (9, 20, 26) {real, imag} */,
  {32'hbca36cb9, 32'hbd185782} /* (9, 20, 25) {real, imag} */,
  {32'h3d70d975, 32'hbcfe95b4} /* (9, 20, 24) {real, imag} */,
  {32'hbdb1277a, 32'hbca1eb88} /* (9, 20, 23) {real, imag} */,
  {32'hbcbab4f0, 32'h3cb4dc10} /* (9, 20, 22) {real, imag} */,
  {32'h3c457a9e, 32'hbdb876e8} /* (9, 20, 21) {real, imag} */,
  {32'hbbb67292, 32'hbd0135f2} /* (9, 20, 20) {real, imag} */,
  {32'h3dca447d, 32'h3c0c0460} /* (9, 20, 19) {real, imag} */,
  {32'h3c5ef817, 32'hbd3ffeea} /* (9, 20, 18) {real, imag} */,
  {32'h39a718c0, 32'h3d06ff5f} /* (9, 20, 17) {real, imag} */,
  {32'h3dbb0d3a, 32'h00000000} /* (9, 20, 16) {real, imag} */,
  {32'h39a718c0, 32'hbd06ff5f} /* (9, 20, 15) {real, imag} */,
  {32'h3c5ef817, 32'h3d3ffeea} /* (9, 20, 14) {real, imag} */,
  {32'h3dca447d, 32'hbc0c0460} /* (9, 20, 13) {real, imag} */,
  {32'hbbb67292, 32'h3d0135f2} /* (9, 20, 12) {real, imag} */,
  {32'h3c457a9e, 32'h3db876e8} /* (9, 20, 11) {real, imag} */,
  {32'hbcbab4f0, 32'hbcb4dc10} /* (9, 20, 10) {real, imag} */,
  {32'hbdb1277a, 32'h3ca1eb88} /* (9, 20, 9) {real, imag} */,
  {32'h3d70d975, 32'h3cfe95b4} /* (9, 20, 8) {real, imag} */,
  {32'hbca36cb9, 32'h3d185782} /* (9, 20, 7) {real, imag} */,
  {32'h3df8b1cc, 32'h3c89f9e3} /* (9, 20, 6) {real, imag} */,
  {32'h3d9fae32, 32'h3d019336} /* (9, 20, 5) {real, imag} */,
  {32'hbe316a45, 32'h3d4c269c} /* (9, 20, 4) {real, imag} */,
  {32'h3c862aa4, 32'hbe16a083} /* (9, 20, 3) {real, imag} */,
  {32'h3efa8a88, 32'h3e772e4f} /* (9, 20, 2) {real, imag} */,
  {32'hbfa37382, 32'hbde5c240} /* (9, 20, 1) {real, imag} */,
  {32'hbf0b07e4, 32'h00000000} /* (9, 20, 0) {real, imag} */,
  {32'hc0272452, 32'h3e3ed0e0} /* (9, 19, 31) {real, imag} */,
  {32'h3f8fe2b7, 32'hbecbe218} /* (9, 19, 30) {real, imag} */,
  {32'hbd567e2a, 32'h3e322659} /* (9, 19, 29) {real, imag} */,
  {32'hbe452e81, 32'h3d27d064} /* (9, 19, 28) {real, imag} */,
  {32'h3e04a652, 32'h3ca8e4e0} /* (9, 19, 27) {real, imag} */,
  {32'h3d88525e, 32'hbdd57f85} /* (9, 19, 26) {real, imag} */,
  {32'hbcb647e4, 32'h3e0e37cc} /* (9, 19, 25) {real, imag} */,
  {32'h3dc87466, 32'hbcc7a30a} /* (9, 19, 24) {real, imag} */,
  {32'h3d901333, 32'hbc47d4f7} /* (9, 19, 23) {real, imag} */,
  {32'h3cc9289c, 32'hbc8b9112} /* (9, 19, 22) {real, imag} */,
  {32'h3c898176, 32'hbda5c2e4} /* (9, 19, 21) {real, imag} */,
  {32'hb9914c20, 32'h3d45e7eb} /* (9, 19, 20) {real, imag} */,
  {32'hbd7063f0, 32'h3b7995c0} /* (9, 19, 19) {real, imag} */,
  {32'h3e020ba5, 32'hbd51f142} /* (9, 19, 18) {real, imag} */,
  {32'hbbdd8d80, 32'hbb9b74e9} /* (9, 19, 17) {real, imag} */,
  {32'hbc0210c1, 32'h00000000} /* (9, 19, 16) {real, imag} */,
  {32'hbbdd8d80, 32'h3b9b74e9} /* (9, 19, 15) {real, imag} */,
  {32'h3e020ba5, 32'h3d51f142} /* (9, 19, 14) {real, imag} */,
  {32'hbd7063f0, 32'hbb7995c0} /* (9, 19, 13) {real, imag} */,
  {32'hb9914c20, 32'hbd45e7eb} /* (9, 19, 12) {real, imag} */,
  {32'h3c898176, 32'h3da5c2e4} /* (9, 19, 11) {real, imag} */,
  {32'h3cc9289c, 32'h3c8b9112} /* (9, 19, 10) {real, imag} */,
  {32'h3d901333, 32'h3c47d4f7} /* (9, 19, 9) {real, imag} */,
  {32'h3dc87466, 32'h3cc7a30a} /* (9, 19, 8) {real, imag} */,
  {32'hbcb647e4, 32'hbe0e37cc} /* (9, 19, 7) {real, imag} */,
  {32'h3d88525e, 32'h3dd57f85} /* (9, 19, 6) {real, imag} */,
  {32'h3e04a652, 32'hbca8e4e0} /* (9, 19, 5) {real, imag} */,
  {32'hbe452e81, 32'hbd27d064} /* (9, 19, 4) {real, imag} */,
  {32'hbd567e2a, 32'hbe322659} /* (9, 19, 3) {real, imag} */,
  {32'h3f8fe2b7, 32'h3ecbe218} /* (9, 19, 2) {real, imag} */,
  {32'hc0272452, 32'hbe3ed0e0} /* (9, 19, 1) {real, imag} */,
  {32'hbfe0c5c5, 32'h00000000} /* (9, 19, 0) {real, imag} */,
  {32'hc066e06f, 32'h3ead142e} /* (9, 18, 31) {real, imag} */,
  {32'h3fa8d5ff, 32'hbeb9d92a} /* (9, 18, 30) {real, imag} */,
  {32'hbd93c72e, 32'h3daa07df} /* (9, 18, 29) {real, imag} */,
  {32'hbe762732, 32'hbc240844} /* (9, 18, 28) {real, imag} */,
  {32'h3e6a8c94, 32'h3d8ce85c} /* (9, 18, 27) {real, imag} */,
  {32'h3dbaeeb1, 32'hbca18c39} /* (9, 18, 26) {real, imag} */,
  {32'hbe0895f8, 32'h3cb3528e} /* (9, 18, 25) {real, imag} */,
  {32'h3da77fe6, 32'hbd116aec} /* (9, 18, 24) {real, imag} */,
  {32'hbdaf005e, 32'h3d12cbd2} /* (9, 18, 23) {real, imag} */,
  {32'h3da5da0c, 32'h3c8db913} /* (9, 18, 22) {real, imag} */,
  {32'hbd999b3b, 32'hbda458ce} /* (9, 18, 21) {real, imag} */,
  {32'h3cb9fdd1, 32'h3b228280} /* (9, 18, 20) {real, imag} */,
  {32'h3d0cbebe, 32'h3c5e2fd2} /* (9, 18, 19) {real, imag} */,
  {32'h3d0ebcfe, 32'hbd41cd1c} /* (9, 18, 18) {real, imag} */,
  {32'hbc16614b, 32'h3d1ce820} /* (9, 18, 17) {real, imag} */,
  {32'h3dda3e37, 32'h00000000} /* (9, 18, 16) {real, imag} */,
  {32'hbc16614b, 32'hbd1ce820} /* (9, 18, 15) {real, imag} */,
  {32'h3d0ebcfe, 32'h3d41cd1c} /* (9, 18, 14) {real, imag} */,
  {32'h3d0cbebe, 32'hbc5e2fd2} /* (9, 18, 13) {real, imag} */,
  {32'h3cb9fdd1, 32'hbb228280} /* (9, 18, 12) {real, imag} */,
  {32'hbd999b3b, 32'h3da458ce} /* (9, 18, 11) {real, imag} */,
  {32'h3da5da0c, 32'hbc8db913} /* (9, 18, 10) {real, imag} */,
  {32'hbdaf005e, 32'hbd12cbd2} /* (9, 18, 9) {real, imag} */,
  {32'h3da77fe6, 32'h3d116aec} /* (9, 18, 8) {real, imag} */,
  {32'hbe0895f8, 32'hbcb3528e} /* (9, 18, 7) {real, imag} */,
  {32'h3dbaeeb1, 32'h3ca18c39} /* (9, 18, 6) {real, imag} */,
  {32'h3e6a8c94, 32'hbd8ce85c} /* (9, 18, 5) {real, imag} */,
  {32'hbe762732, 32'h3c240844} /* (9, 18, 4) {real, imag} */,
  {32'hbd93c72e, 32'hbdaa07df} /* (9, 18, 3) {real, imag} */,
  {32'h3fa8d5ff, 32'h3eb9d92a} /* (9, 18, 2) {real, imag} */,
  {32'hc066e06f, 32'hbead142e} /* (9, 18, 1) {real, imag} */,
  {32'hc01f64db, 32'h00000000} /* (9, 18, 0) {real, imag} */,
  {32'hc084309d, 32'h3eb52f12} /* (9, 17, 31) {real, imag} */,
  {32'h3fba857c, 32'hbe20febc} /* (9, 17, 30) {real, imag} */,
  {32'h3d312796, 32'hbc31789c} /* (9, 17, 29) {real, imag} */,
  {32'hbe6b7fa4, 32'h3cc23568} /* (9, 17, 28) {real, imag} */,
  {32'h3ea03589, 32'hbc7e4fc8} /* (9, 17, 27) {real, imag} */,
  {32'h3e14972c, 32'hbd3584fc} /* (9, 17, 26) {real, imag} */,
  {32'hbdb4fd3c, 32'hbb73e148} /* (9, 17, 25) {real, imag} */,
  {32'h3da37f7a, 32'h3b9c7380} /* (9, 17, 24) {real, imag} */,
  {32'h3d816b0a, 32'hbbac6252} /* (9, 17, 23) {real, imag} */,
  {32'h3dea3f92, 32'h3dd1bd02} /* (9, 17, 22) {real, imag} */,
  {32'hbcc31c2a, 32'hbd145b63} /* (9, 17, 21) {real, imag} */,
  {32'hbda37095, 32'h3d57b479} /* (9, 17, 20) {real, imag} */,
  {32'h3d7ff9d2, 32'h3bf17276} /* (9, 17, 19) {real, imag} */,
  {32'hbcf9906c, 32'hbd2ddc2c} /* (9, 17, 18) {real, imag} */,
  {32'h3ce823e6, 32'h3c178544} /* (9, 17, 17) {real, imag} */,
  {32'hbd8a4bae, 32'h00000000} /* (9, 17, 16) {real, imag} */,
  {32'h3ce823e6, 32'hbc178544} /* (9, 17, 15) {real, imag} */,
  {32'hbcf9906c, 32'h3d2ddc2c} /* (9, 17, 14) {real, imag} */,
  {32'h3d7ff9d2, 32'hbbf17276} /* (9, 17, 13) {real, imag} */,
  {32'hbda37095, 32'hbd57b479} /* (9, 17, 12) {real, imag} */,
  {32'hbcc31c2a, 32'h3d145b63} /* (9, 17, 11) {real, imag} */,
  {32'h3dea3f92, 32'hbdd1bd02} /* (9, 17, 10) {real, imag} */,
  {32'h3d816b0a, 32'h3bac6252} /* (9, 17, 9) {real, imag} */,
  {32'h3da37f7a, 32'hbb9c7380} /* (9, 17, 8) {real, imag} */,
  {32'hbdb4fd3c, 32'h3b73e148} /* (9, 17, 7) {real, imag} */,
  {32'h3e14972c, 32'h3d3584fc} /* (9, 17, 6) {real, imag} */,
  {32'h3ea03589, 32'h3c7e4fc8} /* (9, 17, 5) {real, imag} */,
  {32'hbe6b7fa4, 32'hbcc23568} /* (9, 17, 4) {real, imag} */,
  {32'h3d312796, 32'h3c31789c} /* (9, 17, 3) {real, imag} */,
  {32'h3fba857c, 32'h3e20febc} /* (9, 17, 2) {real, imag} */,
  {32'hc084309d, 32'hbeb52f12} /* (9, 17, 1) {real, imag} */,
  {32'hc04fec68, 32'h00000000} /* (9, 17, 0) {real, imag} */,
  {32'hc089f147, 32'h3eb6035c} /* (9, 16, 31) {real, imag} */,
  {32'h3fc68b90, 32'hbe19f3d0} /* (9, 16, 30) {real, imag} */,
  {32'hbd3a3a3a, 32'h3cec0622} /* (9, 16, 29) {real, imag} */,
  {32'hbd95ea78, 32'h3d185666} /* (9, 16, 28) {real, imag} */,
  {32'h3e80b7cd, 32'hbd8857f2} /* (9, 16, 27) {real, imag} */,
  {32'h3e068dce, 32'hbc90ca5a} /* (9, 16, 26) {real, imag} */,
  {32'hbc33a02c, 32'h3cf2d110} /* (9, 16, 25) {real, imag} */,
  {32'h3da4d2ec, 32'h3ce32173} /* (9, 16, 24) {real, imag} */,
  {32'h3d157c90, 32'h3c548940} /* (9, 16, 23) {real, imag} */,
  {32'h3bcd0af0, 32'hba8fc700} /* (9, 16, 22) {real, imag} */,
  {32'h3da0df65, 32'h3d1d7b33} /* (9, 16, 21) {real, imag} */,
  {32'hbba745a8, 32'hbd5bb5fa} /* (9, 16, 20) {real, imag} */,
  {32'hbceaf7ea, 32'hbdadea93} /* (9, 16, 19) {real, imag} */,
  {32'h3c01b3e1, 32'hbd8734ae} /* (9, 16, 18) {real, imag} */,
  {32'hbcc3a9d6, 32'hbca1dd61} /* (9, 16, 17) {real, imag} */,
  {32'h3c117098, 32'h00000000} /* (9, 16, 16) {real, imag} */,
  {32'hbcc3a9d6, 32'h3ca1dd61} /* (9, 16, 15) {real, imag} */,
  {32'h3c01b3e1, 32'h3d8734ae} /* (9, 16, 14) {real, imag} */,
  {32'hbceaf7ea, 32'h3dadea93} /* (9, 16, 13) {real, imag} */,
  {32'hbba745a8, 32'h3d5bb5fa} /* (9, 16, 12) {real, imag} */,
  {32'h3da0df65, 32'hbd1d7b33} /* (9, 16, 11) {real, imag} */,
  {32'h3bcd0af0, 32'h3a8fc700} /* (9, 16, 10) {real, imag} */,
  {32'h3d157c90, 32'hbc548940} /* (9, 16, 9) {real, imag} */,
  {32'h3da4d2ec, 32'hbce32173} /* (9, 16, 8) {real, imag} */,
  {32'hbc33a02c, 32'hbcf2d110} /* (9, 16, 7) {real, imag} */,
  {32'h3e068dce, 32'h3c90ca5a} /* (9, 16, 6) {real, imag} */,
  {32'h3e80b7cd, 32'h3d8857f2} /* (9, 16, 5) {real, imag} */,
  {32'hbd95ea78, 32'hbd185666} /* (9, 16, 4) {real, imag} */,
  {32'hbd3a3a3a, 32'hbcec0622} /* (9, 16, 3) {real, imag} */,
  {32'h3fc68b90, 32'h3e19f3d0} /* (9, 16, 2) {real, imag} */,
  {32'hc089f147, 32'hbeb6035c} /* (9, 16, 1) {real, imag} */,
  {32'hc057fb42, 32'h00000000} /* (9, 16, 0) {real, imag} */,
  {32'hc0894b6b, 32'h3ea2746e} /* (9, 15, 31) {real, imag} */,
  {32'h3fc30904, 32'hbe51fb8c} /* (9, 15, 30) {real, imag} */,
  {32'h3beaa870, 32'hbc4476dc} /* (9, 15, 29) {real, imag} */,
  {32'hbe5d7316, 32'h3d12ee20} /* (9, 15, 28) {real, imag} */,
  {32'h3e29d75a, 32'hbde9a025} /* (9, 15, 27) {real, imag} */,
  {32'h3dbadbdf, 32'h3cc72a1f} /* (9, 15, 26) {real, imag} */,
  {32'hbd01ec4c, 32'hbc0ff8a6} /* (9, 15, 25) {real, imag} */,
  {32'h3dd1c740, 32'h3ca3ba88} /* (9, 15, 24) {real, imag} */,
  {32'hbcf367ef, 32'h3c6e3deb} /* (9, 15, 23) {real, imag} */,
  {32'hbb9e77f8, 32'hbd5583b0} /* (9, 15, 22) {real, imag} */,
  {32'h3cc90d3c, 32'hbcbc3204} /* (9, 15, 21) {real, imag} */,
  {32'hbd28822e, 32'hbd7f6437} /* (9, 15, 20) {real, imag} */,
  {32'hbd731b4e, 32'hbb8a9446} /* (9, 15, 19) {real, imag} */,
  {32'h3c2e5f21, 32'hbc0b017c} /* (9, 15, 18) {real, imag} */,
  {32'hbd2d4c11, 32'h3d22ede9} /* (9, 15, 17) {real, imag} */,
  {32'hbd3886f0, 32'h00000000} /* (9, 15, 16) {real, imag} */,
  {32'hbd2d4c11, 32'hbd22ede9} /* (9, 15, 15) {real, imag} */,
  {32'h3c2e5f21, 32'h3c0b017c} /* (9, 15, 14) {real, imag} */,
  {32'hbd731b4e, 32'h3b8a9446} /* (9, 15, 13) {real, imag} */,
  {32'hbd28822e, 32'h3d7f6437} /* (9, 15, 12) {real, imag} */,
  {32'h3cc90d3c, 32'h3cbc3204} /* (9, 15, 11) {real, imag} */,
  {32'hbb9e77f8, 32'h3d5583b0} /* (9, 15, 10) {real, imag} */,
  {32'hbcf367ef, 32'hbc6e3deb} /* (9, 15, 9) {real, imag} */,
  {32'h3dd1c740, 32'hbca3ba88} /* (9, 15, 8) {real, imag} */,
  {32'hbd01ec4c, 32'h3c0ff8a6} /* (9, 15, 7) {real, imag} */,
  {32'h3dbadbdf, 32'hbcc72a1f} /* (9, 15, 6) {real, imag} */,
  {32'h3e29d75a, 32'h3de9a025} /* (9, 15, 5) {real, imag} */,
  {32'hbe5d7316, 32'hbd12ee20} /* (9, 15, 4) {real, imag} */,
  {32'h3beaa870, 32'h3c4476dc} /* (9, 15, 3) {real, imag} */,
  {32'h3fc30904, 32'h3e51fb8c} /* (9, 15, 2) {real, imag} */,
  {32'hc0894b6b, 32'hbea2746e} /* (9, 15, 1) {real, imag} */,
  {32'hc04f7f1e, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'hc07884bb, 32'h3eba7cba} /* (9, 14, 31) {real, imag} */,
  {32'h3fb70375, 32'hbe4445cc} /* (9, 14, 30) {real, imag} */,
  {32'h3dcafb5a, 32'h3e05e0ce} /* (9, 14, 29) {real, imag} */,
  {32'hbe8ada2d, 32'hbd958b78} /* (9, 14, 28) {real, imag} */,
  {32'h3e1a1c74, 32'hbdfe884e} /* (9, 14, 27) {real, imag} */,
  {32'hbce173d8, 32'h3d55c078} /* (9, 14, 26) {real, imag} */,
  {32'hbcbf42fc, 32'h3d587d97} /* (9, 14, 25) {real, imag} */,
  {32'h3de626f4, 32'h3d2dbfd4} /* (9, 14, 24) {real, imag} */,
  {32'h3da57774, 32'hbd552b1e} /* (9, 14, 23) {real, imag} */,
  {32'h3deea30e, 32'h3d59d7fe} /* (9, 14, 22) {real, imag} */,
  {32'h3d55ea3a, 32'hbd89da0a} /* (9, 14, 21) {real, imag} */,
  {32'hbb33a5c8, 32'hbd8fc69c} /* (9, 14, 20) {real, imag} */,
  {32'hbd10a58e, 32'h3c9b266b} /* (9, 14, 19) {real, imag} */,
  {32'hbd23ff82, 32'h3be7c3f0} /* (9, 14, 18) {real, imag} */,
  {32'h3c0a5101, 32'h3d73c104} /* (9, 14, 17) {real, imag} */,
  {32'h3d9a0625, 32'h00000000} /* (9, 14, 16) {real, imag} */,
  {32'h3c0a5101, 32'hbd73c104} /* (9, 14, 15) {real, imag} */,
  {32'hbd23ff82, 32'hbbe7c3f0} /* (9, 14, 14) {real, imag} */,
  {32'hbd10a58e, 32'hbc9b266b} /* (9, 14, 13) {real, imag} */,
  {32'hbb33a5c8, 32'h3d8fc69c} /* (9, 14, 12) {real, imag} */,
  {32'h3d55ea3a, 32'h3d89da0a} /* (9, 14, 11) {real, imag} */,
  {32'h3deea30e, 32'hbd59d7fe} /* (9, 14, 10) {real, imag} */,
  {32'h3da57774, 32'h3d552b1e} /* (9, 14, 9) {real, imag} */,
  {32'h3de626f4, 32'hbd2dbfd4} /* (9, 14, 8) {real, imag} */,
  {32'hbcbf42fc, 32'hbd587d97} /* (9, 14, 7) {real, imag} */,
  {32'hbce173d8, 32'hbd55c078} /* (9, 14, 6) {real, imag} */,
  {32'h3e1a1c74, 32'h3dfe884e} /* (9, 14, 5) {real, imag} */,
  {32'hbe8ada2d, 32'h3d958b78} /* (9, 14, 4) {real, imag} */,
  {32'h3dcafb5a, 32'hbe05e0ce} /* (9, 14, 3) {real, imag} */,
  {32'h3fb70375, 32'h3e4445cc} /* (9, 14, 2) {real, imag} */,
  {32'hc07884bb, 32'hbeba7cba} /* (9, 14, 1) {real, imag} */,
  {32'hc03d213d, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hc050853c, 32'h3d69cf40} /* (9, 13, 31) {real, imag} */,
  {32'h3f9f7c6f, 32'hbe07e30f} /* (9, 13, 30) {real, imag} */,
  {32'h3d4d6604, 32'h3d99b7a4} /* (9, 13, 29) {real, imag} */,
  {32'hbe9b4d73, 32'h3caed904} /* (9, 13, 28) {real, imag} */,
  {32'h3e69bf32, 32'hbdd9af50} /* (9, 13, 27) {real, imag} */,
  {32'h3c330bec, 32'h3d3e8036} /* (9, 13, 26) {real, imag} */,
  {32'hbd86f44f, 32'hbccd7898} /* (9, 13, 25) {real, imag} */,
  {32'hbd06940b, 32'h3c6d6244} /* (9, 13, 24) {real, imag} */,
  {32'hbd6da4a6, 32'hbd02a95f} /* (9, 13, 23) {real, imag} */,
  {32'hbdc0fbf9, 32'h3cfeb312} /* (9, 13, 22) {real, imag} */,
  {32'h3c22650b, 32'hbc97f8df} /* (9, 13, 21) {real, imag} */,
  {32'h3cd03ffe, 32'hbc2b8dc0} /* (9, 13, 20) {real, imag} */,
  {32'h3c0d3d02, 32'h3d7d2d06} /* (9, 13, 19) {real, imag} */,
  {32'hbd49ac04, 32'hbe277fbe} /* (9, 13, 18) {real, imag} */,
  {32'hbb8e8c58, 32'hbc877abc} /* (9, 13, 17) {real, imag} */,
  {32'h3d02d54c, 32'h00000000} /* (9, 13, 16) {real, imag} */,
  {32'hbb8e8c58, 32'h3c877abc} /* (9, 13, 15) {real, imag} */,
  {32'hbd49ac04, 32'h3e277fbe} /* (9, 13, 14) {real, imag} */,
  {32'h3c0d3d02, 32'hbd7d2d06} /* (9, 13, 13) {real, imag} */,
  {32'h3cd03ffe, 32'h3c2b8dc0} /* (9, 13, 12) {real, imag} */,
  {32'h3c22650b, 32'h3c97f8df} /* (9, 13, 11) {real, imag} */,
  {32'hbdc0fbf9, 32'hbcfeb312} /* (9, 13, 10) {real, imag} */,
  {32'hbd6da4a6, 32'h3d02a95f} /* (9, 13, 9) {real, imag} */,
  {32'hbd06940b, 32'hbc6d6244} /* (9, 13, 8) {real, imag} */,
  {32'hbd86f44f, 32'h3ccd7898} /* (9, 13, 7) {real, imag} */,
  {32'h3c330bec, 32'hbd3e8036} /* (9, 13, 6) {real, imag} */,
  {32'h3e69bf32, 32'h3dd9af50} /* (9, 13, 5) {real, imag} */,
  {32'hbe9b4d73, 32'hbcaed904} /* (9, 13, 4) {real, imag} */,
  {32'h3d4d6604, 32'hbd99b7a4} /* (9, 13, 3) {real, imag} */,
  {32'h3f9f7c6f, 32'h3e07e30f} /* (9, 13, 2) {real, imag} */,
  {32'hc050853c, 32'hbd69cf40} /* (9, 13, 1) {real, imag} */,
  {32'hc01d934e, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'hc01b21bd, 32'hbe182a20} /* (9, 12, 31) {real, imag} */,
  {32'h3f802ff8, 32'h3ac5e980} /* (9, 12, 30) {real, imag} */,
  {32'h3d5cfbc8, 32'h3daf0064} /* (9, 12, 29) {real, imag} */,
  {32'hbe3a18f3, 32'h3c9018b8} /* (9, 12, 28) {real, imag} */,
  {32'h3e1ba2fd, 32'hbbd548bc} /* (9, 12, 27) {real, imag} */,
  {32'h3cb68cbe, 32'hbbd720eb} /* (9, 12, 26) {real, imag} */,
  {32'hbd8ac006, 32'h3c164af8} /* (9, 12, 25) {real, imag} */,
  {32'h3dea11b2, 32'hbd74ba7c} /* (9, 12, 24) {real, imag} */,
  {32'hbbc936f8, 32'h3d866a7e} /* (9, 12, 23) {real, imag} */,
  {32'hbd53f10c, 32'h3b7a2860} /* (9, 12, 22) {real, imag} */,
  {32'hbcaf45f5, 32'hbdc247c2} /* (9, 12, 21) {real, imag} */,
  {32'h3c61e4b3, 32'hbc5a961f} /* (9, 12, 20) {real, imag} */,
  {32'hbc5d1a08, 32'hbd1859c4} /* (9, 12, 19) {real, imag} */,
  {32'hbc3d7185, 32'h3d9bd703} /* (9, 12, 18) {real, imag} */,
  {32'hbd474adc, 32'hbd8c1302} /* (9, 12, 17) {real, imag} */,
  {32'h3c468bc0, 32'h00000000} /* (9, 12, 16) {real, imag} */,
  {32'hbd474adc, 32'h3d8c1302} /* (9, 12, 15) {real, imag} */,
  {32'hbc3d7185, 32'hbd9bd703} /* (9, 12, 14) {real, imag} */,
  {32'hbc5d1a08, 32'h3d1859c4} /* (9, 12, 13) {real, imag} */,
  {32'h3c61e4b3, 32'h3c5a961f} /* (9, 12, 12) {real, imag} */,
  {32'hbcaf45f5, 32'h3dc247c2} /* (9, 12, 11) {real, imag} */,
  {32'hbd53f10c, 32'hbb7a2860} /* (9, 12, 10) {real, imag} */,
  {32'hbbc936f8, 32'hbd866a7e} /* (9, 12, 9) {real, imag} */,
  {32'h3dea11b2, 32'h3d74ba7c} /* (9, 12, 8) {real, imag} */,
  {32'hbd8ac006, 32'hbc164af8} /* (9, 12, 7) {real, imag} */,
  {32'h3cb68cbe, 32'h3bd720eb} /* (9, 12, 6) {real, imag} */,
  {32'h3e1ba2fd, 32'h3bd548bc} /* (9, 12, 5) {real, imag} */,
  {32'hbe3a18f3, 32'hbc9018b8} /* (9, 12, 4) {real, imag} */,
  {32'h3d5cfbc8, 32'hbdaf0064} /* (9, 12, 3) {real, imag} */,
  {32'h3f802ff8, 32'hbac5e980} /* (9, 12, 2) {real, imag} */,
  {32'hc01b21bd, 32'h3e182a20} /* (9, 12, 1) {real, imag} */,
  {32'hbfd33986, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'hbf8c5114, 32'hbe938701} /* (9, 11, 31) {real, imag} */,
  {32'h3f099b16, 32'h3d3b8b44} /* (9, 11, 30) {real, imag} */,
  {32'hbab67c10, 32'h3cb40ec4} /* (9, 11, 29) {real, imag} */,
  {32'hbe011512, 32'hbe0f88f6} /* (9, 11, 28) {real, imag} */,
  {32'h3d8c9572, 32'hbc8f8462} /* (9, 11, 27) {real, imag} */,
  {32'hbc93d1ae, 32'hbdb1cc2c} /* (9, 11, 26) {real, imag} */,
  {32'h3cf5768c, 32'hbd1f2b26} /* (9, 11, 25) {real, imag} */,
  {32'h3d481aca, 32'h3c4f6468} /* (9, 11, 24) {real, imag} */,
  {32'hbd24a900, 32'hba361ee0} /* (9, 11, 23) {real, imag} */,
  {32'h3dbbea08, 32'hbd4de2d7} /* (9, 11, 22) {real, imag} */,
  {32'h3d9478b3, 32'hbdf45568} /* (9, 11, 21) {real, imag} */,
  {32'hbd1363ae, 32'h3c854b68} /* (9, 11, 20) {real, imag} */,
  {32'h3ca9120f, 32'h3a6fa5c0} /* (9, 11, 19) {real, imag} */,
  {32'h3cbe9340, 32'h3cd07624} /* (9, 11, 18) {real, imag} */,
  {32'hbc497cc1, 32'h3d43a168} /* (9, 11, 17) {real, imag} */,
  {32'h3d62814f, 32'h00000000} /* (9, 11, 16) {real, imag} */,
  {32'hbc497cc1, 32'hbd43a168} /* (9, 11, 15) {real, imag} */,
  {32'h3cbe9340, 32'hbcd07624} /* (9, 11, 14) {real, imag} */,
  {32'h3ca9120f, 32'hba6fa5c0} /* (9, 11, 13) {real, imag} */,
  {32'hbd1363ae, 32'hbc854b68} /* (9, 11, 12) {real, imag} */,
  {32'h3d9478b3, 32'h3df45568} /* (9, 11, 11) {real, imag} */,
  {32'h3dbbea08, 32'h3d4de2d7} /* (9, 11, 10) {real, imag} */,
  {32'hbd24a900, 32'h3a361ee0} /* (9, 11, 9) {real, imag} */,
  {32'h3d481aca, 32'hbc4f6468} /* (9, 11, 8) {real, imag} */,
  {32'h3cf5768c, 32'h3d1f2b26} /* (9, 11, 7) {real, imag} */,
  {32'hbc93d1ae, 32'h3db1cc2c} /* (9, 11, 6) {real, imag} */,
  {32'h3d8c9572, 32'h3c8f8462} /* (9, 11, 5) {real, imag} */,
  {32'hbe011512, 32'h3e0f88f6} /* (9, 11, 4) {real, imag} */,
  {32'hbab67c10, 32'hbcb40ec4} /* (9, 11, 3) {real, imag} */,
  {32'h3f099b16, 32'hbd3b8b44} /* (9, 11, 2) {real, imag} */,
  {32'hbf8c5114, 32'h3e938701} /* (9, 11, 1) {real, imag} */,
  {32'hbeb98164, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h3f2794d0, 32'hbf31adf4} /* (9, 10, 31) {real, imag} */,
  {32'hbe8c58d0, 32'h3e631598} /* (9, 10, 30) {real, imag} */,
  {32'hbd2a1340, 32'hbd32bdca} /* (9, 10, 29) {real, imag} */,
  {32'hbda5390d, 32'hbe7ff851} /* (9, 10, 28) {real, imag} */,
  {32'hbdbe68b2, 32'h3a2a2060} /* (9, 10, 27) {real, imag} */,
  {32'h3df69ab2, 32'h3c589b60} /* (9, 10, 26) {real, imag} */,
  {32'h3d30f37a, 32'hbcb3c6d0} /* (9, 10, 25) {real, imag} */,
  {32'hbbe36392, 32'h3d8a400e} /* (9, 10, 24) {real, imag} */,
  {32'h3cf53065, 32'hbaf15780} /* (9, 10, 23) {real, imag} */,
  {32'h3d8e4de1, 32'h39e48240} /* (9, 10, 22) {real, imag} */,
  {32'hbbc98cf8, 32'hbd4604ff} /* (9, 10, 21) {real, imag} */,
  {32'h3ca76d8e, 32'h3d5d0ec4} /* (9, 10, 20) {real, imag} */,
  {32'h3dd8d4d0, 32'hbdac1d36} /* (9, 10, 19) {real, imag} */,
  {32'hbd49184c, 32'hbd917e4e} /* (9, 10, 18) {real, imag} */,
  {32'h3d03582c, 32'h3d23d38a} /* (9, 10, 17) {real, imag} */,
  {32'hbdf6bf91, 32'h00000000} /* (9, 10, 16) {real, imag} */,
  {32'h3d03582c, 32'hbd23d38a} /* (9, 10, 15) {real, imag} */,
  {32'hbd49184c, 32'h3d917e4e} /* (9, 10, 14) {real, imag} */,
  {32'h3dd8d4d0, 32'h3dac1d36} /* (9, 10, 13) {real, imag} */,
  {32'h3ca76d8e, 32'hbd5d0ec4} /* (9, 10, 12) {real, imag} */,
  {32'hbbc98cf8, 32'h3d4604ff} /* (9, 10, 11) {real, imag} */,
  {32'h3d8e4de1, 32'hb9e48240} /* (9, 10, 10) {real, imag} */,
  {32'h3cf53065, 32'h3af15780} /* (9, 10, 9) {real, imag} */,
  {32'hbbe36392, 32'hbd8a400e} /* (9, 10, 8) {real, imag} */,
  {32'h3d30f37a, 32'h3cb3c6d0} /* (9, 10, 7) {real, imag} */,
  {32'h3df69ab2, 32'hbc589b60} /* (9, 10, 6) {real, imag} */,
  {32'hbdbe68b2, 32'hba2a2060} /* (9, 10, 5) {real, imag} */,
  {32'hbda5390d, 32'h3e7ff851} /* (9, 10, 4) {real, imag} */,
  {32'hbd2a1340, 32'h3d32bdca} /* (9, 10, 3) {real, imag} */,
  {32'hbe8c58d0, 32'hbe631598} /* (9, 10, 2) {real, imag} */,
  {32'h3f2794d0, 32'h3f31adf4} /* (9, 10, 1) {real, imag} */,
  {32'h3f9007bf, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'h40004fee, 32'hbf96357a} /* (9, 9, 31) {real, imag} */,
  {32'hbf47ceac, 32'h3ec96ce2} /* (9, 9, 30) {real, imag} */,
  {32'hbd32fc59, 32'hbd2f1dae} /* (9, 9, 29) {real, imag} */,
  {32'hbd863fa9, 32'hbe47883e} /* (9, 9, 28) {real, imag} */,
  {32'hbe23305e, 32'h3d9f57bc} /* (9, 9, 27) {real, imag} */,
  {32'h3d3ef7d0, 32'hbd46bb24} /* (9, 9, 26) {real, imag} */,
  {32'h3c2983c8, 32'h3dd4505c} /* (9, 9, 25) {real, imag} */,
  {32'hbc8075e5, 32'hbcb3343a} /* (9, 9, 24) {real, imag} */,
  {32'hbd4a1383, 32'hbd46254d} /* (9, 9, 23) {real, imag} */,
  {32'hbbc9b016, 32'h3c7ae2a6} /* (9, 9, 22) {real, imag} */,
  {32'hbc496098, 32'h3a097940} /* (9, 9, 21) {real, imag} */,
  {32'h3d8e516a, 32'h3b9b5580} /* (9, 9, 20) {real, imag} */,
  {32'h3c829270, 32'hbc3498e4} /* (9, 9, 19) {real, imag} */,
  {32'h3c77a500, 32'h3d4f69bc} /* (9, 9, 18) {real, imag} */,
  {32'h3b4cdef0, 32'hbd0dc564} /* (9, 9, 17) {real, imag} */,
  {32'hbd765732, 32'h00000000} /* (9, 9, 16) {real, imag} */,
  {32'h3b4cdef0, 32'h3d0dc564} /* (9, 9, 15) {real, imag} */,
  {32'h3c77a500, 32'hbd4f69bc} /* (9, 9, 14) {real, imag} */,
  {32'h3c829270, 32'h3c3498e4} /* (9, 9, 13) {real, imag} */,
  {32'h3d8e516a, 32'hbb9b5580} /* (9, 9, 12) {real, imag} */,
  {32'hbc496098, 32'hba097940} /* (9, 9, 11) {real, imag} */,
  {32'hbbc9b016, 32'hbc7ae2a6} /* (9, 9, 10) {real, imag} */,
  {32'hbd4a1383, 32'h3d46254d} /* (9, 9, 9) {real, imag} */,
  {32'hbc8075e5, 32'h3cb3343a} /* (9, 9, 8) {real, imag} */,
  {32'h3c2983c8, 32'hbdd4505c} /* (9, 9, 7) {real, imag} */,
  {32'h3d3ef7d0, 32'h3d46bb24} /* (9, 9, 6) {real, imag} */,
  {32'hbe23305e, 32'hbd9f57bc} /* (9, 9, 5) {real, imag} */,
  {32'hbd863fa9, 32'h3e47883e} /* (9, 9, 4) {real, imag} */,
  {32'hbd32fc59, 32'h3d2f1dae} /* (9, 9, 3) {real, imag} */,
  {32'hbf47ceac, 32'hbec96ce2} /* (9, 9, 2) {real, imag} */,
  {32'h40004fee, 32'h3f96357a} /* (9, 9, 1) {real, imag} */,
  {32'h400f9792, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h4034b00a, 32'hbfb8b947} /* (9, 8, 31) {real, imag} */,
  {32'hbf8f078d, 32'h3f0d2a50} /* (9, 8, 30) {real, imag} */,
  {32'hbd90f7b8, 32'hbdfb2505} /* (9, 8, 29) {real, imag} */,
  {32'h3d18ed98, 32'hbe2143fd} /* (9, 8, 28) {real, imag} */,
  {32'hbdfc382a, 32'h3d99327d} /* (9, 8, 27) {real, imag} */,
  {32'hbd87426d, 32'h3d9de48b} /* (9, 8, 26) {real, imag} */,
  {32'h3d413866, 32'h3d26dda8} /* (9, 8, 25) {real, imag} */,
  {32'hbd5bdf2c, 32'hbd4866bc} /* (9, 8, 24) {real, imag} */,
  {32'h3c655bbe, 32'h3c18d644} /* (9, 8, 23) {real, imag} */,
  {32'h3d2c7e88, 32'h3cebeed4} /* (9, 8, 22) {real, imag} */,
  {32'hbd421fcc, 32'h3d037388} /* (9, 8, 21) {real, imag} */,
  {32'h3c969688, 32'hbcbdefac} /* (9, 8, 20) {real, imag} */,
  {32'hbcd44678, 32'hbd76fd0a} /* (9, 8, 19) {real, imag} */,
  {32'hbd6a4a1e, 32'hbc878b84} /* (9, 8, 18) {real, imag} */,
  {32'hbcac05dc, 32'hbd894762} /* (9, 8, 17) {real, imag} */,
  {32'hbd0725b6, 32'h00000000} /* (9, 8, 16) {real, imag} */,
  {32'hbcac05dc, 32'h3d894762} /* (9, 8, 15) {real, imag} */,
  {32'hbd6a4a1e, 32'h3c878b84} /* (9, 8, 14) {real, imag} */,
  {32'hbcd44678, 32'h3d76fd0a} /* (9, 8, 13) {real, imag} */,
  {32'h3c969688, 32'h3cbdefac} /* (9, 8, 12) {real, imag} */,
  {32'hbd421fcc, 32'hbd037388} /* (9, 8, 11) {real, imag} */,
  {32'h3d2c7e88, 32'hbcebeed4} /* (9, 8, 10) {real, imag} */,
  {32'h3c655bbe, 32'hbc18d644} /* (9, 8, 9) {real, imag} */,
  {32'hbd5bdf2c, 32'h3d4866bc} /* (9, 8, 8) {real, imag} */,
  {32'h3d413866, 32'hbd26dda8} /* (9, 8, 7) {real, imag} */,
  {32'hbd87426d, 32'hbd9de48b} /* (9, 8, 6) {real, imag} */,
  {32'hbdfc382a, 32'hbd99327d} /* (9, 8, 5) {real, imag} */,
  {32'h3d18ed98, 32'h3e2143fd} /* (9, 8, 4) {real, imag} */,
  {32'hbd90f7b8, 32'h3dfb2505} /* (9, 8, 3) {real, imag} */,
  {32'hbf8f078d, 32'hbf0d2a50} /* (9, 8, 2) {real, imag} */,
  {32'h4034b00a, 32'h3fb8b947} /* (9, 8, 1) {real, imag} */,
  {32'h405a19f1, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h40564cfd, 32'hbfe449ee} /* (9, 7, 31) {real, imag} */,
  {32'hbf8c9735, 32'h3f4da56b} /* (9, 7, 30) {real, imag} */,
  {32'hbd0349c9, 32'hbdd57579} /* (9, 7, 29) {real, imag} */,
  {32'h3dc55541, 32'hbd8d00ae} /* (9, 7, 28) {real, imag} */,
  {32'hbe5e3930, 32'h3e436732} /* (9, 7, 27) {real, imag} */,
  {32'hb7a7c000, 32'h3c3f0a09} /* (9, 7, 26) {real, imag} */,
  {32'h3dca47b2, 32'h3d0af8d0} /* (9, 7, 25) {real, imag} */,
  {32'hbc819245, 32'h3d6d5eed} /* (9, 7, 24) {real, imag} */,
  {32'h3cad86a3, 32'h3d76d93c} /* (9, 7, 23) {real, imag} */,
  {32'h3d63bac5, 32'h3a46c780} /* (9, 7, 22) {real, imag} */,
  {32'hbd689952, 32'h3cca84cf} /* (9, 7, 21) {real, imag} */,
  {32'hbd0c6e9e, 32'hbd3e1232} /* (9, 7, 20) {real, imag} */,
  {32'hbd89f0eb, 32'hbcb2549a} /* (9, 7, 19) {real, imag} */,
  {32'h3d1cb390, 32'hbd266042} /* (9, 7, 18) {real, imag} */,
  {32'hbb943d26, 32'h3c9bb0cd} /* (9, 7, 17) {real, imag} */,
  {32'h3d5fa17a, 32'h00000000} /* (9, 7, 16) {real, imag} */,
  {32'hbb943d26, 32'hbc9bb0cd} /* (9, 7, 15) {real, imag} */,
  {32'h3d1cb390, 32'h3d266042} /* (9, 7, 14) {real, imag} */,
  {32'hbd89f0eb, 32'h3cb2549a} /* (9, 7, 13) {real, imag} */,
  {32'hbd0c6e9e, 32'h3d3e1232} /* (9, 7, 12) {real, imag} */,
  {32'hbd689952, 32'hbcca84cf} /* (9, 7, 11) {real, imag} */,
  {32'h3d63bac5, 32'hba46c780} /* (9, 7, 10) {real, imag} */,
  {32'h3cad86a3, 32'hbd76d93c} /* (9, 7, 9) {real, imag} */,
  {32'hbc819245, 32'hbd6d5eed} /* (9, 7, 8) {real, imag} */,
  {32'h3dca47b2, 32'hbd0af8d0} /* (9, 7, 7) {real, imag} */,
  {32'hb7a7c000, 32'hbc3f0a09} /* (9, 7, 6) {real, imag} */,
  {32'hbe5e3930, 32'hbe436732} /* (9, 7, 5) {real, imag} */,
  {32'h3dc55541, 32'h3d8d00ae} /* (9, 7, 4) {real, imag} */,
  {32'hbd0349c9, 32'h3dd57579} /* (9, 7, 3) {real, imag} */,
  {32'hbf8c9735, 32'hbf4da56b} /* (9, 7, 2) {real, imag} */,
  {32'h40564cfd, 32'h3fe449ee} /* (9, 7, 1) {real, imag} */,
  {32'h40845442, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h4062b082, 32'hc0150e2e} /* (9, 6, 31) {real, imag} */,
  {32'hbf6c602d, 32'h3f84e77d} /* (9, 6, 30) {real, imag} */,
  {32'hbcc81b89, 32'hbc474bd0} /* (9, 6, 29) {real, imag} */,
  {32'h3d3b0b1e, 32'hbdb2d53e} /* (9, 6, 28) {real, imag} */,
  {32'hbe3a53f2, 32'h3d3518b2} /* (9, 6, 27) {real, imag} */,
  {32'h3d5b1e4c, 32'h3dae7a2d} /* (9, 6, 26) {real, imag} */,
  {32'h3e06bac6, 32'h3df7ca74} /* (9, 6, 25) {real, imag} */,
  {32'h3cf1715c, 32'h3db5601f} /* (9, 6, 24) {real, imag} */,
  {32'hbd1de3ba, 32'hbc2152f1} /* (9, 6, 23) {real, imag} */,
  {32'hbc9a3c35, 32'h3d3758a0} /* (9, 6, 22) {real, imag} */,
  {32'h37acf000, 32'hbd6b3009} /* (9, 6, 21) {real, imag} */,
  {32'h3b00a1d4, 32'hbd31df62} /* (9, 6, 20) {real, imag} */,
  {32'h3caad3da, 32'hbd4f4764} /* (9, 6, 19) {real, imag} */,
  {32'h3d52dc52, 32'h3dd403d9} /* (9, 6, 18) {real, imag} */,
  {32'hbd7aa253, 32'h3d193a38} /* (9, 6, 17) {real, imag} */,
  {32'hbdbaeaf4, 32'h00000000} /* (9, 6, 16) {real, imag} */,
  {32'hbd7aa253, 32'hbd193a38} /* (9, 6, 15) {real, imag} */,
  {32'h3d52dc52, 32'hbdd403d9} /* (9, 6, 14) {real, imag} */,
  {32'h3caad3da, 32'h3d4f4764} /* (9, 6, 13) {real, imag} */,
  {32'h3b00a1d4, 32'h3d31df62} /* (9, 6, 12) {real, imag} */,
  {32'h37acf000, 32'h3d6b3009} /* (9, 6, 11) {real, imag} */,
  {32'hbc9a3c35, 32'hbd3758a0} /* (9, 6, 10) {real, imag} */,
  {32'hbd1de3ba, 32'h3c2152f1} /* (9, 6, 9) {real, imag} */,
  {32'h3cf1715c, 32'hbdb5601f} /* (9, 6, 8) {real, imag} */,
  {32'h3e06bac6, 32'hbdf7ca74} /* (9, 6, 7) {real, imag} */,
  {32'h3d5b1e4c, 32'hbdae7a2d} /* (9, 6, 6) {real, imag} */,
  {32'hbe3a53f2, 32'hbd3518b2} /* (9, 6, 5) {real, imag} */,
  {32'h3d3b0b1e, 32'h3db2d53e} /* (9, 6, 4) {real, imag} */,
  {32'hbcc81b89, 32'h3c474bd0} /* (9, 6, 3) {real, imag} */,
  {32'hbf6c602d, 32'hbf84e77d} /* (9, 6, 2) {real, imag} */,
  {32'h4062b082, 32'h40150e2e} /* (9, 6, 1) {real, imag} */,
  {32'h40960f59, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'h405ab55d, 32'hc0423622} /* (9, 5, 31) {real, imag} */,
  {32'hbebf16b0, 32'h3f9f2cf6} /* (9, 5, 30) {real, imag} */,
  {32'hbdc725ab, 32'h3c9f7c46} /* (9, 5, 29) {real, imag} */,
  {32'h3c01e020, 32'h3d335bf8} /* (9, 5, 28) {real, imag} */,
  {32'hbd6e26eb, 32'h3da3ed8d} /* (9, 5, 27) {real, imag} */,
  {32'h3dfb3226, 32'h3dad268c} /* (9, 5, 26) {real, imag} */,
  {32'h3d55bf41, 32'hbb5a6bc0} /* (9, 5, 25) {real, imag} */,
  {32'hbce4cbb7, 32'h3e00563b} /* (9, 5, 24) {real, imag} */,
  {32'hbdad3a05, 32'hbdc4d508} /* (9, 5, 23) {real, imag} */,
  {32'h3dec3cf2, 32'h3d801e58} /* (9, 5, 22) {real, imag} */,
  {32'h3d854d29, 32'hbdccf716} /* (9, 5, 21) {real, imag} */,
  {32'hbc2dd86a, 32'h3c4ce108} /* (9, 5, 20) {real, imag} */,
  {32'h3d3e7e1d, 32'h3dce61c2} /* (9, 5, 19) {real, imag} */,
  {32'hbdc5acf6, 32'h3def20f2} /* (9, 5, 18) {real, imag} */,
  {32'h3c15b5dc, 32'h3cfb4ea1} /* (9, 5, 17) {real, imag} */,
  {32'h3d02c51d, 32'h00000000} /* (9, 5, 16) {real, imag} */,
  {32'h3c15b5dc, 32'hbcfb4ea1} /* (9, 5, 15) {real, imag} */,
  {32'hbdc5acf6, 32'hbdef20f2} /* (9, 5, 14) {real, imag} */,
  {32'h3d3e7e1d, 32'hbdce61c2} /* (9, 5, 13) {real, imag} */,
  {32'hbc2dd86a, 32'hbc4ce108} /* (9, 5, 12) {real, imag} */,
  {32'h3d854d29, 32'h3dccf716} /* (9, 5, 11) {real, imag} */,
  {32'h3dec3cf2, 32'hbd801e58} /* (9, 5, 10) {real, imag} */,
  {32'hbdad3a05, 32'h3dc4d508} /* (9, 5, 9) {real, imag} */,
  {32'hbce4cbb7, 32'hbe00563b} /* (9, 5, 8) {real, imag} */,
  {32'h3d55bf41, 32'h3b5a6bc0} /* (9, 5, 7) {real, imag} */,
  {32'h3dfb3226, 32'hbdad268c} /* (9, 5, 6) {real, imag} */,
  {32'hbd6e26eb, 32'hbda3ed8d} /* (9, 5, 5) {real, imag} */,
  {32'h3c01e020, 32'hbd335bf8} /* (9, 5, 4) {real, imag} */,
  {32'hbdc725ab, 32'hbc9f7c46} /* (9, 5, 3) {real, imag} */,
  {32'hbebf16b0, 32'hbf9f2cf6} /* (9, 5, 2) {real, imag} */,
  {32'h405ab55d, 32'h40423622} /* (9, 5, 1) {real, imag} */,
  {32'h40a93d4c, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'h4055c031, 32'hc06785f7} /* (9, 4, 31) {real, imag} */,
  {32'hbc684300, 32'h3f94cf60} /* (9, 4, 30) {real, imag} */,
  {32'hbdb3a628, 32'hbd2d1e07} /* (9, 4, 29) {real, imag} */,
  {32'hbd7ff010, 32'h3e7bf1c4} /* (9, 4, 28) {real, imag} */,
  {32'hbdf82f00, 32'h3df981fd} /* (9, 4, 27) {real, imag} */,
  {32'hbc5eadf4, 32'hbd9595c4} /* (9, 4, 26) {real, imag} */,
  {32'h3e17f305, 32'hbdbac1f6} /* (9, 4, 25) {real, imag} */,
  {32'hbb810372, 32'hbb93cdea} /* (9, 4, 24) {real, imag} */,
  {32'hbce8ba76, 32'hbc649b28} /* (9, 4, 23) {real, imag} */,
  {32'h3cc6f99a, 32'h3e095548} /* (9, 4, 22) {real, imag} */,
  {32'hbd318527, 32'hbd3be2c9} /* (9, 4, 21) {real, imag} */,
  {32'h3d1aab88, 32'hbc3fc873} /* (9, 4, 20) {real, imag} */,
  {32'h3d70faa8, 32'hbda6643a} /* (9, 4, 19) {real, imag} */,
  {32'h3c9009ce, 32'hbd97856e} /* (9, 4, 18) {real, imag} */,
  {32'hbca660e6, 32'h3d374277} /* (9, 4, 17) {real, imag} */,
  {32'hbc93fedc, 32'h00000000} /* (9, 4, 16) {real, imag} */,
  {32'hbca660e6, 32'hbd374277} /* (9, 4, 15) {real, imag} */,
  {32'h3c9009ce, 32'h3d97856e} /* (9, 4, 14) {real, imag} */,
  {32'h3d70faa8, 32'h3da6643a} /* (9, 4, 13) {real, imag} */,
  {32'h3d1aab88, 32'h3c3fc873} /* (9, 4, 12) {real, imag} */,
  {32'hbd318527, 32'h3d3be2c9} /* (9, 4, 11) {real, imag} */,
  {32'h3cc6f99a, 32'hbe095548} /* (9, 4, 10) {real, imag} */,
  {32'hbce8ba76, 32'h3c649b28} /* (9, 4, 9) {real, imag} */,
  {32'hbb810372, 32'h3b93cdea} /* (9, 4, 8) {real, imag} */,
  {32'h3e17f305, 32'h3dbac1f6} /* (9, 4, 7) {real, imag} */,
  {32'hbc5eadf4, 32'h3d9595c4} /* (9, 4, 6) {real, imag} */,
  {32'hbdf82f00, 32'hbdf981fd} /* (9, 4, 5) {real, imag} */,
  {32'hbd7ff010, 32'hbe7bf1c4} /* (9, 4, 4) {real, imag} */,
  {32'hbdb3a628, 32'h3d2d1e07} /* (9, 4, 3) {real, imag} */,
  {32'hbc684300, 32'hbf94cf60} /* (9, 4, 2) {real, imag} */,
  {32'h4055c031, 32'h406785f7} /* (9, 4, 1) {real, imag} */,
  {32'h40b017fc, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'h404f4f16, 32'hc07c4646} /* (9, 3, 31) {real, imag} */,
  {32'h3e9fdaac, 32'h3f94d3fe} /* (9, 3, 30) {real, imag} */,
  {32'hbddd6987, 32'h3de0ea11} /* (9, 3, 29) {real, imag} */,
  {32'hbd831a84, 32'h3e8b0ab6} /* (9, 3, 28) {real, imag} */,
  {32'hbdc47331, 32'h3cff5061} /* (9, 3, 27) {real, imag} */,
  {32'hbd5414f7, 32'hbd80938a} /* (9, 3, 26) {real, imag} */,
  {32'h3dda9a8f, 32'h3c963374} /* (9, 3, 25) {real, imag} */,
  {32'h3c5211ab, 32'h3e35bb5c} /* (9, 3, 24) {real, imag} */,
  {32'hbd5f4b0b, 32'h3c75f3aa} /* (9, 3, 23) {real, imag} */,
  {32'h3d666fc2, 32'h3dd24c2a} /* (9, 3, 22) {real, imag} */,
  {32'hbbac11c8, 32'h3d80fec6} /* (9, 3, 21) {real, imag} */,
  {32'h3d287f36, 32'h3cfa3cf4} /* (9, 3, 20) {real, imag} */,
  {32'h3ced4479, 32'h3d814574} /* (9, 3, 19) {real, imag} */,
  {32'h3ccf821b, 32'h3cef474f} /* (9, 3, 18) {real, imag} */,
  {32'hbd946d96, 32'hbd2dd8f0} /* (9, 3, 17) {real, imag} */,
  {32'h3cf2f514, 32'h00000000} /* (9, 3, 16) {real, imag} */,
  {32'hbd946d96, 32'h3d2dd8f0} /* (9, 3, 15) {real, imag} */,
  {32'h3ccf821b, 32'hbcef474f} /* (9, 3, 14) {real, imag} */,
  {32'h3ced4479, 32'hbd814574} /* (9, 3, 13) {real, imag} */,
  {32'h3d287f36, 32'hbcfa3cf4} /* (9, 3, 12) {real, imag} */,
  {32'hbbac11c8, 32'hbd80fec6} /* (9, 3, 11) {real, imag} */,
  {32'h3d666fc2, 32'hbdd24c2a} /* (9, 3, 10) {real, imag} */,
  {32'hbd5f4b0b, 32'hbc75f3aa} /* (9, 3, 9) {real, imag} */,
  {32'h3c5211ab, 32'hbe35bb5c} /* (9, 3, 8) {real, imag} */,
  {32'h3dda9a8f, 32'hbc963374} /* (9, 3, 7) {real, imag} */,
  {32'hbd5414f7, 32'h3d80938a} /* (9, 3, 6) {real, imag} */,
  {32'hbdc47331, 32'hbcff5061} /* (9, 3, 5) {real, imag} */,
  {32'hbd831a84, 32'hbe8b0ab6} /* (9, 3, 4) {real, imag} */,
  {32'hbddd6987, 32'hbde0ea11} /* (9, 3, 3) {real, imag} */,
  {32'h3e9fdaac, 32'hbf94d3fe} /* (9, 3, 2) {real, imag} */,
  {32'h404f4f16, 32'h407c4646} /* (9, 3, 1) {real, imag} */,
  {32'h40b2f865, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'h40440347, 32'hc07b92e6} /* (9, 2, 31) {real, imag} */,
  {32'h3eb803f1, 32'h3f893b88} /* (9, 2, 30) {real, imag} */,
  {32'hbe5e44bc, 32'h3e2aa7a6} /* (9, 2, 29) {real, imag} */,
  {32'hbc9cb78c, 32'h3e971dd4} /* (9, 2, 28) {real, imag} */,
  {32'hbdb9fc36, 32'hbe56e856} /* (9, 2, 27) {real, imag} */,
  {32'hbdf845ae, 32'hbd1959d0} /* (9, 2, 26) {real, imag} */,
  {32'h3c36eeaa, 32'hbc897cc6} /* (9, 2, 25) {real, imag} */,
  {32'h3da746d9, 32'h3de9171a} /* (9, 2, 24) {real, imag} */,
  {32'hbc18ce58, 32'h3b15f2b2} /* (9, 2, 23) {real, imag} */,
  {32'hbde0d2d1, 32'h3d3f2510} /* (9, 2, 22) {real, imag} */,
  {32'hbdecaffe, 32'hbdb67f2a} /* (9, 2, 21) {real, imag} */,
  {32'h3d3885f4, 32'h3d379a7a} /* (9, 2, 20) {real, imag} */,
  {32'h3d3d7be2, 32'hbdac1ade} /* (9, 2, 19) {real, imag} */,
  {32'hbc6a9578, 32'h3cf84ce4} /* (9, 2, 18) {real, imag} */,
  {32'hbb996587, 32'h3ce05a3a} /* (9, 2, 17) {real, imag} */,
  {32'h3d20d688, 32'h00000000} /* (9, 2, 16) {real, imag} */,
  {32'hbb996587, 32'hbce05a3a} /* (9, 2, 15) {real, imag} */,
  {32'hbc6a9578, 32'hbcf84ce4} /* (9, 2, 14) {real, imag} */,
  {32'h3d3d7be2, 32'h3dac1ade} /* (9, 2, 13) {real, imag} */,
  {32'h3d3885f4, 32'hbd379a7a} /* (9, 2, 12) {real, imag} */,
  {32'hbdecaffe, 32'h3db67f2a} /* (9, 2, 11) {real, imag} */,
  {32'hbde0d2d1, 32'hbd3f2510} /* (9, 2, 10) {real, imag} */,
  {32'hbc18ce58, 32'hbb15f2b2} /* (9, 2, 9) {real, imag} */,
  {32'h3da746d9, 32'hbde9171a} /* (9, 2, 8) {real, imag} */,
  {32'h3c36eeaa, 32'h3c897cc6} /* (9, 2, 7) {real, imag} */,
  {32'hbdf845ae, 32'h3d1959d0} /* (9, 2, 6) {real, imag} */,
  {32'hbdb9fc36, 32'h3e56e856} /* (9, 2, 5) {real, imag} */,
  {32'hbc9cb78c, 32'hbe971dd4} /* (9, 2, 4) {real, imag} */,
  {32'hbe5e44bc, 32'hbe2aa7a6} /* (9, 2, 3) {real, imag} */,
  {32'h3eb803f1, 32'hbf893b88} /* (9, 2, 2) {real, imag} */,
  {32'h40440347, 32'h407b92e6} /* (9, 2, 1) {real, imag} */,
  {32'h40b61095, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'h404fb855, 32'hc06a1c71} /* (9, 1, 31) {real, imag} */,
  {32'h3e87ba5c, 32'h3f7f7470} /* (9, 1, 30) {real, imag} */,
  {32'hbe9f3bc5, 32'h3d2be16b} /* (9, 1, 29) {real, imag} */,
  {32'h3bf1e3c8, 32'h3ea60387} /* (9, 1, 28) {real, imag} */,
  {32'hbe234561, 32'hbe303336} /* (9, 1, 27) {real, imag} */,
  {32'hbcefc840, 32'h3d1ed080} /* (9, 1, 26) {real, imag} */,
  {32'h3c4d7d12, 32'h3c73f18a} /* (9, 1, 25) {real, imag} */,
  {32'h3d7f6b28, 32'h3d897cae} /* (9, 1, 24) {real, imag} */,
  {32'h3d333654, 32'hbccaba62} /* (9, 1, 23) {real, imag} */,
  {32'hbd9b90f2, 32'hbab9dba8} /* (9, 1, 22) {real, imag} */,
  {32'hbd91280c, 32'hba8b0100} /* (9, 1, 21) {real, imag} */,
  {32'h3c9c0964, 32'h3da4a1b2} /* (9, 1, 20) {real, imag} */,
  {32'h3dc1a4ae, 32'hbdb80ef8} /* (9, 1, 19) {real, imag} */,
  {32'hbd017487, 32'h3cc1a182} /* (9, 1, 18) {real, imag} */,
  {32'hbbc71a93, 32'hbd0693f4} /* (9, 1, 17) {real, imag} */,
  {32'hbcd820bf, 32'h00000000} /* (9, 1, 16) {real, imag} */,
  {32'hbbc71a93, 32'h3d0693f4} /* (9, 1, 15) {real, imag} */,
  {32'hbd017487, 32'hbcc1a182} /* (9, 1, 14) {real, imag} */,
  {32'h3dc1a4ae, 32'h3db80ef8} /* (9, 1, 13) {real, imag} */,
  {32'h3c9c0964, 32'hbda4a1b2} /* (9, 1, 12) {real, imag} */,
  {32'hbd91280c, 32'h3a8b0100} /* (9, 1, 11) {real, imag} */,
  {32'hbd9b90f2, 32'h3ab9dba8} /* (9, 1, 10) {real, imag} */,
  {32'h3d333654, 32'h3ccaba62} /* (9, 1, 9) {real, imag} */,
  {32'h3d7f6b28, 32'hbd897cae} /* (9, 1, 8) {real, imag} */,
  {32'h3c4d7d12, 32'hbc73f18a} /* (9, 1, 7) {real, imag} */,
  {32'hbcefc840, 32'hbd1ed080} /* (9, 1, 6) {real, imag} */,
  {32'hbe234561, 32'h3e303336} /* (9, 1, 5) {real, imag} */,
  {32'h3bf1e3c8, 32'hbea60387} /* (9, 1, 4) {real, imag} */,
  {32'hbe9f3bc5, 32'hbd2be16b} /* (9, 1, 3) {real, imag} */,
  {32'h3e87ba5c, 32'hbf7f7470} /* (9, 1, 2) {real, imag} */,
  {32'h404fb855, 32'h406a1c71} /* (9, 1, 1) {real, imag} */,
  {32'h40b359c9, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'h405d1b56, 32'hc03c6bd6} /* (9, 0, 31) {real, imag} */,
  {32'hbe163e04, 32'h3f57a754} /* (9, 0, 30) {real, imag} */,
  {32'hbe43f42c, 32'h3d82e6e4} /* (9, 0, 29) {real, imag} */,
  {32'h3d623904, 32'h3e134cf0} /* (9, 0, 28) {real, imag} */,
  {32'hbdde8181, 32'hbdb3078c} /* (9, 0, 27) {real, imag} */,
  {32'h3ce772b8, 32'hbcedf8c6} /* (9, 0, 26) {real, imag} */,
  {32'h3cb94da8, 32'h3b856962} /* (9, 0, 25) {real, imag} */,
  {32'hba664840, 32'hbcdf6d81} /* (9, 0, 24) {real, imag} */,
  {32'h3c1bf2e4, 32'hbd3ad7d2} /* (9, 0, 23) {real, imag} */,
  {32'hbd597e8b, 32'hbc07d0e0} /* (9, 0, 22) {real, imag} */,
  {32'hbcc73cb8, 32'h3d34c8f7} /* (9, 0, 21) {real, imag} */,
  {32'hbd0a114d, 32'h3cc4ea0f} /* (9, 0, 20) {real, imag} */,
  {32'hbd3ba99d, 32'h3d35328a} /* (9, 0, 19) {real, imag} */,
  {32'h3c6ee83d, 32'h3ce5c313} /* (9, 0, 18) {real, imag} */,
  {32'hbcb105f2, 32'hbcded6a3} /* (9, 0, 17) {real, imag} */,
  {32'h3d993aa9, 32'h00000000} /* (9, 0, 16) {real, imag} */,
  {32'hbcb105f2, 32'h3cded6a3} /* (9, 0, 15) {real, imag} */,
  {32'h3c6ee83d, 32'hbce5c313} /* (9, 0, 14) {real, imag} */,
  {32'hbd3ba99d, 32'hbd35328a} /* (9, 0, 13) {real, imag} */,
  {32'hbd0a114d, 32'hbcc4ea0f} /* (9, 0, 12) {real, imag} */,
  {32'hbcc73cb8, 32'hbd34c8f7} /* (9, 0, 11) {real, imag} */,
  {32'hbd597e8b, 32'h3c07d0e0} /* (9, 0, 10) {real, imag} */,
  {32'h3c1bf2e4, 32'h3d3ad7d2} /* (9, 0, 9) {real, imag} */,
  {32'hba664840, 32'h3cdf6d81} /* (9, 0, 8) {real, imag} */,
  {32'h3cb94da8, 32'hbb856962} /* (9, 0, 7) {real, imag} */,
  {32'h3ce772b8, 32'h3cedf8c6} /* (9, 0, 6) {real, imag} */,
  {32'hbdde8181, 32'h3db3078c} /* (9, 0, 5) {real, imag} */,
  {32'h3d623904, 32'hbe134cf0} /* (9, 0, 4) {real, imag} */,
  {32'hbe43f42c, 32'hbd82e6e4} /* (9, 0, 3) {real, imag} */,
  {32'hbe163e04, 32'hbf57a754} /* (9, 0, 2) {real, imag} */,
  {32'h405d1b56, 32'h403c6bd6} /* (9, 0, 1) {real, imag} */,
  {32'h40a8b349, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h4062e33d, 32'hbffb271c} /* (8, 31, 31) {real, imag} */,
  {32'hbf3667ba, 32'h3f0b375e} /* (8, 31, 30) {real, imag} */,
  {32'hbd37a3d2, 32'hbcfb6b58} /* (8, 31, 29) {real, imag} */,
  {32'h3cb90f2e, 32'h3dc57365} /* (8, 31, 28) {real, imag} */,
  {32'hbe03a102, 32'h3b45dea0} /* (8, 31, 27) {real, imag} */,
  {32'h3be687ec, 32'hb98a67c0} /* (8, 31, 26) {real, imag} */,
  {32'h3d7baa56, 32'hb9e9c680} /* (8, 31, 25) {real, imag} */,
  {32'hbdc699a0, 32'h3cb8d2eb} /* (8, 31, 24) {real, imag} */,
  {32'h3d94bc9e, 32'hbc5de536} /* (8, 31, 23) {real, imag} */,
  {32'h3dba5c88, 32'h3c5acaa4} /* (8, 31, 22) {real, imag} */,
  {32'hbd5094f3, 32'h3d8f8234} /* (8, 31, 21) {real, imag} */,
  {32'hbd38766b, 32'hbd3ae02e} /* (8, 31, 20) {real, imag} */,
  {32'h3d581694, 32'hbd09cc5c} /* (8, 31, 19) {real, imag} */,
  {32'hbd2ac209, 32'h3d10e7d9} /* (8, 31, 18) {real, imag} */,
  {32'hbce21969, 32'hbd81f6d5} /* (8, 31, 17) {real, imag} */,
  {32'h3d3e4c6f, 32'h00000000} /* (8, 31, 16) {real, imag} */,
  {32'hbce21969, 32'h3d81f6d5} /* (8, 31, 15) {real, imag} */,
  {32'hbd2ac209, 32'hbd10e7d9} /* (8, 31, 14) {real, imag} */,
  {32'h3d581694, 32'h3d09cc5c} /* (8, 31, 13) {real, imag} */,
  {32'hbd38766b, 32'h3d3ae02e} /* (8, 31, 12) {real, imag} */,
  {32'hbd5094f3, 32'hbd8f8234} /* (8, 31, 11) {real, imag} */,
  {32'h3dba5c88, 32'hbc5acaa4} /* (8, 31, 10) {real, imag} */,
  {32'h3d94bc9e, 32'h3c5de536} /* (8, 31, 9) {real, imag} */,
  {32'hbdc699a0, 32'hbcb8d2eb} /* (8, 31, 8) {real, imag} */,
  {32'h3d7baa56, 32'h39e9c680} /* (8, 31, 7) {real, imag} */,
  {32'h3be687ec, 32'h398a67c0} /* (8, 31, 6) {real, imag} */,
  {32'hbe03a102, 32'hbb45dea0} /* (8, 31, 5) {real, imag} */,
  {32'h3cb90f2e, 32'hbdc57365} /* (8, 31, 4) {real, imag} */,
  {32'hbd37a3d2, 32'h3cfb6b58} /* (8, 31, 3) {real, imag} */,
  {32'hbf3667ba, 32'hbf0b375e} /* (8, 31, 2) {real, imag} */,
  {32'h4062e33d, 32'h3ffb271c} /* (8, 31, 1) {real, imag} */,
  {32'h40a28aaf, 32'h00000000} /* (8, 31, 0) {real, imag} */,
  {32'h4082e612, 32'hbfc58433} /* (8, 30, 31) {real, imag} */,
  {32'hbf88f4f1, 32'h3f03e919} /* (8, 30, 30) {real, imag} */,
  {32'h3aa73080, 32'h3d2c57f6} /* (8, 30, 29) {real, imag} */,
  {32'h3d491036, 32'h3b7c5680} /* (8, 30, 28) {real, imag} */,
  {32'hbe2a107a, 32'h3d994a9a} /* (8, 30, 27) {real, imag} */,
  {32'h3dd608e8, 32'h3cc813c5} /* (8, 30, 26) {real, imag} */,
  {32'h3d9ddf37, 32'hbc85a42e} /* (8, 30, 25) {real, imag} */,
  {32'hbdb81ea0, 32'h3e242dfc} /* (8, 30, 24) {real, imag} */,
  {32'h3d9090aa, 32'hbcded204} /* (8, 30, 23) {real, imag} */,
  {32'hbe03626a, 32'h3b348a00} /* (8, 30, 22) {real, imag} */,
  {32'hbe1da687, 32'h3d50b30c} /* (8, 30, 21) {real, imag} */,
  {32'hbd5266d0, 32'hbc4a75cc} /* (8, 30, 20) {real, imag} */,
  {32'h3daa3318, 32'h3be15f00} /* (8, 30, 19) {real, imag} */,
  {32'hbd6ae84e, 32'h3d9db482} /* (8, 30, 18) {real, imag} */,
  {32'hbd0ac3c9, 32'hbb679340} /* (8, 30, 17) {real, imag} */,
  {32'hbca8afa8, 32'h00000000} /* (8, 30, 16) {real, imag} */,
  {32'hbd0ac3c9, 32'h3b679340} /* (8, 30, 15) {real, imag} */,
  {32'hbd6ae84e, 32'hbd9db482} /* (8, 30, 14) {real, imag} */,
  {32'h3daa3318, 32'hbbe15f00} /* (8, 30, 13) {real, imag} */,
  {32'hbd5266d0, 32'h3c4a75cc} /* (8, 30, 12) {real, imag} */,
  {32'hbe1da687, 32'hbd50b30c} /* (8, 30, 11) {real, imag} */,
  {32'hbe03626a, 32'hbb348a00} /* (8, 30, 10) {real, imag} */,
  {32'h3d9090aa, 32'h3cded204} /* (8, 30, 9) {real, imag} */,
  {32'hbdb81ea0, 32'hbe242dfc} /* (8, 30, 8) {real, imag} */,
  {32'h3d9ddf37, 32'h3c85a42e} /* (8, 30, 7) {real, imag} */,
  {32'h3dd608e8, 32'hbcc813c5} /* (8, 30, 6) {real, imag} */,
  {32'hbe2a107a, 32'hbd994a9a} /* (8, 30, 5) {real, imag} */,
  {32'h3d491036, 32'hbb7c5680} /* (8, 30, 4) {real, imag} */,
  {32'h3aa73080, 32'hbd2c57f6} /* (8, 30, 3) {real, imag} */,
  {32'hbf88f4f1, 32'hbf03e919} /* (8, 30, 2) {real, imag} */,
  {32'h4082e612, 32'h3fc58433} /* (8, 30, 1) {real, imag} */,
  {32'h40a839b4, 32'h00000000} /* (8, 30, 0) {real, imag} */,
  {32'h408d906c, 32'hbf93c068} /* (8, 29, 31) {real, imag} */,
  {32'hbf9012aa, 32'h3f028db4} /* (8, 29, 30) {real, imag} */,
  {32'h3dcf5cd2, 32'h3da3ab9c} /* (8, 29, 29) {real, imag} */,
  {32'h3e472fce, 32'hbd685edc} /* (8, 29, 28) {real, imag} */,
  {32'hbe7033c6, 32'h3da73851} /* (8, 29, 27) {real, imag} */,
  {32'h3cca5b3c, 32'hba3e5e00} /* (8, 29, 26) {real, imag} */,
  {32'h3c9b9c30, 32'hbdb569d1} /* (8, 29, 25) {real, imag} */,
  {32'hbde2d9fb, 32'h3d9d1f3a} /* (8, 29, 24) {real, imag} */,
  {32'hbd17088d, 32'h3cf0026a} /* (8, 29, 23) {real, imag} */,
  {32'hbd5beb76, 32'hbc984a82} /* (8, 29, 22) {real, imag} */,
  {32'hbe060289, 32'h3d4113ee} /* (8, 29, 21) {real, imag} */,
  {32'hbb89e7a0, 32'h3c327023} /* (8, 29, 20) {real, imag} */,
  {32'hbbcf79f0, 32'hbd1410b1} /* (8, 29, 19) {real, imag} */,
  {32'hbcf45e70, 32'h3de0a1de} /* (8, 29, 18) {real, imag} */,
  {32'hbc710870, 32'hbd0a2d3d} /* (8, 29, 17) {real, imag} */,
  {32'hbc9444a8, 32'h00000000} /* (8, 29, 16) {real, imag} */,
  {32'hbc710870, 32'h3d0a2d3d} /* (8, 29, 15) {real, imag} */,
  {32'hbcf45e70, 32'hbde0a1de} /* (8, 29, 14) {real, imag} */,
  {32'hbbcf79f0, 32'h3d1410b1} /* (8, 29, 13) {real, imag} */,
  {32'hbb89e7a0, 32'hbc327023} /* (8, 29, 12) {real, imag} */,
  {32'hbe060289, 32'hbd4113ee} /* (8, 29, 11) {real, imag} */,
  {32'hbd5beb76, 32'h3c984a82} /* (8, 29, 10) {real, imag} */,
  {32'hbd17088d, 32'hbcf0026a} /* (8, 29, 9) {real, imag} */,
  {32'hbde2d9fb, 32'hbd9d1f3a} /* (8, 29, 8) {real, imag} */,
  {32'h3c9b9c30, 32'h3db569d1} /* (8, 29, 7) {real, imag} */,
  {32'h3cca5b3c, 32'h3a3e5e00} /* (8, 29, 6) {real, imag} */,
  {32'hbe7033c6, 32'hbda73851} /* (8, 29, 5) {real, imag} */,
  {32'h3e472fce, 32'h3d685edc} /* (8, 29, 4) {real, imag} */,
  {32'h3dcf5cd2, 32'hbda3ab9c} /* (8, 29, 3) {real, imag} */,
  {32'hbf9012aa, 32'hbf028db4} /* (8, 29, 2) {real, imag} */,
  {32'h408d906c, 32'h3f93c068} /* (8, 29, 1) {real, imag} */,
  {32'h40a1f8d5, 32'h00000000} /* (8, 29, 0) {real, imag} */,
  {32'h408f57ae, 32'hbf7a587e} /* (8, 28, 31) {real, imag} */,
  {32'hbfabf274, 32'h3f149a39} /* (8, 28, 30) {real, imag} */,
  {32'h3bd99c80, 32'hbb9f6960} /* (8, 28, 29) {real, imag} */,
  {32'h3e5bad6c, 32'hb95af000} /* (8, 28, 28) {real, imag} */,
  {32'hbe687df2, 32'h3c09b428} /* (8, 28, 27) {real, imag} */,
  {32'hbd44a29c, 32'hbd696e54} /* (8, 28, 26) {real, imag} */,
  {32'hbd90b664, 32'hbe06073f} /* (8, 28, 25) {real, imag} */,
  {32'hbd50ddb6, 32'h3da89302} /* (8, 28, 24) {real, imag} */,
  {32'hbd9db5a2, 32'h3d96d644} /* (8, 28, 23) {real, imag} */,
  {32'hbcf8e43e, 32'hbceed1f8} /* (8, 28, 22) {real, imag} */,
  {32'h3c60ad34, 32'h3c5dc080} /* (8, 28, 21) {real, imag} */,
  {32'hbd2565c7, 32'hbcf0b88c} /* (8, 28, 20) {real, imag} */,
  {32'h3d3775fa, 32'h3a41baa0} /* (8, 28, 19) {real, imag} */,
  {32'hbd0b8600, 32'h3cd401d4} /* (8, 28, 18) {real, imag} */,
  {32'h3dd1f7fe, 32'hbdf95b36} /* (8, 28, 17) {real, imag} */,
  {32'h3d7f3cb4, 32'h00000000} /* (8, 28, 16) {real, imag} */,
  {32'h3dd1f7fe, 32'h3df95b36} /* (8, 28, 15) {real, imag} */,
  {32'hbd0b8600, 32'hbcd401d4} /* (8, 28, 14) {real, imag} */,
  {32'h3d3775fa, 32'hba41baa0} /* (8, 28, 13) {real, imag} */,
  {32'hbd2565c7, 32'h3cf0b88c} /* (8, 28, 12) {real, imag} */,
  {32'h3c60ad34, 32'hbc5dc080} /* (8, 28, 11) {real, imag} */,
  {32'hbcf8e43e, 32'h3ceed1f8} /* (8, 28, 10) {real, imag} */,
  {32'hbd9db5a2, 32'hbd96d644} /* (8, 28, 9) {real, imag} */,
  {32'hbd50ddb6, 32'hbda89302} /* (8, 28, 8) {real, imag} */,
  {32'hbd90b664, 32'h3e06073f} /* (8, 28, 7) {real, imag} */,
  {32'hbd44a29c, 32'h3d696e54} /* (8, 28, 6) {real, imag} */,
  {32'hbe687df2, 32'hbc09b428} /* (8, 28, 5) {real, imag} */,
  {32'h3e5bad6c, 32'h395af000} /* (8, 28, 4) {real, imag} */,
  {32'h3bd99c80, 32'h3b9f6960} /* (8, 28, 3) {real, imag} */,
  {32'hbfabf274, 32'hbf149a39} /* (8, 28, 2) {real, imag} */,
  {32'h408f57ae, 32'h3f7a587e} /* (8, 28, 1) {real, imag} */,
  {32'h409dec2e, 32'h00000000} /* (8, 28, 0) {real, imag} */,
  {32'h40926426, 32'hbf43dd94} /* (8, 27, 31) {real, imag} */,
  {32'hbfcb6a58, 32'h3eef2ebd} /* (8, 27, 30) {real, imag} */,
  {32'h3ddab9de, 32'h3a9ec760} /* (8, 27, 29) {real, imag} */,
  {32'h3e21aeb5, 32'hbd44ce2a} /* (8, 27, 28) {real, imag} */,
  {32'hbe1aa9e8, 32'h3cc18861} /* (8, 27, 27) {real, imag} */,
  {32'hbd28affa, 32'hbde193d8} /* (8, 27, 26) {real, imag} */,
  {32'h3dbac754, 32'hbda941cc} /* (8, 27, 25) {real, imag} */,
  {32'h3dc181d6, 32'h3ca34e02} /* (8, 27, 24) {real, imag} */,
  {32'h3c50b5b1, 32'h3d5f1546} /* (8, 27, 23) {real, imag} */,
  {32'hbb2c4d20, 32'h3dd0277e} /* (8, 27, 22) {real, imag} */,
  {32'hbace3380, 32'h3d7e1b1c} /* (8, 27, 21) {real, imag} */,
  {32'hbdd56215, 32'hbde34ea8} /* (8, 27, 20) {real, imag} */,
  {32'hbdefafc3, 32'h3d745136} /* (8, 27, 19) {real, imag} */,
  {32'h3dad3704, 32'h3cd9d4c4} /* (8, 27, 18) {real, imag} */,
  {32'h3d6cd9a8, 32'h3c2d8d80} /* (8, 27, 17) {real, imag} */,
  {32'h3d0f557c, 32'h00000000} /* (8, 27, 16) {real, imag} */,
  {32'h3d6cd9a8, 32'hbc2d8d80} /* (8, 27, 15) {real, imag} */,
  {32'h3dad3704, 32'hbcd9d4c4} /* (8, 27, 14) {real, imag} */,
  {32'hbdefafc3, 32'hbd745136} /* (8, 27, 13) {real, imag} */,
  {32'hbdd56215, 32'h3de34ea8} /* (8, 27, 12) {real, imag} */,
  {32'hbace3380, 32'hbd7e1b1c} /* (8, 27, 11) {real, imag} */,
  {32'hbb2c4d20, 32'hbdd0277e} /* (8, 27, 10) {real, imag} */,
  {32'h3c50b5b1, 32'hbd5f1546} /* (8, 27, 9) {real, imag} */,
  {32'h3dc181d6, 32'hbca34e02} /* (8, 27, 8) {real, imag} */,
  {32'h3dbac754, 32'h3da941cc} /* (8, 27, 7) {real, imag} */,
  {32'hbd28affa, 32'h3de193d8} /* (8, 27, 6) {real, imag} */,
  {32'hbe1aa9e8, 32'hbcc18861} /* (8, 27, 5) {real, imag} */,
  {32'h3e21aeb5, 32'h3d44ce2a} /* (8, 27, 4) {real, imag} */,
  {32'h3ddab9de, 32'hba9ec760} /* (8, 27, 3) {real, imag} */,
  {32'hbfcb6a58, 32'hbeef2ebd} /* (8, 27, 2) {real, imag} */,
  {32'h40926426, 32'h3f43dd94} /* (8, 27, 1) {real, imag} */,
  {32'h409f0b34, 32'h00000000} /* (8, 27, 0) {real, imag} */,
  {32'h408e900d, 32'hbf133d16} /* (8, 26, 31) {real, imag} */,
  {32'hbfce6715, 32'h3e9d6402} /* (8, 26, 30) {real, imag} */,
  {32'h3ac35770, 32'hbce862d7} /* (8, 26, 29) {real, imag} */,
  {32'h3e7108c8, 32'h3cb71eee} /* (8, 26, 28) {real, imag} */,
  {32'hbe2a3011, 32'h3d466871} /* (8, 26, 27) {real, imag} */,
  {32'hbd369201, 32'hbcfea270} /* (8, 26, 26) {real, imag} */,
  {32'h3cb06d1c, 32'hbde2e991} /* (8, 26, 25) {real, imag} */,
  {32'h3d7d9324, 32'h3d3341e9} /* (8, 26, 24) {real, imag} */,
  {32'h3c322cc9, 32'h3da9e579} /* (8, 26, 23) {real, imag} */,
  {32'h3d44881e, 32'hbc930950} /* (8, 26, 22) {real, imag} */,
  {32'hbd9293ae, 32'h3c59b358} /* (8, 26, 21) {real, imag} */,
  {32'hbe20668e, 32'hbd8ea0d0} /* (8, 26, 20) {real, imag} */,
  {32'hbd172654, 32'hbd0cb08a} /* (8, 26, 19) {real, imag} */,
  {32'hbbecf8f2, 32'h3ca6966e} /* (8, 26, 18) {real, imag} */,
  {32'hbbf59810, 32'hbd2f8614} /* (8, 26, 17) {real, imag} */,
  {32'h3d128d78, 32'h00000000} /* (8, 26, 16) {real, imag} */,
  {32'hbbf59810, 32'h3d2f8614} /* (8, 26, 15) {real, imag} */,
  {32'hbbecf8f2, 32'hbca6966e} /* (8, 26, 14) {real, imag} */,
  {32'hbd172654, 32'h3d0cb08a} /* (8, 26, 13) {real, imag} */,
  {32'hbe20668e, 32'h3d8ea0d0} /* (8, 26, 12) {real, imag} */,
  {32'hbd9293ae, 32'hbc59b358} /* (8, 26, 11) {real, imag} */,
  {32'h3d44881e, 32'h3c930950} /* (8, 26, 10) {real, imag} */,
  {32'h3c322cc9, 32'hbda9e579} /* (8, 26, 9) {real, imag} */,
  {32'h3d7d9324, 32'hbd3341e9} /* (8, 26, 8) {real, imag} */,
  {32'h3cb06d1c, 32'h3de2e991} /* (8, 26, 7) {real, imag} */,
  {32'hbd369201, 32'h3cfea270} /* (8, 26, 6) {real, imag} */,
  {32'hbe2a3011, 32'hbd466871} /* (8, 26, 5) {real, imag} */,
  {32'h3e7108c8, 32'hbcb71eee} /* (8, 26, 4) {real, imag} */,
  {32'h3ac35770, 32'h3ce862d7} /* (8, 26, 3) {real, imag} */,
  {32'hbfce6715, 32'hbe9d6402} /* (8, 26, 2) {real, imag} */,
  {32'h408e900d, 32'h3f133d16} /* (8, 26, 1) {real, imag} */,
  {32'h40963245, 32'h00000000} /* (8, 26, 0) {real, imag} */,
  {32'h4083c709, 32'hbeef5d8c} /* (8, 25, 31) {real, imag} */,
  {32'hbfbc878c, 32'h3e75822e} /* (8, 25, 30) {real, imag} */,
  {32'hbd7d9ad1, 32'hbd8f8c47} /* (8, 25, 29) {real, imag} */,
  {32'h3e564962, 32'hbba6bcd0} /* (8, 25, 28) {real, imag} */,
  {32'hbe699dc4, 32'hbc057c30} /* (8, 25, 27) {real, imag} */,
  {32'h3d2fa309, 32'h3cbff562} /* (8, 25, 26) {real, imag} */,
  {32'hbc6ab85c, 32'hbdb8861e} /* (8, 25, 25) {real, imag} */,
  {32'h3d99ab00, 32'h3d90883c} /* (8, 25, 24) {real, imag} */,
  {32'h3cba017c, 32'h3d635a5a} /* (8, 25, 23) {real, imag} */,
  {32'hbc7ad758, 32'h3be05556} /* (8, 25, 22) {real, imag} */,
  {32'hbd823736, 32'h3d969b11} /* (8, 25, 21) {real, imag} */,
  {32'hbd900dea, 32'hbbfe9368} /* (8, 25, 20) {real, imag} */,
  {32'h3d3de1aa, 32'hbcb44361} /* (8, 25, 19) {real, imag} */,
  {32'h3d6397f8, 32'h3cef4196} /* (8, 25, 18) {real, imag} */,
  {32'h3a133840, 32'h3c6c3efa} /* (8, 25, 17) {real, imag} */,
  {32'hbc151663, 32'h00000000} /* (8, 25, 16) {real, imag} */,
  {32'h3a133840, 32'hbc6c3efa} /* (8, 25, 15) {real, imag} */,
  {32'h3d6397f8, 32'hbcef4196} /* (8, 25, 14) {real, imag} */,
  {32'h3d3de1aa, 32'h3cb44361} /* (8, 25, 13) {real, imag} */,
  {32'hbd900dea, 32'h3bfe9368} /* (8, 25, 12) {real, imag} */,
  {32'hbd823736, 32'hbd969b11} /* (8, 25, 11) {real, imag} */,
  {32'hbc7ad758, 32'hbbe05556} /* (8, 25, 10) {real, imag} */,
  {32'h3cba017c, 32'hbd635a5a} /* (8, 25, 9) {real, imag} */,
  {32'h3d99ab00, 32'hbd90883c} /* (8, 25, 8) {real, imag} */,
  {32'hbc6ab85c, 32'h3db8861e} /* (8, 25, 7) {real, imag} */,
  {32'h3d2fa309, 32'hbcbff562} /* (8, 25, 6) {real, imag} */,
  {32'hbe699dc4, 32'h3c057c30} /* (8, 25, 5) {real, imag} */,
  {32'h3e564962, 32'h3ba6bcd0} /* (8, 25, 4) {real, imag} */,
  {32'hbd7d9ad1, 32'h3d8f8c47} /* (8, 25, 3) {real, imag} */,
  {32'hbfbc878c, 32'hbe75822e} /* (8, 25, 2) {real, imag} */,
  {32'h4083c709, 32'h3eef5d8c} /* (8, 25, 1) {real, imag} */,
  {32'h40897753, 32'h00000000} /* (8, 25, 0) {real, imag} */,
  {32'h406d9426, 32'hbec3ce30} /* (8, 24, 31) {real, imag} */,
  {32'hbfb7431a, 32'h3e22aa0a} /* (8, 24, 30) {real, imag} */,
  {32'hbdc3779d, 32'hbd91a886} /* (8, 24, 29) {real, imag} */,
  {32'h3e101ed8, 32'h3d861a28} /* (8, 24, 28) {real, imag} */,
  {32'hbe62aa3a, 32'h3ddf470a} /* (8, 24, 27) {real, imag} */,
  {32'h3e20199c, 32'h3ce4be22} /* (8, 24, 26) {real, imag} */,
  {32'hbcd5d98a, 32'hbd8445f8} /* (8, 24, 25) {real, imag} */,
  {32'hbd12654b, 32'h3dcdb43e} /* (8, 24, 24) {real, imag} */,
  {32'h3cdf0b14, 32'hbdc3e2ff} /* (8, 24, 23) {real, imag} */,
  {32'h3be21b00, 32'h3d1ac8b2} /* (8, 24, 22) {real, imag} */,
  {32'hbd9c8a2b, 32'h3d236375} /* (8, 24, 21) {real, imag} */,
  {32'hbda91fba, 32'h3d93f1ff} /* (8, 24, 20) {real, imag} */,
  {32'hbdb0074c, 32'h3d787344} /* (8, 24, 19) {real, imag} */,
  {32'hbbeb1ba0, 32'h3c6e0586} /* (8, 24, 18) {real, imag} */,
  {32'hbd6c0b18, 32'h3d4eaed7} /* (8, 24, 17) {real, imag} */,
  {32'h3df380fb, 32'h00000000} /* (8, 24, 16) {real, imag} */,
  {32'hbd6c0b18, 32'hbd4eaed7} /* (8, 24, 15) {real, imag} */,
  {32'hbbeb1ba0, 32'hbc6e0586} /* (8, 24, 14) {real, imag} */,
  {32'hbdb0074c, 32'hbd787344} /* (8, 24, 13) {real, imag} */,
  {32'hbda91fba, 32'hbd93f1ff} /* (8, 24, 12) {real, imag} */,
  {32'hbd9c8a2b, 32'hbd236375} /* (8, 24, 11) {real, imag} */,
  {32'h3be21b00, 32'hbd1ac8b2} /* (8, 24, 10) {real, imag} */,
  {32'h3cdf0b14, 32'h3dc3e2ff} /* (8, 24, 9) {real, imag} */,
  {32'hbd12654b, 32'hbdcdb43e} /* (8, 24, 8) {real, imag} */,
  {32'hbcd5d98a, 32'h3d8445f8} /* (8, 24, 7) {real, imag} */,
  {32'h3e20199c, 32'hbce4be22} /* (8, 24, 6) {real, imag} */,
  {32'hbe62aa3a, 32'hbddf470a} /* (8, 24, 5) {real, imag} */,
  {32'h3e101ed8, 32'hbd861a28} /* (8, 24, 4) {real, imag} */,
  {32'hbdc3779d, 32'h3d91a886} /* (8, 24, 3) {real, imag} */,
  {32'hbfb7431a, 32'hbe22aa0a} /* (8, 24, 2) {real, imag} */,
  {32'h406d9426, 32'h3ec3ce30} /* (8, 24, 1) {real, imag} */,
  {32'h407d9060, 32'h00000000} /* (8, 24, 0) {real, imag} */,
  {32'h403f86a7, 32'hbe9a5e50} /* (8, 23, 31) {real, imag} */,
  {32'hbf965d1b, 32'h3e536c6a} /* (8, 23, 30) {real, imag} */,
  {32'hbe3d6b04, 32'hbe4f408f} /* (8, 23, 29) {real, imag} */,
  {32'h3e23f0a0, 32'hbd266b3e} /* (8, 23, 28) {real, imag} */,
  {32'hbeaeab77, 32'h3db3c34e} /* (8, 23, 27) {real, imag} */,
  {32'hbbd40878, 32'hba87c2a8} /* (8, 23, 26) {real, imag} */,
  {32'hbd018419, 32'hbd728cf9} /* (8, 23, 25) {real, imag} */,
  {32'hbdca7b9f, 32'h3cd813ca} /* (8, 23, 24) {real, imag} */,
  {32'h3c5ac8ee, 32'hbd1e6d9f} /* (8, 23, 23) {real, imag} */,
  {32'hbd79f0c2, 32'hbcaf3978} /* (8, 23, 22) {real, imag} */,
  {32'hbb06d3c0, 32'h3d423347} /* (8, 23, 21) {real, imag} */,
  {32'hbda21edc, 32'h3c2efd8e} /* (8, 23, 20) {real, imag} */,
  {32'hbba584e4, 32'hbd2c3626} /* (8, 23, 19) {real, imag} */,
  {32'h3dec5c23, 32'h3d3725e1} /* (8, 23, 18) {real, imag} */,
  {32'h3d4b559e, 32'h3dbcffb6} /* (8, 23, 17) {real, imag} */,
  {32'hbd493156, 32'h00000000} /* (8, 23, 16) {real, imag} */,
  {32'h3d4b559e, 32'hbdbcffb6} /* (8, 23, 15) {real, imag} */,
  {32'h3dec5c23, 32'hbd3725e1} /* (8, 23, 14) {real, imag} */,
  {32'hbba584e4, 32'h3d2c3626} /* (8, 23, 13) {real, imag} */,
  {32'hbda21edc, 32'hbc2efd8e} /* (8, 23, 12) {real, imag} */,
  {32'hbb06d3c0, 32'hbd423347} /* (8, 23, 11) {real, imag} */,
  {32'hbd79f0c2, 32'h3caf3978} /* (8, 23, 10) {real, imag} */,
  {32'h3c5ac8ee, 32'h3d1e6d9f} /* (8, 23, 9) {real, imag} */,
  {32'hbdca7b9f, 32'hbcd813ca} /* (8, 23, 8) {real, imag} */,
  {32'hbd018419, 32'h3d728cf9} /* (8, 23, 7) {real, imag} */,
  {32'hbbd40878, 32'h3a87c2a8} /* (8, 23, 6) {real, imag} */,
  {32'hbeaeab77, 32'hbdb3c34e} /* (8, 23, 5) {real, imag} */,
  {32'h3e23f0a0, 32'h3d266b3e} /* (8, 23, 4) {real, imag} */,
  {32'hbe3d6b04, 32'h3e4f408f} /* (8, 23, 3) {real, imag} */,
  {32'hbf965d1b, 32'hbe536c6a} /* (8, 23, 2) {real, imag} */,
  {32'h403f86a7, 32'h3e9a5e50} /* (8, 23, 1) {real, imag} */,
  {32'h405029f0, 32'h00000000} /* (8, 23, 0) {real, imag} */,
  {32'h3ff2dfe7, 32'hbe8a0bee} /* (8, 22, 31) {real, imag} */,
  {32'hbf5dce94, 32'h3e0a52dc} /* (8, 22, 30) {real, imag} */,
  {32'hbd228a52, 32'hbd6e7806} /* (8, 22, 29) {real, imag} */,
  {32'h3dd44344, 32'hbd86a816} /* (8, 22, 28) {real, imag} */,
  {32'hbe88edec, 32'h3d5a2813} /* (8, 22, 27) {real, imag} */,
  {32'h3ba59012, 32'hbc130f04} /* (8, 22, 26) {real, imag} */,
  {32'hbda83cb9, 32'h3d090a9d} /* (8, 22, 25) {real, imag} */,
  {32'hbdb6871a, 32'h3d209efc} /* (8, 22, 24) {real, imag} */,
  {32'hbc99e9dd, 32'hbc9a9dfd} /* (8, 22, 23) {real, imag} */,
  {32'h3daa5720, 32'h3d729757} /* (8, 22, 22) {real, imag} */,
  {32'h3d432115, 32'h3dc4e3d3} /* (8, 22, 21) {real, imag} */,
  {32'h3d34050a, 32'hbe12a789} /* (8, 22, 20) {real, imag} */,
  {32'h3da07604, 32'hbcb5853e} /* (8, 22, 19) {real, imag} */,
  {32'hbc967d2a, 32'h3ceb2d66} /* (8, 22, 18) {real, imag} */,
  {32'hbd907f48, 32'h38f29600} /* (8, 22, 17) {real, imag} */,
  {32'hbdb94f5a, 32'h00000000} /* (8, 22, 16) {real, imag} */,
  {32'hbd907f48, 32'hb8f29600} /* (8, 22, 15) {real, imag} */,
  {32'hbc967d2a, 32'hbceb2d66} /* (8, 22, 14) {real, imag} */,
  {32'h3da07604, 32'h3cb5853e} /* (8, 22, 13) {real, imag} */,
  {32'h3d34050a, 32'h3e12a789} /* (8, 22, 12) {real, imag} */,
  {32'h3d432115, 32'hbdc4e3d3} /* (8, 22, 11) {real, imag} */,
  {32'h3daa5720, 32'hbd729757} /* (8, 22, 10) {real, imag} */,
  {32'hbc99e9dd, 32'h3c9a9dfd} /* (8, 22, 9) {real, imag} */,
  {32'hbdb6871a, 32'hbd209efc} /* (8, 22, 8) {real, imag} */,
  {32'hbda83cb9, 32'hbd090a9d} /* (8, 22, 7) {real, imag} */,
  {32'h3ba59012, 32'h3c130f04} /* (8, 22, 6) {real, imag} */,
  {32'hbe88edec, 32'hbd5a2813} /* (8, 22, 5) {real, imag} */,
  {32'h3dd44344, 32'h3d86a816} /* (8, 22, 4) {real, imag} */,
  {32'hbd228a52, 32'h3d6e7806} /* (8, 22, 3) {real, imag} */,
  {32'hbf5dce94, 32'hbe0a52dc} /* (8, 22, 2) {real, imag} */,
  {32'h3ff2dfe7, 32'h3e8a0bee} /* (8, 22, 1) {real, imag} */,
  {32'h401792bc, 32'h00000000} /* (8, 22, 0) {real, imag} */,
  {32'h3f05f0de, 32'hbd86b03c} /* (8, 21, 31) {real, imag} */,
  {32'hbe81fd60, 32'hbdd929df} /* (8, 21, 30) {real, imag} */,
  {32'h3c9b3e60, 32'hbae14ca0} /* (8, 21, 29) {real, imag} */,
  {32'hbcf1efc8, 32'hbca25594} /* (8, 21, 28) {real, imag} */,
  {32'hbdfb794d, 32'h3ce617c9} /* (8, 21, 27) {real, imag} */,
  {32'h3c93478b, 32'hbce65904} /* (8, 21, 26) {real, imag} */,
  {32'hbdb940aa, 32'hbcdfb664} /* (8, 21, 25) {real, imag} */,
  {32'hbc4184c0, 32'h3d251674} /* (8, 21, 24) {real, imag} */,
  {32'hbcb70b0c, 32'hbd7f0e8e} /* (8, 21, 23) {real, imag} */,
  {32'hbbe7ba70, 32'hbd25104b} /* (8, 21, 22) {real, imag} */,
  {32'h3d2343c4, 32'h3dabde5a} /* (8, 21, 21) {real, imag} */,
  {32'hbd524248, 32'hbd09f6d6} /* (8, 21, 20) {real, imag} */,
  {32'h3d66f966, 32'h3dded1c0} /* (8, 21, 19) {real, imag} */,
  {32'hbd67093e, 32'h3cb69c24} /* (8, 21, 18) {real, imag} */,
  {32'hbd68c700, 32'h3a8e9600} /* (8, 21, 17) {real, imag} */,
  {32'hbd82930a, 32'h00000000} /* (8, 21, 16) {real, imag} */,
  {32'hbd68c700, 32'hba8e9600} /* (8, 21, 15) {real, imag} */,
  {32'hbd67093e, 32'hbcb69c24} /* (8, 21, 14) {real, imag} */,
  {32'h3d66f966, 32'hbdded1c0} /* (8, 21, 13) {real, imag} */,
  {32'hbd524248, 32'h3d09f6d6} /* (8, 21, 12) {real, imag} */,
  {32'h3d2343c4, 32'hbdabde5a} /* (8, 21, 11) {real, imag} */,
  {32'hbbe7ba70, 32'h3d25104b} /* (8, 21, 10) {real, imag} */,
  {32'hbcb70b0c, 32'h3d7f0e8e} /* (8, 21, 9) {real, imag} */,
  {32'hbc4184c0, 32'hbd251674} /* (8, 21, 8) {real, imag} */,
  {32'hbdb940aa, 32'h3cdfb664} /* (8, 21, 7) {real, imag} */,
  {32'h3c93478b, 32'h3ce65904} /* (8, 21, 6) {real, imag} */,
  {32'hbdfb794d, 32'hbce617c9} /* (8, 21, 5) {real, imag} */,
  {32'hbcf1efc8, 32'h3ca25594} /* (8, 21, 4) {real, imag} */,
  {32'h3c9b3e60, 32'h3ae14ca0} /* (8, 21, 3) {real, imag} */,
  {32'hbe81fd60, 32'h3dd929df} /* (8, 21, 2) {real, imag} */,
  {32'h3f05f0de, 32'h3d86b03c} /* (8, 21, 1) {real, imag} */,
  {32'h3f7ab9b4, 32'h00000000} /* (8, 21, 0) {real, imag} */,
  {32'hbfa34c60, 32'h3caffb80} /* (8, 20, 31) {real, imag} */,
  {32'h3f0eea07, 32'hbe945a7a} /* (8, 20, 30) {real, imag} */,
  {32'hbaddfd80, 32'h3d1b33d9} /* (8, 20, 29) {real, imag} */,
  {32'hbdb4af84, 32'h3d7136a0} /* (8, 20, 28) {real, imag} */,
  {32'h3d8d4bd2, 32'hbd70b464} /* (8, 20, 27) {real, imag} */,
  {32'h3c88e11f, 32'h3d7ad1e0} /* (8, 20, 26) {real, imag} */,
  {32'hbce82178, 32'h3b3134b0} /* (8, 20, 25) {real, imag} */,
  {32'h3d7237fa, 32'h3d094aac} /* (8, 20, 24) {real, imag} */,
  {32'h3d4ddb83, 32'hbdd3595f} /* (8, 20, 23) {real, imag} */,
  {32'h3dac1b22, 32'hbe04b744} /* (8, 20, 22) {real, imag} */,
  {32'h3d8701fe, 32'hbd8bdbdc} /* (8, 20, 21) {real, imag} */,
  {32'hbafd6650, 32'h3ba64bc2} /* (8, 20, 20) {real, imag} */,
  {32'hbc9b0e97, 32'h3c2317f4} /* (8, 20, 19) {real, imag} */,
  {32'hbd60c151, 32'hbc1fcf5c} /* (8, 20, 18) {real, imag} */,
  {32'h3c1428f8, 32'h3cd21a66} /* (8, 20, 17) {real, imag} */,
  {32'hbd9e21b3, 32'h00000000} /* (8, 20, 16) {real, imag} */,
  {32'h3c1428f8, 32'hbcd21a66} /* (8, 20, 15) {real, imag} */,
  {32'hbd60c151, 32'h3c1fcf5c} /* (8, 20, 14) {real, imag} */,
  {32'hbc9b0e97, 32'hbc2317f4} /* (8, 20, 13) {real, imag} */,
  {32'hbafd6650, 32'hbba64bc2} /* (8, 20, 12) {real, imag} */,
  {32'h3d8701fe, 32'h3d8bdbdc} /* (8, 20, 11) {real, imag} */,
  {32'h3dac1b22, 32'h3e04b744} /* (8, 20, 10) {real, imag} */,
  {32'h3d4ddb83, 32'h3dd3595f} /* (8, 20, 9) {real, imag} */,
  {32'h3d7237fa, 32'hbd094aac} /* (8, 20, 8) {real, imag} */,
  {32'hbce82178, 32'hbb3134b0} /* (8, 20, 7) {real, imag} */,
  {32'h3c88e11f, 32'hbd7ad1e0} /* (8, 20, 6) {real, imag} */,
  {32'h3d8d4bd2, 32'h3d70b464} /* (8, 20, 5) {real, imag} */,
  {32'hbdb4af84, 32'hbd7136a0} /* (8, 20, 4) {real, imag} */,
  {32'hbaddfd80, 32'hbd1b33d9} /* (8, 20, 3) {real, imag} */,
  {32'h3f0eea07, 32'h3e945a7a} /* (8, 20, 2) {real, imag} */,
  {32'hbfa34c60, 32'hbcaffb80} /* (8, 20, 1) {real, imag} */,
  {32'hbf018449, 32'h00000000} /* (8, 20, 0) {real, imag} */,
  {32'hc01ed520, 32'h3d08f0d0} /* (8, 19, 31) {real, imag} */,
  {32'h3f85f5cf, 32'hbe8bc138} /* (8, 19, 30) {real, imag} */,
  {32'h3c2af2c4, 32'h3cf9035c} /* (8, 19, 29) {real, imag} */,
  {32'hbe65cfd4, 32'hbe040507} /* (8, 19, 28) {real, imag} */,
  {32'h3e8209fd, 32'hbdf4d9f5} /* (8, 19, 27) {real, imag} */,
  {32'h3dbd0016, 32'hbcf7bacf} /* (8, 19, 26) {real, imag} */,
  {32'h3d457aa4, 32'h3e0fca82} /* (8, 19, 25) {real, imag} */,
  {32'h3c350af8, 32'hbd1acf42} /* (8, 19, 24) {real, imag} */,
  {32'hbd81a2e2, 32'hbd95e9f8} /* (8, 19, 23) {real, imag} */,
  {32'h3d063657, 32'h3e336a9b} /* (8, 19, 22) {real, imag} */,
  {32'hbdf8d02c, 32'hbcb9aa5c} /* (8, 19, 21) {real, imag} */,
  {32'h3cf0407c, 32'hbc39bbab} /* (8, 19, 20) {real, imag} */,
  {32'h3dca2482, 32'h3d294082} /* (8, 19, 19) {real, imag} */,
  {32'hbdc67553, 32'hbd73e9d0} /* (8, 19, 18) {real, imag} */,
  {32'h3ce5bfb0, 32'hbc5bb05a} /* (8, 19, 17) {real, imag} */,
  {32'hbbf9d920, 32'h00000000} /* (8, 19, 16) {real, imag} */,
  {32'h3ce5bfb0, 32'h3c5bb05a} /* (8, 19, 15) {real, imag} */,
  {32'hbdc67553, 32'h3d73e9d0} /* (8, 19, 14) {real, imag} */,
  {32'h3dca2482, 32'hbd294082} /* (8, 19, 13) {real, imag} */,
  {32'h3cf0407c, 32'h3c39bbab} /* (8, 19, 12) {real, imag} */,
  {32'hbdf8d02c, 32'h3cb9aa5c} /* (8, 19, 11) {real, imag} */,
  {32'h3d063657, 32'hbe336a9b} /* (8, 19, 10) {real, imag} */,
  {32'hbd81a2e2, 32'h3d95e9f8} /* (8, 19, 9) {real, imag} */,
  {32'h3c350af8, 32'h3d1acf42} /* (8, 19, 8) {real, imag} */,
  {32'h3d457aa4, 32'hbe0fca82} /* (8, 19, 7) {real, imag} */,
  {32'h3dbd0016, 32'h3cf7bacf} /* (8, 19, 6) {real, imag} */,
  {32'h3e8209fd, 32'h3df4d9f5} /* (8, 19, 5) {real, imag} */,
  {32'hbe65cfd4, 32'h3e040507} /* (8, 19, 4) {real, imag} */,
  {32'h3c2af2c4, 32'hbcf9035c} /* (8, 19, 3) {real, imag} */,
  {32'h3f85f5cf, 32'h3e8bc138} /* (8, 19, 2) {real, imag} */,
  {32'hc01ed520, 32'hbd08f0d0} /* (8, 19, 1) {real, imag} */,
  {32'hbfb7bdc0, 32'h00000000} /* (8, 19, 0) {real, imag} */,
  {32'hc0579699, 32'h3e878570} /* (8, 18, 31) {real, imag} */,
  {32'h3f9ee1d2, 32'hbe8db865} /* (8, 18, 30) {real, imag} */,
  {32'hbe190cfe, 32'hbde475e3} /* (8, 18, 29) {real, imag} */,
  {32'hbea72d34, 32'hbd6841af} /* (8, 18, 28) {real, imag} */,
  {32'h3e832f86, 32'h3d8e0b5c} /* (8, 18, 27) {real, imag} */,
  {32'h3d6b41f6, 32'hbdc7c270} /* (8, 18, 26) {real, imag} */,
  {32'hbb5978c8, 32'h3dba53d6} /* (8, 18, 25) {real, imag} */,
  {32'h3e1f32f2, 32'h3d814065} /* (8, 18, 24) {real, imag} */,
  {32'hbd00a6d4, 32'h3d1d6c46} /* (8, 18, 23) {real, imag} */,
  {32'hbd13eae4, 32'hbd9c30a3} /* (8, 18, 22) {real, imag} */,
  {32'h3d3e2998, 32'hbd44b0a1} /* (8, 18, 21) {real, imag} */,
  {32'hbd37540e, 32'h3d08d3e8} /* (8, 18, 20) {real, imag} */,
  {32'hbbdc9f34, 32'hbdc8f57a} /* (8, 18, 19) {real, imag} */,
  {32'h3d60a8a0, 32'hbce9acf6} /* (8, 18, 18) {real, imag} */,
  {32'hbc0e23a4, 32'h3ccbf776} /* (8, 18, 17) {real, imag} */,
  {32'h3b88b3ae, 32'h00000000} /* (8, 18, 16) {real, imag} */,
  {32'hbc0e23a4, 32'hbccbf776} /* (8, 18, 15) {real, imag} */,
  {32'h3d60a8a0, 32'h3ce9acf6} /* (8, 18, 14) {real, imag} */,
  {32'hbbdc9f34, 32'h3dc8f57a} /* (8, 18, 13) {real, imag} */,
  {32'hbd37540e, 32'hbd08d3e8} /* (8, 18, 12) {real, imag} */,
  {32'h3d3e2998, 32'h3d44b0a1} /* (8, 18, 11) {real, imag} */,
  {32'hbd13eae4, 32'h3d9c30a3} /* (8, 18, 10) {real, imag} */,
  {32'hbd00a6d4, 32'hbd1d6c46} /* (8, 18, 9) {real, imag} */,
  {32'h3e1f32f2, 32'hbd814065} /* (8, 18, 8) {real, imag} */,
  {32'hbb5978c8, 32'hbdba53d6} /* (8, 18, 7) {real, imag} */,
  {32'h3d6b41f6, 32'h3dc7c270} /* (8, 18, 6) {real, imag} */,
  {32'h3e832f86, 32'hbd8e0b5c} /* (8, 18, 5) {real, imag} */,
  {32'hbea72d34, 32'h3d6841af} /* (8, 18, 4) {real, imag} */,
  {32'hbe190cfe, 32'h3de475e3} /* (8, 18, 3) {real, imag} */,
  {32'h3f9ee1d2, 32'h3e8db865} /* (8, 18, 2) {real, imag} */,
  {32'hc0579699, 32'hbe878570} /* (8, 18, 1) {real, imag} */,
  {32'hc00e7556, 32'h00000000} /* (8, 18, 0) {real, imag} */,
  {32'hc071653b, 32'h3e8f8c82} /* (8, 17, 31) {real, imag} */,
  {32'h3f9fcc1b, 32'hbe4fb7cc} /* (8, 17, 30) {real, imag} */,
  {32'hbd40b305, 32'hbd4e54db} /* (8, 17, 29) {real, imag} */,
  {32'hbe003335, 32'h3dac0ae9} /* (8, 17, 28) {real, imag} */,
  {32'h3e89ea8e, 32'h3e013104} /* (8, 17, 27) {real, imag} */,
  {32'h3e654d4a, 32'hbd97b235} /* (8, 17, 26) {real, imag} */,
  {32'hbd066266, 32'h3c3476e6} /* (8, 17, 25) {real, imag} */,
  {32'h3da29442, 32'h3deea609} /* (8, 17, 24) {real, imag} */,
  {32'h3d9b117f, 32'hbd2d5714} /* (8, 17, 23) {real, imag} */,
  {32'h3c883e7c, 32'hbd4c013d} /* (8, 17, 22) {real, imag} */,
  {32'hbd0cabcd, 32'hbcbfc788} /* (8, 17, 21) {real, imag} */,
  {32'hbbcd283e, 32'hbda3dc1b} /* (8, 17, 20) {real, imag} */,
  {32'hbcb87d95, 32'hbdb7cfd8} /* (8, 17, 19) {real, imag} */,
  {32'h3d44dbc2, 32'hbcc6d26e} /* (8, 17, 18) {real, imag} */,
  {32'hbd0210be, 32'h3d183892} /* (8, 17, 17) {real, imag} */,
  {32'h3cb0330e, 32'h00000000} /* (8, 17, 16) {real, imag} */,
  {32'hbd0210be, 32'hbd183892} /* (8, 17, 15) {real, imag} */,
  {32'h3d44dbc2, 32'h3cc6d26e} /* (8, 17, 14) {real, imag} */,
  {32'hbcb87d95, 32'h3db7cfd8} /* (8, 17, 13) {real, imag} */,
  {32'hbbcd283e, 32'h3da3dc1b} /* (8, 17, 12) {real, imag} */,
  {32'hbd0cabcd, 32'h3cbfc788} /* (8, 17, 11) {real, imag} */,
  {32'h3c883e7c, 32'h3d4c013d} /* (8, 17, 10) {real, imag} */,
  {32'h3d9b117f, 32'h3d2d5714} /* (8, 17, 9) {real, imag} */,
  {32'h3da29442, 32'hbdeea609} /* (8, 17, 8) {real, imag} */,
  {32'hbd066266, 32'hbc3476e6} /* (8, 17, 7) {real, imag} */,
  {32'h3e654d4a, 32'h3d97b235} /* (8, 17, 6) {real, imag} */,
  {32'h3e89ea8e, 32'hbe013104} /* (8, 17, 5) {real, imag} */,
  {32'hbe003335, 32'hbdac0ae9} /* (8, 17, 4) {real, imag} */,
  {32'hbd40b305, 32'h3d4e54db} /* (8, 17, 3) {real, imag} */,
  {32'h3f9fcc1b, 32'h3e4fb7cc} /* (8, 17, 2) {real, imag} */,
  {32'hc071653b, 32'hbe8f8c82} /* (8, 17, 1) {real, imag} */,
  {32'hc0425110, 32'h00000000} /* (8, 17, 0) {real, imag} */,
  {32'hc0811c96, 32'h3e886fac} /* (8, 16, 31) {real, imag} */,
  {32'h3fa9c94a, 32'hbe78ac38} /* (8, 16, 30) {real, imag} */,
  {32'hbd9d1317, 32'hbcf5597a} /* (8, 16, 29) {real, imag} */,
  {32'hbdf68f38, 32'h3c6c4778} /* (8, 16, 28) {real, imag} */,
  {32'h3e8d6641, 32'hbcd2e4c4} /* (8, 16, 27) {real, imag} */,
  {32'h3db40e88, 32'hbcda9e40} /* (8, 16, 26) {real, imag} */,
  {32'hbb3ed030, 32'h3d037256} /* (8, 16, 25) {real, imag} */,
  {32'h3d460e9c, 32'h3bfa766a} /* (8, 16, 24) {real, imag} */,
  {32'h3db72d22, 32'hbcced608} /* (8, 16, 23) {real, imag} */,
  {32'h3d749520, 32'hbc09e570} /* (8, 16, 22) {real, imag} */,
  {32'h3d5ca64b, 32'hbcfd2f61} /* (8, 16, 21) {real, imag} */,
  {32'hbcab1208, 32'hbe030d39} /* (8, 16, 20) {real, imag} */,
  {32'h3d5bbb82, 32'hbd021b83} /* (8, 16, 19) {real, imag} */,
  {32'hbd60f8d9, 32'hbca4bc00} /* (8, 16, 18) {real, imag} */,
  {32'h3c7c8118, 32'h3d1372fa} /* (8, 16, 17) {real, imag} */,
  {32'hbd46b56b, 32'h00000000} /* (8, 16, 16) {real, imag} */,
  {32'h3c7c8118, 32'hbd1372fa} /* (8, 16, 15) {real, imag} */,
  {32'hbd60f8d9, 32'h3ca4bc00} /* (8, 16, 14) {real, imag} */,
  {32'h3d5bbb82, 32'h3d021b83} /* (8, 16, 13) {real, imag} */,
  {32'hbcab1208, 32'h3e030d39} /* (8, 16, 12) {real, imag} */,
  {32'h3d5ca64b, 32'h3cfd2f61} /* (8, 16, 11) {real, imag} */,
  {32'h3d749520, 32'h3c09e570} /* (8, 16, 10) {real, imag} */,
  {32'h3db72d22, 32'h3cced608} /* (8, 16, 9) {real, imag} */,
  {32'h3d460e9c, 32'hbbfa766a} /* (8, 16, 8) {real, imag} */,
  {32'hbb3ed030, 32'hbd037256} /* (8, 16, 7) {real, imag} */,
  {32'h3db40e88, 32'h3cda9e40} /* (8, 16, 6) {real, imag} */,
  {32'h3e8d6641, 32'h3cd2e4c4} /* (8, 16, 5) {real, imag} */,
  {32'hbdf68f38, 32'hbc6c4778} /* (8, 16, 4) {real, imag} */,
  {32'hbd9d1317, 32'h3cf5597a} /* (8, 16, 3) {real, imag} */,
  {32'h3fa9c94a, 32'h3e78ac38} /* (8, 16, 2) {real, imag} */,
  {32'hc0811c96, 32'hbe886fac} /* (8, 16, 1) {real, imag} */,
  {32'hc0409f22, 32'h00000000} /* (8, 16, 0) {real, imag} */,
  {32'hc080454e, 32'h3e7d90bc} /* (8, 15, 31) {real, imag} */,
  {32'h3fb2f205, 32'hbe50d6f0} /* (8, 15, 30) {real, imag} */,
  {32'hbccfc082, 32'h3d95221a} /* (8, 15, 29) {real, imag} */,
  {32'hbe72be83, 32'h3dac21cf} /* (8, 15, 28) {real, imag} */,
  {32'h3e1f3267, 32'hbbfa0a70} /* (8, 15, 27) {real, imag} */,
  {32'h3e3097d2, 32'h3a23dd80} /* (8, 15, 26) {real, imag} */,
  {32'h3dbb905f, 32'hbd7d819c} /* (8, 15, 25) {real, imag} */,
  {32'h3db0e452, 32'h3dabdd71} /* (8, 15, 24) {real, imag} */,
  {32'hbc5ba306, 32'hbc836ae3} /* (8, 15, 23) {real, imag} */,
  {32'hbd48b4fa, 32'hbc925292} /* (8, 15, 22) {real, imag} */,
  {32'h3d7ecdf1, 32'hbd8e622e} /* (8, 15, 21) {real, imag} */,
  {32'hbc880e70, 32'h3d646a86} /* (8, 15, 20) {real, imag} */,
  {32'h3ca30c23, 32'h3d8f98f4} /* (8, 15, 19) {real, imag} */,
  {32'h3d2adcc6, 32'hbd425131} /* (8, 15, 18) {real, imag} */,
  {32'hbce3287b, 32'hbb571618} /* (8, 15, 17) {real, imag} */,
  {32'hba2f8f00, 32'h00000000} /* (8, 15, 16) {real, imag} */,
  {32'hbce3287b, 32'h3b571618} /* (8, 15, 15) {real, imag} */,
  {32'h3d2adcc6, 32'h3d425131} /* (8, 15, 14) {real, imag} */,
  {32'h3ca30c23, 32'hbd8f98f4} /* (8, 15, 13) {real, imag} */,
  {32'hbc880e70, 32'hbd646a86} /* (8, 15, 12) {real, imag} */,
  {32'h3d7ecdf1, 32'h3d8e622e} /* (8, 15, 11) {real, imag} */,
  {32'hbd48b4fa, 32'h3c925292} /* (8, 15, 10) {real, imag} */,
  {32'hbc5ba306, 32'h3c836ae3} /* (8, 15, 9) {real, imag} */,
  {32'h3db0e452, 32'hbdabdd71} /* (8, 15, 8) {real, imag} */,
  {32'h3dbb905f, 32'h3d7d819c} /* (8, 15, 7) {real, imag} */,
  {32'h3e3097d2, 32'hba23dd80} /* (8, 15, 6) {real, imag} */,
  {32'h3e1f3267, 32'h3bfa0a70} /* (8, 15, 5) {real, imag} */,
  {32'hbe72be83, 32'hbdac21cf} /* (8, 15, 4) {real, imag} */,
  {32'hbccfc082, 32'hbd95221a} /* (8, 15, 3) {real, imag} */,
  {32'h3fb2f205, 32'h3e50d6f0} /* (8, 15, 2) {real, imag} */,
  {32'hc080454e, 32'hbe7d90bc} /* (8, 15, 1) {real, imag} */,
  {32'hc03a4a9c, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'hc05d6df3, 32'h3e68b670} /* (8, 14, 31) {real, imag} */,
  {32'h3fac3086, 32'hbe6beda2} /* (8, 14, 30) {real, imag} */,
  {32'h3d64d451, 32'h3d1de046} /* (8, 14, 29) {real, imag} */,
  {32'hbe8c91e0, 32'h3d23a5d3} /* (8, 14, 28) {real, imag} */,
  {32'h3da9658a, 32'hbe71507c} /* (8, 14, 27) {real, imag} */,
  {32'h3d47a3f2, 32'hbd29a2b0} /* (8, 14, 26) {real, imag} */,
  {32'hbbd12b04, 32'h3d91fe7e} /* (8, 14, 25) {real, imag} */,
  {32'h3c426fa0, 32'hbc96a348} /* (8, 14, 24) {real, imag} */,
  {32'hbcf6b77b, 32'hbddff245} /* (8, 14, 23) {real, imag} */,
  {32'hbd8722e4, 32'h3d824e55} /* (8, 14, 22) {real, imag} */,
  {32'h3d196234, 32'hbd12aaa3} /* (8, 14, 21) {real, imag} */,
  {32'h3d41930a, 32'hbd894843} /* (8, 14, 20) {real, imag} */,
  {32'hbc816407, 32'hbbdb3de0} /* (8, 14, 19) {real, imag} */,
  {32'hbd8db9e7, 32'hbcf4b7ba} /* (8, 14, 18) {real, imag} */,
  {32'hbc2621b0, 32'hbbb30ad8} /* (8, 14, 17) {real, imag} */,
  {32'hbca0b2c2, 32'h00000000} /* (8, 14, 16) {real, imag} */,
  {32'hbc2621b0, 32'h3bb30ad8} /* (8, 14, 15) {real, imag} */,
  {32'hbd8db9e7, 32'h3cf4b7ba} /* (8, 14, 14) {real, imag} */,
  {32'hbc816407, 32'h3bdb3de0} /* (8, 14, 13) {real, imag} */,
  {32'h3d41930a, 32'h3d894843} /* (8, 14, 12) {real, imag} */,
  {32'h3d196234, 32'h3d12aaa3} /* (8, 14, 11) {real, imag} */,
  {32'hbd8722e4, 32'hbd824e55} /* (8, 14, 10) {real, imag} */,
  {32'hbcf6b77b, 32'h3ddff245} /* (8, 14, 9) {real, imag} */,
  {32'h3c426fa0, 32'h3c96a348} /* (8, 14, 8) {real, imag} */,
  {32'hbbd12b04, 32'hbd91fe7e} /* (8, 14, 7) {real, imag} */,
  {32'h3d47a3f2, 32'h3d29a2b0} /* (8, 14, 6) {real, imag} */,
  {32'h3da9658a, 32'h3e71507c} /* (8, 14, 5) {real, imag} */,
  {32'hbe8c91e0, 32'hbd23a5d3} /* (8, 14, 4) {real, imag} */,
  {32'h3d64d451, 32'hbd1de046} /* (8, 14, 3) {real, imag} */,
  {32'h3fac3086, 32'h3e6beda2} /* (8, 14, 2) {real, imag} */,
  {32'hc05d6df3, 32'hbe68b670} /* (8, 14, 1) {real, imag} */,
  {32'hc039979a, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'hc03ebcd2, 32'h3debc4f8} /* (8, 13, 31) {real, imag} */,
  {32'h3f9b1285, 32'hbe9d436e} /* (8, 13, 30) {real, imag} */,
  {32'h3d8ce678, 32'h3d1fa31a} /* (8, 13, 29) {real, imag} */,
  {32'hbe50a666, 32'h3d54890c} /* (8, 13, 28) {real, imag} */,
  {32'h3df44dad, 32'hbdf545cd} /* (8, 13, 27) {real, imag} */,
  {32'hbd08f5e8, 32'hbc975e9f} /* (8, 13, 26) {real, imag} */,
  {32'hbe1fea79, 32'h3d055f43} /* (8, 13, 25) {real, imag} */,
  {32'h3e42b19e, 32'hbe08451c} /* (8, 13, 24) {real, imag} */,
  {32'h3d52ec00, 32'hbc357d0c} /* (8, 13, 23) {real, imag} */,
  {32'h3d5db003, 32'h3d05d38c} /* (8, 13, 22) {real, imag} */,
  {32'h3dac2ad8, 32'hbd2269d4} /* (8, 13, 21) {real, imag} */,
  {32'hbd74b2bc, 32'hbccfeb82} /* (8, 13, 20) {real, imag} */,
  {32'hbc4f22a0, 32'h3caf514c} /* (8, 13, 19) {real, imag} */,
  {32'h3d157ed2, 32'hbd03d4fe} /* (8, 13, 18) {real, imag} */,
  {32'h3b0d499c, 32'h3a8368d0} /* (8, 13, 17) {real, imag} */,
  {32'hbd638cf8, 32'h00000000} /* (8, 13, 16) {real, imag} */,
  {32'h3b0d499c, 32'hba8368d0} /* (8, 13, 15) {real, imag} */,
  {32'h3d157ed2, 32'h3d03d4fe} /* (8, 13, 14) {real, imag} */,
  {32'hbc4f22a0, 32'hbcaf514c} /* (8, 13, 13) {real, imag} */,
  {32'hbd74b2bc, 32'h3ccfeb82} /* (8, 13, 12) {real, imag} */,
  {32'h3dac2ad8, 32'h3d2269d4} /* (8, 13, 11) {real, imag} */,
  {32'h3d5db003, 32'hbd05d38c} /* (8, 13, 10) {real, imag} */,
  {32'h3d52ec00, 32'h3c357d0c} /* (8, 13, 9) {real, imag} */,
  {32'h3e42b19e, 32'h3e08451c} /* (8, 13, 8) {real, imag} */,
  {32'hbe1fea79, 32'hbd055f43} /* (8, 13, 7) {real, imag} */,
  {32'hbd08f5e8, 32'h3c975e9f} /* (8, 13, 6) {real, imag} */,
  {32'h3df44dad, 32'h3df545cd} /* (8, 13, 5) {real, imag} */,
  {32'hbe50a666, 32'hbd54890c} /* (8, 13, 4) {real, imag} */,
  {32'h3d8ce678, 32'hbd1fa31a} /* (8, 13, 3) {real, imag} */,
  {32'h3f9b1285, 32'h3e9d436e} /* (8, 13, 2) {real, imag} */,
  {32'hc03ebcd2, 32'hbdebc4f8} /* (8, 13, 1) {real, imag} */,
  {32'hc0126c5e, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'hc00a6992, 32'hbda0b9c0} /* (8, 12, 31) {real, imag} */,
  {32'h3f835d8c, 32'hbcdddec8} /* (8, 12, 30) {real, imag} */,
  {32'h3e5e046c, 32'h3c09a210} /* (8, 12, 29) {real, imag} */,
  {32'hbd825480, 32'hbe0cb669} /* (8, 12, 28) {real, imag} */,
  {32'h3df1625a, 32'hbd4e6cac} /* (8, 12, 27) {real, imag} */,
  {32'h3d946556, 32'hbd1095e8} /* (8, 12, 26) {real, imag} */,
  {32'hbe07d481, 32'h3d56f749} /* (8, 12, 25) {real, imag} */,
  {32'h3d22d340, 32'hbd88b8e3} /* (8, 12, 24) {real, imag} */,
  {32'hbd0d145f, 32'h3d54e256} /* (8, 12, 23) {real, imag} */,
  {32'hbd642af4, 32'h3dc362c4} /* (8, 12, 22) {real, imag} */,
  {32'hbb4e3a90, 32'hbd581d1e} /* (8, 12, 21) {real, imag} */,
  {32'hbca86ff3, 32'hbcffdbc4} /* (8, 12, 20) {real, imag} */,
  {32'h3d80116c, 32'h3b87b114} /* (8, 12, 19) {real, imag} */,
  {32'hbd8ae7de, 32'hbd6e8f3b} /* (8, 12, 18) {real, imag} */,
  {32'hbac0ec40, 32'hbc174f10} /* (8, 12, 17) {real, imag} */,
  {32'h3b3f5a80, 32'h00000000} /* (8, 12, 16) {real, imag} */,
  {32'hbac0ec40, 32'h3c174f10} /* (8, 12, 15) {real, imag} */,
  {32'hbd8ae7de, 32'h3d6e8f3b} /* (8, 12, 14) {real, imag} */,
  {32'h3d80116c, 32'hbb87b114} /* (8, 12, 13) {real, imag} */,
  {32'hbca86ff3, 32'h3cffdbc4} /* (8, 12, 12) {real, imag} */,
  {32'hbb4e3a90, 32'h3d581d1e} /* (8, 12, 11) {real, imag} */,
  {32'hbd642af4, 32'hbdc362c4} /* (8, 12, 10) {real, imag} */,
  {32'hbd0d145f, 32'hbd54e256} /* (8, 12, 9) {real, imag} */,
  {32'h3d22d340, 32'h3d88b8e3} /* (8, 12, 8) {real, imag} */,
  {32'hbe07d481, 32'hbd56f749} /* (8, 12, 7) {real, imag} */,
  {32'h3d946556, 32'h3d1095e8} /* (8, 12, 6) {real, imag} */,
  {32'h3df1625a, 32'h3d4e6cac} /* (8, 12, 5) {real, imag} */,
  {32'hbd825480, 32'h3e0cb669} /* (8, 12, 4) {real, imag} */,
  {32'h3e5e046c, 32'hbc09a210} /* (8, 12, 3) {real, imag} */,
  {32'h3f835d8c, 32'h3cdddec8} /* (8, 12, 2) {real, imag} */,
  {32'hc00a6992, 32'h3da0b9c0} /* (8, 12, 1) {real, imag} */,
  {32'hbfc2b7bc, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'hbf8464ef, 32'hbe92aaf1} /* (8, 11, 31) {real, imag} */,
  {32'h3f05441e, 32'h3c6e43b8} /* (8, 11, 30) {real, imag} */,
  {32'h3e50db9c, 32'h3d995d98} /* (8, 11, 29) {real, imag} */,
  {32'hbe18f5bd, 32'hbe329e7a} /* (8, 11, 28) {real, imag} */,
  {32'h3bf190f0, 32'hbd9e444a} /* (8, 11, 27) {real, imag} */,
  {32'h3cda9917, 32'hbdd6f2c7} /* (8, 11, 26) {real, imag} */,
  {32'hbe0980cd, 32'hbe21e178} /* (8, 11, 25) {real, imag} */,
  {32'hbc1099f0, 32'hbdf24d0e} /* (8, 11, 24) {real, imag} */,
  {32'h3db010e9, 32'h3d640bbe} /* (8, 11, 23) {real, imag} */,
  {32'h3dcc92ef, 32'h3d50b86b} /* (8, 11, 22) {real, imag} */,
  {32'hbc9ea28f, 32'hbc4f1948} /* (8, 11, 21) {real, imag} */,
  {32'h3b519000, 32'hbd2d2436} /* (8, 11, 20) {real, imag} */,
  {32'hbd60e786, 32'h3cab9788} /* (8, 11, 19) {real, imag} */,
  {32'h3d2ef5d2, 32'hbd426368} /* (8, 11, 18) {real, imag} */,
  {32'h3cda2d9b, 32'hbb8428f0} /* (8, 11, 17) {real, imag} */,
  {32'hbda7ea3c, 32'h00000000} /* (8, 11, 16) {real, imag} */,
  {32'h3cda2d9b, 32'h3b8428f0} /* (8, 11, 15) {real, imag} */,
  {32'h3d2ef5d2, 32'h3d426368} /* (8, 11, 14) {real, imag} */,
  {32'hbd60e786, 32'hbcab9788} /* (8, 11, 13) {real, imag} */,
  {32'h3b519000, 32'h3d2d2436} /* (8, 11, 12) {real, imag} */,
  {32'hbc9ea28f, 32'h3c4f1948} /* (8, 11, 11) {real, imag} */,
  {32'h3dcc92ef, 32'hbd50b86b} /* (8, 11, 10) {real, imag} */,
  {32'h3db010e9, 32'hbd640bbe} /* (8, 11, 9) {real, imag} */,
  {32'hbc1099f0, 32'h3df24d0e} /* (8, 11, 8) {real, imag} */,
  {32'hbe0980cd, 32'h3e21e178} /* (8, 11, 7) {real, imag} */,
  {32'h3cda9917, 32'h3dd6f2c7} /* (8, 11, 6) {real, imag} */,
  {32'h3bf190f0, 32'h3d9e444a} /* (8, 11, 5) {real, imag} */,
  {32'hbe18f5bd, 32'h3e329e7a} /* (8, 11, 4) {real, imag} */,
  {32'h3e50db9c, 32'hbd995d98} /* (8, 11, 3) {real, imag} */,
  {32'h3f05441e, 32'hbc6e43b8} /* (8, 11, 2) {real, imag} */,
  {32'hbf8464ef, 32'h3e92aaf1} /* (8, 11, 1) {real, imag} */,
  {32'hbf1bb374, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h3f0b928a, 32'hbf2ea12a} /* (8, 10, 31) {real, imag} */,
  {32'hbe8df841, 32'h3e46f7c4} /* (8, 10, 30) {real, imag} */,
  {32'h3de3e56b, 32'h3d3a578a} /* (8, 10, 29) {real, imag} */,
  {32'hbd5e8920, 32'hbe2be61f} /* (8, 10, 28) {real, imag} */,
  {32'hbde9966a, 32'h3e179a77} /* (8, 10, 27) {real, imag} */,
  {32'hbbb42f72, 32'hbca3c336} /* (8, 10, 26) {real, imag} */,
  {32'h3cb53f08, 32'hbe0a3e6b} /* (8, 10, 25) {real, imag} */,
  {32'h3db2c1b6, 32'hbdd1224a} /* (8, 10, 24) {real, imag} */,
  {32'hbd0b3a12, 32'hbc86e6b9} /* (8, 10, 23) {real, imag} */,
  {32'h3d765901, 32'h3d8e588e} /* (8, 10, 22) {real, imag} */,
  {32'h3b21b4c0, 32'h3cf4542c} /* (8, 10, 21) {real, imag} */,
  {32'hbd54ce52, 32'h3d30abdc} /* (8, 10, 20) {real, imag} */,
  {32'hbab116a0, 32'h3db5a9a2} /* (8, 10, 19) {real, imag} */,
  {32'h3d8a8e8a, 32'h3ce01086} /* (8, 10, 18) {real, imag} */,
  {32'hbc1192ee, 32'hbd9faf14} /* (8, 10, 17) {real, imag} */,
  {32'hbbc0a2f8, 32'h00000000} /* (8, 10, 16) {real, imag} */,
  {32'hbc1192ee, 32'h3d9faf14} /* (8, 10, 15) {real, imag} */,
  {32'h3d8a8e8a, 32'hbce01086} /* (8, 10, 14) {real, imag} */,
  {32'hbab116a0, 32'hbdb5a9a2} /* (8, 10, 13) {real, imag} */,
  {32'hbd54ce52, 32'hbd30abdc} /* (8, 10, 12) {real, imag} */,
  {32'h3b21b4c0, 32'hbcf4542c} /* (8, 10, 11) {real, imag} */,
  {32'h3d765901, 32'hbd8e588e} /* (8, 10, 10) {real, imag} */,
  {32'hbd0b3a12, 32'h3c86e6b9} /* (8, 10, 9) {real, imag} */,
  {32'h3db2c1b6, 32'h3dd1224a} /* (8, 10, 8) {real, imag} */,
  {32'h3cb53f08, 32'h3e0a3e6b} /* (8, 10, 7) {real, imag} */,
  {32'hbbb42f72, 32'h3ca3c336} /* (8, 10, 6) {real, imag} */,
  {32'hbde9966a, 32'hbe179a77} /* (8, 10, 5) {real, imag} */,
  {32'hbd5e8920, 32'h3e2be61f} /* (8, 10, 4) {real, imag} */,
  {32'h3de3e56b, 32'hbd3a578a} /* (8, 10, 3) {real, imag} */,
  {32'hbe8df841, 32'hbe46f7c4} /* (8, 10, 2) {real, imag} */,
  {32'h3f0b928a, 32'h3f2ea12a} /* (8, 10, 1) {real, imag} */,
  {32'h3f72eb51, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'h3ff30a1e, 32'hbf7e1134} /* (8, 9, 31) {real, imag} */,
  {32'hbf48360a, 32'h3ee03f2d} /* (8, 9, 30) {real, imag} */,
  {32'h3d40d132, 32'hbe125491} /* (8, 9, 29) {real, imag} */,
  {32'h3e087d6a, 32'hbdd388db} /* (8, 9, 28) {real, imag} */,
  {32'hbe2cc492, 32'h3dae83ea} /* (8, 9, 27) {real, imag} */,
  {32'h3d7db2c1, 32'h3c098261} /* (8, 9, 26) {real, imag} */,
  {32'hbd6e9df5, 32'h3d33ad71} /* (8, 9, 25) {real, imag} */,
  {32'h3dc595b1, 32'h3cbb661e} /* (8, 9, 24) {real, imag} */,
  {32'h3d845f5d, 32'h3d31de7f} /* (8, 9, 23) {real, imag} */,
  {32'hbd97d28b, 32'h3d5409e0} /* (8, 9, 22) {real, imag} */,
  {32'h3d492d84, 32'hbdb97c72} /* (8, 9, 21) {real, imag} */,
  {32'hbd1dfd75, 32'h3d71ded4} /* (8, 9, 20) {real, imag} */,
  {32'h3d544936, 32'hbd5a9da6} /* (8, 9, 19) {real, imag} */,
  {32'h3d9e2af1, 32'h3b75f770} /* (8, 9, 18) {real, imag} */,
  {32'hbd46f674, 32'hbc067604} /* (8, 9, 17) {real, imag} */,
  {32'hbca5cfc0, 32'h00000000} /* (8, 9, 16) {real, imag} */,
  {32'hbd46f674, 32'h3c067604} /* (8, 9, 15) {real, imag} */,
  {32'h3d9e2af1, 32'hbb75f770} /* (8, 9, 14) {real, imag} */,
  {32'h3d544936, 32'h3d5a9da6} /* (8, 9, 13) {real, imag} */,
  {32'hbd1dfd75, 32'hbd71ded4} /* (8, 9, 12) {real, imag} */,
  {32'h3d492d84, 32'h3db97c72} /* (8, 9, 11) {real, imag} */,
  {32'hbd97d28b, 32'hbd5409e0} /* (8, 9, 10) {real, imag} */,
  {32'h3d845f5d, 32'hbd31de7f} /* (8, 9, 9) {real, imag} */,
  {32'h3dc595b1, 32'hbcbb661e} /* (8, 9, 8) {real, imag} */,
  {32'hbd6e9df5, 32'hbd33ad71} /* (8, 9, 7) {real, imag} */,
  {32'h3d7db2c1, 32'hbc098261} /* (8, 9, 6) {real, imag} */,
  {32'hbe2cc492, 32'hbdae83ea} /* (8, 9, 5) {real, imag} */,
  {32'h3e087d6a, 32'h3dd388db} /* (8, 9, 4) {real, imag} */,
  {32'h3d40d132, 32'h3e125491} /* (8, 9, 3) {real, imag} */,
  {32'hbf48360a, 32'hbee03f2d} /* (8, 9, 2) {real, imag} */,
  {32'h3ff30a1e, 32'h3f7e1134} /* (8, 9, 1) {real, imag} */,
  {32'h4006bc5c, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'h402d34cc, 32'hbfaca5d2} /* (8, 8, 31) {real, imag} */,
  {32'hbf8695ba, 32'h3f02ea10} /* (8, 8, 30) {real, imag} */,
  {32'h3dd0de17, 32'hbd2cec0f} /* (8, 8, 29) {real, imag} */,
  {32'h3e00a73c, 32'hbdc220a0} /* (8, 8, 28) {real, imag} */,
  {32'hbe20c182, 32'hbd1ed40c} /* (8, 8, 27) {real, imag} */,
  {32'h3d437d9e, 32'hbccbaaf6} /* (8, 8, 26) {real, imag} */,
  {32'h3c8f8c10, 32'hbc02431c} /* (8, 8, 25) {real, imag} */,
  {32'hbc38b123, 32'h3ce27e42} /* (8, 8, 24) {real, imag} */,
  {32'hbd6aa5cc, 32'hbcda669c} /* (8, 8, 23) {real, imag} */,
  {32'h3da69046, 32'hbc55ec56} /* (8, 8, 22) {real, imag} */,
  {32'h3d1f8678, 32'h3cec45be} /* (8, 8, 21) {real, imag} */,
  {32'h3cd3645f, 32'hbd4cea2a} /* (8, 8, 20) {real, imag} */,
  {32'hbd96def2, 32'hbd553bec} /* (8, 8, 19) {real, imag} */,
  {32'hbe055c53, 32'hbcdb169d} /* (8, 8, 18) {real, imag} */,
  {32'hbd0f2ee8, 32'hbc974ffa} /* (8, 8, 17) {real, imag} */,
  {32'h3ddfdead, 32'h00000000} /* (8, 8, 16) {real, imag} */,
  {32'hbd0f2ee8, 32'h3c974ffa} /* (8, 8, 15) {real, imag} */,
  {32'hbe055c53, 32'h3cdb169d} /* (8, 8, 14) {real, imag} */,
  {32'hbd96def2, 32'h3d553bec} /* (8, 8, 13) {real, imag} */,
  {32'h3cd3645f, 32'h3d4cea2a} /* (8, 8, 12) {real, imag} */,
  {32'h3d1f8678, 32'hbcec45be} /* (8, 8, 11) {real, imag} */,
  {32'h3da69046, 32'h3c55ec56} /* (8, 8, 10) {real, imag} */,
  {32'hbd6aa5cc, 32'h3cda669c} /* (8, 8, 9) {real, imag} */,
  {32'hbc38b123, 32'hbce27e42} /* (8, 8, 8) {real, imag} */,
  {32'h3c8f8c10, 32'h3c02431c} /* (8, 8, 7) {real, imag} */,
  {32'h3d437d9e, 32'h3ccbaaf6} /* (8, 8, 6) {real, imag} */,
  {32'hbe20c182, 32'h3d1ed40c} /* (8, 8, 5) {real, imag} */,
  {32'h3e00a73c, 32'h3dc220a0} /* (8, 8, 4) {real, imag} */,
  {32'h3dd0de17, 32'h3d2cec0f} /* (8, 8, 3) {real, imag} */,
  {32'hbf8695ba, 32'hbf02ea10} /* (8, 8, 2) {real, imag} */,
  {32'h402d34cc, 32'h3faca5d2} /* (8, 8, 1) {real, imag} */,
  {32'h4041489c, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h404f2c10, 32'hbfca0631} /* (8, 7, 31) {real, imag} */,
  {32'hbf8e6964, 32'h3f24ef50} /* (8, 7, 30) {real, imag} */,
  {32'h3e03aa3f, 32'hbd99b6c7} /* (8, 7, 29) {real, imag} */,
  {32'h3e161424, 32'hbe019e10} /* (8, 7, 28) {real, imag} */,
  {32'hbe83fd4a, 32'h3e2d89f1} /* (8, 7, 27) {real, imag} */,
  {32'hbde68484, 32'h3d7e8cdf} /* (8, 7, 26) {real, imag} */,
  {32'h3dc57f8a, 32'hbd8890be} /* (8, 7, 25) {real, imag} */,
  {32'h3d9b7c12, 32'h3dfca390} /* (8, 7, 24) {real, imag} */,
  {32'h3d0da715, 32'h3d69acba} /* (8, 7, 23) {real, imag} */,
  {32'h3cbe6300, 32'h3cbab8e4} /* (8, 7, 22) {real, imag} */,
  {32'h3ce72e96, 32'h3d09f32c} /* (8, 7, 21) {real, imag} */,
  {32'h3dc3679e, 32'h3ce61694} /* (8, 7, 20) {real, imag} */,
  {32'h3dcbce5b, 32'hbd2fa8bc} /* (8, 7, 19) {real, imag} */,
  {32'hbcbc1ed0, 32'h3cf52536} /* (8, 7, 18) {real, imag} */,
  {32'hbd9e2878, 32'hbd61e02c} /* (8, 7, 17) {real, imag} */,
  {32'h3c9219c4, 32'h00000000} /* (8, 7, 16) {real, imag} */,
  {32'hbd9e2878, 32'h3d61e02c} /* (8, 7, 15) {real, imag} */,
  {32'hbcbc1ed0, 32'hbcf52536} /* (8, 7, 14) {real, imag} */,
  {32'h3dcbce5b, 32'h3d2fa8bc} /* (8, 7, 13) {real, imag} */,
  {32'h3dc3679e, 32'hbce61694} /* (8, 7, 12) {real, imag} */,
  {32'h3ce72e96, 32'hbd09f32c} /* (8, 7, 11) {real, imag} */,
  {32'h3cbe6300, 32'hbcbab8e4} /* (8, 7, 10) {real, imag} */,
  {32'h3d0da715, 32'hbd69acba} /* (8, 7, 9) {real, imag} */,
  {32'h3d9b7c12, 32'hbdfca390} /* (8, 7, 8) {real, imag} */,
  {32'h3dc57f8a, 32'h3d8890be} /* (8, 7, 7) {real, imag} */,
  {32'hbde68484, 32'hbd7e8cdf} /* (8, 7, 6) {real, imag} */,
  {32'hbe83fd4a, 32'hbe2d89f1} /* (8, 7, 5) {real, imag} */,
  {32'h3e161424, 32'h3e019e10} /* (8, 7, 4) {real, imag} */,
  {32'h3e03aa3f, 32'h3d99b6c7} /* (8, 7, 3) {real, imag} */,
  {32'hbf8e6964, 32'hbf24ef50} /* (8, 7, 2) {real, imag} */,
  {32'h404f2c10, 32'h3fca0631} /* (8, 7, 1) {real, imag} */,
  {32'h406bc8bf, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h405a8070, 32'hc0036202} /* (8, 6, 31) {real, imag} */,
  {32'hbf6cddba, 32'h3f59f31d} /* (8, 6, 30) {real, imag} */,
  {32'h3b844aec, 32'hbcc25c5f} /* (8, 6, 29) {real, imag} */,
  {32'h3dd8a4ec, 32'h3c07c7a4} /* (8, 6, 28) {real, imag} */,
  {32'hbe586115, 32'h3defd4d4} /* (8, 6, 27) {real, imag} */,
  {32'h3bd35428, 32'h3d2f071e} /* (8, 6, 26) {real, imag} */,
  {32'hbca27d38, 32'hbd41f7ce} /* (8, 6, 25) {real, imag} */,
  {32'hbd9cac5a, 32'h3d4bb047} /* (8, 6, 24) {real, imag} */,
  {32'hbb78288c, 32'hbd34f296} /* (8, 6, 23) {real, imag} */,
  {32'hbd81d17c, 32'hbd01f455} /* (8, 6, 22) {real, imag} */,
  {32'h3d6cc484, 32'hbce235ac} /* (8, 6, 21) {real, imag} */,
  {32'h3c5e70a8, 32'hbd6a8daf} /* (8, 6, 20) {real, imag} */,
  {32'hbca1e41b, 32'h3c9a6c05} /* (8, 6, 19) {real, imag} */,
  {32'hbbaf089a, 32'hbcc7cb5e} /* (8, 6, 18) {real, imag} */,
  {32'h3d75cffa, 32'hbcd8219d} /* (8, 6, 17) {real, imag} */,
  {32'h3dbe4cce, 32'h00000000} /* (8, 6, 16) {real, imag} */,
  {32'h3d75cffa, 32'h3cd8219d} /* (8, 6, 15) {real, imag} */,
  {32'hbbaf089a, 32'h3cc7cb5e} /* (8, 6, 14) {real, imag} */,
  {32'hbca1e41b, 32'hbc9a6c05} /* (8, 6, 13) {real, imag} */,
  {32'h3c5e70a8, 32'h3d6a8daf} /* (8, 6, 12) {real, imag} */,
  {32'h3d6cc484, 32'h3ce235ac} /* (8, 6, 11) {real, imag} */,
  {32'hbd81d17c, 32'h3d01f455} /* (8, 6, 10) {real, imag} */,
  {32'hbb78288c, 32'h3d34f296} /* (8, 6, 9) {real, imag} */,
  {32'hbd9cac5a, 32'hbd4bb047} /* (8, 6, 8) {real, imag} */,
  {32'hbca27d38, 32'h3d41f7ce} /* (8, 6, 7) {real, imag} */,
  {32'h3bd35428, 32'hbd2f071e} /* (8, 6, 6) {real, imag} */,
  {32'hbe586115, 32'hbdefd4d4} /* (8, 6, 5) {real, imag} */,
  {32'h3dd8a4ec, 32'hbc07c7a4} /* (8, 6, 4) {real, imag} */,
  {32'h3b844aec, 32'h3cc25c5f} /* (8, 6, 3) {real, imag} */,
  {32'hbf6cddba, 32'hbf59f31d} /* (8, 6, 2) {real, imag} */,
  {32'h405a8070, 32'h40036202} /* (8, 6, 1) {real, imag} */,
  {32'h408310c7, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'h404e6375, 32'hc036f323} /* (8, 5, 31) {real, imag} */,
  {32'hbec06df4, 32'h3f868fe3} /* (8, 5, 30) {real, imag} */,
  {32'h3d7a81ed, 32'hbd4a82ef} /* (8, 5, 29) {real, imag} */,
  {32'h3a721d00, 32'h3e456a7a} /* (8, 5, 28) {real, imag} */,
  {32'hbd6ff3a6, 32'h3d1114e8} /* (8, 5, 27) {real, imag} */,
  {32'h3db0765f, 32'h3dc4a23a} /* (8, 5, 26) {real, imag} */,
  {32'h3d9679f0, 32'hbc478370} /* (8, 5, 25) {real, imag} */,
  {32'h3d9b35e2, 32'h3d803424} /* (8, 5, 24) {real, imag} */,
  {32'h3c13b33d, 32'h3df9cd01} /* (8, 5, 23) {real, imag} */,
  {32'h3d1e2012, 32'h3d422c13} /* (8, 5, 22) {real, imag} */,
  {32'hbdc80992, 32'hbce2755c} /* (8, 5, 21) {real, imag} */,
  {32'hbd5ded4a, 32'hbd0a5384} /* (8, 5, 20) {real, imag} */,
  {32'h3dc047a7, 32'hbdb447d3} /* (8, 5, 19) {real, imag} */,
  {32'h3cb50e9f, 32'h3c187b41} /* (8, 5, 18) {real, imag} */,
  {32'hbd112556, 32'h3dc6dcc5} /* (8, 5, 17) {real, imag} */,
  {32'hbda9a751, 32'h00000000} /* (8, 5, 16) {real, imag} */,
  {32'hbd112556, 32'hbdc6dcc5} /* (8, 5, 15) {real, imag} */,
  {32'h3cb50e9f, 32'hbc187b41} /* (8, 5, 14) {real, imag} */,
  {32'h3dc047a7, 32'h3db447d3} /* (8, 5, 13) {real, imag} */,
  {32'hbd5ded4a, 32'h3d0a5384} /* (8, 5, 12) {real, imag} */,
  {32'hbdc80992, 32'h3ce2755c} /* (8, 5, 11) {real, imag} */,
  {32'h3d1e2012, 32'hbd422c13} /* (8, 5, 10) {real, imag} */,
  {32'h3c13b33d, 32'hbdf9cd01} /* (8, 5, 9) {real, imag} */,
  {32'h3d9b35e2, 32'hbd803424} /* (8, 5, 8) {real, imag} */,
  {32'h3d9679f0, 32'h3c478370} /* (8, 5, 7) {real, imag} */,
  {32'h3db0765f, 32'hbdc4a23a} /* (8, 5, 6) {real, imag} */,
  {32'hbd6ff3a6, 32'hbd1114e8} /* (8, 5, 5) {real, imag} */,
  {32'h3a721d00, 32'hbe456a7a} /* (8, 5, 4) {real, imag} */,
  {32'h3d7a81ed, 32'h3d4a82ef} /* (8, 5, 3) {real, imag} */,
  {32'hbec06df4, 32'hbf868fe3} /* (8, 5, 2) {real, imag} */,
  {32'h404e6375, 32'h4036f323} /* (8, 5, 1) {real, imag} */,
  {32'h4099ba1a, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'h403bcf36, 32'hc04f89b0} /* (8, 4, 31) {real, imag} */,
  {32'h3d4a4ff0, 32'h3f93e68e} /* (8, 4, 30) {real, imag} */,
  {32'hbd44aa1c, 32'h3d2c56cb} /* (8, 4, 29) {real, imag} */,
  {32'hbdc6b56c, 32'h3e4dcf19} /* (8, 4, 28) {real, imag} */,
  {32'hbe044de0, 32'h3dc42dc3} /* (8, 4, 27) {real, imag} */,
  {32'h3da22480, 32'h3dab28a2} /* (8, 4, 26) {real, imag} */,
  {32'h3d98dba4, 32'hbde59b20} /* (8, 4, 25) {real, imag} */,
  {32'hbb85c380, 32'h3d0438cb} /* (8, 4, 24) {real, imag} */,
  {32'hbd31a829, 32'hbdeae782} /* (8, 4, 23) {real, imag} */,
  {32'hbce8163a, 32'h3dc53832} /* (8, 4, 22) {real, imag} */,
  {32'hbe05124d, 32'h3c938314} /* (8, 4, 21) {real, imag} */,
  {32'h3d2812bd, 32'h3d59e0e4} /* (8, 4, 20) {real, imag} */,
  {32'h3d8e14e5, 32'h3cd3e8e4} /* (8, 4, 19) {real, imag} */,
  {32'h3d0b8b30, 32'h3b0ae638} /* (8, 4, 18) {real, imag} */,
  {32'hbd4235cf, 32'h3ce12ee8} /* (8, 4, 17) {real, imag} */,
  {32'hb8eb3c00, 32'h00000000} /* (8, 4, 16) {real, imag} */,
  {32'hbd4235cf, 32'hbce12ee8} /* (8, 4, 15) {real, imag} */,
  {32'h3d0b8b30, 32'hbb0ae638} /* (8, 4, 14) {real, imag} */,
  {32'h3d8e14e5, 32'hbcd3e8e4} /* (8, 4, 13) {real, imag} */,
  {32'h3d2812bd, 32'hbd59e0e4} /* (8, 4, 12) {real, imag} */,
  {32'hbe05124d, 32'hbc938314} /* (8, 4, 11) {real, imag} */,
  {32'hbce8163a, 32'hbdc53832} /* (8, 4, 10) {real, imag} */,
  {32'hbd31a829, 32'h3deae782} /* (8, 4, 9) {real, imag} */,
  {32'hbb85c380, 32'hbd0438cb} /* (8, 4, 8) {real, imag} */,
  {32'h3d98dba4, 32'h3de59b20} /* (8, 4, 7) {real, imag} */,
  {32'h3da22480, 32'hbdab28a2} /* (8, 4, 6) {real, imag} */,
  {32'hbe044de0, 32'hbdc42dc3} /* (8, 4, 5) {real, imag} */,
  {32'hbdc6b56c, 32'hbe4dcf19} /* (8, 4, 4) {real, imag} */,
  {32'hbd44aa1c, 32'hbd2c56cb} /* (8, 4, 3) {real, imag} */,
  {32'h3d4a4ff0, 32'hbf93e68e} /* (8, 4, 2) {real, imag} */,
  {32'h403bcf36, 32'h404f89b0} /* (8, 4, 1) {real, imag} */,
  {32'h40a36678, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'h40376d5e, 32'hc063b414} /* (8, 3, 31) {real, imag} */,
  {32'h3e72fcb0, 32'h3f898a86} /* (8, 3, 30) {real, imag} */,
  {32'hbd930fd8, 32'h3dc6ccb0} /* (8, 3, 29) {real, imag} */,
  {32'hbd379860, 32'h3e9e024e} /* (8, 3, 28) {real, imag} */,
  {32'hbe1a1852, 32'hbd6c987e} /* (8, 3, 27) {real, imag} */,
  {32'hbda6b8dc, 32'hbe21c094} /* (8, 3, 26) {real, imag} */,
  {32'h3cb0a260, 32'h3d781dd6} /* (8, 3, 25) {real, imag} */,
  {32'hbcdc41a4, 32'h3cd020f7} /* (8, 3, 24) {real, imag} */,
  {32'h3dcb902c, 32'h3cc86c4c} /* (8, 3, 23) {real, imag} */,
  {32'hbd62d00c, 32'h3db6c78c} /* (8, 3, 22) {real, imag} */,
  {32'hbd7f660d, 32'hbac06680} /* (8, 3, 21) {real, imag} */,
  {32'h3e102309, 32'h3bb834fa} /* (8, 3, 20) {real, imag} */,
  {32'hbdb2b26f, 32'h3bc16870} /* (8, 3, 19) {real, imag} */,
  {32'hbd4daa98, 32'h3d04e9f5} /* (8, 3, 18) {real, imag} */,
  {32'hbce0302c, 32'h3c41bb44} /* (8, 3, 17) {real, imag} */,
  {32'hbd966662, 32'h00000000} /* (8, 3, 16) {real, imag} */,
  {32'hbce0302c, 32'hbc41bb44} /* (8, 3, 15) {real, imag} */,
  {32'hbd4daa98, 32'hbd04e9f5} /* (8, 3, 14) {real, imag} */,
  {32'hbdb2b26f, 32'hbbc16870} /* (8, 3, 13) {real, imag} */,
  {32'h3e102309, 32'hbbb834fa} /* (8, 3, 12) {real, imag} */,
  {32'hbd7f660d, 32'h3ac06680} /* (8, 3, 11) {real, imag} */,
  {32'hbd62d00c, 32'hbdb6c78c} /* (8, 3, 10) {real, imag} */,
  {32'h3dcb902c, 32'hbcc86c4c} /* (8, 3, 9) {real, imag} */,
  {32'hbcdc41a4, 32'hbcd020f7} /* (8, 3, 8) {real, imag} */,
  {32'h3cb0a260, 32'hbd781dd6} /* (8, 3, 7) {real, imag} */,
  {32'hbda6b8dc, 32'h3e21c094} /* (8, 3, 6) {real, imag} */,
  {32'hbe1a1852, 32'h3d6c987e} /* (8, 3, 5) {real, imag} */,
  {32'hbd379860, 32'hbe9e024e} /* (8, 3, 4) {real, imag} */,
  {32'hbd930fd8, 32'hbdc6ccb0} /* (8, 3, 3) {real, imag} */,
  {32'h3e72fcb0, 32'hbf898a86} /* (8, 3, 2) {real, imag} */,
  {32'h40376d5e, 32'h4063b414} /* (8, 3, 1) {real, imag} */,
  {32'h40a4409b, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'h403c7398, 32'hc066e3be} /* (8, 2, 31) {real, imag} */,
  {32'h3ed12c91, 32'h3f904aaa} /* (8, 2, 30) {real, imag} */,
  {32'hbe524b9b, 32'h3e83b49d} /* (8, 2, 29) {real, imag} */,
  {32'hbdca7ed7, 32'h3e8cfafb} /* (8, 2, 28) {real, imag} */,
  {32'hbe207806, 32'hbe317201} /* (8, 2, 27) {real, imag} */,
  {32'hbd30fabc, 32'hbc99d881} /* (8, 2, 26) {real, imag} */,
  {32'h3bfcd010, 32'h3d58de1d} /* (8, 2, 25) {real, imag} */,
  {32'h3ddf1424, 32'h3cff4c00} /* (8, 2, 24) {real, imag} */,
  {32'hbd79b024, 32'h3e0fc2f4} /* (8, 2, 23) {real, imag} */,
  {32'hbd8f6b3e, 32'h3dced0cd} /* (8, 2, 22) {real, imag} */,
  {32'hbdbd0b64, 32'hbdd47202} /* (8, 2, 21) {real, imag} */,
  {32'h3c28d906, 32'hbd8bea5e} /* (8, 2, 20) {real, imag} */,
  {32'h3d1a0d26, 32'hbd8fe42c} /* (8, 2, 19) {real, imag} */,
  {32'h3cad108f, 32'h3ddbd03e} /* (8, 2, 18) {real, imag} */,
  {32'hbc14b2bf, 32'h3d3d1a2e} /* (8, 2, 17) {real, imag} */,
  {32'hbd9ec37e, 32'h00000000} /* (8, 2, 16) {real, imag} */,
  {32'hbc14b2bf, 32'hbd3d1a2e} /* (8, 2, 15) {real, imag} */,
  {32'h3cad108f, 32'hbddbd03e} /* (8, 2, 14) {real, imag} */,
  {32'h3d1a0d26, 32'h3d8fe42c} /* (8, 2, 13) {real, imag} */,
  {32'h3c28d906, 32'h3d8bea5e} /* (8, 2, 12) {real, imag} */,
  {32'hbdbd0b64, 32'h3dd47202} /* (8, 2, 11) {real, imag} */,
  {32'hbd8f6b3e, 32'hbdced0cd} /* (8, 2, 10) {real, imag} */,
  {32'hbd79b024, 32'hbe0fc2f4} /* (8, 2, 9) {real, imag} */,
  {32'h3ddf1424, 32'hbcff4c00} /* (8, 2, 8) {real, imag} */,
  {32'h3bfcd010, 32'hbd58de1d} /* (8, 2, 7) {real, imag} */,
  {32'hbd30fabc, 32'h3c99d881} /* (8, 2, 6) {real, imag} */,
  {32'hbe207806, 32'h3e317201} /* (8, 2, 5) {real, imag} */,
  {32'hbdca7ed7, 32'hbe8cfafb} /* (8, 2, 4) {real, imag} */,
  {32'hbe524b9b, 32'hbe83b49d} /* (8, 2, 3) {real, imag} */,
  {32'h3ed12c91, 32'hbf904aaa} /* (8, 2, 2) {real, imag} */,
  {32'h403c7398, 32'h4066e3be} /* (8, 2, 1) {real, imag} */,
  {32'h40aa85c8, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'h403e08cb, 32'hc053afb8} /* (8, 1, 31) {real, imag} */,
  {32'h3e555dd2, 32'h3f6477b2} /* (8, 1, 30) {real, imag} */,
  {32'hbe767c2c, 32'h3e46b20d} /* (8, 1, 29) {real, imag} */,
  {32'hbd6b0f6b, 32'h3ea55397} /* (8, 1, 28) {real, imag} */,
  {32'hbdca4b50, 32'hbdf60fc3} /* (8, 1, 27) {real, imag} */,
  {32'h3b41ac28, 32'hbd35718a} /* (8, 1, 26) {real, imag} */,
  {32'hbda4cb13, 32'h3d844bea} /* (8, 1, 25) {real, imag} */,
  {32'h3da07628, 32'hbce3e90b} /* (8, 1, 24) {real, imag} */,
  {32'hbc2ca7a2, 32'hbd15d356} /* (8, 1, 23) {real, imag} */,
  {32'h3b7a3a40, 32'h3db809a4} /* (8, 1, 22) {real, imag} */,
  {32'hbd80baea, 32'hbab5ce20} /* (8, 1, 21) {real, imag} */,
  {32'h3da1bb28, 32'hbdd3f0b1} /* (8, 1, 20) {real, imag} */,
  {32'h3cbbb750, 32'h3db21b4e} /* (8, 1, 19) {real, imag} */,
  {32'hbc10fc1c, 32'hbc9248a6} /* (8, 1, 18) {real, imag} */,
  {32'hbca7f013, 32'hbd05877a} /* (8, 1, 17) {real, imag} */,
  {32'hbcac4d0a, 32'h00000000} /* (8, 1, 16) {real, imag} */,
  {32'hbca7f013, 32'h3d05877a} /* (8, 1, 15) {real, imag} */,
  {32'hbc10fc1c, 32'h3c9248a6} /* (8, 1, 14) {real, imag} */,
  {32'h3cbbb750, 32'hbdb21b4e} /* (8, 1, 13) {real, imag} */,
  {32'h3da1bb28, 32'h3dd3f0b1} /* (8, 1, 12) {real, imag} */,
  {32'hbd80baea, 32'h3ab5ce20} /* (8, 1, 11) {real, imag} */,
  {32'h3b7a3a40, 32'hbdb809a4} /* (8, 1, 10) {real, imag} */,
  {32'hbc2ca7a2, 32'h3d15d356} /* (8, 1, 9) {real, imag} */,
  {32'h3da07628, 32'h3ce3e90b} /* (8, 1, 8) {real, imag} */,
  {32'hbda4cb13, 32'hbd844bea} /* (8, 1, 7) {real, imag} */,
  {32'h3b41ac28, 32'h3d35718a} /* (8, 1, 6) {real, imag} */,
  {32'hbdca4b50, 32'h3df60fc3} /* (8, 1, 5) {real, imag} */,
  {32'hbd6b0f6b, 32'hbea55397} /* (8, 1, 4) {real, imag} */,
  {32'hbe767c2c, 32'hbe46b20d} /* (8, 1, 3) {real, imag} */,
  {32'h3e555dd2, 32'hbf6477b2} /* (8, 1, 2) {real, imag} */,
  {32'h403e08cb, 32'h4053afb8} /* (8, 1, 1) {real, imag} */,
  {32'h40a7271f, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'h404677d7, 32'hc02ede9a} /* (8, 0, 31) {real, imag} */,
  {32'hbda4bcc8, 32'h3f3c6c82} /* (8, 0, 30) {real, imag} */,
  {32'hbe5dafcc, 32'h3db2c60e} /* (8, 0, 29) {real, imag} */,
  {32'h3bebb548, 32'h3e77fc34} /* (8, 0, 28) {real, imag} */,
  {32'hbda01cdc, 32'hbdd6c1f9} /* (8, 0, 27) {real, imag} */,
  {32'hbcfde1b8, 32'h3d08944c} /* (8, 0, 26) {real, imag} */,
  {32'hbd845720, 32'hb9f4f340} /* (8, 0, 25) {real, imag} */,
  {32'h3c904328, 32'h3c85d1ce} /* (8, 0, 24) {real, imag} */,
  {32'h37aa2800, 32'h3c46b4c0} /* (8, 0, 23) {real, imag} */,
  {32'hbcbfd260, 32'hbd2b460f} /* (8, 0, 22) {real, imag} */,
  {32'h3d1bd0ff, 32'h3d8d58b7} /* (8, 0, 21) {real, imag} */,
  {32'h3df23c2e, 32'h3bcc47c0} /* (8, 0, 20) {real, imag} */,
  {32'hb8da0d00, 32'hbca4a8a2} /* (8, 0, 19) {real, imag} */,
  {32'hbd0a9f6b, 32'hbd420cbc} /* (8, 0, 18) {real, imag} */,
  {32'h3c81a0e6, 32'h3d4038b4} /* (8, 0, 17) {real, imag} */,
  {32'hbd4c8d7d, 32'h00000000} /* (8, 0, 16) {real, imag} */,
  {32'h3c81a0e6, 32'hbd4038b4} /* (8, 0, 15) {real, imag} */,
  {32'hbd0a9f6b, 32'h3d420cbc} /* (8, 0, 14) {real, imag} */,
  {32'hb8da0d00, 32'h3ca4a8a2} /* (8, 0, 13) {real, imag} */,
  {32'h3df23c2e, 32'hbbcc47c0} /* (8, 0, 12) {real, imag} */,
  {32'h3d1bd0ff, 32'hbd8d58b7} /* (8, 0, 11) {real, imag} */,
  {32'hbcbfd260, 32'h3d2b460f} /* (8, 0, 10) {real, imag} */,
  {32'h37aa2800, 32'hbc46b4c0} /* (8, 0, 9) {real, imag} */,
  {32'h3c904328, 32'hbc85d1ce} /* (8, 0, 8) {real, imag} */,
  {32'hbd845720, 32'h39f4f340} /* (8, 0, 7) {real, imag} */,
  {32'hbcfde1b8, 32'hbd08944c} /* (8, 0, 6) {real, imag} */,
  {32'hbda01cdc, 32'h3dd6c1f9} /* (8, 0, 5) {real, imag} */,
  {32'h3bebb548, 32'hbe77fc34} /* (8, 0, 4) {real, imag} */,
  {32'hbe5dafcc, 32'hbdb2c60e} /* (8, 0, 3) {real, imag} */,
  {32'hbda4bcc8, 32'hbf3c6c82} /* (8, 0, 2) {real, imag} */,
  {32'h404677d7, 32'h402ede9a} /* (8, 0, 1) {real, imag} */,
  {32'h40a025b5, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h4040025a, 32'hbfccfbe4} /* (7, 31, 31) {real, imag} */,
  {32'hbeec3489, 32'h3ec0bdeb} /* (7, 31, 30) {real, imag} */,
  {32'hbdb4f2fb, 32'h3beaf3d0} /* (7, 31, 29) {real, imag} */,
  {32'h3e12c268, 32'h3ceb6df0} /* (7, 31, 28) {real, imag} */,
  {32'hbddb0233, 32'h3d377c51} /* (7, 31, 27) {real, imag} */,
  {32'h3b2d1100, 32'h3d168f05} /* (7, 31, 26) {real, imag} */,
  {32'h3c17efad, 32'h3d37c9c9} /* (7, 31, 25) {real, imag} */,
  {32'hbde83951, 32'h3d2a9963} /* (7, 31, 24) {real, imag} */,
  {32'h3d63eb56, 32'hbd35ff9b} /* (7, 31, 23) {real, imag} */,
  {32'h3da164a9, 32'h3d9577e8} /* (7, 31, 22) {real, imag} */,
  {32'hbdb53de8, 32'h3d8863c6} /* (7, 31, 21) {real, imag} */,
  {32'hbce2382a, 32'hbd1800f8} /* (7, 31, 20) {real, imag} */,
  {32'h3c975308, 32'hbc8544ab} /* (7, 31, 19) {real, imag} */,
  {32'h3cd69e92, 32'h3d4437a9} /* (7, 31, 18) {real, imag} */,
  {32'hbcc38a32, 32'h3c9082b2} /* (7, 31, 17) {real, imag} */,
  {32'hbdb7ead1, 32'h00000000} /* (7, 31, 16) {real, imag} */,
  {32'hbcc38a32, 32'hbc9082b2} /* (7, 31, 15) {real, imag} */,
  {32'h3cd69e92, 32'hbd4437a9} /* (7, 31, 14) {real, imag} */,
  {32'h3c975308, 32'h3c8544ab} /* (7, 31, 13) {real, imag} */,
  {32'hbce2382a, 32'h3d1800f8} /* (7, 31, 12) {real, imag} */,
  {32'hbdb53de8, 32'hbd8863c6} /* (7, 31, 11) {real, imag} */,
  {32'h3da164a9, 32'hbd9577e8} /* (7, 31, 10) {real, imag} */,
  {32'h3d63eb56, 32'h3d35ff9b} /* (7, 31, 9) {real, imag} */,
  {32'hbde83951, 32'hbd2a9963} /* (7, 31, 8) {real, imag} */,
  {32'h3c17efad, 32'hbd37c9c9} /* (7, 31, 7) {real, imag} */,
  {32'h3b2d1100, 32'hbd168f05} /* (7, 31, 6) {real, imag} */,
  {32'hbddb0233, 32'hbd377c51} /* (7, 31, 5) {real, imag} */,
  {32'h3e12c268, 32'hbceb6df0} /* (7, 31, 4) {real, imag} */,
  {32'hbdb4f2fb, 32'hbbeaf3d0} /* (7, 31, 3) {real, imag} */,
  {32'hbeec3489, 32'hbec0bdeb} /* (7, 31, 2) {real, imag} */,
  {32'h4040025a, 32'h3fccfbe4} /* (7, 31, 1) {real, imag} */,
  {32'h408c1258, 32'h00000000} /* (7, 31, 0) {real, imag} */,
  {32'h4066b534, 32'hbf9a89d2} /* (7, 30, 31) {real, imag} */,
  {32'hbf55c914, 32'h3ed71557} /* (7, 30, 30) {real, imag} */,
  {32'hbce77864, 32'h3daaa002} /* (7, 30, 29) {real, imag} */,
  {32'h3e24195a, 32'hbe012400} /* (7, 30, 28) {real, imag} */,
  {32'hbe84f0dd, 32'h3da43f2e} /* (7, 30, 27) {real, imag} */,
  {32'hbd28bcbf, 32'h3e2ace48} /* (7, 30, 26) {real, imag} */,
  {32'h3dc944b6, 32'hbcb6d44a} /* (7, 30, 25) {real, imag} */,
  {32'hbdf09a0e, 32'h3d4c3864} /* (7, 30, 24) {real, imag} */,
  {32'hba8171e0, 32'h3d833542} /* (7, 30, 23) {real, imag} */,
  {32'hbc3646ea, 32'hbbeb80a8} /* (7, 30, 22) {real, imag} */,
  {32'hbda241c0, 32'h3b689c40} /* (7, 30, 21) {real, imag} */,
  {32'hbd748f62, 32'hbd0c0e6c} /* (7, 30, 20) {real, imag} */,
  {32'hbc38de26, 32'hbc986310} /* (7, 30, 19) {real, imag} */,
  {32'hbd1c8da4, 32'hbceaddf0} /* (7, 30, 18) {real, imag} */,
  {32'h3d6a5251, 32'hbdc1e4b8} /* (7, 30, 17) {real, imag} */,
  {32'h3c465dce, 32'h00000000} /* (7, 30, 16) {real, imag} */,
  {32'h3d6a5251, 32'h3dc1e4b8} /* (7, 30, 15) {real, imag} */,
  {32'hbd1c8da4, 32'h3ceaddf0} /* (7, 30, 14) {real, imag} */,
  {32'hbc38de26, 32'h3c986310} /* (7, 30, 13) {real, imag} */,
  {32'hbd748f62, 32'h3d0c0e6c} /* (7, 30, 12) {real, imag} */,
  {32'hbda241c0, 32'hbb689c40} /* (7, 30, 11) {real, imag} */,
  {32'hbc3646ea, 32'h3beb80a8} /* (7, 30, 10) {real, imag} */,
  {32'hba8171e0, 32'hbd833542} /* (7, 30, 9) {real, imag} */,
  {32'hbdf09a0e, 32'hbd4c3864} /* (7, 30, 8) {real, imag} */,
  {32'h3dc944b6, 32'h3cb6d44a} /* (7, 30, 7) {real, imag} */,
  {32'hbd28bcbf, 32'hbe2ace48} /* (7, 30, 6) {real, imag} */,
  {32'hbe84f0dd, 32'hbda43f2e} /* (7, 30, 5) {real, imag} */,
  {32'h3e24195a, 32'h3e012400} /* (7, 30, 4) {real, imag} */,
  {32'hbce77864, 32'hbdaaa002} /* (7, 30, 3) {real, imag} */,
  {32'hbf55c914, 32'hbed71557} /* (7, 30, 2) {real, imag} */,
  {32'h4066b534, 32'h3f9a89d2} /* (7, 30, 1) {real, imag} */,
  {32'h408b44fc, 32'h00000000} /* (7, 30, 0) {real, imag} */,
  {32'h4072cff6, 32'hbf40404c} /* (7, 29, 31) {real, imag} */,
  {32'hbf77c517, 32'h3eeae323} /* (7, 29, 30) {real, imag} */,
  {32'hbd511e34, 32'h3d645fce} /* (7, 29, 29) {real, imag} */,
  {32'h3e25b38e, 32'hbc89ccf8} /* (7, 29, 28) {real, imag} */,
  {32'hbe87f5f2, 32'h3d98ad13} /* (7, 29, 27) {real, imag} */,
  {32'h3c87c220, 32'h3d48adfe} /* (7, 29, 26) {real, imag} */,
  {32'h3d4804fc, 32'hbda3b22e} /* (7, 29, 25) {real, imag} */,
  {32'hbdd521b9, 32'h3e0b633c} /* (7, 29, 24) {real, imag} */,
  {32'h3c92e01a, 32'h3cd09525} /* (7, 29, 23) {real, imag} */,
  {32'hbcfefcc0, 32'hbdf88288} /* (7, 29, 22) {real, imag} */,
  {32'hbd1fa45a, 32'h3d0b30a7} /* (7, 29, 21) {real, imag} */,
  {32'h3dcb71f2, 32'hbd5d91c4} /* (7, 29, 20) {real, imag} */,
  {32'hbcb90438, 32'hbbe1c160} /* (7, 29, 19) {real, imag} */,
  {32'h3d2acae6, 32'h3db169dc} /* (7, 29, 18) {real, imag} */,
  {32'h3d384e3f, 32'hbd84bdd8} /* (7, 29, 17) {real, imag} */,
  {32'hbcf75012, 32'h00000000} /* (7, 29, 16) {real, imag} */,
  {32'h3d384e3f, 32'h3d84bdd8} /* (7, 29, 15) {real, imag} */,
  {32'h3d2acae6, 32'hbdb169dc} /* (7, 29, 14) {real, imag} */,
  {32'hbcb90438, 32'h3be1c160} /* (7, 29, 13) {real, imag} */,
  {32'h3dcb71f2, 32'h3d5d91c4} /* (7, 29, 12) {real, imag} */,
  {32'hbd1fa45a, 32'hbd0b30a7} /* (7, 29, 11) {real, imag} */,
  {32'hbcfefcc0, 32'h3df88288} /* (7, 29, 10) {real, imag} */,
  {32'h3c92e01a, 32'hbcd09525} /* (7, 29, 9) {real, imag} */,
  {32'hbdd521b9, 32'hbe0b633c} /* (7, 29, 8) {real, imag} */,
  {32'h3d4804fc, 32'h3da3b22e} /* (7, 29, 7) {real, imag} */,
  {32'h3c87c220, 32'hbd48adfe} /* (7, 29, 6) {real, imag} */,
  {32'hbe87f5f2, 32'hbd98ad13} /* (7, 29, 5) {real, imag} */,
  {32'h3e25b38e, 32'h3c89ccf8} /* (7, 29, 4) {real, imag} */,
  {32'hbd511e34, 32'hbd645fce} /* (7, 29, 3) {real, imag} */,
  {32'hbf77c517, 32'hbeeae323} /* (7, 29, 2) {real, imag} */,
  {32'h4072cff6, 32'h3f40404c} /* (7, 29, 1) {real, imag} */,
  {32'h408b4dfb, 32'h00000000} /* (7, 29, 0) {real, imag} */,
  {32'h4068e901, 32'hbf27cc3c} /* (7, 28, 31) {real, imag} */,
  {32'hbf87abe7, 32'h3ed434c7} /* (7, 28, 30) {real, imag} */,
  {32'hbce5e9b0, 32'hbdac738f} /* (7, 28, 29) {real, imag} */,
  {32'h3d9a17c3, 32'hbdf52f09} /* (7, 28, 28) {real, imag} */,
  {32'hbe473112, 32'h3d61971a} /* (7, 28, 27) {real, imag} */,
  {32'hbd55064d, 32'h3ceab5f4} /* (7, 28, 26) {real, imag} */,
  {32'hbd338e4c, 32'hbbf79f20} /* (7, 28, 25) {real, imag} */,
  {32'h3d93d0be, 32'hbc44ab5e} /* (7, 28, 24) {real, imag} */,
  {32'h3d188fc4, 32'hbcca0def} /* (7, 28, 23) {real, imag} */,
  {32'h3d9e6f4e, 32'hbd5dbb3e} /* (7, 28, 22) {real, imag} */,
  {32'hbd127367, 32'hbc362100} /* (7, 28, 21) {real, imag} */,
  {32'hbd452726, 32'hbcd67d66} /* (7, 28, 20) {real, imag} */,
  {32'hbd307b57, 32'hbd5909e5} /* (7, 28, 19) {real, imag} */,
  {32'h3d966db5, 32'h3d8151f0} /* (7, 28, 18) {real, imag} */,
  {32'hbc885d8c, 32'h3dc529dc} /* (7, 28, 17) {real, imag} */,
  {32'hbd32e5bc, 32'h00000000} /* (7, 28, 16) {real, imag} */,
  {32'hbc885d8c, 32'hbdc529dc} /* (7, 28, 15) {real, imag} */,
  {32'h3d966db5, 32'hbd8151f0} /* (7, 28, 14) {real, imag} */,
  {32'hbd307b57, 32'h3d5909e5} /* (7, 28, 13) {real, imag} */,
  {32'hbd452726, 32'h3cd67d66} /* (7, 28, 12) {real, imag} */,
  {32'hbd127367, 32'h3c362100} /* (7, 28, 11) {real, imag} */,
  {32'h3d9e6f4e, 32'h3d5dbb3e} /* (7, 28, 10) {real, imag} */,
  {32'h3d188fc4, 32'h3cca0def} /* (7, 28, 9) {real, imag} */,
  {32'h3d93d0be, 32'h3c44ab5e} /* (7, 28, 8) {real, imag} */,
  {32'hbd338e4c, 32'h3bf79f20} /* (7, 28, 7) {real, imag} */,
  {32'hbd55064d, 32'hbceab5f4} /* (7, 28, 6) {real, imag} */,
  {32'hbe473112, 32'hbd61971a} /* (7, 28, 5) {real, imag} */,
  {32'h3d9a17c3, 32'h3df52f09} /* (7, 28, 4) {real, imag} */,
  {32'hbce5e9b0, 32'h3dac738f} /* (7, 28, 3) {real, imag} */,
  {32'hbf87abe7, 32'hbed434c7} /* (7, 28, 2) {real, imag} */,
  {32'h4068e901, 32'h3f27cc3c} /* (7, 28, 1) {real, imag} */,
  {32'h408b3e54, 32'h00000000} /* (7, 28, 0) {real, imag} */,
  {32'h406b4ea4, 32'hbf181e02} /* (7, 27, 31) {real, imag} */,
  {32'hbf9be5a2, 32'h3ebbb596} /* (7, 27, 30) {real, imag} */,
  {32'hbbd8bfbc, 32'hbce5ec5d} /* (7, 27, 29) {real, imag} */,
  {32'h3e2cf618, 32'hbe0d2dca} /* (7, 27, 28) {real, imag} */,
  {32'hbe41356e, 32'h3d8900da} /* (7, 27, 27) {real, imag} */,
  {32'hbd0e69cb, 32'hbcb0c138} /* (7, 27, 26) {real, imag} */,
  {32'h3e080b78, 32'hbd8e0415} /* (7, 27, 25) {real, imag} */,
  {32'h38d1e200, 32'hbb8b5bb0} /* (7, 27, 24) {real, imag} */,
  {32'h3cadebfa, 32'hbd525cdc} /* (7, 27, 23) {real, imag} */,
  {32'hbc14885e, 32'hbc1fe0ae} /* (7, 27, 22) {real, imag} */,
  {32'hbcf08534, 32'h3d9b34b4} /* (7, 27, 21) {real, imag} */,
  {32'hbc591ec2, 32'hbd80e4ed} /* (7, 27, 20) {real, imag} */,
  {32'hbcf26f8e, 32'hbd918150} /* (7, 27, 19) {real, imag} */,
  {32'hbcecbb64, 32'h3da83bce} /* (7, 27, 18) {real, imag} */,
  {32'hbb89822c, 32'h3d17f8f1} /* (7, 27, 17) {real, imag} */,
  {32'hbc512d1a, 32'h00000000} /* (7, 27, 16) {real, imag} */,
  {32'hbb89822c, 32'hbd17f8f1} /* (7, 27, 15) {real, imag} */,
  {32'hbcecbb64, 32'hbda83bce} /* (7, 27, 14) {real, imag} */,
  {32'hbcf26f8e, 32'h3d918150} /* (7, 27, 13) {real, imag} */,
  {32'hbc591ec2, 32'h3d80e4ed} /* (7, 27, 12) {real, imag} */,
  {32'hbcf08534, 32'hbd9b34b4} /* (7, 27, 11) {real, imag} */,
  {32'hbc14885e, 32'h3c1fe0ae} /* (7, 27, 10) {real, imag} */,
  {32'h3cadebfa, 32'h3d525cdc} /* (7, 27, 9) {real, imag} */,
  {32'h38d1e200, 32'h3b8b5bb0} /* (7, 27, 8) {real, imag} */,
  {32'h3e080b78, 32'h3d8e0415} /* (7, 27, 7) {real, imag} */,
  {32'hbd0e69cb, 32'h3cb0c138} /* (7, 27, 6) {real, imag} */,
  {32'hbe41356e, 32'hbd8900da} /* (7, 27, 5) {real, imag} */,
  {32'h3e2cf618, 32'h3e0d2dca} /* (7, 27, 4) {real, imag} */,
  {32'hbbd8bfbc, 32'h3ce5ec5d} /* (7, 27, 3) {real, imag} */,
  {32'hbf9be5a2, 32'hbebbb596} /* (7, 27, 2) {real, imag} */,
  {32'h406b4ea4, 32'h3f181e02} /* (7, 27, 1) {real, imag} */,
  {32'h4084142f, 32'h00000000} /* (7, 27, 0) {real, imag} */,
  {32'h40635b62, 32'hbf1e0339} /* (7, 26, 31) {real, imag} */,
  {32'hbfa7e94e, 32'h3e62ae04} /* (7, 26, 30) {real, imag} */,
  {32'h3d855c09, 32'hbda3a92e} /* (7, 26, 29) {real, imag} */,
  {32'h3dddb3c7, 32'h3d40f13b} /* (7, 26, 28) {real, imag} */,
  {32'hbe3f86f9, 32'h3d7ab970} /* (7, 26, 27) {real, imag} */,
  {32'h3d47156c, 32'h3c1a5070} /* (7, 26, 26) {real, imag} */,
  {32'h3db71dfb, 32'hbce55240} /* (7, 26, 25) {real, imag} */,
  {32'h3c904280, 32'h3dc8635a} /* (7, 26, 24) {real, imag} */,
  {32'h3dedfa52, 32'h3d311cbf} /* (7, 26, 23) {real, imag} */,
  {32'h3b949020, 32'hbcc7f18c} /* (7, 26, 22) {real, imag} */,
  {32'h3d90585e, 32'h3d542a37} /* (7, 26, 21) {real, imag} */,
  {32'h3bd19c18, 32'h3c11f58a} /* (7, 26, 20) {real, imag} */,
  {32'h3d25fe36, 32'hbc8472c1} /* (7, 26, 19) {real, imag} */,
  {32'h3c191008, 32'h3c767270} /* (7, 26, 18) {real, imag} */,
  {32'h3c481f9a, 32'h3c6ab9c8} /* (7, 26, 17) {real, imag} */,
  {32'hbd761b5a, 32'h00000000} /* (7, 26, 16) {real, imag} */,
  {32'h3c481f9a, 32'hbc6ab9c8} /* (7, 26, 15) {real, imag} */,
  {32'h3c191008, 32'hbc767270} /* (7, 26, 14) {real, imag} */,
  {32'h3d25fe36, 32'h3c8472c1} /* (7, 26, 13) {real, imag} */,
  {32'h3bd19c18, 32'hbc11f58a} /* (7, 26, 12) {real, imag} */,
  {32'h3d90585e, 32'hbd542a37} /* (7, 26, 11) {real, imag} */,
  {32'h3b949020, 32'h3cc7f18c} /* (7, 26, 10) {real, imag} */,
  {32'h3dedfa52, 32'hbd311cbf} /* (7, 26, 9) {real, imag} */,
  {32'h3c904280, 32'hbdc8635a} /* (7, 26, 8) {real, imag} */,
  {32'h3db71dfb, 32'h3ce55240} /* (7, 26, 7) {real, imag} */,
  {32'h3d47156c, 32'hbc1a5070} /* (7, 26, 6) {real, imag} */,
  {32'hbe3f86f9, 32'hbd7ab970} /* (7, 26, 5) {real, imag} */,
  {32'h3dddb3c7, 32'hbd40f13b} /* (7, 26, 4) {real, imag} */,
  {32'h3d855c09, 32'h3da3a92e} /* (7, 26, 3) {real, imag} */,
  {32'hbfa7e94e, 32'hbe62ae04} /* (7, 26, 2) {real, imag} */,
  {32'h40635b62, 32'h3f1e0339} /* (7, 26, 1) {real, imag} */,
  {32'h407ea796, 32'h00000000} /* (7, 26, 0) {real, imag} */,
  {32'h4052f8ef, 32'hbf0d4b01} /* (7, 25, 31) {real, imag} */,
  {32'hbfaa006c, 32'h3e532284} /* (7, 25, 30) {real, imag} */,
  {32'hbcb37b88, 32'hbdf19597} /* (7, 25, 29) {real, imag} */,
  {32'h3e41f538, 32'hbc7e0be8} /* (7, 25, 28) {real, imag} */,
  {32'hbe4a75f3, 32'h3de9cf4c} /* (7, 25, 27) {real, imag} */,
  {32'h3cb92754, 32'hbcb49783} /* (7, 25, 26) {real, imag} */,
  {32'h3c6a8085, 32'hbe0f02cc} /* (7, 25, 25) {real, imag} */,
  {32'hbc87c573, 32'h3d16c24f} /* (7, 25, 24) {real, imag} */,
  {32'hbd478511, 32'hbd300a7a} /* (7, 25, 23) {real, imag} */,
  {32'h3b2ddea8, 32'h3d01d1d5} /* (7, 25, 22) {real, imag} */,
  {32'hbc4e7c3a, 32'h3d0f2556} /* (7, 25, 21) {real, imag} */,
  {32'hbc5acfde, 32'hbe2254f5} /* (7, 25, 20) {real, imag} */,
  {32'h3ce65905, 32'h3de66013} /* (7, 25, 19) {real, imag} */,
  {32'hbddff83e, 32'hbda5b1d5} /* (7, 25, 18) {real, imag} */,
  {32'hbc220340, 32'h3c84ebc4} /* (7, 25, 17) {real, imag} */,
  {32'hbbd87890, 32'h00000000} /* (7, 25, 16) {real, imag} */,
  {32'hbc220340, 32'hbc84ebc4} /* (7, 25, 15) {real, imag} */,
  {32'hbddff83e, 32'h3da5b1d5} /* (7, 25, 14) {real, imag} */,
  {32'h3ce65905, 32'hbde66013} /* (7, 25, 13) {real, imag} */,
  {32'hbc5acfde, 32'h3e2254f5} /* (7, 25, 12) {real, imag} */,
  {32'hbc4e7c3a, 32'hbd0f2556} /* (7, 25, 11) {real, imag} */,
  {32'h3b2ddea8, 32'hbd01d1d5} /* (7, 25, 10) {real, imag} */,
  {32'hbd478511, 32'h3d300a7a} /* (7, 25, 9) {real, imag} */,
  {32'hbc87c573, 32'hbd16c24f} /* (7, 25, 8) {real, imag} */,
  {32'h3c6a8085, 32'h3e0f02cc} /* (7, 25, 7) {real, imag} */,
  {32'h3cb92754, 32'h3cb49783} /* (7, 25, 6) {real, imag} */,
  {32'hbe4a75f3, 32'hbde9cf4c} /* (7, 25, 5) {real, imag} */,
  {32'h3e41f538, 32'h3c7e0be8} /* (7, 25, 4) {real, imag} */,
  {32'hbcb37b88, 32'h3df19597} /* (7, 25, 3) {real, imag} */,
  {32'hbfaa006c, 32'hbe532284} /* (7, 25, 2) {real, imag} */,
  {32'h4052f8ef, 32'h3f0d4b01} /* (7, 25, 1) {real, imag} */,
  {32'h406cb6e8, 32'h00000000} /* (7, 25, 0) {real, imag} */,
  {32'h403e5a3c, 32'hbf0cd597} /* (7, 24, 31) {real, imag} */,
  {32'hbfa5062a, 32'h3e894126} /* (7, 24, 30) {real, imag} */,
  {32'hbb947940, 32'hbdccac0b} /* (7, 24, 29) {real, imag} */,
  {32'h3e5304f9, 32'h3cbcc8d4} /* (7, 24, 28) {real, imag} */,
  {32'hbe76e830, 32'h3db75c64} /* (7, 24, 27) {real, imag} */,
  {32'hbd3f0673, 32'hbcc92ea0} /* (7, 24, 26) {real, imag} */,
  {32'h3cb95561, 32'hbd921ff0} /* (7, 24, 25) {real, imag} */,
  {32'hbdda6491, 32'hbd05d5fc} /* (7, 24, 24) {real, imag} */,
  {32'hbb177ad0, 32'h3c0945a8} /* (7, 24, 23) {real, imag} */,
  {32'hbd62c36c, 32'hbe11474e} /* (7, 24, 22) {real, imag} */,
  {32'hbc7cf000, 32'hbc00bbde} /* (7, 24, 21) {real, imag} */,
  {32'hbc5e6c6e, 32'h3e2c8900} /* (7, 24, 20) {real, imag} */,
  {32'hbd2ac1bb, 32'hbdd8ae27} /* (7, 24, 19) {real, imag} */,
  {32'h3dc16f9f, 32'h3d305ab0} /* (7, 24, 18) {real, imag} */,
  {32'h3bc5da5e, 32'hbcc03034} /* (7, 24, 17) {real, imag} */,
  {32'hbc8ccc17, 32'h00000000} /* (7, 24, 16) {real, imag} */,
  {32'h3bc5da5e, 32'h3cc03034} /* (7, 24, 15) {real, imag} */,
  {32'h3dc16f9f, 32'hbd305ab0} /* (7, 24, 14) {real, imag} */,
  {32'hbd2ac1bb, 32'h3dd8ae27} /* (7, 24, 13) {real, imag} */,
  {32'hbc5e6c6e, 32'hbe2c8900} /* (7, 24, 12) {real, imag} */,
  {32'hbc7cf000, 32'h3c00bbde} /* (7, 24, 11) {real, imag} */,
  {32'hbd62c36c, 32'h3e11474e} /* (7, 24, 10) {real, imag} */,
  {32'hbb177ad0, 32'hbc0945a8} /* (7, 24, 9) {real, imag} */,
  {32'hbdda6491, 32'h3d05d5fc} /* (7, 24, 8) {real, imag} */,
  {32'h3cb95561, 32'h3d921ff0} /* (7, 24, 7) {real, imag} */,
  {32'hbd3f0673, 32'h3cc92ea0} /* (7, 24, 6) {real, imag} */,
  {32'hbe76e830, 32'hbdb75c64} /* (7, 24, 5) {real, imag} */,
  {32'h3e5304f9, 32'hbcbcc8d4} /* (7, 24, 4) {real, imag} */,
  {32'hbb947940, 32'h3dccac0b} /* (7, 24, 3) {real, imag} */,
  {32'hbfa5062a, 32'hbe894126} /* (7, 24, 2) {real, imag} */,
  {32'h403e5a3c, 32'h3f0cd597} /* (7, 24, 1) {real, imag} */,
  {32'h405728b6, 32'h00000000} /* (7, 24, 0) {real, imag} */,
  {32'h401615f4, 32'hbedffe5a} /* (7, 23, 31) {real, imag} */,
  {32'hbf8b8830, 32'h3e5403ee} /* (7, 23, 30) {real, imag} */,
  {32'hbe37449a, 32'hbe2a93d2} /* (7, 23, 29) {real, imag} */,
  {32'h3de3b5ba, 32'hbcff1904} /* (7, 23, 28) {real, imag} */,
  {32'hbe025bdf, 32'h3d97ef0a} /* (7, 23, 27) {real, imag} */,
  {32'h3dcda87b, 32'h3c9c31a2} /* (7, 23, 26) {real, imag} */,
  {32'hbc35771c, 32'hbbb64912} /* (7, 23, 25) {real, imag} */,
  {32'hbd9e7f8d, 32'hbd119360} /* (7, 23, 24) {real, imag} */,
  {32'hbd89866f, 32'h3d88b392} /* (7, 23, 23) {real, imag} */,
  {32'hbcfa7dc2, 32'hbd024b2f} /* (7, 23, 22) {real, imag} */,
  {32'h3d83a163, 32'h3c56b792} /* (7, 23, 21) {real, imag} */,
  {32'h3ca3aacd, 32'h3d33dac8} /* (7, 23, 20) {real, imag} */,
  {32'h3b4562d8, 32'hbc3813c2} /* (7, 23, 19) {real, imag} */,
  {32'h3ced6a9a, 32'h3c91dd31} /* (7, 23, 18) {real, imag} */,
  {32'hbc3fb4a2, 32'hbd29c6e0} /* (7, 23, 17) {real, imag} */,
  {32'hbb9abfdc, 32'h00000000} /* (7, 23, 16) {real, imag} */,
  {32'hbc3fb4a2, 32'h3d29c6e0} /* (7, 23, 15) {real, imag} */,
  {32'h3ced6a9a, 32'hbc91dd31} /* (7, 23, 14) {real, imag} */,
  {32'h3b4562d8, 32'h3c3813c2} /* (7, 23, 13) {real, imag} */,
  {32'h3ca3aacd, 32'hbd33dac8} /* (7, 23, 12) {real, imag} */,
  {32'h3d83a163, 32'hbc56b792} /* (7, 23, 11) {real, imag} */,
  {32'hbcfa7dc2, 32'h3d024b2f} /* (7, 23, 10) {real, imag} */,
  {32'hbd89866f, 32'hbd88b392} /* (7, 23, 9) {real, imag} */,
  {32'hbd9e7f8d, 32'h3d119360} /* (7, 23, 8) {real, imag} */,
  {32'hbc35771c, 32'h3bb64912} /* (7, 23, 7) {real, imag} */,
  {32'h3dcda87b, 32'hbc9c31a2} /* (7, 23, 6) {real, imag} */,
  {32'hbe025bdf, 32'hbd97ef0a} /* (7, 23, 5) {real, imag} */,
  {32'h3de3b5ba, 32'h3cff1904} /* (7, 23, 4) {real, imag} */,
  {32'hbe37449a, 32'h3e2a93d2} /* (7, 23, 3) {real, imag} */,
  {32'hbf8b8830, 32'hbe5403ee} /* (7, 23, 2) {real, imag} */,
  {32'h401615f4, 32'h3edffe5a} /* (7, 23, 1) {real, imag} */,
  {32'h4039a5ac, 32'h00000000} /* (7, 23, 0) {real, imag} */,
  {32'h3fc5234c, 32'hbe9ed4b8} /* (7, 22, 31) {real, imag} */,
  {32'hbf6db420, 32'h3e1a86c0} /* (7, 22, 30) {real, imag} */,
  {32'hbe4eb3a0, 32'hbe5382fa} /* (7, 22, 29) {real, imag} */,
  {32'h3e0d5be6, 32'hbcde9d36} /* (7, 22, 28) {real, imag} */,
  {32'hbe1bf16d, 32'h3e24122b} /* (7, 22, 27) {real, imag} */,
  {32'h3ac6ab00, 32'h3d955aca} /* (7, 22, 26) {real, imag} */,
  {32'h3dafc747, 32'hbd80da0a} /* (7, 22, 25) {real, imag} */,
  {32'hbde22e2e, 32'h3b57fa90} /* (7, 22, 24) {real, imag} */,
  {32'h3d4cfb04, 32'h38404800} /* (7, 22, 23) {real, imag} */,
  {32'hbdca76a7, 32'hbd473338} /* (7, 22, 22) {real, imag} */,
  {32'hbcd038e0, 32'hbd6be4b2} /* (7, 22, 21) {real, imag} */,
  {32'h3ba36798, 32'hbd8904d5} /* (7, 22, 20) {real, imag} */,
  {32'h3e1c96e5, 32'h3d844691} /* (7, 22, 19) {real, imag} */,
  {32'hbd1e80e6, 32'hbd9b7893} /* (7, 22, 18) {real, imag} */,
  {32'h3954d780, 32'hbbc97988} /* (7, 22, 17) {real, imag} */,
  {32'hbbaf4cda, 32'h00000000} /* (7, 22, 16) {real, imag} */,
  {32'h3954d780, 32'h3bc97988} /* (7, 22, 15) {real, imag} */,
  {32'hbd1e80e6, 32'h3d9b7893} /* (7, 22, 14) {real, imag} */,
  {32'h3e1c96e5, 32'hbd844691} /* (7, 22, 13) {real, imag} */,
  {32'h3ba36798, 32'h3d8904d5} /* (7, 22, 12) {real, imag} */,
  {32'hbcd038e0, 32'h3d6be4b2} /* (7, 22, 11) {real, imag} */,
  {32'hbdca76a7, 32'h3d473338} /* (7, 22, 10) {real, imag} */,
  {32'h3d4cfb04, 32'hb8404800} /* (7, 22, 9) {real, imag} */,
  {32'hbde22e2e, 32'hbb57fa90} /* (7, 22, 8) {real, imag} */,
  {32'h3dafc747, 32'h3d80da0a} /* (7, 22, 7) {real, imag} */,
  {32'h3ac6ab00, 32'hbd955aca} /* (7, 22, 6) {real, imag} */,
  {32'hbe1bf16d, 32'hbe24122b} /* (7, 22, 5) {real, imag} */,
  {32'h3e0d5be6, 32'h3cde9d36} /* (7, 22, 4) {real, imag} */,
  {32'hbe4eb3a0, 32'h3e5382fa} /* (7, 22, 3) {real, imag} */,
  {32'hbf6db420, 32'hbe1a86c0} /* (7, 22, 2) {real, imag} */,
  {32'h3fc5234c, 32'h3e9ed4b8} /* (7, 22, 1) {real, imag} */,
  {32'h400d3684, 32'h00000000} /* (7, 22, 0) {real, imag} */,
  {32'h3ee38668, 32'hbe442e3e} /* (7, 21, 31) {real, imag} */,
  {32'hbe993d1b, 32'hbe3ea792} /* (7, 21, 30) {real, imag} */,
  {32'hbdeed2ed, 32'hbe0d0030} /* (7, 21, 29) {real, imag} */,
  {32'h3ddf90a3, 32'h3d79cd54} /* (7, 21, 28) {real, imag} */,
  {32'hbe0414d0, 32'h3dff32e4} /* (7, 21, 27) {real, imag} */,
  {32'hbc32da22, 32'h3d605948} /* (7, 21, 26) {real, imag} */,
  {32'h3d3d21d0, 32'hbdd255fa} /* (7, 21, 25) {real, imag} */,
  {32'hbd923c1a, 32'hbd759ad7} /* (7, 21, 24) {real, imag} */,
  {32'hbd24d22e, 32'h3af0b328} /* (7, 21, 23) {real, imag} */,
  {32'h3d11f378, 32'h3d5d0e27} /* (7, 21, 22) {real, imag} */,
  {32'hbdbcd9bc, 32'h3d6d7de1} /* (7, 21, 21) {real, imag} */,
  {32'h3d260fb0, 32'h3cb36750} /* (7, 21, 20) {real, imag} */,
  {32'hbc7df13c, 32'h3d03fab4} /* (7, 21, 19) {real, imag} */,
  {32'h3dd41fae, 32'hbce1427a} /* (7, 21, 18) {real, imag} */,
  {32'h3d01ae96, 32'hbcf30e64} /* (7, 21, 17) {real, imag} */,
  {32'hbdbd2f0d, 32'h00000000} /* (7, 21, 16) {real, imag} */,
  {32'h3d01ae96, 32'h3cf30e64} /* (7, 21, 15) {real, imag} */,
  {32'h3dd41fae, 32'h3ce1427a} /* (7, 21, 14) {real, imag} */,
  {32'hbc7df13c, 32'hbd03fab4} /* (7, 21, 13) {real, imag} */,
  {32'h3d260fb0, 32'hbcb36750} /* (7, 21, 12) {real, imag} */,
  {32'hbdbcd9bc, 32'hbd6d7de1} /* (7, 21, 11) {real, imag} */,
  {32'h3d11f378, 32'hbd5d0e27} /* (7, 21, 10) {real, imag} */,
  {32'hbd24d22e, 32'hbaf0b328} /* (7, 21, 9) {real, imag} */,
  {32'hbd923c1a, 32'h3d759ad7} /* (7, 21, 8) {real, imag} */,
  {32'h3d3d21d0, 32'h3dd255fa} /* (7, 21, 7) {real, imag} */,
  {32'hbc32da22, 32'hbd605948} /* (7, 21, 6) {real, imag} */,
  {32'hbe0414d0, 32'hbdff32e4} /* (7, 21, 5) {real, imag} */,
  {32'h3ddf90a3, 32'hbd79cd54} /* (7, 21, 4) {real, imag} */,
  {32'hbdeed2ed, 32'h3e0d0030} /* (7, 21, 3) {real, imag} */,
  {32'hbe993d1b, 32'h3e3ea792} /* (7, 21, 2) {real, imag} */,
  {32'h3ee38668, 32'h3e442e3e} /* (7, 21, 1) {real, imag} */,
  {32'h3f9be120, 32'h00000000} /* (7, 21, 0) {real, imag} */,
  {32'hbf828468, 32'hbbf4bc80} /* (7, 20, 31) {real, imag} */,
  {32'h3ef964bc, 32'hbeaad63d} /* (7, 20, 30) {real, imag} */,
  {32'hbe1f2986, 32'hbdf38038} /* (7, 20, 29) {real, imag} */,
  {32'hbe006c99, 32'h3dbd086b} /* (7, 20, 28) {real, imag} */,
  {32'h3e399d10, 32'hbdbc72c8} /* (7, 20, 27) {real, imag} */,
  {32'h3cdcd04e, 32'hbd40d529} /* (7, 20, 26) {real, imag} */,
  {32'h3d1677a8, 32'hbc9175b8} /* (7, 20, 25) {real, imag} */,
  {32'h3b828ec8, 32'hbcc445cc} /* (7, 20, 24) {real, imag} */,
  {32'h3d0df310, 32'hbd29b2b6} /* (7, 20, 23) {real, imag} */,
  {32'hbe0e09d6, 32'h3c2f7444} /* (7, 20, 22) {real, imag} */,
  {32'hbd50de3c, 32'hbc713562} /* (7, 20, 21) {real, imag} */,
  {32'hbc971ab4, 32'hbcb143c2} /* (7, 20, 20) {real, imag} */,
  {32'h3b399690, 32'hbce8863f} /* (7, 20, 19) {real, imag} */,
  {32'h3dc3e7ce, 32'h3d186284} /* (7, 20, 18) {real, imag} */,
  {32'h3c458735, 32'hbc322812} /* (7, 20, 17) {real, imag} */,
  {32'h3d2f06c7, 32'h00000000} /* (7, 20, 16) {real, imag} */,
  {32'h3c458735, 32'h3c322812} /* (7, 20, 15) {real, imag} */,
  {32'h3dc3e7ce, 32'hbd186284} /* (7, 20, 14) {real, imag} */,
  {32'h3b399690, 32'h3ce8863f} /* (7, 20, 13) {real, imag} */,
  {32'hbc971ab4, 32'h3cb143c2} /* (7, 20, 12) {real, imag} */,
  {32'hbd50de3c, 32'h3c713562} /* (7, 20, 11) {real, imag} */,
  {32'hbe0e09d6, 32'hbc2f7444} /* (7, 20, 10) {real, imag} */,
  {32'h3d0df310, 32'h3d29b2b6} /* (7, 20, 9) {real, imag} */,
  {32'h3b828ec8, 32'h3cc445cc} /* (7, 20, 8) {real, imag} */,
  {32'h3d1677a8, 32'h3c9175b8} /* (7, 20, 7) {real, imag} */,
  {32'h3cdcd04e, 32'h3d40d529} /* (7, 20, 6) {real, imag} */,
  {32'h3e399d10, 32'h3dbc72c8} /* (7, 20, 5) {real, imag} */,
  {32'hbe006c99, 32'hbdbd086b} /* (7, 20, 4) {real, imag} */,
  {32'hbe1f2986, 32'h3df38038} /* (7, 20, 3) {real, imag} */,
  {32'h3ef964bc, 32'h3eaad63d} /* (7, 20, 2) {real, imag} */,
  {32'hbf828468, 32'h3bf4bc80} /* (7, 20, 1) {real, imag} */,
  {32'hbe9662c2, 32'h00000000} /* (7, 20, 0) {real, imag} */,
  {32'hc00413f1, 32'h3e0355e8} /* (7, 19, 31) {real, imag} */,
  {32'h3f7ae556, 32'hbe948bc9} /* (7, 19, 30) {real, imag} */,
  {32'hbe78a950, 32'hbdea6319} /* (7, 19, 29) {real, imag} */,
  {32'hbe233889, 32'hbd61a246} /* (7, 19, 28) {real, imag} */,
  {32'h3e4910c9, 32'hbdebb60c} /* (7, 19, 27) {real, imag} */,
  {32'h3d0ddc60, 32'hbc63666d} /* (7, 19, 26) {real, imag} */,
  {32'hbd2eba4d, 32'h3d74ca4c} /* (7, 19, 25) {real, imag} */,
  {32'h3b0c0f68, 32'h3c9a073c} /* (7, 19, 24) {real, imag} */,
  {32'hbb224b90, 32'hbdc84baa} /* (7, 19, 23) {real, imag} */,
  {32'hbcf2b706, 32'hbcb1a0a6} /* (7, 19, 22) {real, imag} */,
  {32'h3db155e5, 32'h3d86252c} /* (7, 19, 21) {real, imag} */,
  {32'h3c6abc52, 32'h3d1f471e} /* (7, 19, 20) {real, imag} */,
  {32'hbc8617d0, 32'hbd95c002} /* (7, 19, 19) {real, imag} */,
  {32'h3da1b958, 32'hbd169c82} /* (7, 19, 18) {real, imag} */,
  {32'h3bad6bcd, 32'h3d5e07e8} /* (7, 19, 17) {real, imag} */,
  {32'hbdcebd75, 32'h00000000} /* (7, 19, 16) {real, imag} */,
  {32'h3bad6bcd, 32'hbd5e07e8} /* (7, 19, 15) {real, imag} */,
  {32'h3da1b958, 32'h3d169c82} /* (7, 19, 14) {real, imag} */,
  {32'hbc8617d0, 32'h3d95c002} /* (7, 19, 13) {real, imag} */,
  {32'h3c6abc52, 32'hbd1f471e} /* (7, 19, 12) {real, imag} */,
  {32'h3db155e5, 32'hbd86252c} /* (7, 19, 11) {real, imag} */,
  {32'hbcf2b706, 32'h3cb1a0a6} /* (7, 19, 10) {real, imag} */,
  {32'hbb224b90, 32'h3dc84baa} /* (7, 19, 9) {real, imag} */,
  {32'h3b0c0f68, 32'hbc9a073c} /* (7, 19, 8) {real, imag} */,
  {32'hbd2eba4d, 32'hbd74ca4c} /* (7, 19, 7) {real, imag} */,
  {32'h3d0ddc60, 32'h3c63666d} /* (7, 19, 6) {real, imag} */,
  {32'h3e4910c9, 32'h3debb60c} /* (7, 19, 5) {real, imag} */,
  {32'hbe233889, 32'h3d61a246} /* (7, 19, 4) {real, imag} */,
  {32'hbe78a950, 32'h3dea6319} /* (7, 19, 3) {real, imag} */,
  {32'h3f7ae556, 32'h3e948bc9} /* (7, 19, 2) {real, imag} */,
  {32'hc00413f1, 32'hbe0355e8} /* (7, 19, 1) {real, imag} */,
  {32'hbf7730ad, 32'h00000000} /* (7, 19, 0) {real, imag} */,
  {32'hc0332d74, 32'h3e87144d} /* (7, 18, 31) {real, imag} */,
  {32'h3f925f32, 32'hbe9a345a} /* (7, 18, 30) {real, imag} */,
  {32'hbe39f1dc, 32'hbd02e0cd} /* (7, 18, 29) {real, imag} */,
  {32'hbde6ab1b, 32'hbc8dc118} /* (7, 18, 28) {real, imag} */,
  {32'h3dd87f34, 32'hbbd3c380} /* (7, 18, 27) {real, imag} */,
  {32'h3e15d629, 32'h3c6c8256} /* (7, 18, 26) {real, imag} */,
  {32'hbd83cbac, 32'h3b780dac} /* (7, 18, 25) {real, imag} */,
  {32'h3d19a0be, 32'h3d4c5edf} /* (7, 18, 24) {real, imag} */,
  {32'h3d681c90, 32'hbdedcfbe} /* (7, 18, 23) {real, imag} */,
  {32'h3d16de82, 32'h3dd590dc} /* (7, 18, 22) {real, imag} */,
  {32'hbd254cb8, 32'hbe42ec8f} /* (7, 18, 21) {real, imag} */,
  {32'hbd003f76, 32'h3c01dbac} /* (7, 18, 20) {real, imag} */,
  {32'hbc402f5a, 32'hbd647d76} /* (7, 18, 19) {real, imag} */,
  {32'h3be5f51c, 32'hbbc1b570} /* (7, 18, 18) {real, imag} */,
  {32'h3c919d0e, 32'hbc3975d4} /* (7, 18, 17) {real, imag} */,
  {32'hbd3e2680, 32'h00000000} /* (7, 18, 16) {real, imag} */,
  {32'h3c919d0e, 32'h3c3975d4} /* (7, 18, 15) {real, imag} */,
  {32'h3be5f51c, 32'h3bc1b570} /* (7, 18, 14) {real, imag} */,
  {32'hbc402f5a, 32'h3d647d76} /* (7, 18, 13) {real, imag} */,
  {32'hbd003f76, 32'hbc01dbac} /* (7, 18, 12) {real, imag} */,
  {32'hbd254cb8, 32'h3e42ec8f} /* (7, 18, 11) {real, imag} */,
  {32'h3d16de82, 32'hbdd590dc} /* (7, 18, 10) {real, imag} */,
  {32'h3d681c90, 32'h3dedcfbe} /* (7, 18, 9) {real, imag} */,
  {32'h3d19a0be, 32'hbd4c5edf} /* (7, 18, 8) {real, imag} */,
  {32'hbd83cbac, 32'hbb780dac} /* (7, 18, 7) {real, imag} */,
  {32'h3e15d629, 32'hbc6c8256} /* (7, 18, 6) {real, imag} */,
  {32'h3dd87f34, 32'h3bd3c380} /* (7, 18, 5) {real, imag} */,
  {32'hbde6ab1b, 32'h3c8dc118} /* (7, 18, 4) {real, imag} */,
  {32'hbe39f1dc, 32'h3d02e0cd} /* (7, 18, 3) {real, imag} */,
  {32'h3f925f32, 32'h3e9a345a} /* (7, 18, 2) {real, imag} */,
  {32'hc0332d74, 32'hbe87144d} /* (7, 18, 1) {real, imag} */,
  {32'hbfcd2b7f, 32'h00000000} /* (7, 18, 0) {real, imag} */,
  {32'hc049cf34, 32'h3e93a56d} /* (7, 17, 31) {real, imag} */,
  {32'h3f919d4a, 32'hbe9f6a7e} /* (7, 17, 30) {real, imag} */,
  {32'hbd741a9c, 32'hbd372b08} /* (7, 17, 29) {real, imag} */,
  {32'hbe24bf63, 32'hbcebeb36} /* (7, 17, 28) {real, imag} */,
  {32'h3e5837d6, 32'h3da348ae} /* (7, 17, 27) {real, imag} */,
  {32'h3db5cc6c, 32'h3d6c9fe5} /* (7, 17, 26) {real, imag} */,
  {32'h3d9b8e89, 32'h3d38e983} /* (7, 17, 25) {real, imag} */,
  {32'h3d24891b, 32'hbd242e3f} /* (7, 17, 24) {real, imag} */,
  {32'h3d9d6d7d, 32'h3e0276aa} /* (7, 17, 23) {real, imag} */,
  {32'h3c3f56d6, 32'hbcec7159} /* (7, 17, 22) {real, imag} */,
  {32'h3d948902, 32'hbdc6ea42} /* (7, 17, 21) {real, imag} */,
  {32'hbe04631c, 32'hbd30c80a} /* (7, 17, 20) {real, imag} */,
  {32'h3bb08e42, 32'hbd48f26c} /* (7, 17, 19) {real, imag} */,
  {32'hbb18b218, 32'h3d164830} /* (7, 17, 18) {real, imag} */,
  {32'h3d026ed4, 32'hbb134cf0} /* (7, 17, 17) {real, imag} */,
  {32'hbcdb1b78, 32'h00000000} /* (7, 17, 16) {real, imag} */,
  {32'h3d026ed4, 32'h3b134cf0} /* (7, 17, 15) {real, imag} */,
  {32'hbb18b218, 32'hbd164830} /* (7, 17, 14) {real, imag} */,
  {32'h3bb08e42, 32'h3d48f26c} /* (7, 17, 13) {real, imag} */,
  {32'hbe04631c, 32'h3d30c80a} /* (7, 17, 12) {real, imag} */,
  {32'h3d948902, 32'h3dc6ea42} /* (7, 17, 11) {real, imag} */,
  {32'h3c3f56d6, 32'h3cec7159} /* (7, 17, 10) {real, imag} */,
  {32'h3d9d6d7d, 32'hbe0276aa} /* (7, 17, 9) {real, imag} */,
  {32'h3d24891b, 32'h3d242e3f} /* (7, 17, 8) {real, imag} */,
  {32'h3d9b8e89, 32'hbd38e983} /* (7, 17, 7) {real, imag} */,
  {32'h3db5cc6c, 32'hbd6c9fe5} /* (7, 17, 6) {real, imag} */,
  {32'h3e5837d6, 32'hbda348ae} /* (7, 17, 5) {real, imag} */,
  {32'hbe24bf63, 32'h3cebeb36} /* (7, 17, 4) {real, imag} */,
  {32'hbd741a9c, 32'h3d372b08} /* (7, 17, 3) {real, imag} */,
  {32'h3f919d4a, 32'h3e9f6a7e} /* (7, 17, 2) {real, imag} */,
  {32'hc049cf34, 32'hbe93a56d} /* (7, 17, 1) {real, imag} */,
  {32'hc00c5fad, 32'h00000000} /* (7, 17, 0) {real, imag} */,
  {32'hc0505974, 32'h3e90c12e} /* (7, 16, 31) {real, imag} */,
  {32'h3f98c566, 32'hbe158007} /* (7, 16, 30) {real, imag} */,
  {32'hbd93f79b, 32'hbe13a01b} /* (7, 16, 29) {real, imag} */,
  {32'hbe233d27, 32'h3d83031d} /* (7, 16, 28) {real, imag} */,
  {32'h3dec9800, 32'hbd355008} /* (7, 16, 27) {real, imag} */,
  {32'h3d364e96, 32'hbdac5477} /* (7, 16, 26) {real, imag} */,
  {32'h3dd18db2, 32'hbda4fd44} /* (7, 16, 25) {real, imag} */,
  {32'h3d95bb40, 32'hbd9546eb} /* (7, 16, 24) {real, imag} */,
  {32'h3d773028, 32'h3d066969} /* (7, 16, 23) {real, imag} */,
  {32'hbcc9f1c3, 32'h3d8bbe1c} /* (7, 16, 22) {real, imag} */,
  {32'h3dc67c44, 32'hbd2adb1e} /* (7, 16, 21) {real, imag} */,
  {32'h3d09e67f, 32'hbdb615be} /* (7, 16, 20) {real, imag} */,
  {32'hbdb4953a, 32'hbd07478d} /* (7, 16, 19) {real, imag} */,
  {32'h3c0c26a8, 32'h3cb328ee} /* (7, 16, 18) {real, imag} */,
  {32'hbc3a7fb7, 32'h3c9c1dc5} /* (7, 16, 17) {real, imag} */,
  {32'hbda7055e, 32'h00000000} /* (7, 16, 16) {real, imag} */,
  {32'hbc3a7fb7, 32'hbc9c1dc5} /* (7, 16, 15) {real, imag} */,
  {32'h3c0c26a8, 32'hbcb328ee} /* (7, 16, 14) {real, imag} */,
  {32'hbdb4953a, 32'h3d07478d} /* (7, 16, 13) {real, imag} */,
  {32'h3d09e67f, 32'h3db615be} /* (7, 16, 12) {real, imag} */,
  {32'h3dc67c44, 32'h3d2adb1e} /* (7, 16, 11) {real, imag} */,
  {32'hbcc9f1c3, 32'hbd8bbe1c} /* (7, 16, 10) {real, imag} */,
  {32'h3d773028, 32'hbd066969} /* (7, 16, 9) {real, imag} */,
  {32'h3d95bb40, 32'h3d9546eb} /* (7, 16, 8) {real, imag} */,
  {32'h3dd18db2, 32'h3da4fd44} /* (7, 16, 7) {real, imag} */,
  {32'h3d364e96, 32'h3dac5477} /* (7, 16, 6) {real, imag} */,
  {32'h3dec9800, 32'h3d355008} /* (7, 16, 5) {real, imag} */,
  {32'hbe233d27, 32'hbd83031d} /* (7, 16, 4) {real, imag} */,
  {32'hbd93f79b, 32'h3e13a01b} /* (7, 16, 3) {real, imag} */,
  {32'h3f98c566, 32'h3e158007} /* (7, 16, 2) {real, imag} */,
  {32'hc0505974, 32'hbe90c12e} /* (7, 16, 1) {real, imag} */,
  {32'hc0197b68, 32'h00000000} /* (7, 16, 0) {real, imag} */,
  {32'hc053f368, 32'h3ea9c467} /* (7, 15, 31) {real, imag} */,
  {32'h3f9e8c36, 32'hbdde9443} /* (7, 15, 30) {real, imag} */,
  {32'hbc176d30, 32'hbdd463cc} /* (7, 15, 29) {real, imag} */,
  {32'hbe1bd419, 32'hbe04a3af} /* (7, 15, 28) {real, imag} */,
  {32'h3df68160, 32'hbe35d0d1} /* (7, 15, 27) {real, imag} */,
  {32'h3d190144, 32'hbdd8b540} /* (7, 15, 26) {real, imag} */,
  {32'hbda49f63, 32'hbd65f4dd} /* (7, 15, 25) {real, imag} */,
  {32'h3df9e6cc, 32'hbd293335} /* (7, 15, 24) {real, imag} */,
  {32'hbd315bc6, 32'hbdfb2225} /* (7, 15, 23) {real, imag} */,
  {32'hbc5e5a56, 32'h3d26ec78} /* (7, 15, 22) {real, imag} */,
  {32'h3cfcae10, 32'hbb976c28} /* (7, 15, 21) {real, imag} */,
  {32'h3d8b6378, 32'hbdbdc789} /* (7, 15, 20) {real, imag} */,
  {32'h3d09bd06, 32'h3d373384} /* (7, 15, 19) {real, imag} */,
  {32'h3d119c24, 32'h3d4097fc} /* (7, 15, 18) {real, imag} */,
  {32'h3d238870, 32'hbd5bbe63} /* (7, 15, 17) {real, imag} */,
  {32'h3c3e0b90, 32'h00000000} /* (7, 15, 16) {real, imag} */,
  {32'h3d238870, 32'h3d5bbe63} /* (7, 15, 15) {real, imag} */,
  {32'h3d119c24, 32'hbd4097fc} /* (7, 15, 14) {real, imag} */,
  {32'h3d09bd06, 32'hbd373384} /* (7, 15, 13) {real, imag} */,
  {32'h3d8b6378, 32'h3dbdc789} /* (7, 15, 12) {real, imag} */,
  {32'h3cfcae10, 32'h3b976c28} /* (7, 15, 11) {real, imag} */,
  {32'hbc5e5a56, 32'hbd26ec78} /* (7, 15, 10) {real, imag} */,
  {32'hbd315bc6, 32'h3dfb2225} /* (7, 15, 9) {real, imag} */,
  {32'h3df9e6cc, 32'h3d293335} /* (7, 15, 8) {real, imag} */,
  {32'hbda49f63, 32'h3d65f4dd} /* (7, 15, 7) {real, imag} */,
  {32'h3d190144, 32'h3dd8b540} /* (7, 15, 6) {real, imag} */,
  {32'h3df68160, 32'h3e35d0d1} /* (7, 15, 5) {real, imag} */,
  {32'hbe1bd419, 32'h3e04a3af} /* (7, 15, 4) {real, imag} */,
  {32'hbc176d30, 32'h3dd463cc} /* (7, 15, 3) {real, imag} */,
  {32'h3f9e8c36, 32'h3dde9443} /* (7, 15, 2) {real, imag} */,
  {32'hc053f368, 32'hbea9c467} /* (7, 15, 1) {real, imag} */,
  {32'hc0265e19, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'hc03b27fc, 32'h3dfd296c} /* (7, 14, 31) {real, imag} */,
  {32'h3f9d6130, 32'hbe763dd0} /* (7, 14, 30) {real, imag} */,
  {32'h3d6ebc26, 32'h3c84287a} /* (7, 14, 29) {real, imag} */,
  {32'hbe4c12ba, 32'hbde061d0} /* (7, 14, 28) {real, imag} */,
  {32'h3e02ba9b, 32'hbdd03ede} /* (7, 14, 27) {real, imag} */,
  {32'h3d86d5d2, 32'hbd5dee3e} /* (7, 14, 26) {real, imag} */,
  {32'hbd35ee4c, 32'h3cd58690} /* (7, 14, 25) {real, imag} */,
  {32'h3c03c7c6, 32'hbcc3cee2} /* (7, 14, 24) {real, imag} */,
  {32'hbdae5360, 32'hbc647700} /* (7, 14, 23) {real, imag} */,
  {32'h3d888a1b, 32'hbd32c840} /* (7, 14, 22) {real, imag} */,
  {32'h3d962e15, 32'hbc9e2db8} /* (7, 14, 21) {real, imag} */,
  {32'h3d608ac2, 32'hbdabfbe2} /* (7, 14, 20) {real, imag} */,
  {32'h3d1df9a6, 32'h3bf87be0} /* (7, 14, 19) {real, imag} */,
  {32'hbd660df0, 32'hbd40a1f4} /* (7, 14, 18) {real, imag} */,
  {32'h3d6c4569, 32'h3d1c87fe} /* (7, 14, 17) {real, imag} */,
  {32'h3dde0812, 32'h00000000} /* (7, 14, 16) {real, imag} */,
  {32'h3d6c4569, 32'hbd1c87fe} /* (7, 14, 15) {real, imag} */,
  {32'hbd660df0, 32'h3d40a1f4} /* (7, 14, 14) {real, imag} */,
  {32'h3d1df9a6, 32'hbbf87be0} /* (7, 14, 13) {real, imag} */,
  {32'h3d608ac2, 32'h3dabfbe2} /* (7, 14, 12) {real, imag} */,
  {32'h3d962e15, 32'h3c9e2db8} /* (7, 14, 11) {real, imag} */,
  {32'h3d888a1b, 32'h3d32c840} /* (7, 14, 10) {real, imag} */,
  {32'hbdae5360, 32'h3c647700} /* (7, 14, 9) {real, imag} */,
  {32'h3c03c7c6, 32'h3cc3cee2} /* (7, 14, 8) {real, imag} */,
  {32'hbd35ee4c, 32'hbcd58690} /* (7, 14, 7) {real, imag} */,
  {32'h3d86d5d2, 32'h3d5dee3e} /* (7, 14, 6) {real, imag} */,
  {32'h3e02ba9b, 32'h3dd03ede} /* (7, 14, 5) {real, imag} */,
  {32'hbe4c12ba, 32'h3de061d0} /* (7, 14, 4) {real, imag} */,
  {32'h3d6ebc26, 32'hbc84287a} /* (7, 14, 3) {real, imag} */,
  {32'h3f9d6130, 32'h3e763dd0} /* (7, 14, 2) {real, imag} */,
  {32'hc03b27fc, 32'hbdfd296c} /* (7, 14, 1) {real, imag} */,
  {32'hc01f5728, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hc01e1ab5, 32'h3c09a200} /* (7, 13, 31) {real, imag} */,
  {32'h3f8c36a5, 32'hbe10f7f6} /* (7, 13, 30) {real, imag} */,
  {32'h3d227c7e, 32'hbd4c774a} /* (7, 13, 29) {real, imag} */,
  {32'hbe06e433, 32'h3b1615e0} /* (7, 13, 28) {real, imag} */,
  {32'h3e61dd67, 32'hbd748a98} /* (7, 13, 27) {real, imag} */,
  {32'h3d93c8bc, 32'h3c8975be} /* (7, 13, 26) {real, imag} */,
  {32'hbe130b55, 32'h3dabe742} /* (7, 13, 25) {real, imag} */,
  {32'h3d03474e, 32'hbe20956a} /* (7, 13, 24) {real, imag} */,
  {32'h3de55b92, 32'hbc8e4b4e} /* (7, 13, 23) {real, imag} */,
  {32'hbbdb7a48, 32'h3d4774cf} /* (7, 13, 22) {real, imag} */,
  {32'hbd7c53ca, 32'h3c8dda16} /* (7, 13, 21) {real, imag} */,
  {32'h3cb6eceb, 32'hbd70d65a} /* (7, 13, 20) {real, imag} */,
  {32'hbc920586, 32'hbc2c9b18} /* (7, 13, 19) {real, imag} */,
  {32'h3c83a464, 32'h3c44d2f0} /* (7, 13, 18) {real, imag} */,
  {32'h3c0be1fe, 32'hbd98aa40} /* (7, 13, 17) {real, imag} */,
  {32'h3da3c4ab, 32'h00000000} /* (7, 13, 16) {real, imag} */,
  {32'h3c0be1fe, 32'h3d98aa40} /* (7, 13, 15) {real, imag} */,
  {32'h3c83a464, 32'hbc44d2f0} /* (7, 13, 14) {real, imag} */,
  {32'hbc920586, 32'h3c2c9b18} /* (7, 13, 13) {real, imag} */,
  {32'h3cb6eceb, 32'h3d70d65a} /* (7, 13, 12) {real, imag} */,
  {32'hbd7c53ca, 32'hbc8dda16} /* (7, 13, 11) {real, imag} */,
  {32'hbbdb7a48, 32'hbd4774cf} /* (7, 13, 10) {real, imag} */,
  {32'h3de55b92, 32'h3c8e4b4e} /* (7, 13, 9) {real, imag} */,
  {32'h3d03474e, 32'h3e20956a} /* (7, 13, 8) {real, imag} */,
  {32'hbe130b55, 32'hbdabe742} /* (7, 13, 7) {real, imag} */,
  {32'h3d93c8bc, 32'hbc8975be} /* (7, 13, 6) {real, imag} */,
  {32'h3e61dd67, 32'h3d748a98} /* (7, 13, 5) {real, imag} */,
  {32'hbe06e433, 32'hbb1615e0} /* (7, 13, 4) {real, imag} */,
  {32'h3d227c7e, 32'h3d4c774a} /* (7, 13, 3) {real, imag} */,
  {32'h3f8c36a5, 32'h3e10f7f6} /* (7, 13, 2) {real, imag} */,
  {32'hc01e1ab5, 32'hbc09a200} /* (7, 13, 1) {real, imag} */,
  {32'hc0073d23, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'hbfe195a4, 32'h3c6daf40} /* (7, 12, 31) {real, imag} */,
  {32'h3f6f9e1c, 32'hbd4fc0f8} /* (7, 12, 30) {real, imag} */,
  {32'h3e951847, 32'h3d9c81e4} /* (7, 12, 29) {real, imag} */,
  {32'hbe0e20a3, 32'hbd48967a} /* (7, 12, 28) {real, imag} */,
  {32'h3d0db572, 32'hbc4a7640} /* (7, 12, 27) {real, imag} */,
  {32'h3d446cd1, 32'hbd39ff35} /* (7, 12, 26) {real, imag} */,
  {32'hbdc2a158, 32'hbe224fcf} /* (7, 12, 25) {real, imag} */,
  {32'hbc74d86c, 32'hbe0b8d42} /* (7, 12, 24) {real, imag} */,
  {32'h3a1892a0, 32'h3d731caa} /* (7, 12, 23) {real, imag} */,
  {32'hbd07b78f, 32'h3da591ce} /* (7, 12, 22) {real, imag} */,
  {32'h3d2d8ae0, 32'hbd44d710} /* (7, 12, 21) {real, imag} */,
  {32'h3bf44a52, 32'hbd9063a6} /* (7, 12, 20) {real, imag} */,
  {32'h3d8ba7b4, 32'h3d06774a} /* (7, 12, 19) {real, imag} */,
  {32'hbd2d2ff3, 32'hbacbe4f0} /* (7, 12, 18) {real, imag} */,
  {32'hbc79fee5, 32'h3cc86843} /* (7, 12, 17) {real, imag} */,
  {32'hbc98301e, 32'h00000000} /* (7, 12, 16) {real, imag} */,
  {32'hbc79fee5, 32'hbcc86843} /* (7, 12, 15) {real, imag} */,
  {32'hbd2d2ff3, 32'h3acbe4f0} /* (7, 12, 14) {real, imag} */,
  {32'h3d8ba7b4, 32'hbd06774a} /* (7, 12, 13) {real, imag} */,
  {32'h3bf44a52, 32'h3d9063a6} /* (7, 12, 12) {real, imag} */,
  {32'h3d2d8ae0, 32'h3d44d710} /* (7, 12, 11) {real, imag} */,
  {32'hbd07b78f, 32'hbda591ce} /* (7, 12, 10) {real, imag} */,
  {32'h3a1892a0, 32'hbd731caa} /* (7, 12, 9) {real, imag} */,
  {32'hbc74d86c, 32'h3e0b8d42} /* (7, 12, 8) {real, imag} */,
  {32'hbdc2a158, 32'h3e224fcf} /* (7, 12, 7) {real, imag} */,
  {32'h3d446cd1, 32'h3d39ff35} /* (7, 12, 6) {real, imag} */,
  {32'h3d0db572, 32'h3c4a7640} /* (7, 12, 5) {real, imag} */,
  {32'hbe0e20a3, 32'h3d48967a} /* (7, 12, 4) {real, imag} */,
  {32'h3e951847, 32'hbd9c81e4} /* (7, 12, 3) {real, imag} */,
  {32'h3f6f9e1c, 32'h3d4fc0f8} /* (7, 12, 2) {real, imag} */,
  {32'hbfe195a4, 32'hbc6daf40} /* (7, 12, 1) {real, imag} */,
  {32'hbfbe5c64, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'hbf64e748, 32'hbe80fdb5} /* (7, 11, 31) {real, imag} */,
  {32'h3f00e71c, 32'hbd901873} /* (7, 11, 30) {real, imag} */,
  {32'h3e30d081, 32'h3da989a3} /* (7, 11, 29) {real, imag} */,
  {32'hbe2789b0, 32'hbde08dce} /* (7, 11, 28) {real, imag} */,
  {32'h3c813b60, 32'hbd0f3d49} /* (7, 11, 27) {real, imag} */,
  {32'hbd8e3941, 32'h3ca694ef} /* (7, 11, 26) {real, imag} */,
  {32'hbd5f1294, 32'hbd47f0f0} /* (7, 11, 25) {real, imag} */,
  {32'h3e03a5c3, 32'hbe2326f7} /* (7, 11, 24) {real, imag} */,
  {32'hbc938fbf, 32'h3ca78a4c} /* (7, 11, 23) {real, imag} */,
  {32'hbcc068a3, 32'h3bf8a818} /* (7, 11, 22) {real, imag} */,
  {32'h3d561bf5, 32'hbd38f143} /* (7, 11, 21) {real, imag} */,
  {32'hbd1e10a8, 32'hbd0a8a5c} /* (7, 11, 20) {real, imag} */,
  {32'hbdd892be, 32'hbd8ddf68} /* (7, 11, 19) {real, imag} */,
  {32'h3c46ead0, 32'hbd54f02f} /* (7, 11, 18) {real, imag} */,
  {32'h3b60d150, 32'h3d427b80} /* (7, 11, 17) {real, imag} */,
  {32'h3d71f0e6, 32'h00000000} /* (7, 11, 16) {real, imag} */,
  {32'h3b60d150, 32'hbd427b80} /* (7, 11, 15) {real, imag} */,
  {32'h3c46ead0, 32'h3d54f02f} /* (7, 11, 14) {real, imag} */,
  {32'hbdd892be, 32'h3d8ddf68} /* (7, 11, 13) {real, imag} */,
  {32'hbd1e10a8, 32'h3d0a8a5c} /* (7, 11, 12) {real, imag} */,
  {32'h3d561bf5, 32'h3d38f143} /* (7, 11, 11) {real, imag} */,
  {32'hbcc068a3, 32'hbbf8a818} /* (7, 11, 10) {real, imag} */,
  {32'hbc938fbf, 32'hbca78a4c} /* (7, 11, 9) {real, imag} */,
  {32'h3e03a5c3, 32'h3e2326f7} /* (7, 11, 8) {real, imag} */,
  {32'hbd5f1294, 32'h3d47f0f0} /* (7, 11, 7) {real, imag} */,
  {32'hbd8e3941, 32'hbca694ef} /* (7, 11, 6) {real, imag} */,
  {32'h3c813b60, 32'h3d0f3d49} /* (7, 11, 5) {real, imag} */,
  {32'hbe2789b0, 32'h3de08dce} /* (7, 11, 4) {real, imag} */,
  {32'h3e30d081, 32'hbda989a3} /* (7, 11, 3) {real, imag} */,
  {32'h3f00e71c, 32'h3d901873} /* (7, 11, 2) {real, imag} */,
  {32'hbf64e748, 32'h3e80fdb5} /* (7, 11, 1) {real, imag} */,
  {32'hbef6881e, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'h3f1e5e48, 32'hbf10f856} /* (7, 10, 31) {real, imag} */,
  {32'hbe78054a, 32'h3e42b4d4} /* (7, 10, 30) {real, imag} */,
  {32'h3e0e95a4, 32'hbca2d124} /* (7, 10, 29) {real, imag} */,
  {32'h3b97e1d0, 32'hbe0224a4} /* (7, 10, 28) {real, imag} */,
  {32'h3d858e82, 32'h3d94be94} /* (7, 10, 27) {real, imag} */,
  {32'hbdb29482, 32'h3c83c408} /* (7, 10, 26) {real, imag} */,
  {32'h3e0ffbcc, 32'h3ca16df9} /* (7, 10, 25) {real, imag} */,
  {32'hbd4bffeb, 32'h3c8a43da} /* (7, 10, 24) {real, imag} */,
  {32'h3cbcb0b0, 32'hbddf3d0a} /* (7, 10, 23) {real, imag} */,
  {32'hbd20efee, 32'h3bce0da4} /* (7, 10, 22) {real, imag} */,
  {32'h3ab67a88, 32'h3d5df7f4} /* (7, 10, 21) {real, imag} */,
  {32'hbd16beb5, 32'hbdbd9a1b} /* (7, 10, 20) {real, imag} */,
  {32'h3dab8612, 32'h3c458d6a} /* (7, 10, 19) {real, imag} */,
  {32'hbb979a20, 32'h3d256a30} /* (7, 10, 18) {real, imag} */,
  {32'h3d008d66, 32'hbbb50f48} /* (7, 10, 17) {real, imag} */,
  {32'hbc98bb92, 32'h00000000} /* (7, 10, 16) {real, imag} */,
  {32'h3d008d66, 32'h3bb50f48} /* (7, 10, 15) {real, imag} */,
  {32'hbb979a20, 32'hbd256a30} /* (7, 10, 14) {real, imag} */,
  {32'h3dab8612, 32'hbc458d6a} /* (7, 10, 13) {real, imag} */,
  {32'hbd16beb5, 32'h3dbd9a1b} /* (7, 10, 12) {real, imag} */,
  {32'h3ab67a88, 32'hbd5df7f4} /* (7, 10, 11) {real, imag} */,
  {32'hbd20efee, 32'hbbce0da4} /* (7, 10, 10) {real, imag} */,
  {32'h3cbcb0b0, 32'h3ddf3d0a} /* (7, 10, 9) {real, imag} */,
  {32'hbd4bffeb, 32'hbc8a43da} /* (7, 10, 8) {real, imag} */,
  {32'h3e0ffbcc, 32'hbca16df9} /* (7, 10, 7) {real, imag} */,
  {32'hbdb29482, 32'hbc83c408} /* (7, 10, 6) {real, imag} */,
  {32'h3d858e82, 32'hbd94be94} /* (7, 10, 5) {real, imag} */,
  {32'h3b97e1d0, 32'h3e0224a4} /* (7, 10, 4) {real, imag} */,
  {32'h3e0e95a4, 32'h3ca2d124} /* (7, 10, 3) {real, imag} */,
  {32'hbe78054a, 32'hbe42b4d4} /* (7, 10, 2) {real, imag} */,
  {32'h3f1e5e48, 32'h3f10f856} /* (7, 10, 1) {real, imag} */,
  {32'h3f2e2e40, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'h3fd51beb, 32'hbf69e8dd} /* (7, 9, 31) {real, imag} */,
  {32'hbf27d1aa, 32'h3ec91f53} /* (7, 9, 30) {real, imag} */,
  {32'h3e8fc30e, 32'h3da17e23} /* (7, 9, 29) {real, imag} */,
  {32'h3e1cb173, 32'hbe4c04be} /* (7, 9, 28) {real, imag} */,
  {32'h3a7ea100, 32'h3e36f827} /* (7, 9, 27) {real, imag} */,
  {32'hbd9d4a23, 32'hbbcbaff2} /* (7, 9, 26) {real, imag} */,
  {32'hbd6bde71, 32'h3c8af294} /* (7, 9, 25) {real, imag} */,
  {32'hbd4432c6, 32'hbbf91134} /* (7, 9, 24) {real, imag} */,
  {32'h3dea5aa5, 32'h3c055b18} /* (7, 9, 23) {real, imag} */,
  {32'hbdd4a7de, 32'hbcf41596} /* (7, 9, 22) {real, imag} */,
  {32'hbda705d5, 32'h3cdf1dcf} /* (7, 9, 21) {real, imag} */,
  {32'h3b8bc9d4, 32'h3d93b578} /* (7, 9, 20) {real, imag} */,
  {32'h3c6e64da, 32'hbc19b566} /* (7, 9, 19) {real, imag} */,
  {32'hbc8e301e, 32'h3d99fc66} /* (7, 9, 18) {real, imag} */,
  {32'hbd5bbe38, 32'hbc9d48b3} /* (7, 9, 17) {real, imag} */,
  {32'hbc27b3b8, 32'h00000000} /* (7, 9, 16) {real, imag} */,
  {32'hbd5bbe38, 32'h3c9d48b3} /* (7, 9, 15) {real, imag} */,
  {32'hbc8e301e, 32'hbd99fc66} /* (7, 9, 14) {real, imag} */,
  {32'h3c6e64da, 32'h3c19b566} /* (7, 9, 13) {real, imag} */,
  {32'h3b8bc9d4, 32'hbd93b578} /* (7, 9, 12) {real, imag} */,
  {32'hbda705d5, 32'hbcdf1dcf} /* (7, 9, 11) {real, imag} */,
  {32'hbdd4a7de, 32'h3cf41596} /* (7, 9, 10) {real, imag} */,
  {32'h3dea5aa5, 32'hbc055b18} /* (7, 9, 9) {real, imag} */,
  {32'hbd4432c6, 32'h3bf91134} /* (7, 9, 8) {real, imag} */,
  {32'hbd6bde71, 32'hbc8af294} /* (7, 9, 7) {real, imag} */,
  {32'hbd9d4a23, 32'h3bcbaff2} /* (7, 9, 6) {real, imag} */,
  {32'h3a7ea100, 32'hbe36f827} /* (7, 9, 5) {real, imag} */,
  {32'h3e1cb173, 32'h3e4c04be} /* (7, 9, 4) {real, imag} */,
  {32'h3e8fc30e, 32'hbda17e23} /* (7, 9, 3) {real, imag} */,
  {32'hbf27d1aa, 32'hbec91f53} /* (7, 9, 2) {real, imag} */,
  {32'h3fd51beb, 32'h3f69e8dd} /* (7, 9, 1) {real, imag} */,
  {32'h3ffd1d40, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'h400f6040, 32'hbf85f3d4} /* (7, 8, 31) {real, imag} */,
  {32'hbf43b66b, 32'h3ee2279e} /* (7, 8, 30) {real, imag} */,
  {32'h3e4067a8, 32'h3e0ff5c6} /* (7, 8, 29) {real, imag} */,
  {32'h3e30a681, 32'hbe21128a} /* (7, 8, 28) {real, imag} */,
  {32'hbe3613fa, 32'h3e114998} /* (7, 8, 27) {real, imag} */,
  {32'hbcaa397e, 32'h3d9df706} /* (7, 8, 26) {real, imag} */,
  {32'h3c6702fa, 32'hbd29cdbc} /* (7, 8, 25) {real, imag} */,
  {32'hbccbb234, 32'hbd4b179a} /* (7, 8, 24) {real, imag} */,
  {32'hbce1171e, 32'h3e187a20} /* (7, 8, 23) {real, imag} */,
  {32'h3d9d354a, 32'h3c83eaa0} /* (7, 8, 22) {real, imag} */,
  {32'hbe08d8ca, 32'hbd55b398} /* (7, 8, 21) {real, imag} */,
  {32'hbd87273b, 32'h3cdd8efc} /* (7, 8, 20) {real, imag} */,
  {32'h3ceeef6a, 32'hbcfd35e4} /* (7, 8, 19) {real, imag} */,
  {32'h3d487d3e, 32'h3cf1ed50} /* (7, 8, 18) {real, imag} */,
  {32'h3cbc38a6, 32'h3d38895c} /* (7, 8, 17) {real, imag} */,
  {32'h3d3e575c, 32'h00000000} /* (7, 8, 16) {real, imag} */,
  {32'h3cbc38a6, 32'hbd38895c} /* (7, 8, 15) {real, imag} */,
  {32'h3d487d3e, 32'hbcf1ed50} /* (7, 8, 14) {real, imag} */,
  {32'h3ceeef6a, 32'h3cfd35e4} /* (7, 8, 13) {real, imag} */,
  {32'hbd87273b, 32'hbcdd8efc} /* (7, 8, 12) {real, imag} */,
  {32'hbe08d8ca, 32'h3d55b398} /* (7, 8, 11) {real, imag} */,
  {32'h3d9d354a, 32'hbc83eaa0} /* (7, 8, 10) {real, imag} */,
  {32'hbce1171e, 32'hbe187a20} /* (7, 8, 9) {real, imag} */,
  {32'hbccbb234, 32'h3d4b179a} /* (7, 8, 8) {real, imag} */,
  {32'h3c6702fa, 32'h3d29cdbc} /* (7, 8, 7) {real, imag} */,
  {32'hbcaa397e, 32'hbd9df706} /* (7, 8, 6) {real, imag} */,
  {32'hbe3613fa, 32'hbe114998} /* (7, 8, 5) {real, imag} */,
  {32'h3e30a681, 32'h3e21128a} /* (7, 8, 4) {real, imag} */,
  {32'h3e4067a8, 32'hbe0ff5c6} /* (7, 8, 3) {real, imag} */,
  {32'hbf43b66b, 32'hbee2279e} /* (7, 8, 2) {real, imag} */,
  {32'h400f6040, 32'h3f85f3d4} /* (7, 8, 1) {real, imag} */,
  {32'h40251cf6, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'h402ace2f, 32'hbfa448a8} /* (7, 7, 31) {real, imag} */,
  {32'hbf5eb0d8, 32'h3f15bcda} /* (7, 7, 30) {real, imag} */,
  {32'h3e522ad9, 32'hbce46f64} /* (7, 7, 29) {real, imag} */,
  {32'h3e27e850, 32'hbe19646c} /* (7, 7, 28) {real, imag} */,
  {32'hbe87944f, 32'h3cd55cae} /* (7, 7, 27) {real, imag} */,
  {32'hbdd3748d, 32'hbc826621} /* (7, 7, 26) {real, imag} */,
  {32'h3ca1568e, 32'hbe1910fa} /* (7, 7, 25) {real, imag} */,
  {32'hbc93eb8d, 32'hbcda1842} /* (7, 7, 24) {real, imag} */,
  {32'hbd1c5d0b, 32'hbd5323dc} /* (7, 7, 23) {real, imag} */,
  {32'hbc93d93b, 32'h3d88d5d0} /* (7, 7, 22) {real, imag} */,
  {32'hbd3a1746, 32'h3de67e9f} /* (7, 7, 21) {real, imag} */,
  {32'h3ca6e131, 32'h3d515d20} /* (7, 7, 20) {real, imag} */,
  {32'h3d9f38b9, 32'h3d255b6a} /* (7, 7, 19) {real, imag} */,
  {32'hbe09b509, 32'h3cf7b273} /* (7, 7, 18) {real, imag} */,
  {32'hbba149e0, 32'hbb806778} /* (7, 7, 17) {real, imag} */,
  {32'h3d23b238, 32'h00000000} /* (7, 7, 16) {real, imag} */,
  {32'hbba149e0, 32'h3b806778} /* (7, 7, 15) {real, imag} */,
  {32'hbe09b509, 32'hbcf7b273} /* (7, 7, 14) {real, imag} */,
  {32'h3d9f38b9, 32'hbd255b6a} /* (7, 7, 13) {real, imag} */,
  {32'h3ca6e131, 32'hbd515d20} /* (7, 7, 12) {real, imag} */,
  {32'hbd3a1746, 32'hbde67e9f} /* (7, 7, 11) {real, imag} */,
  {32'hbc93d93b, 32'hbd88d5d0} /* (7, 7, 10) {real, imag} */,
  {32'hbd1c5d0b, 32'h3d5323dc} /* (7, 7, 9) {real, imag} */,
  {32'hbc93eb8d, 32'h3cda1842} /* (7, 7, 8) {real, imag} */,
  {32'h3ca1568e, 32'h3e1910fa} /* (7, 7, 7) {real, imag} */,
  {32'hbdd3748d, 32'h3c826621} /* (7, 7, 6) {real, imag} */,
  {32'hbe87944f, 32'hbcd55cae} /* (7, 7, 5) {real, imag} */,
  {32'h3e27e850, 32'h3e19646c} /* (7, 7, 4) {real, imag} */,
  {32'h3e522ad9, 32'h3ce46f64} /* (7, 7, 3) {real, imag} */,
  {32'hbf5eb0d8, 32'hbf15bcda} /* (7, 7, 2) {real, imag} */,
  {32'h402ace2f, 32'h3fa448a8} /* (7, 7, 1) {real, imag} */,
  {32'h4044dd04, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'h403b5b46, 32'hbfd8e070} /* (7, 6, 31) {real, imag} */,
  {32'hbf27463a, 32'h3f2accd4} /* (7, 6, 30) {real, imag} */,
  {32'h3d6e7b9a, 32'h3d2a3c49} /* (7, 6, 29) {real, imag} */,
  {32'h3e0b6dd0, 32'hbc755c7c} /* (7, 6, 28) {real, imag} */,
  {32'hbe23a93d, 32'h3e000f8f} /* (7, 6, 27) {real, imag} */,
  {32'hbd810422, 32'h3d0d501c} /* (7, 6, 26) {real, imag} */,
  {32'h3db4e455, 32'hbe09f206} /* (7, 6, 25) {real, imag} */,
  {32'hbdd70235, 32'h3e1de345} /* (7, 6, 24) {real, imag} */,
  {32'hbd26c020, 32'h3e2a6504} /* (7, 6, 23) {real, imag} */,
  {32'hbe0729be, 32'hbd8ae391} /* (7, 6, 22) {real, imag} */,
  {32'hbd734d79, 32'h3da70938} /* (7, 6, 21) {real, imag} */,
  {32'h3dc8eb9e, 32'hbbaf78a4} /* (7, 6, 20) {real, imag} */,
  {32'h3d1bd222, 32'h3d0b7bf0} /* (7, 6, 19) {real, imag} */,
  {32'hbda913e2, 32'h3da9fa87} /* (7, 6, 18) {real, imag} */,
  {32'hbcffd13d, 32'hbd6b25d2} /* (7, 6, 17) {real, imag} */,
  {32'h3dd8db93, 32'h00000000} /* (7, 6, 16) {real, imag} */,
  {32'hbcffd13d, 32'h3d6b25d2} /* (7, 6, 15) {real, imag} */,
  {32'hbda913e2, 32'hbda9fa87} /* (7, 6, 14) {real, imag} */,
  {32'h3d1bd222, 32'hbd0b7bf0} /* (7, 6, 13) {real, imag} */,
  {32'h3dc8eb9e, 32'h3baf78a4} /* (7, 6, 12) {real, imag} */,
  {32'hbd734d79, 32'hbda70938} /* (7, 6, 11) {real, imag} */,
  {32'hbe0729be, 32'h3d8ae391} /* (7, 6, 10) {real, imag} */,
  {32'hbd26c020, 32'hbe2a6504} /* (7, 6, 9) {real, imag} */,
  {32'hbdd70235, 32'hbe1de345} /* (7, 6, 8) {real, imag} */,
  {32'h3db4e455, 32'h3e09f206} /* (7, 6, 7) {real, imag} */,
  {32'hbd810422, 32'hbd0d501c} /* (7, 6, 6) {real, imag} */,
  {32'hbe23a93d, 32'hbe000f8f} /* (7, 6, 5) {real, imag} */,
  {32'h3e0b6dd0, 32'h3c755c7c} /* (7, 6, 4) {real, imag} */,
  {32'h3d6e7b9a, 32'hbd2a3c49} /* (7, 6, 3) {real, imag} */,
  {32'hbf27463a, 32'hbf2accd4} /* (7, 6, 2) {real, imag} */,
  {32'h403b5b46, 32'h3fd8e070} /* (7, 6, 1) {real, imag} */,
  {32'h406cdce6, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'h4031bf90, 32'hc0101f84} /* (7, 5, 31) {real, imag} */,
  {32'hbe9f5ff6, 32'h3f67f14d} /* (7, 5, 30) {real, imag} */,
  {32'h3be35324, 32'h3ceafb1b} /* (7, 5, 29) {real, imag} */,
  {32'h3c3c38e8, 32'h3e6c70ea} /* (7, 5, 28) {real, imag} */,
  {32'hbe3ef250, 32'h3cc033c6} /* (7, 5, 27) {real, imag} */,
  {32'h3db75ee0, 32'h3dced9aa} /* (7, 5, 26) {real, imag} */,
  {32'h3e0204cc, 32'hbbb96390} /* (7, 5, 25) {real, imag} */,
  {32'h3c428424, 32'h3e005dce} /* (7, 5, 24) {real, imag} */,
  {32'hbd7b44f3, 32'h3d603d14} /* (7, 5, 23) {real, imag} */,
  {32'hbd5c88b6, 32'h3b336670} /* (7, 5, 22) {real, imag} */,
  {32'hbe37a06c, 32'hbd142ad3} /* (7, 5, 21) {real, imag} */,
  {32'hbbed1794, 32'hbc30bfe8} /* (7, 5, 20) {real, imag} */,
  {32'hbd56416d, 32'h3b404340} /* (7, 5, 19) {real, imag} */,
  {32'hbd570efe, 32'hbda1312e} /* (7, 5, 18) {real, imag} */,
  {32'hbc85fd9d, 32'hbd8723b0} /* (7, 5, 17) {real, imag} */,
  {32'hbd8a443d, 32'h00000000} /* (7, 5, 16) {real, imag} */,
  {32'hbc85fd9d, 32'h3d8723b0} /* (7, 5, 15) {real, imag} */,
  {32'hbd570efe, 32'h3da1312e} /* (7, 5, 14) {real, imag} */,
  {32'hbd56416d, 32'hbb404340} /* (7, 5, 13) {real, imag} */,
  {32'hbbed1794, 32'h3c30bfe8} /* (7, 5, 12) {real, imag} */,
  {32'hbe37a06c, 32'h3d142ad3} /* (7, 5, 11) {real, imag} */,
  {32'hbd5c88b6, 32'hbb336670} /* (7, 5, 10) {real, imag} */,
  {32'hbd7b44f3, 32'hbd603d14} /* (7, 5, 9) {real, imag} */,
  {32'h3c428424, 32'hbe005dce} /* (7, 5, 8) {real, imag} */,
  {32'h3e0204cc, 32'h3bb96390} /* (7, 5, 7) {real, imag} */,
  {32'h3db75ee0, 32'hbdced9aa} /* (7, 5, 6) {real, imag} */,
  {32'hbe3ef250, 32'hbcc033c6} /* (7, 5, 5) {real, imag} */,
  {32'h3c3c38e8, 32'hbe6c70ea} /* (7, 5, 4) {real, imag} */,
  {32'h3be35324, 32'hbceafb1b} /* (7, 5, 3) {real, imag} */,
  {32'hbe9f5ff6, 32'hbf67f14d} /* (7, 5, 2) {real, imag} */,
  {32'h4031bf90, 32'h40101f84} /* (7, 5, 1) {real, imag} */,
  {32'h407d8496, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'h401caacd, 32'hc02bc1e5} /* (7, 4, 31) {real, imag} */,
  {32'h3d7e3898, 32'h3f789206} /* (7, 4, 30) {real, imag} */,
  {32'h3d661948, 32'hbd1d02fa} /* (7, 4, 29) {real, imag} */,
  {32'h3cfbf98c, 32'h3e6557c6} /* (7, 4, 28) {real, imag} */,
  {32'hbddfb7d4, 32'hbccd9a85} /* (7, 4, 27) {real, imag} */,
  {32'hbcc0f0ae, 32'h3de56e25} /* (7, 4, 26) {real, imag} */,
  {32'h3d069f8e, 32'hbe0aa1af} /* (7, 4, 25) {real, imag} */,
  {32'hbd9095fe, 32'h3ccbe277} /* (7, 4, 24) {real, imag} */,
  {32'hbc839185, 32'hbda07816} /* (7, 4, 23) {real, imag} */,
  {32'h3cefd774, 32'h3dc55de5} /* (7, 4, 22) {real, imag} */,
  {32'hbcc6f3b2, 32'h3db0a12c} /* (7, 4, 21) {real, imag} */,
  {32'hbc9e5294, 32'h3d37d13b} /* (7, 4, 20) {real, imag} */,
  {32'hbcf4312a, 32'h3d917c0b} /* (7, 4, 19) {real, imag} */,
  {32'h3dce7d43, 32'h3db9d9e2} /* (7, 4, 18) {real, imag} */,
  {32'hbccd77c8, 32'h3b7bb850} /* (7, 4, 17) {real, imag} */,
  {32'hbd59296c, 32'h00000000} /* (7, 4, 16) {real, imag} */,
  {32'hbccd77c8, 32'hbb7bb850} /* (7, 4, 15) {real, imag} */,
  {32'h3dce7d43, 32'hbdb9d9e2} /* (7, 4, 14) {real, imag} */,
  {32'hbcf4312a, 32'hbd917c0b} /* (7, 4, 13) {real, imag} */,
  {32'hbc9e5294, 32'hbd37d13b} /* (7, 4, 12) {real, imag} */,
  {32'hbcc6f3b2, 32'hbdb0a12c} /* (7, 4, 11) {real, imag} */,
  {32'h3cefd774, 32'hbdc55de5} /* (7, 4, 10) {real, imag} */,
  {32'hbc839185, 32'h3da07816} /* (7, 4, 9) {real, imag} */,
  {32'hbd9095fe, 32'hbccbe277} /* (7, 4, 8) {real, imag} */,
  {32'h3d069f8e, 32'h3e0aa1af} /* (7, 4, 7) {real, imag} */,
  {32'hbcc0f0ae, 32'hbde56e25} /* (7, 4, 6) {real, imag} */,
  {32'hbddfb7d4, 32'h3ccd9a85} /* (7, 4, 5) {real, imag} */,
  {32'h3cfbf98c, 32'hbe6557c6} /* (7, 4, 4) {real, imag} */,
  {32'h3d661948, 32'h3d1d02fa} /* (7, 4, 3) {real, imag} */,
  {32'h3d7e3898, 32'hbf789206} /* (7, 4, 2) {real, imag} */,
  {32'h401caacd, 32'h402bc1e5} /* (7, 4, 1) {real, imag} */,
  {32'h4088a70c, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'h4018a76c, 32'hc0386a85} /* (7, 3, 31) {real, imag} */,
  {32'h3e96b5ea, 32'h3f682ee4} /* (7, 3, 30) {real, imag} */,
  {32'h3d33fb28, 32'h3e3ed196} /* (7, 3, 29) {real, imag} */,
  {32'hbd9b4001, 32'h3eb2ec00} /* (7, 3, 28) {real, imag} */,
  {32'hbe5fa46d, 32'hbdbb76fd} /* (7, 3, 27) {real, imag} */,
  {32'hbd4961bc, 32'hbd060d38} /* (7, 3, 26) {real, imag} */,
  {32'h397c1e00, 32'hbdc82882} /* (7, 3, 25) {real, imag} */,
  {32'hbd0f2fd2, 32'h3d258dfa} /* (7, 3, 24) {real, imag} */,
  {32'hbd8edd9a, 32'hbd02e7b0} /* (7, 3, 23) {real, imag} */,
  {32'hbde740a8, 32'hbd26f8a5} /* (7, 3, 22) {real, imag} */,
  {32'h3db38e71, 32'h3ced8afe} /* (7, 3, 21) {real, imag} */,
  {32'h3de630ea, 32'hbd15d968} /* (7, 3, 20) {real, imag} */,
  {32'hbbab5398, 32'h3ccc5fcc} /* (7, 3, 19) {real, imag} */,
  {32'h3cff37e0, 32'h3d979880} /* (7, 3, 18) {real, imag} */,
  {32'hbcad162a, 32'h3c829ea9} /* (7, 3, 17) {real, imag} */,
  {32'h3da8be9c, 32'h00000000} /* (7, 3, 16) {real, imag} */,
  {32'hbcad162a, 32'hbc829ea9} /* (7, 3, 15) {real, imag} */,
  {32'h3cff37e0, 32'hbd979880} /* (7, 3, 14) {real, imag} */,
  {32'hbbab5398, 32'hbccc5fcc} /* (7, 3, 13) {real, imag} */,
  {32'h3de630ea, 32'h3d15d968} /* (7, 3, 12) {real, imag} */,
  {32'h3db38e71, 32'hbced8afe} /* (7, 3, 11) {real, imag} */,
  {32'hbde740a8, 32'h3d26f8a5} /* (7, 3, 10) {real, imag} */,
  {32'hbd8edd9a, 32'h3d02e7b0} /* (7, 3, 9) {real, imag} */,
  {32'hbd0f2fd2, 32'hbd258dfa} /* (7, 3, 8) {real, imag} */,
  {32'h397c1e00, 32'h3dc82882} /* (7, 3, 7) {real, imag} */,
  {32'hbd4961bc, 32'h3d060d38} /* (7, 3, 6) {real, imag} */,
  {32'hbe5fa46d, 32'h3dbb76fd} /* (7, 3, 5) {real, imag} */,
  {32'hbd9b4001, 32'hbeb2ec00} /* (7, 3, 4) {real, imag} */,
  {32'h3d33fb28, 32'hbe3ed196} /* (7, 3, 3) {real, imag} */,
  {32'h3e96b5ea, 32'hbf682ee4} /* (7, 3, 2) {real, imag} */,
  {32'h4018a76c, 32'h40386a85} /* (7, 3, 1) {real, imag} */,
  {32'h408d17b5, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'h40133db4, 32'hc03d396b} /* (7, 2, 31) {real, imag} */,
  {32'h3ec6cedf, 32'h3f5c5274} /* (7, 2, 30) {real, imag} */,
  {32'h3c66ce38, 32'h3ded423a} /* (7, 2, 29) {real, imag} */,
  {32'hbe081f06, 32'h3e93de68} /* (7, 2, 28) {real, imag} */,
  {32'hbe1e5fe1, 32'hbcd29aa0} /* (7, 2, 27) {real, imag} */,
  {32'h3cb5c24e, 32'hbd6904ac} /* (7, 2, 26) {real, imag} */,
  {32'hbc9a70d0, 32'hbd58734f} /* (7, 2, 25) {real, imag} */,
  {32'h3ccf0098, 32'h3df011be} /* (7, 2, 24) {real, imag} */,
  {32'h3d81e300, 32'h3d8fb5e8} /* (7, 2, 23) {real, imag} */,
  {32'h3cb478d5, 32'h3d32f42d} /* (7, 2, 22) {real, imag} */,
  {32'hbbdac8f0, 32'h3d362d2c} /* (7, 2, 21) {real, imag} */,
  {32'h3bb5aaf4, 32'hbd25ac0e} /* (7, 2, 20) {real, imag} */,
  {32'hbca98e05, 32'hbb986130} /* (7, 2, 19) {real, imag} */,
  {32'hbc735eec, 32'hbb44b824} /* (7, 2, 18) {real, imag} */,
  {32'h3c93ec3e, 32'hbd3c1fc0} /* (7, 2, 17) {real, imag} */,
  {32'h3d4137c0, 32'h00000000} /* (7, 2, 16) {real, imag} */,
  {32'h3c93ec3e, 32'h3d3c1fc0} /* (7, 2, 15) {real, imag} */,
  {32'hbc735eec, 32'h3b44b824} /* (7, 2, 14) {real, imag} */,
  {32'hbca98e05, 32'h3b986130} /* (7, 2, 13) {real, imag} */,
  {32'h3bb5aaf4, 32'h3d25ac0e} /* (7, 2, 12) {real, imag} */,
  {32'hbbdac8f0, 32'hbd362d2c} /* (7, 2, 11) {real, imag} */,
  {32'h3cb478d5, 32'hbd32f42d} /* (7, 2, 10) {real, imag} */,
  {32'h3d81e300, 32'hbd8fb5e8} /* (7, 2, 9) {real, imag} */,
  {32'h3ccf0098, 32'hbdf011be} /* (7, 2, 8) {real, imag} */,
  {32'hbc9a70d0, 32'h3d58734f} /* (7, 2, 7) {real, imag} */,
  {32'h3cb5c24e, 32'h3d6904ac} /* (7, 2, 6) {real, imag} */,
  {32'hbe1e5fe1, 32'h3cd29aa0} /* (7, 2, 5) {real, imag} */,
  {32'hbe081f06, 32'hbe93de68} /* (7, 2, 4) {real, imag} */,
  {32'h3c66ce38, 32'hbded423a} /* (7, 2, 3) {real, imag} */,
  {32'h3ec6cedf, 32'hbf5c5274} /* (7, 2, 2) {real, imag} */,
  {32'h40133db4, 32'h403d396b} /* (7, 2, 1) {real, imag} */,
  {32'h409434b6, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'h40154b8e, 32'hc02ee45c} /* (7, 1, 31) {real, imag} */,
  {32'h3eb56681, 32'h3f43c58a} /* (7, 1, 30) {real, imag} */,
  {32'hbe2cd73e, 32'h3d8cab81} /* (7, 1, 29) {real, imag} */,
  {32'hbdcca31b, 32'h3e388af0} /* (7, 1, 28) {real, imag} */,
  {32'hbd8079a1, 32'h3c96f4fa} /* (7, 1, 27) {real, imag} */,
  {32'hbde7b6f2, 32'h3d4a9bb1} /* (7, 1, 26) {real, imag} */,
  {32'hbc937076, 32'hbd913bc8} /* (7, 1, 25) {real, imag} */,
  {32'h3d595d16, 32'h3d9da270} /* (7, 1, 24) {real, imag} */,
  {32'h3da7a8bb, 32'hbdc922b6} /* (7, 1, 23) {real, imag} */,
  {32'h3d798ebe, 32'h3cdfe301} /* (7, 1, 22) {real, imag} */,
  {32'h3d61867c, 32'h3e04374f} /* (7, 1, 21) {real, imag} */,
  {32'hbd920d88, 32'h3d14743c} /* (7, 1, 20) {real, imag} */,
  {32'hbd896140, 32'h3d71a35a} /* (7, 1, 19) {real, imag} */,
  {32'h3da5bc08, 32'h3caed796} /* (7, 1, 18) {real, imag} */,
  {32'hbccc8bb6, 32'hbc843b46} /* (7, 1, 17) {real, imag} */,
  {32'h3a883a40, 32'h00000000} /* (7, 1, 16) {real, imag} */,
  {32'hbccc8bb6, 32'h3c843b46} /* (7, 1, 15) {real, imag} */,
  {32'h3da5bc08, 32'hbcaed796} /* (7, 1, 14) {real, imag} */,
  {32'hbd896140, 32'hbd71a35a} /* (7, 1, 13) {real, imag} */,
  {32'hbd920d88, 32'hbd14743c} /* (7, 1, 12) {real, imag} */,
  {32'h3d61867c, 32'hbe04374f} /* (7, 1, 11) {real, imag} */,
  {32'h3d798ebe, 32'hbcdfe301} /* (7, 1, 10) {real, imag} */,
  {32'h3da7a8bb, 32'h3dc922b6} /* (7, 1, 9) {real, imag} */,
  {32'h3d595d16, 32'hbd9da270} /* (7, 1, 8) {real, imag} */,
  {32'hbc937076, 32'h3d913bc8} /* (7, 1, 7) {real, imag} */,
  {32'hbde7b6f2, 32'hbd4a9bb1} /* (7, 1, 6) {real, imag} */,
  {32'hbd8079a1, 32'hbc96f4fa} /* (7, 1, 5) {real, imag} */,
  {32'hbdcca31b, 32'hbe388af0} /* (7, 1, 4) {real, imag} */,
  {32'hbe2cd73e, 32'hbd8cab81} /* (7, 1, 3) {real, imag} */,
  {32'h3eb56681, 32'hbf43c58a} /* (7, 1, 2) {real, imag} */,
  {32'h40154b8e, 32'h402ee45c} /* (7, 1, 1) {real, imag} */,
  {32'h4091cf8c, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'h4021c640, 32'hc00853a3} /* (7, 0, 31) {real, imag} */,
  {32'h3c52cc00, 32'h3f1aec3c} /* (7, 0, 30) {real, imag} */,
  {32'hbe11e958, 32'hbd903db2} /* (7, 0, 29) {real, imag} */,
  {32'h3c411650, 32'h3e1d1a94} /* (7, 0, 28) {real, imag} */,
  {32'hbb7d2590, 32'hbbe0b57c} /* (7, 0, 27) {real, imag} */,
  {32'h3c89cc67, 32'hbcd15864} /* (7, 0, 26) {real, imag} */,
  {32'hbd326228, 32'hbd45f4a4} /* (7, 0, 25) {real, imag} */,
  {32'hbd9e2388, 32'hbd41cefc} /* (7, 0, 24) {real, imag} */,
  {32'hbcd44d30, 32'hbd77891d} /* (7, 0, 23) {real, imag} */,
  {32'h3d5d487e, 32'hbc5965b0} /* (7, 0, 22) {real, imag} */,
  {32'h3ccbb25e, 32'hbcc87834} /* (7, 0, 21) {real, imag} */,
  {32'h3ce7edce, 32'hbb739290} /* (7, 0, 20) {real, imag} */,
  {32'h3cc511ca, 32'h3dd96f08} /* (7, 0, 19) {real, imag} */,
  {32'hbdbde81b, 32'hbc245c25} /* (7, 0, 18) {real, imag} */,
  {32'hbaf9cb68, 32'hbc0c02b4} /* (7, 0, 17) {real, imag} */,
  {32'hbbe95fa8, 32'h00000000} /* (7, 0, 16) {real, imag} */,
  {32'hbaf9cb68, 32'h3c0c02b4} /* (7, 0, 15) {real, imag} */,
  {32'hbdbde81b, 32'h3c245c25} /* (7, 0, 14) {real, imag} */,
  {32'h3cc511ca, 32'hbdd96f08} /* (7, 0, 13) {real, imag} */,
  {32'h3ce7edce, 32'h3b739290} /* (7, 0, 12) {real, imag} */,
  {32'h3ccbb25e, 32'h3cc87834} /* (7, 0, 11) {real, imag} */,
  {32'h3d5d487e, 32'h3c5965b0} /* (7, 0, 10) {real, imag} */,
  {32'hbcd44d30, 32'h3d77891d} /* (7, 0, 9) {real, imag} */,
  {32'hbd9e2388, 32'h3d41cefc} /* (7, 0, 8) {real, imag} */,
  {32'hbd326228, 32'h3d45f4a4} /* (7, 0, 7) {real, imag} */,
  {32'h3c89cc67, 32'h3cd15864} /* (7, 0, 6) {real, imag} */,
  {32'hbb7d2590, 32'h3be0b57c} /* (7, 0, 5) {real, imag} */,
  {32'h3c411650, 32'hbe1d1a94} /* (7, 0, 4) {real, imag} */,
  {32'hbe11e958, 32'h3d903db2} /* (7, 0, 3) {real, imag} */,
  {32'h3c52cc00, 32'hbf1aec3c} /* (7, 0, 2) {real, imag} */,
  {32'h4021c640, 32'h400853a3} /* (7, 0, 1) {real, imag} */,
  {32'h4087a5ea, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h4007a6e6, 32'hbf8fed82} /* (6, 31, 31) {real, imag} */,
  {32'hbe86a740, 32'h3e1164a8} /* (6, 31, 30) {real, imag} */,
  {32'h3d001704, 32'h3c6c2b28} /* (6, 31, 29) {real, imag} */,
  {32'h3db85e80, 32'h3d1a0173} /* (6, 31, 28) {real, imag} */,
  {32'hbd560a4d, 32'h3bbf46fc} /* (6, 31, 27) {real, imag} */,
  {32'hbc693588, 32'hbc0d4ede} /* (6, 31, 26) {real, imag} */,
  {32'h3ced11ed, 32'h3c6412f4} /* (6, 31, 25) {real, imag} */,
  {32'h3be527cc, 32'h3d57d07e} /* (6, 31, 24) {real, imag} */,
  {32'h3d05cea3, 32'hbc708582} /* (6, 31, 23) {real, imag} */,
  {32'h3c9220aa, 32'hbd00c528} /* (6, 31, 22) {real, imag} */,
  {32'h3c9b7db9, 32'h3cda3f03} /* (6, 31, 21) {real, imag} */,
  {32'hbc0faa60, 32'h3bd52054} /* (6, 31, 20) {real, imag} */,
  {32'h3d0251b2, 32'h3dd0e25c} /* (6, 31, 19) {real, imag} */,
  {32'hbcd4102d, 32'h3d9ff183} /* (6, 31, 18) {real, imag} */,
  {32'h3d0795f0, 32'hbb4c6eda} /* (6, 31, 17) {real, imag} */,
  {32'h3d225610, 32'h00000000} /* (6, 31, 16) {real, imag} */,
  {32'h3d0795f0, 32'h3b4c6eda} /* (6, 31, 15) {real, imag} */,
  {32'hbcd4102d, 32'hbd9ff183} /* (6, 31, 14) {real, imag} */,
  {32'h3d0251b2, 32'hbdd0e25c} /* (6, 31, 13) {real, imag} */,
  {32'hbc0faa60, 32'hbbd52054} /* (6, 31, 12) {real, imag} */,
  {32'h3c9b7db9, 32'hbcda3f03} /* (6, 31, 11) {real, imag} */,
  {32'h3c9220aa, 32'h3d00c528} /* (6, 31, 10) {real, imag} */,
  {32'h3d05cea3, 32'h3c708582} /* (6, 31, 9) {real, imag} */,
  {32'h3be527cc, 32'hbd57d07e} /* (6, 31, 8) {real, imag} */,
  {32'h3ced11ed, 32'hbc6412f4} /* (6, 31, 7) {real, imag} */,
  {32'hbc693588, 32'h3c0d4ede} /* (6, 31, 6) {real, imag} */,
  {32'hbd560a4d, 32'hbbbf46fc} /* (6, 31, 5) {real, imag} */,
  {32'h3db85e80, 32'hbd1a0173} /* (6, 31, 4) {real, imag} */,
  {32'h3d001704, 32'hbc6c2b28} /* (6, 31, 3) {real, imag} */,
  {32'hbe86a740, 32'hbe1164a8} /* (6, 31, 2) {real, imag} */,
  {32'h4007a6e6, 32'h3f8fed82} /* (6, 31, 1) {real, imag} */,
  {32'h4057527f, 32'h00000000} /* (6, 31, 0) {real, imag} */,
  {32'h40295e30, 32'hbf76467d} /* (6, 30, 31) {real, imag} */,
  {32'hbeec2662, 32'h3e088662} /* (6, 30, 30) {real, imag} */,
  {32'h3da4aab3, 32'h3b0843a0} /* (6, 30, 29) {real, imag} */,
  {32'h3dc68b46, 32'hb9491b00} /* (6, 30, 28) {real, imag} */,
  {32'hbe5c9ccc, 32'hbd36eb61} /* (6, 30, 27) {real, imag} */,
  {32'h3c8dbdac, 32'h3df91df3} /* (6, 30, 26) {real, imag} */,
  {32'hbd998ecc, 32'hbd517a26} /* (6, 30, 25) {real, imag} */,
  {32'hbda1e0fb, 32'h3cd9127c} /* (6, 30, 24) {real, imag} */,
  {32'hbc8b5eca, 32'h3db45621} /* (6, 30, 23) {real, imag} */,
  {32'h3daee690, 32'hbdb6ca9d} /* (6, 30, 22) {real, imag} */,
  {32'hbdf0cad9, 32'h3e0919b8} /* (6, 30, 21) {real, imag} */,
  {32'h3ce25432, 32'hbd84478e} /* (6, 30, 20) {real, imag} */,
  {32'h3d50a25b, 32'h3d211fc4} /* (6, 30, 19) {real, imag} */,
  {32'hbd802adb, 32'h3d328ec9} /* (6, 30, 18) {real, imag} */,
  {32'h3c4d827c, 32'h3d2d7af1} /* (6, 30, 17) {real, imag} */,
  {32'hbbf05aa4, 32'h00000000} /* (6, 30, 16) {real, imag} */,
  {32'h3c4d827c, 32'hbd2d7af1} /* (6, 30, 15) {real, imag} */,
  {32'hbd802adb, 32'hbd328ec9} /* (6, 30, 14) {real, imag} */,
  {32'h3d50a25b, 32'hbd211fc4} /* (6, 30, 13) {real, imag} */,
  {32'h3ce25432, 32'h3d84478e} /* (6, 30, 12) {real, imag} */,
  {32'hbdf0cad9, 32'hbe0919b8} /* (6, 30, 11) {real, imag} */,
  {32'h3daee690, 32'h3db6ca9d} /* (6, 30, 10) {real, imag} */,
  {32'hbc8b5eca, 32'hbdb45621} /* (6, 30, 9) {real, imag} */,
  {32'hbda1e0fb, 32'hbcd9127c} /* (6, 30, 8) {real, imag} */,
  {32'hbd998ecc, 32'h3d517a26} /* (6, 30, 7) {real, imag} */,
  {32'h3c8dbdac, 32'hbdf91df3} /* (6, 30, 6) {real, imag} */,
  {32'hbe5c9ccc, 32'h3d36eb61} /* (6, 30, 5) {real, imag} */,
  {32'h3dc68b46, 32'h39491b00} /* (6, 30, 4) {real, imag} */,
  {32'h3da4aab3, 32'hbb0843a0} /* (6, 30, 3) {real, imag} */,
  {32'hbeec2662, 32'hbe088662} /* (6, 30, 2) {real, imag} */,
  {32'h40295e30, 32'h3f76467d} /* (6, 30, 1) {real, imag} */,
  {32'h40598b5d, 32'h00000000} /* (6, 30, 0) {real, imag} */,
  {32'h401e9cf1, 32'hbf1abd58} /* (6, 29, 31) {real, imag} */,
  {32'hbf23c16e, 32'h3e568192} /* (6, 29, 30) {real, imag} */,
  {32'h3d91ece8, 32'hbe2beecb} /* (6, 29, 29) {real, imag} */,
  {32'h3e1d2241, 32'hbe1d2b62} /* (6, 29, 28) {real, imag} */,
  {32'hbe2ead86, 32'h3d536a97} /* (6, 29, 27) {real, imag} */,
  {32'h3d580b5f, 32'h3ccefed1} /* (6, 29, 26) {real, imag} */,
  {32'h3d2f233e, 32'hbd24b671} /* (6, 29, 25) {real, imag} */,
  {32'h3cc3718c, 32'h3cdc216b} /* (6, 29, 24) {real, imag} */,
  {32'hbd321a4c, 32'h3dafc5bc} /* (6, 29, 23) {real, imag} */,
  {32'hbcde2b13, 32'h3c7bccf2} /* (6, 29, 22) {real, imag} */,
  {32'hbb9410f8, 32'h3db1cfdd} /* (6, 29, 21) {real, imag} */,
  {32'hbca3ef76, 32'h3ba24c14} /* (6, 29, 20) {real, imag} */,
  {32'hbd8c93f6, 32'hbd4a31d4} /* (6, 29, 19) {real, imag} */,
  {32'hbd976432, 32'h3d45b8d1} /* (6, 29, 18) {real, imag} */,
  {32'h3cba205e, 32'hbc9299dc} /* (6, 29, 17) {real, imag} */,
  {32'h3d2ea4b2, 32'h00000000} /* (6, 29, 16) {real, imag} */,
  {32'h3cba205e, 32'h3c9299dc} /* (6, 29, 15) {real, imag} */,
  {32'hbd976432, 32'hbd45b8d1} /* (6, 29, 14) {real, imag} */,
  {32'hbd8c93f6, 32'h3d4a31d4} /* (6, 29, 13) {real, imag} */,
  {32'hbca3ef76, 32'hbba24c14} /* (6, 29, 12) {real, imag} */,
  {32'hbb9410f8, 32'hbdb1cfdd} /* (6, 29, 11) {real, imag} */,
  {32'hbcde2b13, 32'hbc7bccf2} /* (6, 29, 10) {real, imag} */,
  {32'hbd321a4c, 32'hbdafc5bc} /* (6, 29, 9) {real, imag} */,
  {32'h3cc3718c, 32'hbcdc216b} /* (6, 29, 8) {real, imag} */,
  {32'h3d2f233e, 32'h3d24b671} /* (6, 29, 7) {real, imag} */,
  {32'h3d580b5f, 32'hbccefed1} /* (6, 29, 6) {real, imag} */,
  {32'hbe2ead86, 32'hbd536a97} /* (6, 29, 5) {real, imag} */,
  {32'h3e1d2241, 32'h3e1d2b62} /* (6, 29, 4) {real, imag} */,
  {32'h3d91ece8, 32'h3e2beecb} /* (6, 29, 3) {real, imag} */,
  {32'hbf23c16e, 32'hbe568192} /* (6, 29, 2) {real, imag} */,
  {32'h401e9cf1, 32'h3f1abd58} /* (6, 29, 1) {real, imag} */,
  {32'h406062f0, 32'h00000000} /* (6, 29, 0) {real, imag} */,
  {32'h401eac1b, 32'hbeb0abd8} /* (6, 28, 31) {real, imag} */,
  {32'hbf4a4f73, 32'h3e945340} /* (6, 28, 30) {real, imag} */,
  {32'h3d98c8d9, 32'hbd482dee} /* (6, 28, 29) {real, imag} */,
  {32'h3dc8e183, 32'hbd92c458} /* (6, 28, 28) {real, imag} */,
  {32'hbea14ad2, 32'h3d840d9c} /* (6, 28, 27) {real, imag} */,
  {32'hbca9018e, 32'hbcd428a0} /* (6, 28, 26) {real, imag} */,
  {32'h3d1fe9e1, 32'hbd7fe680} /* (6, 28, 25) {real, imag} */,
  {32'hbca4982d, 32'h3ca71362} /* (6, 28, 24) {real, imag} */,
  {32'hbd6e63f0, 32'hbd23232c} /* (6, 28, 23) {real, imag} */,
  {32'h3cb98a2a, 32'hbd8ac41b} /* (6, 28, 22) {real, imag} */,
  {32'hbcf3cf87, 32'h3dcb9d6a} /* (6, 28, 21) {real, imag} */,
  {32'h3da71ce8, 32'hbd4c8e66} /* (6, 28, 20) {real, imag} */,
  {32'h3cd3e400, 32'hbc185e2c} /* (6, 28, 19) {real, imag} */,
  {32'h3c31d91b, 32'h3db5e0b9} /* (6, 28, 18) {real, imag} */,
  {32'h3bd9fa38, 32'hbd017ea6} /* (6, 28, 17) {real, imag} */,
  {32'hbca25595, 32'h00000000} /* (6, 28, 16) {real, imag} */,
  {32'h3bd9fa38, 32'h3d017ea6} /* (6, 28, 15) {real, imag} */,
  {32'h3c31d91b, 32'hbdb5e0b9} /* (6, 28, 14) {real, imag} */,
  {32'h3cd3e400, 32'h3c185e2c} /* (6, 28, 13) {real, imag} */,
  {32'h3da71ce8, 32'h3d4c8e66} /* (6, 28, 12) {real, imag} */,
  {32'hbcf3cf87, 32'hbdcb9d6a} /* (6, 28, 11) {real, imag} */,
  {32'h3cb98a2a, 32'h3d8ac41b} /* (6, 28, 10) {real, imag} */,
  {32'hbd6e63f0, 32'h3d23232c} /* (6, 28, 9) {real, imag} */,
  {32'hbca4982d, 32'hbca71362} /* (6, 28, 8) {real, imag} */,
  {32'h3d1fe9e1, 32'h3d7fe680} /* (6, 28, 7) {real, imag} */,
  {32'hbca9018e, 32'h3cd428a0} /* (6, 28, 6) {real, imag} */,
  {32'hbea14ad2, 32'hbd840d9c} /* (6, 28, 5) {real, imag} */,
  {32'h3dc8e183, 32'h3d92c458} /* (6, 28, 4) {real, imag} */,
  {32'h3d98c8d9, 32'h3d482dee} /* (6, 28, 3) {real, imag} */,
  {32'hbf4a4f73, 32'hbe945340} /* (6, 28, 2) {real, imag} */,
  {32'h401eac1b, 32'h3eb0abd8} /* (6, 28, 1) {real, imag} */,
  {32'h405c4b3a, 32'h00000000} /* (6, 28, 0) {real, imag} */,
  {32'h401c98cc, 32'hbededa76} /* (6, 27, 31) {real, imag} */,
  {32'hbf57b72d, 32'h3e964a55} /* (6, 27, 30) {real, imag} */,
  {32'h3d956521, 32'h3d0fd121} /* (6, 27, 29) {real, imag} */,
  {32'h3e1fae8e, 32'hbe2f11cd} /* (6, 27, 28) {real, imag} */,
  {32'hbe51da10, 32'h3d4ab146} /* (6, 27, 27) {real, imag} */,
  {32'h3db63638, 32'h3d47e9ca} /* (6, 27, 26) {real, imag} */,
  {32'h3c3136e8, 32'h3beeb6a0} /* (6, 27, 25) {real, imag} */,
  {32'hbd570b66, 32'hbd0d2c24} /* (6, 27, 24) {real, imag} */,
  {32'h3d341264, 32'hbc3b7c1c} /* (6, 27, 23) {real, imag} */,
  {32'hbd1fa8bc, 32'h3caebeaa} /* (6, 27, 22) {real, imag} */,
  {32'hbcf7b278, 32'h3bde8634} /* (6, 27, 21) {real, imag} */,
  {32'h3d8a3ad4, 32'hbab11ab8} /* (6, 27, 20) {real, imag} */,
  {32'h3d278daa, 32'hbcee31b9} /* (6, 27, 19) {real, imag} */,
  {32'hbdbac404, 32'h3df68ff2} /* (6, 27, 18) {real, imag} */,
  {32'hba3776c0, 32'hbcce3278} /* (6, 27, 17) {real, imag} */,
  {32'h3d1ac9e2, 32'h00000000} /* (6, 27, 16) {real, imag} */,
  {32'hba3776c0, 32'h3cce3278} /* (6, 27, 15) {real, imag} */,
  {32'hbdbac404, 32'hbdf68ff2} /* (6, 27, 14) {real, imag} */,
  {32'h3d278daa, 32'h3cee31b9} /* (6, 27, 13) {real, imag} */,
  {32'h3d8a3ad4, 32'h3ab11ab8} /* (6, 27, 12) {real, imag} */,
  {32'hbcf7b278, 32'hbbde8634} /* (6, 27, 11) {real, imag} */,
  {32'hbd1fa8bc, 32'hbcaebeaa} /* (6, 27, 10) {real, imag} */,
  {32'h3d341264, 32'h3c3b7c1c} /* (6, 27, 9) {real, imag} */,
  {32'hbd570b66, 32'h3d0d2c24} /* (6, 27, 8) {real, imag} */,
  {32'h3c3136e8, 32'hbbeeb6a0} /* (6, 27, 7) {real, imag} */,
  {32'h3db63638, 32'hbd47e9ca} /* (6, 27, 6) {real, imag} */,
  {32'hbe51da10, 32'hbd4ab146} /* (6, 27, 5) {real, imag} */,
  {32'h3e1fae8e, 32'h3e2f11cd} /* (6, 27, 4) {real, imag} */,
  {32'h3d956521, 32'hbd0fd121} /* (6, 27, 3) {real, imag} */,
  {32'hbf57b72d, 32'hbe964a55} /* (6, 27, 2) {real, imag} */,
  {32'h401c98cc, 32'h3ededa76} /* (6, 27, 1) {real, imag} */,
  {32'h404fb75b, 32'h00000000} /* (6, 27, 0) {real, imag} */,
  {32'h40130850, 32'hbe94ad76} /* (6, 26, 31) {real, imag} */,
  {32'hbf5be24a, 32'h3e13e0a5} /* (6, 26, 30) {real, imag} */,
  {32'hbc8775c4, 32'hbe0f3216} /* (6, 26, 29) {real, imag} */,
  {32'h3dffeb5f, 32'hbdd07310} /* (6, 26, 28) {real, imag} */,
  {32'hbe3dee41, 32'h3df23e8b} /* (6, 26, 27) {real, imag} */,
  {32'h3dfc02bb, 32'hbd3ce964} /* (6, 26, 26) {real, imag} */,
  {32'h3ccdb46c, 32'h3cf4a6b6} /* (6, 26, 25) {real, imag} */,
  {32'hb9675700, 32'h3d932393} /* (6, 26, 24) {real, imag} */,
  {32'hbc9b6c2a, 32'h3d9d693a} /* (6, 26, 23) {real, imag} */,
  {32'h3c6f4852, 32'hbd2c7cba} /* (6, 26, 22) {real, imag} */,
  {32'h3bbe7c10, 32'h3d536000} /* (6, 26, 21) {real, imag} */,
  {32'hbd14c0b8, 32'hbce07dce} /* (6, 26, 20) {real, imag} */,
  {32'hbc7b55ae, 32'hbdc1c18c} /* (6, 26, 19) {real, imag} */,
  {32'hbd3541d3, 32'h3d5e4f2c} /* (6, 26, 18) {real, imag} */,
  {32'hbd6312ce, 32'hbc9f73a8} /* (6, 26, 17) {real, imag} */,
  {32'hbc1f38cd, 32'h00000000} /* (6, 26, 16) {real, imag} */,
  {32'hbd6312ce, 32'h3c9f73a8} /* (6, 26, 15) {real, imag} */,
  {32'hbd3541d3, 32'hbd5e4f2c} /* (6, 26, 14) {real, imag} */,
  {32'hbc7b55ae, 32'h3dc1c18c} /* (6, 26, 13) {real, imag} */,
  {32'hbd14c0b8, 32'h3ce07dce} /* (6, 26, 12) {real, imag} */,
  {32'h3bbe7c10, 32'hbd536000} /* (6, 26, 11) {real, imag} */,
  {32'h3c6f4852, 32'h3d2c7cba} /* (6, 26, 10) {real, imag} */,
  {32'hbc9b6c2a, 32'hbd9d693a} /* (6, 26, 9) {real, imag} */,
  {32'hb9675700, 32'hbd932393} /* (6, 26, 8) {real, imag} */,
  {32'h3ccdb46c, 32'hbcf4a6b6} /* (6, 26, 7) {real, imag} */,
  {32'h3dfc02bb, 32'h3d3ce964} /* (6, 26, 6) {real, imag} */,
  {32'hbe3dee41, 32'hbdf23e8b} /* (6, 26, 5) {real, imag} */,
  {32'h3dffeb5f, 32'h3dd07310} /* (6, 26, 4) {real, imag} */,
  {32'hbc8775c4, 32'h3e0f3216} /* (6, 26, 3) {real, imag} */,
  {32'hbf5be24a, 32'hbe13e0a5} /* (6, 26, 2) {real, imag} */,
  {32'h40130850, 32'h3e94ad76} /* (6, 26, 1) {real, imag} */,
  {32'h403f8da8, 32'h00000000} /* (6, 26, 0) {real, imag} */,
  {32'h4008a9c1, 32'hbe91dd51} /* (6, 25, 31) {real, imag} */,
  {32'hbf4e24e9, 32'h3e07fecb} /* (6, 25, 30) {real, imag} */,
  {32'h3d56c334, 32'hbdbf78e6} /* (6, 25, 29) {real, imag} */,
  {32'h3d955817, 32'hbc846be6} /* (6, 25, 28) {real, imag} */,
  {32'hbda90ea2, 32'h3db3923a} /* (6, 25, 27) {real, imag} */,
  {32'h3d43d390, 32'hbe0e3216} /* (6, 25, 26) {real, imag} */,
  {32'hbbc84e6a, 32'h3d1d610f} /* (6, 25, 25) {real, imag} */,
  {32'hbe21f48a, 32'h3d838bce} /* (6, 25, 24) {real, imag} */,
  {32'hbda78e64, 32'h3ce0aa84} /* (6, 25, 23) {real, imag} */,
  {32'h3c97e22e, 32'h3b925e58} /* (6, 25, 22) {real, imag} */,
  {32'hbd9ce3d1, 32'h3d153494} /* (6, 25, 21) {real, imag} */,
  {32'h3d125ea4, 32'hbcb9c8ea} /* (6, 25, 20) {real, imag} */,
  {32'hbda8c309, 32'hbc39d3e2} /* (6, 25, 19) {real, imag} */,
  {32'h3d082859, 32'h3d71c919} /* (6, 25, 18) {real, imag} */,
  {32'hbc6fc424, 32'h3d9bf61c} /* (6, 25, 17) {real, imag} */,
  {32'hbc164408, 32'h00000000} /* (6, 25, 16) {real, imag} */,
  {32'hbc6fc424, 32'hbd9bf61c} /* (6, 25, 15) {real, imag} */,
  {32'h3d082859, 32'hbd71c919} /* (6, 25, 14) {real, imag} */,
  {32'hbda8c309, 32'h3c39d3e2} /* (6, 25, 13) {real, imag} */,
  {32'h3d125ea4, 32'h3cb9c8ea} /* (6, 25, 12) {real, imag} */,
  {32'hbd9ce3d1, 32'hbd153494} /* (6, 25, 11) {real, imag} */,
  {32'h3c97e22e, 32'hbb925e58} /* (6, 25, 10) {real, imag} */,
  {32'hbda78e64, 32'hbce0aa84} /* (6, 25, 9) {real, imag} */,
  {32'hbe21f48a, 32'hbd838bce} /* (6, 25, 8) {real, imag} */,
  {32'hbbc84e6a, 32'hbd1d610f} /* (6, 25, 7) {real, imag} */,
  {32'h3d43d390, 32'h3e0e3216} /* (6, 25, 6) {real, imag} */,
  {32'hbda90ea2, 32'hbdb3923a} /* (6, 25, 5) {real, imag} */,
  {32'h3d955817, 32'h3c846be6} /* (6, 25, 4) {real, imag} */,
  {32'h3d56c334, 32'h3dbf78e6} /* (6, 25, 3) {real, imag} */,
  {32'hbf4e24e9, 32'hbe07fecb} /* (6, 25, 2) {real, imag} */,
  {32'h4008a9c1, 32'h3e91dd51} /* (6, 25, 1) {real, imag} */,
  {32'h4032e6f2, 32'h00000000} /* (6, 25, 0) {real, imag} */,
  {32'h3feb9357, 32'hbe98fd54} /* (6, 24, 31) {real, imag} */,
  {32'hbf3f40c5, 32'h3e01d44c} /* (6, 24, 30) {real, imag} */,
  {32'h3ca99b68, 32'hbd1434b1} /* (6, 24, 29) {real, imag} */,
  {32'h3af62340, 32'hbd030883} /* (6, 24, 28) {real, imag} */,
  {32'hbddb7584, 32'h3d493860} /* (6, 24, 27) {real, imag} */,
  {32'hbbe49d90, 32'hbd15fccc} /* (6, 24, 26) {real, imag} */,
  {32'h3dbce716, 32'h3c29a5c0} /* (6, 24, 25) {real, imag} */,
  {32'hbdb1db51, 32'h3d7558a2} /* (6, 24, 24) {real, imag} */,
  {32'hbc8fcd6d, 32'hbcdfb8ec} /* (6, 24, 23) {real, imag} */,
  {32'hbdc756ca, 32'hbc4c0efa} /* (6, 24, 22) {real, imag} */,
  {32'hbcc8324e, 32'h3d7548b2} /* (6, 24, 21) {real, imag} */,
  {32'h3d4857b6, 32'hbe1f4774} /* (6, 24, 20) {real, imag} */,
  {32'h3daf3eb6, 32'h3db9317a} /* (6, 24, 19) {real, imag} */,
  {32'h3ce7a0a7, 32'h3d3d1ba7} /* (6, 24, 18) {real, imag} */,
  {32'h3c869b98, 32'hbbf7f894} /* (6, 24, 17) {real, imag} */,
  {32'h3d05c26f, 32'h00000000} /* (6, 24, 16) {real, imag} */,
  {32'h3c869b98, 32'h3bf7f894} /* (6, 24, 15) {real, imag} */,
  {32'h3ce7a0a7, 32'hbd3d1ba7} /* (6, 24, 14) {real, imag} */,
  {32'h3daf3eb6, 32'hbdb9317a} /* (6, 24, 13) {real, imag} */,
  {32'h3d4857b6, 32'h3e1f4774} /* (6, 24, 12) {real, imag} */,
  {32'hbcc8324e, 32'hbd7548b2} /* (6, 24, 11) {real, imag} */,
  {32'hbdc756ca, 32'h3c4c0efa} /* (6, 24, 10) {real, imag} */,
  {32'hbc8fcd6d, 32'h3cdfb8ec} /* (6, 24, 9) {real, imag} */,
  {32'hbdb1db51, 32'hbd7558a2} /* (6, 24, 8) {real, imag} */,
  {32'h3dbce716, 32'hbc29a5c0} /* (6, 24, 7) {real, imag} */,
  {32'hbbe49d90, 32'h3d15fccc} /* (6, 24, 6) {real, imag} */,
  {32'hbddb7584, 32'hbd493860} /* (6, 24, 5) {real, imag} */,
  {32'h3af62340, 32'h3d030883} /* (6, 24, 4) {real, imag} */,
  {32'h3ca99b68, 32'h3d1434b1} /* (6, 24, 3) {real, imag} */,
  {32'hbf3f40c5, 32'hbe01d44c} /* (6, 24, 2) {real, imag} */,
  {32'h3feb9357, 32'h3e98fd54} /* (6, 24, 1) {real, imag} */,
  {32'h4026973a, 32'h00000000} /* (6, 24, 0) {real, imag} */,
  {32'h3fafb9df, 32'hbecad4d7} /* (6, 23, 31) {real, imag} */,
  {32'hbf236a69, 32'h3d808a6a} /* (6, 23, 30) {real, imag} */,
  {32'h3d29cce3, 32'hbdeb0f83} /* (6, 23, 29) {real, imag} */,
  {32'h3d6166c0, 32'hbd2a60d8} /* (6, 23, 28) {real, imag} */,
  {32'hbd861237, 32'h3b552a80} /* (6, 23, 27) {real, imag} */,
  {32'hbc858e1b, 32'hbda6bbd3} /* (6, 23, 26) {real, imag} */,
  {32'hbcb0a85e, 32'hbd75a488} /* (6, 23, 25) {real, imag} */,
  {32'hbd947597, 32'hbd4f47ac} /* (6, 23, 24) {real, imag} */,
  {32'h3ca6671f, 32'h3dac1d82} /* (6, 23, 23) {real, imag} */,
  {32'hbd8a109c, 32'h3be8103c} /* (6, 23, 22) {real, imag} */,
  {32'hbc7e0140, 32'h3d5c7e48} /* (6, 23, 21) {real, imag} */,
  {32'h3b71cba8, 32'hbd09665e} /* (6, 23, 20) {real, imag} */,
  {32'h3ce03829, 32'h3d436d68} /* (6, 23, 19) {real, imag} */,
  {32'hbd6b5fc3, 32'hbd5f12bc} /* (6, 23, 18) {real, imag} */,
  {32'h3cffc7a4, 32'hbd13352c} /* (6, 23, 17) {real, imag} */,
  {32'h3c890fde, 32'h00000000} /* (6, 23, 16) {real, imag} */,
  {32'h3cffc7a4, 32'h3d13352c} /* (6, 23, 15) {real, imag} */,
  {32'hbd6b5fc3, 32'h3d5f12bc} /* (6, 23, 14) {real, imag} */,
  {32'h3ce03829, 32'hbd436d68} /* (6, 23, 13) {real, imag} */,
  {32'h3b71cba8, 32'h3d09665e} /* (6, 23, 12) {real, imag} */,
  {32'hbc7e0140, 32'hbd5c7e48} /* (6, 23, 11) {real, imag} */,
  {32'hbd8a109c, 32'hbbe8103c} /* (6, 23, 10) {real, imag} */,
  {32'h3ca6671f, 32'hbdac1d82} /* (6, 23, 9) {real, imag} */,
  {32'hbd947597, 32'h3d4f47ac} /* (6, 23, 8) {real, imag} */,
  {32'hbcb0a85e, 32'h3d75a488} /* (6, 23, 7) {real, imag} */,
  {32'hbc858e1b, 32'h3da6bbd3} /* (6, 23, 6) {real, imag} */,
  {32'hbd861237, 32'hbb552a80} /* (6, 23, 5) {real, imag} */,
  {32'h3d6166c0, 32'h3d2a60d8} /* (6, 23, 4) {real, imag} */,
  {32'h3d29cce3, 32'h3deb0f83} /* (6, 23, 3) {real, imag} */,
  {32'hbf236a69, 32'hbd808a6a} /* (6, 23, 2) {real, imag} */,
  {32'h3fafb9df, 32'h3ecad4d7} /* (6, 23, 1) {real, imag} */,
  {32'h400ecaa4, 32'h00000000} /* (6, 23, 0) {real, imag} */,
  {32'h3f6f0367, 32'hbeae6fd2} /* (6, 22, 31) {real, imag} */,
  {32'hbf331620, 32'h3d7a5af4} /* (6, 22, 30) {real, imag} */,
  {32'hbd9be178, 32'hbe245b78} /* (6, 22, 29) {real, imag} */,
  {32'h3e17eae2, 32'hbcda1ce8} /* (6, 22, 28) {real, imag} */,
  {32'hbd81b8e6, 32'h3e0144be} /* (6, 22, 27) {real, imag} */,
  {32'h3d3f465c, 32'h3c9e4972} /* (6, 22, 26) {real, imag} */,
  {32'h3de99ec8, 32'hbd4866d4} /* (6, 22, 25) {real, imag} */,
  {32'hbda92df8, 32'h3b909f00} /* (6, 22, 24) {real, imag} */,
  {32'hbdec15fb, 32'hbc66bb22} /* (6, 22, 23) {real, imag} */,
  {32'h3da5fceb, 32'hbd195e46} /* (6, 22, 22) {real, imag} */,
  {32'hba8d3180, 32'h3bb14948} /* (6, 22, 21) {real, imag} */,
  {32'h3cb9e0f8, 32'hbc6c9798} /* (6, 22, 20) {real, imag} */,
  {32'hbd9b49be, 32'h3d7352cb} /* (6, 22, 19) {real, imag} */,
  {32'h3c95f6e8, 32'h3d388fe2} /* (6, 22, 18) {real, imag} */,
  {32'hbc88c223, 32'hbc94b424} /* (6, 22, 17) {real, imag} */,
  {32'hbd03f83a, 32'h00000000} /* (6, 22, 16) {real, imag} */,
  {32'hbc88c223, 32'h3c94b424} /* (6, 22, 15) {real, imag} */,
  {32'h3c95f6e8, 32'hbd388fe2} /* (6, 22, 14) {real, imag} */,
  {32'hbd9b49be, 32'hbd7352cb} /* (6, 22, 13) {real, imag} */,
  {32'h3cb9e0f8, 32'h3c6c9798} /* (6, 22, 12) {real, imag} */,
  {32'hba8d3180, 32'hbbb14948} /* (6, 22, 11) {real, imag} */,
  {32'h3da5fceb, 32'h3d195e46} /* (6, 22, 10) {real, imag} */,
  {32'hbdec15fb, 32'h3c66bb22} /* (6, 22, 9) {real, imag} */,
  {32'hbda92df8, 32'hbb909f00} /* (6, 22, 8) {real, imag} */,
  {32'h3de99ec8, 32'h3d4866d4} /* (6, 22, 7) {real, imag} */,
  {32'h3d3f465c, 32'hbc9e4972} /* (6, 22, 6) {real, imag} */,
  {32'hbd81b8e6, 32'hbe0144be} /* (6, 22, 5) {real, imag} */,
  {32'h3e17eae2, 32'h3cda1ce8} /* (6, 22, 4) {real, imag} */,
  {32'hbd9be178, 32'h3e245b78} /* (6, 22, 3) {real, imag} */,
  {32'hbf331620, 32'hbd7a5af4} /* (6, 22, 2) {real, imag} */,
  {32'h3f6f0367, 32'h3eae6fd2} /* (6, 22, 1) {real, imag} */,
  {32'h3fe755a4, 32'h00000000} /* (6, 22, 0) {real, imag} */,
  {32'h3e967708, 32'hbe3b7084} /* (6, 21, 31) {real, imag} */,
  {32'hbeb67964, 32'hbe10441f} /* (6, 21, 30) {real, imag} */,
  {32'hbe431ff5, 32'hbe3963b1} /* (6, 21, 29) {real, imag} */,
  {32'hbc71daf6, 32'h3d7944e3} /* (6, 21, 28) {real, imag} */,
  {32'h3d5b2c3e, 32'h3d938c87} /* (6, 21, 27) {real, imag} */,
  {32'hbd0b347c, 32'h3dd0d68b} /* (6, 21, 26) {real, imag} */,
  {32'h3d8a7dc8, 32'h3dbdc1d4} /* (6, 21, 25) {real, imag} */,
  {32'hbd4cd535, 32'h3cd0372b} /* (6, 21, 24) {real, imag} */,
  {32'h3d27bcc6, 32'hbab33d00} /* (6, 21, 23) {real, imag} */,
  {32'hbd02514b, 32'hbd86d99f} /* (6, 21, 22) {real, imag} */,
  {32'hbd596e28, 32'h3d07d484} /* (6, 21, 21) {real, imag} */,
  {32'h3cf3288a, 32'h3d812890} /* (6, 21, 20) {real, imag} */,
  {32'h3d09811e, 32'h3d8f08ed} /* (6, 21, 19) {real, imag} */,
  {32'hbc952762, 32'h3c8eab61} /* (6, 21, 18) {real, imag} */,
  {32'hbcc792ba, 32'hbe073cb8} /* (6, 21, 17) {real, imag} */,
  {32'h3d9d553a, 32'h00000000} /* (6, 21, 16) {real, imag} */,
  {32'hbcc792ba, 32'h3e073cb8} /* (6, 21, 15) {real, imag} */,
  {32'hbc952762, 32'hbc8eab61} /* (6, 21, 14) {real, imag} */,
  {32'h3d09811e, 32'hbd8f08ed} /* (6, 21, 13) {real, imag} */,
  {32'h3cf3288a, 32'hbd812890} /* (6, 21, 12) {real, imag} */,
  {32'hbd596e28, 32'hbd07d484} /* (6, 21, 11) {real, imag} */,
  {32'hbd02514b, 32'h3d86d99f} /* (6, 21, 10) {real, imag} */,
  {32'h3d27bcc6, 32'h3ab33d00} /* (6, 21, 9) {real, imag} */,
  {32'hbd4cd535, 32'hbcd0372b} /* (6, 21, 8) {real, imag} */,
  {32'h3d8a7dc8, 32'hbdbdc1d4} /* (6, 21, 7) {real, imag} */,
  {32'hbd0b347c, 32'hbdd0d68b} /* (6, 21, 6) {real, imag} */,
  {32'h3d5b2c3e, 32'hbd938c87} /* (6, 21, 5) {real, imag} */,
  {32'hbc71daf6, 32'hbd7944e3} /* (6, 21, 4) {real, imag} */,
  {32'hbe431ff5, 32'h3e3963b1} /* (6, 21, 3) {real, imag} */,
  {32'hbeb67964, 32'h3e10441f} /* (6, 21, 2) {real, imag} */,
  {32'h3e967708, 32'h3e3b7084} /* (6, 21, 1) {real, imag} */,
  {32'h3fa009c0, 32'h00000000} /* (6, 21, 0) {real, imag} */,
  {32'hbf430f92, 32'hbe08aaf8} /* (6, 20, 31) {real, imag} */,
  {32'h3eb9985c, 32'hbe386c8d} /* (6, 20, 30) {real, imag} */,
  {32'hbe323e9c, 32'hbe15ee62} /* (6, 20, 29) {real, imag} */,
  {32'hbe0bc4da, 32'hbd374b98} /* (6, 20, 28) {real, imag} */,
  {32'h3ddedf7b, 32'hbadd2ca0} /* (6, 20, 27) {real, imag} */,
  {32'hbc86b3fe, 32'h3d1c4327} /* (6, 20, 26) {real, imag} */,
  {32'h3ceacfa2, 32'h3ba1e330} /* (6, 20, 25) {real, imag} */,
  {32'h3cf75bcc, 32'hbb7be8c8} /* (6, 20, 24) {real, imag} */,
  {32'hbd6af5bf, 32'h3d077cdd} /* (6, 20, 23) {real, imag} */,
  {32'hbdc40b66, 32'hbca6d29c} /* (6, 20, 22) {real, imag} */,
  {32'h3d5817c0, 32'hbd51c0ea} /* (6, 20, 21) {real, imag} */,
  {32'h3d2e0f3c, 32'hbb0a0c20} /* (6, 20, 20) {real, imag} */,
  {32'hbc9a01b4, 32'hbd2f39b4} /* (6, 20, 19) {real, imag} */,
  {32'h3c21a3f2, 32'hbc79ebbc} /* (6, 20, 18) {real, imag} */,
  {32'h3d68a809, 32'h3d804a90} /* (6, 20, 17) {real, imag} */,
  {32'h3dbc1498, 32'h00000000} /* (6, 20, 16) {real, imag} */,
  {32'h3d68a809, 32'hbd804a90} /* (6, 20, 15) {real, imag} */,
  {32'h3c21a3f2, 32'h3c79ebbc} /* (6, 20, 14) {real, imag} */,
  {32'hbc9a01b4, 32'h3d2f39b4} /* (6, 20, 13) {real, imag} */,
  {32'h3d2e0f3c, 32'h3b0a0c20} /* (6, 20, 12) {real, imag} */,
  {32'h3d5817c0, 32'h3d51c0ea} /* (6, 20, 11) {real, imag} */,
  {32'hbdc40b66, 32'h3ca6d29c} /* (6, 20, 10) {real, imag} */,
  {32'hbd6af5bf, 32'hbd077cdd} /* (6, 20, 9) {real, imag} */,
  {32'h3cf75bcc, 32'h3b7be8c8} /* (6, 20, 8) {real, imag} */,
  {32'h3ceacfa2, 32'hbba1e330} /* (6, 20, 7) {real, imag} */,
  {32'hbc86b3fe, 32'hbd1c4327} /* (6, 20, 6) {real, imag} */,
  {32'h3ddedf7b, 32'h3add2ca0} /* (6, 20, 5) {real, imag} */,
  {32'hbe0bc4da, 32'h3d374b98} /* (6, 20, 4) {real, imag} */,
  {32'hbe323e9c, 32'h3e15ee62} /* (6, 20, 3) {real, imag} */,
  {32'h3eb9985c, 32'h3e386c8d} /* (6, 20, 2) {real, imag} */,
  {32'hbf430f92, 32'h3e08aaf8} /* (6, 20, 1) {real, imag} */,
  {32'h3e4b5c80, 32'h00000000} /* (6, 20, 0) {real, imag} */,
  {32'hbfb0c8e3, 32'h3e53e210} /* (6, 19, 31) {real, imag} */,
  {32'h3f1dffa8, 32'hbdc13162} /* (6, 19, 30) {real, imag} */,
  {32'hbe56c294, 32'hbe9accd6} /* (6, 19, 29) {real, imag} */,
  {32'hbe0185d8, 32'hbd15b02b} /* (6, 19, 28) {real, imag} */,
  {32'h3e02a388, 32'h3bf87104} /* (6, 19, 27) {real, imag} */,
  {32'hbd32f9ba, 32'h3cc2cf7f} /* (6, 19, 26) {real, imag} */,
  {32'hbc709cdc, 32'hbdc72606} /* (6, 19, 25) {real, imag} */,
  {32'h3cec3e48, 32'hbc9daaa5} /* (6, 19, 24) {real, imag} */,
  {32'hbd8b4cba, 32'hbd8bc5b8} /* (6, 19, 23) {real, imag} */,
  {32'h3bf28ab8, 32'hbd9677f5} /* (6, 19, 22) {real, imag} */,
  {32'h3de2bb12, 32'h3c9edd04} /* (6, 19, 21) {real, imag} */,
  {32'hbd97289f, 32'h3d3c8846} /* (6, 19, 20) {real, imag} */,
  {32'hbc5c8512, 32'hbcdcf4b8} /* (6, 19, 19) {real, imag} */,
  {32'h3c3ba174, 32'h3cb91e00} /* (6, 19, 18) {real, imag} */,
  {32'h3ca0c2a0, 32'hbbcdc088} /* (6, 19, 17) {real, imag} */,
  {32'h3d031ea8, 32'h00000000} /* (6, 19, 16) {real, imag} */,
  {32'h3ca0c2a0, 32'h3bcdc088} /* (6, 19, 15) {real, imag} */,
  {32'h3c3ba174, 32'hbcb91e00} /* (6, 19, 14) {real, imag} */,
  {32'hbc5c8512, 32'h3cdcf4b8} /* (6, 19, 13) {real, imag} */,
  {32'hbd97289f, 32'hbd3c8846} /* (6, 19, 12) {real, imag} */,
  {32'h3de2bb12, 32'hbc9edd04} /* (6, 19, 11) {real, imag} */,
  {32'h3bf28ab8, 32'h3d9677f5} /* (6, 19, 10) {real, imag} */,
  {32'hbd8b4cba, 32'h3d8bc5b8} /* (6, 19, 9) {real, imag} */,
  {32'h3cec3e48, 32'h3c9daaa5} /* (6, 19, 8) {real, imag} */,
  {32'hbc709cdc, 32'h3dc72606} /* (6, 19, 7) {real, imag} */,
  {32'hbd32f9ba, 32'hbcc2cf7f} /* (6, 19, 6) {real, imag} */,
  {32'h3e02a388, 32'hbbf87104} /* (6, 19, 5) {real, imag} */,
  {32'hbe0185d8, 32'h3d15b02b} /* (6, 19, 4) {real, imag} */,
  {32'hbe56c294, 32'h3e9accd6} /* (6, 19, 3) {real, imag} */,
  {32'h3f1dffa8, 32'h3dc13162} /* (6, 19, 2) {real, imag} */,
  {32'hbfb0c8e3, 32'hbe53e210} /* (6, 19, 1) {real, imag} */,
  {32'hbed1a462, 32'h00000000} /* (6, 19, 0) {real, imag} */,
  {32'hbfe88566, 32'h3e28dad7} /* (6, 18, 31) {real, imag} */,
  {32'h3f46c93c, 32'hbc9f0ef0} /* (6, 18, 30) {real, imag} */,
  {32'hbe15fa3b, 32'hbe31ab46} /* (6, 18, 29) {real, imag} */,
  {32'hbe2e777b, 32'hbd5f031a} /* (6, 18, 28) {real, imag} */,
  {32'h3e215f31, 32'h3c642d8c} /* (6, 18, 27) {real, imag} */,
  {32'h3d95032a, 32'h3c93dc97} /* (6, 18, 26) {real, imag} */,
  {32'h3c844402, 32'h3cf88235} /* (6, 18, 25) {real, imag} */,
  {32'hbdbd96d6, 32'h3d4c2222} /* (6, 18, 24) {real, imag} */,
  {32'hbd15966d, 32'h3c1ecdd9} /* (6, 18, 23) {real, imag} */,
  {32'h3ddd1f00, 32'h3c314a54} /* (6, 18, 22) {real, imag} */,
  {32'hbd1ae48d, 32'hbda331a6} /* (6, 18, 21) {real, imag} */,
  {32'hbda67722, 32'h3c788cc4} /* (6, 18, 20) {real, imag} */,
  {32'h3d27da53, 32'h3ccc4f72} /* (6, 18, 19) {real, imag} */,
  {32'h3d465e25, 32'hbc494614} /* (6, 18, 18) {real, imag} */,
  {32'h3c3383d6, 32'h3c81d486} /* (6, 18, 17) {real, imag} */,
  {32'hbd8b31d0, 32'h00000000} /* (6, 18, 16) {real, imag} */,
  {32'h3c3383d6, 32'hbc81d486} /* (6, 18, 15) {real, imag} */,
  {32'h3d465e25, 32'h3c494614} /* (6, 18, 14) {real, imag} */,
  {32'h3d27da53, 32'hbccc4f72} /* (6, 18, 13) {real, imag} */,
  {32'hbda67722, 32'hbc788cc4} /* (6, 18, 12) {real, imag} */,
  {32'hbd1ae48d, 32'h3da331a6} /* (6, 18, 11) {real, imag} */,
  {32'h3ddd1f00, 32'hbc314a54} /* (6, 18, 10) {real, imag} */,
  {32'hbd15966d, 32'hbc1ecdd9} /* (6, 18, 9) {real, imag} */,
  {32'hbdbd96d6, 32'hbd4c2222} /* (6, 18, 8) {real, imag} */,
  {32'h3c844402, 32'hbcf88235} /* (6, 18, 7) {real, imag} */,
  {32'h3d95032a, 32'hbc93dc97} /* (6, 18, 6) {real, imag} */,
  {32'h3e215f31, 32'hbc642d8c} /* (6, 18, 5) {real, imag} */,
  {32'hbe2e777b, 32'h3d5f031a} /* (6, 18, 4) {real, imag} */,
  {32'hbe15fa3b, 32'h3e31ab46} /* (6, 18, 3) {real, imag} */,
  {32'h3f46c93c, 32'h3c9f0ef0} /* (6, 18, 2) {real, imag} */,
  {32'hbfe88566, 32'hbe28dad7} /* (6, 18, 1) {real, imag} */,
  {32'hbf3eafb1, 32'h00000000} /* (6, 18, 0) {real, imag} */,
  {32'hc003cdbf, 32'h3e0ad0bb} /* (6, 17, 31) {real, imag} */,
  {32'h3f614028, 32'hbdada668} /* (6, 17, 30) {real, imag} */,
  {32'hbd856265, 32'hbcff83d8} /* (6, 17, 29) {real, imag} */,
  {32'hbdea8e91, 32'hbd3e9df4} /* (6, 17, 28) {real, imag} */,
  {32'h3dd17cd5, 32'h3d948515} /* (6, 17, 27) {real, imag} */,
  {32'h3ba2fb48, 32'h3dbcf1c6} /* (6, 17, 26) {real, imag} */,
  {32'h3c229a86, 32'hbdcb5faa} /* (6, 17, 25) {real, imag} */,
  {32'h3de0791b, 32'hbd470049} /* (6, 17, 24) {real, imag} */,
  {32'hbd6536d3, 32'h3d5b37ec} /* (6, 17, 23) {real, imag} */,
  {32'hbd79c531, 32'h3d62a2ce} /* (6, 17, 22) {real, imag} */,
  {32'h3d1a3b4a, 32'hbda66a24} /* (6, 17, 21) {real, imag} */,
  {32'hbc2475e4, 32'hbd3ccd72} /* (6, 17, 20) {real, imag} */,
  {32'h3d62ff0c, 32'h3c886b07} /* (6, 17, 19) {real, imag} */,
  {32'hbd5c6b0a, 32'h3d254f1e} /* (6, 17, 18) {real, imag} */,
  {32'hbb42e9e4, 32'hbd34bc62} /* (6, 17, 17) {real, imag} */,
  {32'h3d0f8eab, 32'h00000000} /* (6, 17, 16) {real, imag} */,
  {32'hbb42e9e4, 32'h3d34bc62} /* (6, 17, 15) {real, imag} */,
  {32'hbd5c6b0a, 32'hbd254f1e} /* (6, 17, 14) {real, imag} */,
  {32'h3d62ff0c, 32'hbc886b07} /* (6, 17, 13) {real, imag} */,
  {32'hbc2475e4, 32'h3d3ccd72} /* (6, 17, 12) {real, imag} */,
  {32'h3d1a3b4a, 32'h3da66a24} /* (6, 17, 11) {real, imag} */,
  {32'hbd79c531, 32'hbd62a2ce} /* (6, 17, 10) {real, imag} */,
  {32'hbd6536d3, 32'hbd5b37ec} /* (6, 17, 9) {real, imag} */,
  {32'h3de0791b, 32'h3d470049} /* (6, 17, 8) {real, imag} */,
  {32'h3c229a86, 32'h3dcb5faa} /* (6, 17, 7) {real, imag} */,
  {32'h3ba2fb48, 32'hbdbcf1c6} /* (6, 17, 6) {real, imag} */,
  {32'h3dd17cd5, 32'hbd948515} /* (6, 17, 5) {real, imag} */,
  {32'hbdea8e91, 32'h3d3e9df4} /* (6, 17, 4) {real, imag} */,
  {32'hbd856265, 32'h3cff83d8} /* (6, 17, 3) {real, imag} */,
  {32'h3f614028, 32'h3dada668} /* (6, 17, 2) {real, imag} */,
  {32'hc003cdbf, 32'hbe0ad0bb} /* (6, 17, 1) {real, imag} */,
  {32'hbf90a38a, 32'h00000000} /* (6, 17, 0) {real, imag} */,
  {32'hc010a1d4, 32'h3d300420} /* (6, 16, 31) {real, imag} */,
  {32'h3f4892b4, 32'hbe4e9d43} /* (6, 16, 30) {real, imag} */,
  {32'hbdd7b351, 32'hbd226afe} /* (6, 16, 29) {real, imag} */,
  {32'hbd9ea0b0, 32'hbdf2ae3e} /* (6, 16, 28) {real, imag} */,
  {32'h3dba71c6, 32'hbd8af93a} /* (6, 16, 27) {real, imag} */,
  {32'h3cd35f4a, 32'hbe0e6d4e} /* (6, 16, 26) {real, imag} */,
  {32'h3d6b3f88, 32'h3d3f18b0} /* (6, 16, 25) {real, imag} */,
  {32'h3d522916, 32'hbdd1b7ec} /* (6, 16, 24) {real, imag} */,
  {32'hbd77d978, 32'hbd9aaa48} /* (6, 16, 23) {real, imag} */,
  {32'h3c337114, 32'hbe02d09e} /* (6, 16, 22) {real, imag} */,
  {32'h3d94c0f0, 32'hbd52af6e} /* (6, 16, 21) {real, imag} */,
  {32'hbd295c10, 32'hbd3b716e} /* (6, 16, 20) {real, imag} */,
  {32'h3c84664c, 32'h3dadadb4} /* (6, 16, 19) {real, imag} */,
  {32'h3c15e430, 32'hb9a81b00} /* (6, 16, 18) {real, imag} */,
  {32'h3d59dc64, 32'hbd298518} /* (6, 16, 17) {real, imag} */,
  {32'h3cdfd182, 32'h00000000} /* (6, 16, 16) {real, imag} */,
  {32'h3d59dc64, 32'h3d298518} /* (6, 16, 15) {real, imag} */,
  {32'h3c15e430, 32'h39a81b00} /* (6, 16, 14) {real, imag} */,
  {32'h3c84664c, 32'hbdadadb4} /* (6, 16, 13) {real, imag} */,
  {32'hbd295c10, 32'h3d3b716e} /* (6, 16, 12) {real, imag} */,
  {32'h3d94c0f0, 32'h3d52af6e} /* (6, 16, 11) {real, imag} */,
  {32'h3c337114, 32'h3e02d09e} /* (6, 16, 10) {real, imag} */,
  {32'hbd77d978, 32'h3d9aaa48} /* (6, 16, 9) {real, imag} */,
  {32'h3d522916, 32'h3dd1b7ec} /* (6, 16, 8) {real, imag} */,
  {32'h3d6b3f88, 32'hbd3f18b0} /* (6, 16, 7) {real, imag} */,
  {32'h3cd35f4a, 32'h3e0e6d4e} /* (6, 16, 6) {real, imag} */,
  {32'h3dba71c6, 32'h3d8af93a} /* (6, 16, 5) {real, imag} */,
  {32'hbd9ea0b0, 32'h3df2ae3e} /* (6, 16, 4) {real, imag} */,
  {32'hbdd7b351, 32'h3d226afe} /* (6, 16, 3) {real, imag} */,
  {32'h3f4892b4, 32'h3e4e9d43} /* (6, 16, 2) {real, imag} */,
  {32'hc010a1d4, 32'hbd300420} /* (6, 16, 1) {real, imag} */,
  {32'hbfcf5ba8, 32'h00000000} /* (6, 16, 0) {real, imag} */,
  {32'hc00ce4c5, 32'hbc0b8d30} /* (6, 15, 31) {real, imag} */,
  {32'h3f4353c4, 32'hbe0955b8} /* (6, 15, 30) {real, imag} */,
  {32'hbcd1dd54, 32'hbe26253f} /* (6, 15, 29) {real, imag} */,
  {32'hbe175b5d, 32'hbe503e71} /* (6, 15, 28) {real, imag} */,
  {32'h3d9e390f, 32'hbdf664c5} /* (6, 15, 27) {real, imag} */,
  {32'h3df97580, 32'hbe55e289} /* (6, 15, 26) {real, imag} */,
  {32'h3d899bc9, 32'h3d533087} /* (6, 15, 25) {real, imag} */,
  {32'h3d8af1bf, 32'hbd0ebccf} /* (6, 15, 24) {real, imag} */,
  {32'hbd84f549, 32'h3c988f00} /* (6, 15, 23) {real, imag} */,
  {32'h3db6333c, 32'h3cc8ae40} /* (6, 15, 22) {real, imag} */,
  {32'hbb9ece2c, 32'hbd7170c9} /* (6, 15, 21) {real, imag} */,
  {32'h3d46816f, 32'hbdad3c2d} /* (6, 15, 20) {real, imag} */,
  {32'hbd679e70, 32'hbcf33cf5} /* (6, 15, 19) {real, imag} */,
  {32'hbd1ee12a, 32'h3beb7394} /* (6, 15, 18) {real, imag} */,
  {32'hbcb553ac, 32'h3d54ccb2} /* (6, 15, 17) {real, imag} */,
  {32'h3da49848, 32'h00000000} /* (6, 15, 16) {real, imag} */,
  {32'hbcb553ac, 32'hbd54ccb2} /* (6, 15, 15) {real, imag} */,
  {32'hbd1ee12a, 32'hbbeb7394} /* (6, 15, 14) {real, imag} */,
  {32'hbd679e70, 32'h3cf33cf5} /* (6, 15, 13) {real, imag} */,
  {32'h3d46816f, 32'h3dad3c2d} /* (6, 15, 12) {real, imag} */,
  {32'hbb9ece2c, 32'h3d7170c9} /* (6, 15, 11) {real, imag} */,
  {32'h3db6333c, 32'hbcc8ae40} /* (6, 15, 10) {real, imag} */,
  {32'hbd84f549, 32'hbc988f00} /* (6, 15, 9) {real, imag} */,
  {32'h3d8af1bf, 32'h3d0ebccf} /* (6, 15, 8) {real, imag} */,
  {32'h3d899bc9, 32'hbd533087} /* (6, 15, 7) {real, imag} */,
  {32'h3df97580, 32'h3e55e289} /* (6, 15, 6) {real, imag} */,
  {32'h3d9e390f, 32'h3df664c5} /* (6, 15, 5) {real, imag} */,
  {32'hbe175b5d, 32'h3e503e71} /* (6, 15, 4) {real, imag} */,
  {32'hbcd1dd54, 32'h3e26253f} /* (6, 15, 3) {real, imag} */,
  {32'h3f4353c4, 32'h3e0955b8} /* (6, 15, 2) {real, imag} */,
  {32'hc00ce4c5, 32'h3c0b8d30} /* (6, 15, 1) {real, imag} */,
  {32'hbfde820a, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'hbff08f4e, 32'h3d507204} /* (6, 14, 31) {real, imag} */,
  {32'h3f688a4a, 32'hbdf4db34} /* (6, 14, 30) {real, imag} */,
  {32'h3d2c0a00, 32'hbd821ed4} /* (6, 14, 29) {real, imag} */,
  {32'hbe246699, 32'hbe28b4c8} /* (6, 14, 28) {real, imag} */,
  {32'h3e2a79cb, 32'h3d73208f} /* (6, 14, 27) {real, imag} */,
  {32'h3d5e6644, 32'hbd9bbb0a} /* (6, 14, 26) {real, imag} */,
  {32'hbcd95bf6, 32'hbd89642b} /* (6, 14, 25) {real, imag} */,
  {32'h3e393d59, 32'hbb0120d8} /* (6, 14, 24) {real, imag} */,
  {32'h3cf1abaa, 32'h3c93cc44} /* (6, 14, 23) {real, imag} */,
  {32'hbdc3bbcc, 32'h3da9eb26} /* (6, 14, 22) {real, imag} */,
  {32'h3d099933, 32'hbcf0e01a} /* (6, 14, 21) {real, imag} */,
  {32'h3dd0accc, 32'h3dbf06e4} /* (6, 14, 20) {real, imag} */,
  {32'hbd17d167, 32'h3c911622} /* (6, 14, 19) {real, imag} */,
  {32'hbc02c754, 32'hbda4b28e} /* (6, 14, 18) {real, imag} */,
  {32'hbd7c9aa6, 32'h3d936a40} /* (6, 14, 17) {real, imag} */,
  {32'hbb518250, 32'h00000000} /* (6, 14, 16) {real, imag} */,
  {32'hbd7c9aa6, 32'hbd936a40} /* (6, 14, 15) {real, imag} */,
  {32'hbc02c754, 32'h3da4b28e} /* (6, 14, 14) {real, imag} */,
  {32'hbd17d167, 32'hbc911622} /* (6, 14, 13) {real, imag} */,
  {32'h3dd0accc, 32'hbdbf06e4} /* (6, 14, 12) {real, imag} */,
  {32'h3d099933, 32'h3cf0e01a} /* (6, 14, 11) {real, imag} */,
  {32'hbdc3bbcc, 32'hbda9eb26} /* (6, 14, 10) {real, imag} */,
  {32'h3cf1abaa, 32'hbc93cc44} /* (6, 14, 9) {real, imag} */,
  {32'h3e393d59, 32'h3b0120d8} /* (6, 14, 8) {real, imag} */,
  {32'hbcd95bf6, 32'h3d89642b} /* (6, 14, 7) {real, imag} */,
  {32'h3d5e6644, 32'h3d9bbb0a} /* (6, 14, 6) {real, imag} */,
  {32'h3e2a79cb, 32'hbd73208f} /* (6, 14, 5) {real, imag} */,
  {32'hbe246699, 32'h3e28b4c8} /* (6, 14, 4) {real, imag} */,
  {32'h3d2c0a00, 32'h3d821ed4} /* (6, 14, 3) {real, imag} */,
  {32'h3f688a4a, 32'h3df4db34} /* (6, 14, 2) {real, imag} */,
  {32'hbff08f4e, 32'hbd507204} /* (6, 14, 1) {real, imag} */,
  {32'hbfe249ce, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hbfc8675b, 32'hbd26efc0} /* (6, 13, 31) {real, imag} */,
  {32'h3f6f3c68, 32'hbe0a5315} /* (6, 13, 30) {real, imag} */,
  {32'h3d9856bc, 32'h3d0e127c} /* (6, 13, 29) {real, imag} */,
  {32'hbe1521c8, 32'hbda691c4} /* (6, 13, 28) {real, imag} */,
  {32'h3e7711e0, 32'h3c261e4a} /* (6, 13, 27) {real, imag} */,
  {32'h3dfd9317, 32'h3d75c632} /* (6, 13, 26) {real, imag} */,
  {32'hbd0d53f8, 32'hbd7bda43} /* (6, 13, 25) {real, imag} */,
  {32'h3e0bfe43, 32'h3c5d6f2a} /* (6, 13, 24) {real, imag} */,
  {32'hbd2a9a0b, 32'h3e3f31ee} /* (6, 13, 23) {real, imag} */,
  {32'hbdb55da4, 32'h3dab16c1} /* (6, 13, 22) {real, imag} */,
  {32'h3cca123a, 32'hbe545cf4} /* (6, 13, 21) {real, imag} */,
  {32'h3cafb1bc, 32'hbdc2cda5} /* (6, 13, 20) {real, imag} */,
  {32'h3cc499b5, 32'h3e398ed2} /* (6, 13, 19) {real, imag} */,
  {32'hbd6cd3bf, 32'hbde4cf30} /* (6, 13, 18) {real, imag} */,
  {32'h3d83537c, 32'hbc04c20a} /* (6, 13, 17) {real, imag} */,
  {32'h3c74be8e, 32'h00000000} /* (6, 13, 16) {real, imag} */,
  {32'h3d83537c, 32'h3c04c20a} /* (6, 13, 15) {real, imag} */,
  {32'hbd6cd3bf, 32'h3de4cf30} /* (6, 13, 14) {real, imag} */,
  {32'h3cc499b5, 32'hbe398ed2} /* (6, 13, 13) {real, imag} */,
  {32'h3cafb1bc, 32'h3dc2cda5} /* (6, 13, 12) {real, imag} */,
  {32'h3cca123a, 32'h3e545cf4} /* (6, 13, 11) {real, imag} */,
  {32'hbdb55da4, 32'hbdab16c1} /* (6, 13, 10) {real, imag} */,
  {32'hbd2a9a0b, 32'hbe3f31ee} /* (6, 13, 9) {real, imag} */,
  {32'h3e0bfe43, 32'hbc5d6f2a} /* (6, 13, 8) {real, imag} */,
  {32'hbd0d53f8, 32'h3d7bda43} /* (6, 13, 7) {real, imag} */,
  {32'h3dfd9317, 32'hbd75c632} /* (6, 13, 6) {real, imag} */,
  {32'h3e7711e0, 32'hbc261e4a} /* (6, 13, 5) {real, imag} */,
  {32'hbe1521c8, 32'h3da691c4} /* (6, 13, 4) {real, imag} */,
  {32'h3d9856bc, 32'hbd0e127c} /* (6, 13, 3) {real, imag} */,
  {32'h3f6f3c68, 32'h3e0a5315} /* (6, 13, 2) {real, imag} */,
  {32'hbfc8675b, 32'h3d26efc0} /* (6, 13, 1) {real, imag} */,
  {32'hbfcdbb32, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'hbf968af1, 32'hbc4f7500} /* (6, 12, 31) {real, imag} */,
  {32'h3f3475ac, 32'hbe49c0fb} /* (6, 12, 30) {real, imag} */,
  {32'h3e06abee, 32'h3d74799c} /* (6, 12, 29) {real, imag} */,
  {32'hbe45d97a, 32'hbd3df7a4} /* (6, 12, 28) {real, imag} */,
  {32'h3dcb6f61, 32'hbd0627f9} /* (6, 12, 27) {real, imag} */,
  {32'h3d65e1b9, 32'h3e040f20} /* (6, 12, 26) {real, imag} */,
  {32'hbc97494a, 32'hbdaba2b3} /* (6, 12, 25) {real, imag} */,
  {32'h3def2b0b, 32'h3c517aae} /* (6, 12, 24) {real, imag} */,
  {32'hbd3176d3, 32'hbb6f8850} /* (6, 12, 23) {real, imag} */,
  {32'h3e02c4bc, 32'hbd528eaa} /* (6, 12, 22) {real, imag} */,
  {32'hbb534d58, 32'h3c21cb5a} /* (6, 12, 21) {real, imag} */,
  {32'hbdf9d8d6, 32'h3d6f79fb} /* (6, 12, 20) {real, imag} */,
  {32'h3dea3873, 32'hbddc1df2} /* (6, 12, 19) {real, imag} */,
  {32'h3aec5570, 32'h3d07953f} /* (6, 12, 18) {real, imag} */,
  {32'hbd6432eb, 32'h3d05383c} /* (6, 12, 17) {real, imag} */,
  {32'h3c81bf6a, 32'h00000000} /* (6, 12, 16) {real, imag} */,
  {32'hbd6432eb, 32'hbd05383c} /* (6, 12, 15) {real, imag} */,
  {32'h3aec5570, 32'hbd07953f} /* (6, 12, 14) {real, imag} */,
  {32'h3dea3873, 32'h3ddc1df2} /* (6, 12, 13) {real, imag} */,
  {32'hbdf9d8d6, 32'hbd6f79fb} /* (6, 12, 12) {real, imag} */,
  {32'hbb534d58, 32'hbc21cb5a} /* (6, 12, 11) {real, imag} */,
  {32'h3e02c4bc, 32'h3d528eaa} /* (6, 12, 10) {real, imag} */,
  {32'hbd3176d3, 32'h3b6f8850} /* (6, 12, 9) {real, imag} */,
  {32'h3def2b0b, 32'hbc517aae} /* (6, 12, 8) {real, imag} */,
  {32'hbc97494a, 32'h3daba2b3} /* (6, 12, 7) {real, imag} */,
  {32'h3d65e1b9, 32'hbe040f20} /* (6, 12, 6) {real, imag} */,
  {32'h3dcb6f61, 32'h3d0627f9} /* (6, 12, 5) {real, imag} */,
  {32'hbe45d97a, 32'h3d3df7a4} /* (6, 12, 4) {real, imag} */,
  {32'h3e06abee, 32'hbd74799c} /* (6, 12, 3) {real, imag} */,
  {32'h3f3475ac, 32'h3e49c0fb} /* (6, 12, 2) {real, imag} */,
  {32'hbf968af1, 32'h3c4f7500} /* (6, 12, 1) {real, imag} */,
  {32'hbf7a979c, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'hbf2142a8, 32'hbe856d56} /* (6, 11, 31) {real, imag} */,
  {32'h3efe04e8, 32'hbdf136e6} /* (6, 11, 30) {real, imag} */,
  {32'h3e52fe07, 32'h3d94812a} /* (6, 11, 29) {real, imag} */,
  {32'hbb75f668, 32'hbdc18172} /* (6, 11, 28) {real, imag} */,
  {32'h3d8cfd52, 32'hbd8f642b} /* (6, 11, 27) {real, imag} */,
  {32'hbc3068c9, 32'h3d49444e} /* (6, 11, 26) {real, imag} */,
  {32'hbd38edff, 32'hbdbb209e} /* (6, 11, 25) {real, imag} */,
  {32'h3a143080, 32'hbdb240ad} /* (6, 11, 24) {real, imag} */,
  {32'h3cfa6ebc, 32'hbdd4efb7} /* (6, 11, 23) {real, imag} */,
  {32'h3ce96ca6, 32'h3d95bae9} /* (6, 11, 22) {real, imag} */,
  {32'h3b1fb980, 32'hbcfa1210} /* (6, 11, 21) {real, imag} */,
  {32'h3cd9839a, 32'h3d69e704} /* (6, 11, 20) {real, imag} */,
  {32'h3c9f0af5, 32'h3d5dd9fa} /* (6, 11, 19) {real, imag} */,
  {32'h3c3a9dcc, 32'h3d3e08de} /* (6, 11, 18) {real, imag} */,
  {32'hbc66c203, 32'h3d245f7a} /* (6, 11, 17) {real, imag} */,
  {32'h3cdfeaa7, 32'h00000000} /* (6, 11, 16) {real, imag} */,
  {32'hbc66c203, 32'hbd245f7a} /* (6, 11, 15) {real, imag} */,
  {32'h3c3a9dcc, 32'hbd3e08de} /* (6, 11, 14) {real, imag} */,
  {32'h3c9f0af5, 32'hbd5dd9fa} /* (6, 11, 13) {real, imag} */,
  {32'h3cd9839a, 32'hbd69e704} /* (6, 11, 12) {real, imag} */,
  {32'h3b1fb980, 32'h3cfa1210} /* (6, 11, 11) {real, imag} */,
  {32'h3ce96ca6, 32'hbd95bae9} /* (6, 11, 10) {real, imag} */,
  {32'h3cfa6ebc, 32'h3dd4efb7} /* (6, 11, 9) {real, imag} */,
  {32'h3a143080, 32'h3db240ad} /* (6, 11, 8) {real, imag} */,
  {32'hbd38edff, 32'h3dbb209e} /* (6, 11, 7) {real, imag} */,
  {32'hbc3068c9, 32'hbd49444e} /* (6, 11, 6) {real, imag} */,
  {32'h3d8cfd52, 32'h3d8f642b} /* (6, 11, 5) {real, imag} */,
  {32'hbb75f668, 32'h3dc18172} /* (6, 11, 4) {real, imag} */,
  {32'h3e52fe07, 32'hbd94812a} /* (6, 11, 3) {real, imag} */,
  {32'h3efe04e8, 32'h3df136e6} /* (6, 11, 2) {real, imag} */,
  {32'hbf2142a8, 32'h3e856d56} /* (6, 11, 1) {real, imag} */,
  {32'hbf039db1, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h3eecafc6, 32'hbf04e303} /* (6, 10, 31) {real, imag} */,
  {32'hbdda882c, 32'h3d2ee31c} /* (6, 10, 30) {real, imag} */,
  {32'h3d892cb4, 32'h3d7d150a} /* (6, 10, 29) {real, imag} */,
  {32'h3da1f2fd, 32'hbe530961} /* (6, 10, 28) {real, imag} */,
  {32'hbcbbc521, 32'h3d9f5f95} /* (6, 10, 27) {real, imag} */,
  {32'h3cea6280, 32'h3d5cfc03} /* (6, 10, 26) {real, imag} */,
  {32'h3daf1b68, 32'h3c699bc2} /* (6, 10, 25) {real, imag} */,
  {32'h3d29edb7, 32'h3d24974e} /* (6, 10, 24) {real, imag} */,
  {32'h3dd7dcff, 32'hbd20a17e} /* (6, 10, 23) {real, imag} */,
  {32'hbd202838, 32'hbd3a26aa} /* (6, 10, 22) {real, imag} */,
  {32'hbc611298, 32'h3dd2a1f0} /* (6, 10, 21) {real, imag} */,
  {32'hbd7491bc, 32'h3c932658} /* (6, 10, 20) {real, imag} */,
  {32'hbc8c005b, 32'h3d0f45d3} /* (6, 10, 19) {real, imag} */,
  {32'h3d7cea6e, 32'hbd0d1aca} /* (6, 10, 18) {real, imag} */,
  {32'hbc8d68e7, 32'h3d66de1a} /* (6, 10, 17) {real, imag} */,
  {32'h3b428718, 32'h00000000} /* (6, 10, 16) {real, imag} */,
  {32'hbc8d68e7, 32'hbd66de1a} /* (6, 10, 15) {real, imag} */,
  {32'h3d7cea6e, 32'h3d0d1aca} /* (6, 10, 14) {real, imag} */,
  {32'hbc8c005b, 32'hbd0f45d3} /* (6, 10, 13) {real, imag} */,
  {32'hbd7491bc, 32'hbc932658} /* (6, 10, 12) {real, imag} */,
  {32'hbc611298, 32'hbdd2a1f0} /* (6, 10, 11) {real, imag} */,
  {32'hbd202838, 32'h3d3a26aa} /* (6, 10, 10) {real, imag} */,
  {32'h3dd7dcff, 32'h3d20a17e} /* (6, 10, 9) {real, imag} */,
  {32'h3d29edb7, 32'hbd24974e} /* (6, 10, 8) {real, imag} */,
  {32'h3daf1b68, 32'hbc699bc2} /* (6, 10, 7) {real, imag} */,
  {32'h3cea6280, 32'hbd5cfc03} /* (6, 10, 6) {real, imag} */,
  {32'hbcbbc521, 32'hbd9f5f95} /* (6, 10, 5) {real, imag} */,
  {32'h3da1f2fd, 32'h3e530961} /* (6, 10, 4) {real, imag} */,
  {32'h3d892cb4, 32'hbd7d150a} /* (6, 10, 3) {real, imag} */,
  {32'hbdda882c, 32'hbd2ee31c} /* (6, 10, 2) {real, imag} */,
  {32'h3eecafc6, 32'h3f04e303} /* (6, 10, 1) {real, imag} */,
  {32'h3f2b821b, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'h3f9527e9, 32'hbf37bd18} /* (6, 9, 31) {real, imag} */,
  {32'hbee1d09e, 32'h3e56fdd7} /* (6, 9, 30) {real, imag} */,
  {32'h3db389de, 32'h3d887795} /* (6, 9, 29) {real, imag} */,
  {32'h3deb2a1e, 32'hbe81aee9} /* (6, 9, 28) {real, imag} */,
  {32'hbdae70ed, 32'h3e3ce4bf} /* (6, 9, 27) {real, imag} */,
  {32'hbd921251, 32'h3df53e09} /* (6, 9, 26) {real, imag} */,
  {32'h392b4340, 32'hbe4100b6} /* (6, 9, 25) {real, imag} */,
  {32'hbe12707e, 32'hbdd2ca78} /* (6, 9, 24) {real, imag} */,
  {32'hbc786496, 32'h3de1cece} /* (6, 9, 23) {real, imag} */,
  {32'hbd156adb, 32'hbd1b1cce} /* (6, 9, 22) {real, imag} */,
  {32'hbdb2477e, 32'h3e3099b7} /* (6, 9, 21) {real, imag} */,
  {32'h3ce810d3, 32'hbd87e9fc} /* (6, 9, 20) {real, imag} */,
  {32'h3d59e21c, 32'hbbbce324} /* (6, 9, 19) {real, imag} */,
  {32'h3dd1532a, 32'h3cd9d924} /* (6, 9, 18) {real, imag} */,
  {32'hbc5bbc24, 32'hbd9649e8} /* (6, 9, 17) {real, imag} */,
  {32'hbd9a0d0e, 32'h00000000} /* (6, 9, 16) {real, imag} */,
  {32'hbc5bbc24, 32'h3d9649e8} /* (6, 9, 15) {real, imag} */,
  {32'h3dd1532a, 32'hbcd9d924} /* (6, 9, 14) {real, imag} */,
  {32'h3d59e21c, 32'h3bbce324} /* (6, 9, 13) {real, imag} */,
  {32'h3ce810d3, 32'h3d87e9fc} /* (6, 9, 12) {real, imag} */,
  {32'hbdb2477e, 32'hbe3099b7} /* (6, 9, 11) {real, imag} */,
  {32'hbd156adb, 32'h3d1b1cce} /* (6, 9, 10) {real, imag} */,
  {32'hbc786496, 32'hbde1cece} /* (6, 9, 9) {real, imag} */,
  {32'hbe12707e, 32'h3dd2ca78} /* (6, 9, 8) {real, imag} */,
  {32'h392b4340, 32'h3e4100b6} /* (6, 9, 7) {real, imag} */,
  {32'hbd921251, 32'hbdf53e09} /* (6, 9, 6) {real, imag} */,
  {32'hbdae70ed, 32'hbe3ce4bf} /* (6, 9, 5) {real, imag} */,
  {32'h3deb2a1e, 32'h3e81aee9} /* (6, 9, 4) {real, imag} */,
  {32'h3db389de, 32'hbd887795} /* (6, 9, 3) {real, imag} */,
  {32'hbee1d09e, 32'hbe56fdd7} /* (6, 9, 2) {real, imag} */,
  {32'h3f9527e9, 32'h3f37bd18} /* (6, 9, 1) {real, imag} */,
  {32'h3fc6cd63, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'h3fc105c7, 32'hbf3d0352} /* (6, 8, 31) {real, imag} */,
  {32'hbeda60a2, 32'h3ecaf21a} /* (6, 8, 30) {real, imag} */,
  {32'h3e5776f1, 32'hbcbbe80c} /* (6, 8, 29) {real, imag} */,
  {32'h3dbb21a4, 32'hbdeb378a} /* (6, 8, 28) {real, imag} */,
  {32'hbdf0757c, 32'h3da3eb70} /* (6, 8, 27) {real, imag} */,
  {32'hbda3e665, 32'h3daf30b7} /* (6, 8, 26) {real, imag} */,
  {32'hbd554abc, 32'hbde7d9fc} /* (6, 8, 25) {real, imag} */,
  {32'hbdf6aa9b, 32'hbdc0fc9f} /* (6, 8, 24) {real, imag} */,
  {32'h3d083394, 32'h3d82430d} /* (6, 8, 23) {real, imag} */,
  {32'h3ca93342, 32'h3d3c5360} /* (6, 8, 22) {real, imag} */,
  {32'h3d898094, 32'h3dde8655} /* (6, 8, 21) {real, imag} */,
  {32'h3ce3a085, 32'h3c7ff398} /* (6, 8, 20) {real, imag} */,
  {32'h3d923970, 32'h3d255148} /* (6, 8, 19) {real, imag} */,
  {32'hbcbef1f9, 32'h3d43ea45} /* (6, 8, 18) {real, imag} */,
  {32'h3d06fb22, 32'hbc808e35} /* (6, 8, 17) {real, imag} */,
  {32'h3d39fbad, 32'h00000000} /* (6, 8, 16) {real, imag} */,
  {32'h3d06fb22, 32'h3c808e35} /* (6, 8, 15) {real, imag} */,
  {32'hbcbef1f9, 32'hbd43ea45} /* (6, 8, 14) {real, imag} */,
  {32'h3d923970, 32'hbd255148} /* (6, 8, 13) {real, imag} */,
  {32'h3ce3a085, 32'hbc7ff398} /* (6, 8, 12) {real, imag} */,
  {32'h3d898094, 32'hbdde8655} /* (6, 8, 11) {real, imag} */,
  {32'h3ca93342, 32'hbd3c5360} /* (6, 8, 10) {real, imag} */,
  {32'h3d083394, 32'hbd82430d} /* (6, 8, 9) {real, imag} */,
  {32'hbdf6aa9b, 32'h3dc0fc9f} /* (6, 8, 8) {real, imag} */,
  {32'hbd554abc, 32'h3de7d9fc} /* (6, 8, 7) {real, imag} */,
  {32'hbda3e665, 32'hbdaf30b7} /* (6, 8, 6) {real, imag} */,
  {32'hbdf0757c, 32'hbda3eb70} /* (6, 8, 5) {real, imag} */,
  {32'h3dbb21a4, 32'h3deb378a} /* (6, 8, 4) {real, imag} */,
  {32'h3e5776f1, 32'h3cbbe80c} /* (6, 8, 3) {real, imag} */,
  {32'hbeda60a2, 32'hbecaf21a} /* (6, 8, 2) {real, imag} */,
  {32'h3fc105c7, 32'h3f3d0352} /* (6, 8, 1) {real, imag} */,
  {32'h3ff67237, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h3fe54f2f, 32'hbf703c84} /* (6, 7, 31) {real, imag} */,
  {32'hbefea696, 32'h3f1cd6e2} /* (6, 7, 30) {real, imag} */,
  {32'h3e7f176f, 32'hbcc21012} /* (6, 7, 29) {real, imag} */,
  {32'h3d991d3b, 32'h3b349330} /* (6, 7, 28) {real, imag} */,
  {32'hbe2a16d9, 32'h3bd767c0} /* (6, 7, 27) {real, imag} */,
  {32'h3c71361e, 32'h3838d800} /* (6, 7, 26) {real, imag} */,
  {32'h3c2ac34b, 32'hbda865e8} /* (6, 7, 25) {real, imag} */,
  {32'hbd966855, 32'hbc7f2b20} /* (6, 7, 24) {real, imag} */,
  {32'hbcac54c3, 32'h3c21c190} /* (6, 7, 23) {real, imag} */,
  {32'hbdbf9f5e, 32'hbd729fcd} /* (6, 7, 22) {real, imag} */,
  {32'h3cbee6ec, 32'hbd814ed8} /* (6, 7, 21) {real, imag} */,
  {32'h3ce6aff3, 32'hba8e9460} /* (6, 7, 20) {real, imag} */,
  {32'hbd25ea1a, 32'hbc56ff82} /* (6, 7, 19) {real, imag} */,
  {32'hbcbc00a2, 32'h3cd05e46} /* (6, 7, 18) {real, imag} */,
  {32'h3c10c540, 32'hbc24ef00} /* (6, 7, 17) {real, imag} */,
  {32'h3d8b8ef9, 32'h00000000} /* (6, 7, 16) {real, imag} */,
  {32'h3c10c540, 32'h3c24ef00} /* (6, 7, 15) {real, imag} */,
  {32'hbcbc00a2, 32'hbcd05e46} /* (6, 7, 14) {real, imag} */,
  {32'hbd25ea1a, 32'h3c56ff82} /* (6, 7, 13) {real, imag} */,
  {32'h3ce6aff3, 32'h3a8e9460} /* (6, 7, 12) {real, imag} */,
  {32'h3cbee6ec, 32'h3d814ed8} /* (6, 7, 11) {real, imag} */,
  {32'hbdbf9f5e, 32'h3d729fcd} /* (6, 7, 10) {real, imag} */,
  {32'hbcac54c3, 32'hbc21c190} /* (6, 7, 9) {real, imag} */,
  {32'hbd966855, 32'h3c7f2b20} /* (6, 7, 8) {real, imag} */,
  {32'h3c2ac34b, 32'h3da865e8} /* (6, 7, 7) {real, imag} */,
  {32'h3c71361e, 32'hb838d800} /* (6, 7, 6) {real, imag} */,
  {32'hbe2a16d9, 32'hbbd767c0} /* (6, 7, 5) {real, imag} */,
  {32'h3d991d3b, 32'hbb349330} /* (6, 7, 4) {real, imag} */,
  {32'h3e7f176f, 32'h3cc21012} /* (6, 7, 3) {real, imag} */,
  {32'hbefea696, 32'hbf1cd6e2} /* (6, 7, 2) {real, imag} */,
  {32'h3fe54f2f, 32'h3f703c84} /* (6, 7, 1) {real, imag} */,
  {32'h40101a8c, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'h3ffd7eb4, 32'hbf71fe21} /* (6, 6, 31) {real, imag} */,
  {32'hbf04cbee, 32'h3f13635f} /* (6, 6, 30) {real, imag} */,
  {32'h3c87cf68, 32'h3940e800} /* (6, 6, 29) {real, imag} */,
  {32'h3d8c4ba1, 32'hbde171dc} /* (6, 6, 28) {real, imag} */,
  {32'hbe1010e7, 32'hbbf3d2d0} /* (6, 6, 27) {real, imag} */,
  {32'h3d9bf713, 32'hbcfea8a0} /* (6, 6, 26) {real, imag} */,
  {32'h3de6dbdd, 32'h3c82f078} /* (6, 6, 25) {real, imag} */,
  {32'hbdcb7bf4, 32'h3ddd2715} /* (6, 6, 24) {real, imag} */,
  {32'hbd5ed971, 32'h3cdf948b} /* (6, 6, 23) {real, imag} */,
  {32'hbd14b806, 32'h3d9b7b1d} /* (6, 6, 22) {real, imag} */,
  {32'hbdc9930c, 32'h3d2c1ebe} /* (6, 6, 21) {real, imag} */,
  {32'h3e0c35c6, 32'hbd2ad735} /* (6, 6, 20) {real, imag} */,
  {32'h3b6dfad8, 32'hbd50ef7f} /* (6, 6, 19) {real, imag} */,
  {32'hbceb4646, 32'hbc47a23e} /* (6, 6, 18) {real, imag} */,
  {32'h3cafbc5d, 32'hbd052e74} /* (6, 6, 17) {real, imag} */,
  {32'hbbd5005e, 32'h00000000} /* (6, 6, 16) {real, imag} */,
  {32'h3cafbc5d, 32'h3d052e74} /* (6, 6, 15) {real, imag} */,
  {32'hbceb4646, 32'h3c47a23e} /* (6, 6, 14) {real, imag} */,
  {32'h3b6dfad8, 32'h3d50ef7f} /* (6, 6, 13) {real, imag} */,
  {32'h3e0c35c6, 32'h3d2ad735} /* (6, 6, 12) {real, imag} */,
  {32'hbdc9930c, 32'hbd2c1ebe} /* (6, 6, 11) {real, imag} */,
  {32'hbd14b806, 32'hbd9b7b1d} /* (6, 6, 10) {real, imag} */,
  {32'hbd5ed971, 32'hbcdf948b} /* (6, 6, 9) {real, imag} */,
  {32'hbdcb7bf4, 32'hbddd2715} /* (6, 6, 8) {real, imag} */,
  {32'h3de6dbdd, 32'hbc82f078} /* (6, 6, 7) {real, imag} */,
  {32'h3d9bf713, 32'h3cfea8a0} /* (6, 6, 6) {real, imag} */,
  {32'hbe1010e7, 32'h3bf3d2d0} /* (6, 6, 5) {real, imag} */,
  {32'h3d8c4ba1, 32'h3de171dc} /* (6, 6, 4) {real, imag} */,
  {32'h3c87cf68, 32'hb940e800} /* (6, 6, 3) {real, imag} */,
  {32'hbf04cbee, 32'hbf13635f} /* (6, 6, 2) {real, imag} */,
  {32'h3ffd7eb4, 32'h3f71fe21} /* (6, 6, 1) {real, imag} */,
  {32'h4033946c, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'h3fefa338, 32'hbfc32180} /* (6, 5, 31) {real, imag} */,
  {32'hbe1cc9c4, 32'h3f20e3ca} /* (6, 5, 30) {real, imag} */,
  {32'h3ce28a5c, 32'h3d6a9ae3} /* (6, 5, 29) {real, imag} */,
  {32'h3ccab508, 32'h3b95f160} /* (6, 5, 28) {real, imag} */,
  {32'hbdec9173, 32'hbdb9705b} /* (6, 5, 27) {real, imag} */,
  {32'h3d5e7127, 32'hbbbc862c} /* (6, 5, 26) {real, imag} */,
  {32'h3d869de8, 32'hbd9d56c4} /* (6, 5, 25) {real, imag} */,
  {32'hbb9ddfb8, 32'hbc7d5c52} /* (6, 5, 24) {real, imag} */,
  {32'hbdd084f6, 32'hbdf1d38e} /* (6, 5, 23) {real, imag} */,
  {32'h3e131105, 32'hbd2bd33b} /* (6, 5, 22) {real, imag} */,
  {32'hbdb7f392, 32'h3d859a0b} /* (6, 5, 21) {real, imag} */,
  {32'hbddb8334, 32'hbc62fde9} /* (6, 5, 20) {real, imag} */,
  {32'hbd1a8f7a, 32'hbd11d19c} /* (6, 5, 19) {real, imag} */,
  {32'hbba62b98, 32'h3ccadac8} /* (6, 5, 18) {real, imag} */,
  {32'hbcb1462b, 32'hbd472edc} /* (6, 5, 17) {real, imag} */,
  {32'hbd2daaf6, 32'h00000000} /* (6, 5, 16) {real, imag} */,
  {32'hbcb1462b, 32'h3d472edc} /* (6, 5, 15) {real, imag} */,
  {32'hbba62b98, 32'hbccadac8} /* (6, 5, 14) {real, imag} */,
  {32'hbd1a8f7a, 32'h3d11d19c} /* (6, 5, 13) {real, imag} */,
  {32'hbddb8334, 32'h3c62fde9} /* (6, 5, 12) {real, imag} */,
  {32'hbdb7f392, 32'hbd859a0b} /* (6, 5, 11) {real, imag} */,
  {32'h3e131105, 32'h3d2bd33b} /* (6, 5, 10) {real, imag} */,
  {32'hbdd084f6, 32'h3df1d38e} /* (6, 5, 9) {real, imag} */,
  {32'hbb9ddfb8, 32'h3c7d5c52} /* (6, 5, 8) {real, imag} */,
  {32'h3d869de8, 32'h3d9d56c4} /* (6, 5, 7) {real, imag} */,
  {32'h3d5e7127, 32'h3bbc862c} /* (6, 5, 6) {real, imag} */,
  {32'hbdec9173, 32'h3db9705b} /* (6, 5, 5) {real, imag} */,
  {32'h3ccab508, 32'hbb95f160} /* (6, 5, 4) {real, imag} */,
  {32'h3ce28a5c, 32'hbd6a9ae3} /* (6, 5, 3) {real, imag} */,
  {32'hbe1cc9c4, 32'hbf20e3ca} /* (6, 5, 2) {real, imag} */,
  {32'h3fefa338, 32'h3fc32180} /* (6, 5, 1) {real, imag} */,
  {32'h403960f3, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'h3fe797b9, 32'hbfef8c0e} /* (6, 4, 31) {real, imag} */,
  {32'h3e11671c, 32'h3f47635e} /* (6, 4, 30) {real, imag} */,
  {32'h3e15e27c, 32'h3cbe36eb} /* (6, 4, 29) {real, imag} */,
  {32'hbd91d121, 32'h3ea4d910} /* (6, 4, 28) {real, imag} */,
  {32'hbd44f00c, 32'hbde5122e} /* (6, 4, 27) {real, imag} */,
  {32'h3d89ca14, 32'h3d508fce} /* (6, 4, 26) {real, imag} */,
  {32'h3dd563ca, 32'hbde4eccc} /* (6, 4, 25) {real, imag} */,
  {32'h3d81a9bb, 32'h3de454c2} /* (6, 4, 24) {real, imag} */,
  {32'hbd5feae2, 32'hbcfe2db0} /* (6, 4, 23) {real, imag} */,
  {32'h3da7be20, 32'h3ddc00df} /* (6, 4, 22) {real, imag} */,
  {32'hbd6fa3da, 32'h3b548800} /* (6, 4, 21) {real, imag} */,
  {32'hbd271fc8, 32'h3ca57453} /* (6, 4, 20) {real, imag} */,
  {32'hbdd64344, 32'h3d53c715} /* (6, 4, 19) {real, imag} */,
  {32'hbc856f68, 32'hbd55b45e} /* (6, 4, 18) {real, imag} */,
  {32'hbda20b00, 32'h3dd76f4d} /* (6, 4, 17) {real, imag} */,
  {32'h3c6411e2, 32'h00000000} /* (6, 4, 16) {real, imag} */,
  {32'hbda20b00, 32'hbdd76f4d} /* (6, 4, 15) {real, imag} */,
  {32'hbc856f68, 32'h3d55b45e} /* (6, 4, 14) {real, imag} */,
  {32'hbdd64344, 32'hbd53c715} /* (6, 4, 13) {real, imag} */,
  {32'hbd271fc8, 32'hbca57453} /* (6, 4, 12) {real, imag} */,
  {32'hbd6fa3da, 32'hbb548800} /* (6, 4, 11) {real, imag} */,
  {32'h3da7be20, 32'hbddc00df} /* (6, 4, 10) {real, imag} */,
  {32'hbd5feae2, 32'h3cfe2db0} /* (6, 4, 9) {real, imag} */,
  {32'h3d81a9bb, 32'hbde454c2} /* (6, 4, 8) {real, imag} */,
  {32'h3dd563ca, 32'h3de4eccc} /* (6, 4, 7) {real, imag} */,
  {32'h3d89ca14, 32'hbd508fce} /* (6, 4, 6) {real, imag} */,
  {32'hbd44f00c, 32'h3de5122e} /* (6, 4, 5) {real, imag} */,
  {32'hbd91d121, 32'hbea4d910} /* (6, 4, 4) {real, imag} */,
  {32'h3e15e27c, 32'hbcbe36eb} /* (6, 4, 3) {real, imag} */,
  {32'h3e11671c, 32'hbf47635e} /* (6, 4, 2) {real, imag} */,
  {32'h3fe797b9, 32'h3fef8c0e} /* (6, 4, 1) {real, imag} */,
  {32'h403ada56, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'h3fda23ce, 32'hc0027e74} /* (6, 3, 31) {real, imag} */,
  {32'h3e3cf5da, 32'h3f19ee10} /* (6, 3, 30) {real, imag} */,
  {32'h3cf2a142, 32'h3d174284} /* (6, 3, 29) {real, imag} */,
  {32'h3ce1c178, 32'h3e4ded56} /* (6, 3, 28) {real, imag} */,
  {32'hbd9c32e5, 32'hbdc17e00} /* (6, 3, 27) {real, imag} */,
  {32'h3bb885c8, 32'h3c99489b} /* (6, 3, 26) {real, imag} */,
  {32'h3cf1f503, 32'hbd32c329} /* (6, 3, 25) {real, imag} */,
  {32'h3dde13dd, 32'h3cc80881} /* (6, 3, 24) {real, imag} */,
  {32'h3d97fc97, 32'hbb9ccb08} /* (6, 3, 23) {real, imag} */,
  {32'h3c932661, 32'h3cc6eda1} /* (6, 3, 22) {real, imag} */,
  {32'hbdfc0188, 32'h3dd42c55} /* (6, 3, 21) {real, imag} */,
  {32'h3b84cf26, 32'hbbe3e79c} /* (6, 3, 20) {real, imag} */,
  {32'h3d35b681, 32'h3da6d838} /* (6, 3, 19) {real, imag} */,
  {32'hbd46e581, 32'h3b811630} /* (6, 3, 18) {real, imag} */,
  {32'h3ceab584, 32'h3d01b1ce} /* (6, 3, 17) {real, imag} */,
  {32'hbc7b62d6, 32'h00000000} /* (6, 3, 16) {real, imag} */,
  {32'h3ceab584, 32'hbd01b1ce} /* (6, 3, 15) {real, imag} */,
  {32'hbd46e581, 32'hbb811630} /* (6, 3, 14) {real, imag} */,
  {32'h3d35b681, 32'hbda6d838} /* (6, 3, 13) {real, imag} */,
  {32'h3b84cf26, 32'h3be3e79c} /* (6, 3, 12) {real, imag} */,
  {32'hbdfc0188, 32'hbdd42c55} /* (6, 3, 11) {real, imag} */,
  {32'h3c932661, 32'hbcc6eda1} /* (6, 3, 10) {real, imag} */,
  {32'h3d97fc97, 32'h3b9ccb08} /* (6, 3, 9) {real, imag} */,
  {32'h3dde13dd, 32'hbcc80881} /* (6, 3, 8) {real, imag} */,
  {32'h3cf1f503, 32'h3d32c329} /* (6, 3, 7) {real, imag} */,
  {32'h3bb885c8, 32'hbc99489b} /* (6, 3, 6) {real, imag} */,
  {32'hbd9c32e5, 32'h3dc17e00} /* (6, 3, 5) {real, imag} */,
  {32'h3ce1c178, 32'hbe4ded56} /* (6, 3, 4) {real, imag} */,
  {32'h3cf2a142, 32'hbd174284} /* (6, 3, 3) {real, imag} */,
  {32'h3e3cf5da, 32'hbf19ee10} /* (6, 3, 2) {real, imag} */,
  {32'h3fda23ce, 32'h40027e74} /* (6, 3, 1) {real, imag} */,
  {32'h4049922c, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'h3fc70934, 32'hc003bb85} /* (6, 2, 31) {real, imag} */,
  {32'h3e5abc1c, 32'h3f127cd2} /* (6, 2, 30) {real, imag} */,
  {32'h3d00d836, 32'h3d241df4} /* (6, 2, 29) {real, imag} */,
  {32'h3c9bfb3a, 32'h3dcec554} /* (6, 2, 28) {real, imag} */,
  {32'hbe0dad0c, 32'hbbb83828} /* (6, 2, 27) {real, imag} */,
  {32'h3c0132c3, 32'h3d6af036} /* (6, 2, 26) {real, imag} */,
  {32'hbce08e34, 32'hbd809b41} /* (6, 2, 25) {real, imag} */,
  {32'h3cae1a3b, 32'h3de4649b} /* (6, 2, 24) {real, imag} */,
  {32'hbd3139ed, 32'hbdaaa7c9} /* (6, 2, 23) {real, imag} */,
  {32'hbc1dacfc, 32'hbe045306} /* (6, 2, 22) {real, imag} */,
  {32'hbda0cd47, 32'h3b850930} /* (6, 2, 21) {real, imag} */,
  {32'h3d48e245, 32'h3dfdaf0e} /* (6, 2, 20) {real, imag} */,
  {32'h3de1f2c8, 32'hbc4a33a0} /* (6, 2, 19) {real, imag} */,
  {32'h3d467317, 32'hbd1f62ff} /* (6, 2, 18) {real, imag} */,
  {32'h3d379bfc, 32'h3d9a7532} /* (6, 2, 17) {real, imag} */,
  {32'h3d07ee52, 32'h00000000} /* (6, 2, 16) {real, imag} */,
  {32'h3d379bfc, 32'hbd9a7532} /* (6, 2, 15) {real, imag} */,
  {32'h3d467317, 32'h3d1f62ff} /* (6, 2, 14) {real, imag} */,
  {32'h3de1f2c8, 32'h3c4a33a0} /* (6, 2, 13) {real, imag} */,
  {32'h3d48e245, 32'hbdfdaf0e} /* (6, 2, 12) {real, imag} */,
  {32'hbda0cd47, 32'hbb850930} /* (6, 2, 11) {real, imag} */,
  {32'hbc1dacfc, 32'h3e045306} /* (6, 2, 10) {real, imag} */,
  {32'hbd3139ed, 32'h3daaa7c9} /* (6, 2, 9) {real, imag} */,
  {32'h3cae1a3b, 32'hbde4649b} /* (6, 2, 8) {real, imag} */,
  {32'hbce08e34, 32'h3d809b41} /* (6, 2, 7) {real, imag} */,
  {32'h3c0132c3, 32'hbd6af036} /* (6, 2, 6) {real, imag} */,
  {32'hbe0dad0c, 32'h3bb83828} /* (6, 2, 5) {real, imag} */,
  {32'h3c9bfb3a, 32'hbdcec554} /* (6, 2, 4) {real, imag} */,
  {32'h3d00d836, 32'hbd241df4} /* (6, 2, 3) {real, imag} */,
  {32'h3e5abc1c, 32'hbf127cd2} /* (6, 2, 2) {real, imag} */,
  {32'h3fc70934, 32'h4003bb85} /* (6, 2, 1) {real, imag} */,
  {32'h4066f35f, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'h3fce42cf, 32'hbfe521ce} /* (6, 1, 31) {real, imag} */,
  {32'h3e395200, 32'h3ec38656} /* (6, 1, 30) {real, imag} */,
  {32'hbdd6e5a6, 32'h3d499c56} /* (6, 1, 29) {real, imag} */,
  {32'hbb7b6410, 32'h3d584265} /* (6, 1, 28) {real, imag} */,
  {32'hbdcd6ed6, 32'h3cdbf5bf} /* (6, 1, 27) {real, imag} */,
  {32'hbc07f280, 32'hbbdbc8bc} /* (6, 1, 26) {real, imag} */,
  {32'h3d4d197e, 32'hbd3c86c3} /* (6, 1, 25) {real, imag} */,
  {32'hbc87042b, 32'h3da1e0d1} /* (6, 1, 24) {real, imag} */,
  {32'h3d3b410f, 32'hbd133930} /* (6, 1, 23) {real, imag} */,
  {32'hbd7de8bb, 32'hbb5480e0} /* (6, 1, 22) {real, imag} */,
  {32'h3cbfa981, 32'h3bf3352c} /* (6, 1, 21) {real, imag} */,
  {32'hbc9e6778, 32'h3c8f895d} /* (6, 1, 20) {real, imag} */,
  {32'h3d1a9cb6, 32'h3c92eff2} /* (6, 1, 19) {real, imag} */,
  {32'h3ce9c4bd, 32'h3d1f7032} /* (6, 1, 18) {real, imag} */,
  {32'hbdae9402, 32'h3b47a636} /* (6, 1, 17) {real, imag} */,
  {32'hbcb48955, 32'h00000000} /* (6, 1, 16) {real, imag} */,
  {32'hbdae9402, 32'hbb47a636} /* (6, 1, 15) {real, imag} */,
  {32'h3ce9c4bd, 32'hbd1f7032} /* (6, 1, 14) {real, imag} */,
  {32'h3d1a9cb6, 32'hbc92eff2} /* (6, 1, 13) {real, imag} */,
  {32'hbc9e6778, 32'hbc8f895d} /* (6, 1, 12) {real, imag} */,
  {32'h3cbfa981, 32'hbbf3352c} /* (6, 1, 11) {real, imag} */,
  {32'hbd7de8bb, 32'h3b5480e0} /* (6, 1, 10) {real, imag} */,
  {32'h3d3b410f, 32'h3d133930} /* (6, 1, 9) {real, imag} */,
  {32'hbc87042b, 32'hbda1e0d1} /* (6, 1, 8) {real, imag} */,
  {32'h3d4d197e, 32'h3d3c86c3} /* (6, 1, 7) {real, imag} */,
  {32'hbc07f280, 32'h3bdbc8bc} /* (6, 1, 6) {real, imag} */,
  {32'hbdcd6ed6, 32'hbcdbf5bf} /* (6, 1, 5) {real, imag} */,
  {32'hbb7b6410, 32'hbd584265} /* (6, 1, 4) {real, imag} */,
  {32'hbdd6e5a6, 32'hbd499c56} /* (6, 1, 3) {real, imag} */,
  {32'h3e395200, 32'hbec38656} /* (6, 1, 2) {real, imag} */,
  {32'h3fce42cf, 32'h3fe521ce} /* (6, 1, 1) {real, imag} */,
  {32'h405828e7, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'h3fe83bf9, 32'hbfbc41a5} /* (6, 0, 31) {real, imag} */,
  {32'hbc37a1a0, 32'h3e8d1cb4} /* (6, 0, 30) {real, imag} */,
  {32'hbd9c1b6b, 32'h3c2090c2} /* (6, 0, 29) {real, imag} */,
  {32'hbd595b27, 32'h3d98056a} /* (6, 0, 28) {real, imag} */,
  {32'hbd5edc13, 32'h3d064ccd} /* (6, 0, 27) {real, imag} */,
  {32'h3d445293, 32'hbdc82ae4} /* (6, 0, 26) {real, imag} */,
  {32'h3d404f68, 32'hbd64fc60} /* (6, 0, 25) {real, imag} */,
  {32'hbb394200, 32'hbc97a4d0} /* (6, 0, 24) {real, imag} */,
  {32'hbb4cf6f8, 32'hbd8db562} /* (6, 0, 23) {real, imag} */,
  {32'hbde0770e, 32'h3d778b18} /* (6, 0, 22) {real, imag} */,
  {32'hbce326a6, 32'h3cc6ae84} /* (6, 0, 21) {real, imag} */,
  {32'h3d3cc262, 32'h3cd50c1d} /* (6, 0, 20) {real, imag} */,
  {32'h3d08e99a, 32'hbbd06a68} /* (6, 0, 19) {real, imag} */,
  {32'h3d5adc58, 32'hbd56952e} /* (6, 0, 18) {real, imag} */,
  {32'hbd5a8976, 32'hbd8171be} /* (6, 0, 17) {real, imag} */,
  {32'hbd88ab5e, 32'h00000000} /* (6, 0, 16) {real, imag} */,
  {32'hbd5a8976, 32'h3d8171be} /* (6, 0, 15) {real, imag} */,
  {32'h3d5adc58, 32'h3d56952e} /* (6, 0, 14) {real, imag} */,
  {32'h3d08e99a, 32'h3bd06a68} /* (6, 0, 13) {real, imag} */,
  {32'h3d3cc262, 32'hbcd50c1d} /* (6, 0, 12) {real, imag} */,
  {32'hbce326a6, 32'hbcc6ae84} /* (6, 0, 11) {real, imag} */,
  {32'hbde0770e, 32'hbd778b18} /* (6, 0, 10) {real, imag} */,
  {32'hbb4cf6f8, 32'h3d8db562} /* (6, 0, 9) {real, imag} */,
  {32'hbb394200, 32'h3c97a4d0} /* (6, 0, 8) {real, imag} */,
  {32'h3d404f68, 32'h3d64fc60} /* (6, 0, 7) {real, imag} */,
  {32'h3d445293, 32'h3dc82ae4} /* (6, 0, 6) {real, imag} */,
  {32'hbd5edc13, 32'hbd064ccd} /* (6, 0, 5) {real, imag} */,
  {32'hbd595b27, 32'hbd98056a} /* (6, 0, 4) {real, imag} */,
  {32'hbd9c1b6b, 32'hbc2090c2} /* (6, 0, 3) {real, imag} */,
  {32'hbc37a1a0, 32'hbe8d1cb4} /* (6, 0, 2) {real, imag} */,
  {32'h3fe83bf9, 32'h3fbc41a5} /* (6, 0, 1) {real, imag} */,
  {32'h40554f8c, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'h3f5d5fd4, 32'hbf0542d1} /* (5, 31, 31) {real, imag} */,
  {32'h3ca0a4ff, 32'hbdb8b24b} /* (5, 31, 30) {real, imag} */,
  {32'h3db15579, 32'hbdccf1d7} /* (5, 31, 29) {real, imag} */,
  {32'h3cfbc713, 32'hbceba626} /* (5, 31, 28) {real, imag} */,
  {32'h3d27ce59, 32'hbcdabb75} /* (5, 31, 27) {real, imag} */,
  {32'h3d8266b9, 32'h3d189215} /* (5, 31, 26) {real, imag} */,
  {32'h3bcaabcc, 32'h3d23ed12} /* (5, 31, 25) {real, imag} */,
  {32'hbb5345c0, 32'h3d142070} /* (5, 31, 24) {real, imag} */,
  {32'h3d05e63e, 32'h3d0c22d7} /* (5, 31, 23) {real, imag} */,
  {32'h3b3e5e1c, 32'hbccff522} /* (5, 31, 22) {real, imag} */,
  {32'hbd7d151b, 32'h3da2aefd} /* (5, 31, 21) {real, imag} */,
  {32'h3bb43f30, 32'hbd350372} /* (5, 31, 20) {real, imag} */,
  {32'h3c131f70, 32'h3d547f60} /* (5, 31, 19) {real, imag} */,
  {32'h3c3e3374, 32'hbc1ae4b0} /* (5, 31, 18) {real, imag} */,
  {32'h3c9534da, 32'hbc6c3a92} /* (5, 31, 17) {real, imag} */,
  {32'hbd0dbd9e, 32'h00000000} /* (5, 31, 16) {real, imag} */,
  {32'h3c9534da, 32'h3c6c3a92} /* (5, 31, 15) {real, imag} */,
  {32'h3c3e3374, 32'h3c1ae4b0} /* (5, 31, 14) {real, imag} */,
  {32'h3c131f70, 32'hbd547f60} /* (5, 31, 13) {real, imag} */,
  {32'h3bb43f30, 32'h3d350372} /* (5, 31, 12) {real, imag} */,
  {32'hbd7d151b, 32'hbda2aefd} /* (5, 31, 11) {real, imag} */,
  {32'h3b3e5e1c, 32'h3ccff522} /* (5, 31, 10) {real, imag} */,
  {32'h3d05e63e, 32'hbd0c22d7} /* (5, 31, 9) {real, imag} */,
  {32'hbb5345c0, 32'hbd142070} /* (5, 31, 8) {real, imag} */,
  {32'h3bcaabcc, 32'hbd23ed12} /* (5, 31, 7) {real, imag} */,
  {32'h3d8266b9, 32'hbd189215} /* (5, 31, 6) {real, imag} */,
  {32'h3d27ce59, 32'h3cdabb75} /* (5, 31, 5) {real, imag} */,
  {32'h3cfbc713, 32'h3ceba626} /* (5, 31, 4) {real, imag} */,
  {32'h3db15579, 32'h3dccf1d7} /* (5, 31, 3) {real, imag} */,
  {32'h3ca0a4ff, 32'h3db8b24b} /* (5, 31, 2) {real, imag} */,
  {32'h3f5d5fd4, 32'h3f0542d1} /* (5, 31, 1) {real, imag} */,
  {32'h400035c1, 32'h00000000} /* (5, 31, 0) {real, imag} */,
  {32'h3f5d21d9, 32'hbef9f656} /* (5, 30, 31) {real, imag} */,
  {32'h3e35598c, 32'hbd730125} /* (5, 30, 30) {real, imag} */,
  {32'h3e25aaab, 32'hbddf0ab6} /* (5, 30, 29) {real, imag} */,
  {32'h3d804c35, 32'h3ce3f558} /* (5, 30, 28) {real, imag} */,
  {32'hbd1efd91, 32'h3db268f6} /* (5, 30, 27) {real, imag} */,
  {32'hbd4c4d2a, 32'h3d92a631} /* (5, 30, 26) {real, imag} */,
  {32'hbe0d0dd1, 32'hbc2cee08} /* (5, 30, 25) {real, imag} */,
  {32'h3dcd7b9d, 32'hbd3d1f59} /* (5, 30, 24) {real, imag} */,
  {32'h3cf69ad8, 32'hbd4b4842} /* (5, 30, 23) {real, imag} */,
  {32'hbdaabe3d, 32'h3e08fb2d} /* (5, 30, 22) {real, imag} */,
  {32'h3d50d849, 32'h3d92a57b} /* (5, 30, 21) {real, imag} */,
  {32'hbc0ca4ca, 32'hbd62c336} /* (5, 30, 20) {real, imag} */,
  {32'h3d26b186, 32'hbb4abd88} /* (5, 30, 19) {real, imag} */,
  {32'h3d42f6d2, 32'h3cbf35d3} /* (5, 30, 18) {real, imag} */,
  {32'h3c6342a1, 32'hbcaa38ec} /* (5, 30, 17) {real, imag} */,
  {32'hbd846469, 32'h00000000} /* (5, 30, 16) {real, imag} */,
  {32'h3c6342a1, 32'h3caa38ec} /* (5, 30, 15) {real, imag} */,
  {32'h3d42f6d2, 32'hbcbf35d3} /* (5, 30, 14) {real, imag} */,
  {32'h3d26b186, 32'h3b4abd88} /* (5, 30, 13) {real, imag} */,
  {32'hbc0ca4ca, 32'h3d62c336} /* (5, 30, 12) {real, imag} */,
  {32'h3d50d849, 32'hbd92a57b} /* (5, 30, 11) {real, imag} */,
  {32'hbdaabe3d, 32'hbe08fb2d} /* (5, 30, 10) {real, imag} */,
  {32'h3cf69ad8, 32'h3d4b4842} /* (5, 30, 9) {real, imag} */,
  {32'h3dcd7b9d, 32'h3d3d1f59} /* (5, 30, 8) {real, imag} */,
  {32'hbe0d0dd1, 32'h3c2cee08} /* (5, 30, 7) {real, imag} */,
  {32'hbd4c4d2a, 32'hbd92a631} /* (5, 30, 6) {real, imag} */,
  {32'hbd1efd91, 32'hbdb268f6} /* (5, 30, 5) {real, imag} */,
  {32'h3d804c35, 32'hbce3f558} /* (5, 30, 4) {real, imag} */,
  {32'h3e25aaab, 32'h3ddf0ab6} /* (5, 30, 3) {real, imag} */,
  {32'h3e35598c, 32'h3d730125} /* (5, 30, 2) {real, imag} */,
  {32'h3f5d21d9, 32'h3ef9f656} /* (5, 30, 1) {real, imag} */,
  {32'h40040d9a, 32'h00000000} /* (5, 30, 0) {real, imag} */,
  {32'h3f516f18, 32'hbe8871d0} /* (5, 29, 31) {real, imag} */,
  {32'h3e3acb88, 32'h3d3c2968} /* (5, 29, 30) {real, imag} */,
  {32'h3e1f8669, 32'hbcb02f20} /* (5, 29, 29) {real, imag} */,
  {32'h3dcdf156, 32'hbd7ac194} /* (5, 29, 28) {real, imag} */,
  {32'hbc23d76c, 32'h3e2156c8} /* (5, 29, 27) {real, imag} */,
  {32'hbce335cc, 32'h3daa2ffa} /* (5, 29, 26) {real, imag} */,
  {32'hbd182bad, 32'hbdf5db6a} /* (5, 29, 25) {real, imag} */,
  {32'h3e0a2ef5, 32'hbdcfbc2c} /* (5, 29, 24) {real, imag} */,
  {32'h3c8cc474, 32'hbd9cc018} /* (5, 29, 23) {real, imag} */,
  {32'hbe1b1bad, 32'h3b47bc40} /* (5, 29, 22) {real, imag} */,
  {32'hbd98692c, 32'h3bb8db2c} /* (5, 29, 21) {real, imag} */,
  {32'h3d14b246, 32'hbba3fd80} /* (5, 29, 20) {real, imag} */,
  {32'h3d0dd6a5, 32'h3c9d9564} /* (5, 29, 19) {real, imag} */,
  {32'hbd242d0f, 32'h3e14fc16} /* (5, 29, 18) {real, imag} */,
  {32'h3a7b5820, 32'h3d735aef} /* (5, 29, 17) {real, imag} */,
  {32'h3b88efec, 32'h00000000} /* (5, 29, 16) {real, imag} */,
  {32'h3a7b5820, 32'hbd735aef} /* (5, 29, 15) {real, imag} */,
  {32'hbd242d0f, 32'hbe14fc16} /* (5, 29, 14) {real, imag} */,
  {32'h3d0dd6a5, 32'hbc9d9564} /* (5, 29, 13) {real, imag} */,
  {32'h3d14b246, 32'h3ba3fd80} /* (5, 29, 12) {real, imag} */,
  {32'hbd98692c, 32'hbbb8db2c} /* (5, 29, 11) {real, imag} */,
  {32'hbe1b1bad, 32'hbb47bc40} /* (5, 29, 10) {real, imag} */,
  {32'h3c8cc474, 32'h3d9cc018} /* (5, 29, 9) {real, imag} */,
  {32'h3e0a2ef5, 32'h3dcfbc2c} /* (5, 29, 8) {real, imag} */,
  {32'hbd182bad, 32'h3df5db6a} /* (5, 29, 7) {real, imag} */,
  {32'hbce335cc, 32'hbdaa2ffa} /* (5, 29, 6) {real, imag} */,
  {32'hbc23d76c, 32'hbe2156c8} /* (5, 29, 5) {real, imag} */,
  {32'h3dcdf156, 32'h3d7ac194} /* (5, 29, 4) {real, imag} */,
  {32'h3e1f8669, 32'h3cb02f20} /* (5, 29, 3) {real, imag} */,
  {32'h3e3acb88, 32'hbd3c2968} /* (5, 29, 2) {real, imag} */,
  {32'h3f516f18, 32'h3e8871d0} /* (5, 29, 1) {real, imag} */,
  {32'h3fec01a5, 32'h00000000} /* (5, 29, 0) {real, imag} */,
  {32'h3f2bc93a, 32'hbe1148f4} /* (5, 28, 31) {real, imag} */,
  {32'h3ceee107, 32'h3c81cc34} /* (5, 28, 30) {real, imag} */,
  {32'h3e5717bf, 32'h3ceb83b0} /* (5, 28, 29) {real, imag} */,
  {32'hbd982130, 32'h3cc76b33} /* (5, 28, 28) {real, imag} */,
  {32'hbdbae2f4, 32'hbd3bd256} /* (5, 28, 27) {real, imag} */,
  {32'h3e097ac1, 32'h3b431428} /* (5, 28, 26) {real, imag} */,
  {32'h3d5490b0, 32'h3cb1dbf0} /* (5, 28, 25) {real, imag} */,
  {32'h3d8d2998, 32'h3af387d0} /* (5, 28, 24) {real, imag} */,
  {32'h3d4aabb0, 32'hbe04f5b3} /* (5, 28, 23) {real, imag} */,
  {32'hbd46efe6, 32'hbd79a8f0} /* (5, 28, 22) {real, imag} */,
  {32'hbdac6a20, 32'h3dccb767} /* (5, 28, 21) {real, imag} */,
  {32'hbceae2c1, 32'hbd9624f9} /* (5, 28, 20) {real, imag} */,
  {32'h3b0b01a8, 32'hbd41b43b} /* (5, 28, 19) {real, imag} */,
  {32'hbda17fea, 32'h3c00d870} /* (5, 28, 18) {real, imag} */,
  {32'hbd0379f5, 32'hbd703a7f} /* (5, 28, 17) {real, imag} */,
  {32'h3d80cf8d, 32'h00000000} /* (5, 28, 16) {real, imag} */,
  {32'hbd0379f5, 32'h3d703a7f} /* (5, 28, 15) {real, imag} */,
  {32'hbda17fea, 32'hbc00d870} /* (5, 28, 14) {real, imag} */,
  {32'h3b0b01a8, 32'h3d41b43b} /* (5, 28, 13) {real, imag} */,
  {32'hbceae2c1, 32'h3d9624f9} /* (5, 28, 12) {real, imag} */,
  {32'hbdac6a20, 32'hbdccb767} /* (5, 28, 11) {real, imag} */,
  {32'hbd46efe6, 32'h3d79a8f0} /* (5, 28, 10) {real, imag} */,
  {32'h3d4aabb0, 32'h3e04f5b3} /* (5, 28, 9) {real, imag} */,
  {32'h3d8d2998, 32'hbaf387d0} /* (5, 28, 8) {real, imag} */,
  {32'h3d5490b0, 32'hbcb1dbf0} /* (5, 28, 7) {real, imag} */,
  {32'h3e097ac1, 32'hbb431428} /* (5, 28, 6) {real, imag} */,
  {32'hbdbae2f4, 32'h3d3bd256} /* (5, 28, 5) {real, imag} */,
  {32'hbd982130, 32'hbcc76b33} /* (5, 28, 4) {real, imag} */,
  {32'h3e5717bf, 32'hbceb83b0} /* (5, 28, 3) {real, imag} */,
  {32'h3ceee107, 32'hbc81cc34} /* (5, 28, 2) {real, imag} */,
  {32'h3f2bc93a, 32'h3e1148f4} /* (5, 28, 1) {real, imag} */,
  {32'h3fecdf92, 32'h00000000} /* (5, 28, 0) {real, imag} */,
  {32'h3f0aeea5, 32'h3d2fc694} /* (5, 27, 31) {real, imag} */,
  {32'hbc0ec7cc, 32'h3d6607a4} /* (5, 27, 30) {real, imag} */,
  {32'h3e1a1748, 32'hbe209dc6} /* (5, 27, 29) {real, imag} */,
  {32'hbdf55f4a, 32'hbcbc1804} /* (5, 27, 28) {real, imag} */,
  {32'hbc0ac318, 32'h3d248c21} /* (5, 27, 27) {real, imag} */,
  {32'h3de04108, 32'hbcf8242d} /* (5, 27, 26) {real, imag} */,
  {32'hbdd299a6, 32'hbc09e8c8} /* (5, 27, 25) {real, imag} */,
  {32'hbd28d36f, 32'h3d0d0964} /* (5, 27, 24) {real, imag} */,
  {32'h3c112bfc, 32'h3da0abb3} /* (5, 27, 23) {real, imag} */,
  {32'h3d68d25e, 32'hbbb990bc} /* (5, 27, 22) {real, imag} */,
  {32'hbb8184b0, 32'hbda6f3f8} /* (5, 27, 21) {real, imag} */,
  {32'hbd3ec31c, 32'hbd8ccd15} /* (5, 27, 20) {real, imag} */,
  {32'hbdb4d452, 32'h3cbecc44} /* (5, 27, 19) {real, imag} */,
  {32'hbd260dca, 32'hbd49c4bd} /* (5, 27, 18) {real, imag} */,
  {32'h3cb50b3a, 32'hbb5b8250} /* (5, 27, 17) {real, imag} */,
  {32'hbde855b4, 32'h00000000} /* (5, 27, 16) {real, imag} */,
  {32'h3cb50b3a, 32'h3b5b8250} /* (5, 27, 15) {real, imag} */,
  {32'hbd260dca, 32'h3d49c4bd} /* (5, 27, 14) {real, imag} */,
  {32'hbdb4d452, 32'hbcbecc44} /* (5, 27, 13) {real, imag} */,
  {32'hbd3ec31c, 32'h3d8ccd15} /* (5, 27, 12) {real, imag} */,
  {32'hbb8184b0, 32'h3da6f3f8} /* (5, 27, 11) {real, imag} */,
  {32'h3d68d25e, 32'h3bb990bc} /* (5, 27, 10) {real, imag} */,
  {32'h3c112bfc, 32'hbda0abb3} /* (5, 27, 9) {real, imag} */,
  {32'hbd28d36f, 32'hbd0d0964} /* (5, 27, 8) {real, imag} */,
  {32'hbdd299a6, 32'h3c09e8c8} /* (5, 27, 7) {real, imag} */,
  {32'h3de04108, 32'h3cf8242d} /* (5, 27, 6) {real, imag} */,
  {32'hbc0ac318, 32'hbd248c21} /* (5, 27, 5) {real, imag} */,
  {32'hbdf55f4a, 32'h3cbc1804} /* (5, 27, 4) {real, imag} */,
  {32'h3e1a1748, 32'h3e209dc6} /* (5, 27, 3) {real, imag} */,
  {32'hbc0ec7cc, 32'hbd6607a4} /* (5, 27, 2) {real, imag} */,
  {32'h3f0aeea5, 32'hbd2fc694} /* (5, 27, 1) {real, imag} */,
  {32'h3fe23158, 32'h00000000} /* (5, 27, 0) {real, imag} */,
  {32'h3f0edde5, 32'h3c00ea90} /* (5, 26, 31) {real, imag} */,
  {32'h3cdf155a, 32'h3d96c0f8} /* (5, 26, 30) {real, imag} */,
  {32'hbd329850, 32'hbe0f2679} /* (5, 26, 29) {real, imag} */,
  {32'hbd2634c2, 32'hbbaf81a0} /* (5, 26, 28) {real, imag} */,
  {32'h3da36620, 32'h3dd342a2} /* (5, 26, 27) {real, imag} */,
  {32'hbc551341, 32'hbc932b1d} /* (5, 26, 26) {real, imag} */,
  {32'hbbf2cc7c, 32'hbd5a238c} /* (5, 26, 25) {real, imag} */,
  {32'hbd98e7e2, 32'hbd8001c5} /* (5, 26, 24) {real, imag} */,
  {32'hbd229b3e, 32'h3e0b5586} /* (5, 26, 23) {real, imag} */,
  {32'hbd8b51ab, 32'hbccfdfdc} /* (5, 26, 22) {real, imag} */,
  {32'h3d56eae6, 32'h3cca1476} /* (5, 26, 21) {real, imag} */,
  {32'hbdc03bc2, 32'h3b8e9d20} /* (5, 26, 20) {real, imag} */,
  {32'hbcaeb0df, 32'h3c830854} /* (5, 26, 19) {real, imag} */,
  {32'hbad7bb00, 32'hbcbee2e3} /* (5, 26, 18) {real, imag} */,
  {32'hbce4f5c0, 32'hbaefbd78} /* (5, 26, 17) {real, imag} */,
  {32'h3d71ffec, 32'h00000000} /* (5, 26, 16) {real, imag} */,
  {32'hbce4f5c0, 32'h3aefbd78} /* (5, 26, 15) {real, imag} */,
  {32'hbad7bb00, 32'h3cbee2e3} /* (5, 26, 14) {real, imag} */,
  {32'hbcaeb0df, 32'hbc830854} /* (5, 26, 13) {real, imag} */,
  {32'hbdc03bc2, 32'hbb8e9d20} /* (5, 26, 12) {real, imag} */,
  {32'h3d56eae6, 32'hbcca1476} /* (5, 26, 11) {real, imag} */,
  {32'hbd8b51ab, 32'h3ccfdfdc} /* (5, 26, 10) {real, imag} */,
  {32'hbd229b3e, 32'hbe0b5586} /* (5, 26, 9) {real, imag} */,
  {32'hbd98e7e2, 32'h3d8001c5} /* (5, 26, 8) {real, imag} */,
  {32'hbbf2cc7c, 32'h3d5a238c} /* (5, 26, 7) {real, imag} */,
  {32'hbc551341, 32'h3c932b1d} /* (5, 26, 6) {real, imag} */,
  {32'h3da36620, 32'hbdd342a2} /* (5, 26, 5) {real, imag} */,
  {32'hbd2634c2, 32'h3baf81a0} /* (5, 26, 4) {real, imag} */,
  {32'hbd329850, 32'h3e0f2679} /* (5, 26, 3) {real, imag} */,
  {32'h3cdf155a, 32'hbd96c0f8} /* (5, 26, 2) {real, imag} */,
  {32'h3f0edde5, 32'hbc00ea90} /* (5, 26, 1) {real, imag} */,
  {32'h3fdcc66c, 32'h00000000} /* (5, 26, 0) {real, imag} */,
  {32'h3e9266f6, 32'hbba89f20} /* (5, 25, 31) {real, imag} */,
  {32'h3d9fa41c, 32'h3da68e40} /* (5, 25, 30) {real, imag} */,
  {32'hbdb86666, 32'hbdf5fbe1} /* (5, 25, 29) {real, imag} */,
  {32'hbdbff5b6, 32'h3c1d2ee4} /* (5, 25, 28) {real, imag} */,
  {32'h3dd170c6, 32'hbd16cdc4} /* (5, 25, 27) {real, imag} */,
  {32'h3e1be93c, 32'hbd0f2186} /* (5, 25, 26) {real, imag} */,
  {32'h3da7f70f, 32'h3db0e4bc} /* (5, 25, 25) {real, imag} */,
  {32'h3c8591f1, 32'hbcec2308} /* (5, 25, 24) {real, imag} */,
  {32'hbcd1a208, 32'h3cfb1f7e} /* (5, 25, 23) {real, imag} */,
  {32'hbcb08bda, 32'h3d03d854} /* (5, 25, 22) {real, imag} */,
  {32'h3d7e554a, 32'hbd75bcb6} /* (5, 25, 21) {real, imag} */,
  {32'hbe109f66, 32'h3d9a05f8} /* (5, 25, 20) {real, imag} */,
  {32'h3d09010a, 32'hbd3d2028} /* (5, 25, 19) {real, imag} */,
  {32'hbcbb9aa4, 32'hbb3df130} /* (5, 25, 18) {real, imag} */,
  {32'hbd5e73ab, 32'hbbcb92e8} /* (5, 25, 17) {real, imag} */,
  {32'hbda4c52c, 32'h00000000} /* (5, 25, 16) {real, imag} */,
  {32'hbd5e73ab, 32'h3bcb92e8} /* (5, 25, 15) {real, imag} */,
  {32'hbcbb9aa4, 32'h3b3df130} /* (5, 25, 14) {real, imag} */,
  {32'h3d09010a, 32'h3d3d2028} /* (5, 25, 13) {real, imag} */,
  {32'hbe109f66, 32'hbd9a05f8} /* (5, 25, 12) {real, imag} */,
  {32'h3d7e554a, 32'h3d75bcb6} /* (5, 25, 11) {real, imag} */,
  {32'hbcb08bda, 32'hbd03d854} /* (5, 25, 10) {real, imag} */,
  {32'hbcd1a208, 32'hbcfb1f7e} /* (5, 25, 9) {real, imag} */,
  {32'h3c8591f1, 32'h3cec2308} /* (5, 25, 8) {real, imag} */,
  {32'h3da7f70f, 32'hbdb0e4bc} /* (5, 25, 7) {real, imag} */,
  {32'h3e1be93c, 32'h3d0f2186} /* (5, 25, 6) {real, imag} */,
  {32'h3dd170c6, 32'h3d16cdc4} /* (5, 25, 5) {real, imag} */,
  {32'hbdbff5b6, 32'hbc1d2ee4} /* (5, 25, 4) {real, imag} */,
  {32'hbdb86666, 32'h3df5fbe1} /* (5, 25, 3) {real, imag} */,
  {32'h3d9fa41c, 32'hbda68e40} /* (5, 25, 2) {real, imag} */,
  {32'h3e9266f6, 32'h3ba89f20} /* (5, 25, 1) {real, imag} */,
  {32'h3fc13279, 32'h00000000} /* (5, 25, 0) {real, imag} */,
  {32'h3e42172f, 32'hbd95cb1c} /* (5, 24, 31) {real, imag} */,
  {32'h3ca46d98, 32'h3e0b0fa6} /* (5, 24, 30) {real, imag} */,
  {32'h3db89581, 32'hbe0244f8} /* (5, 24, 29) {real, imag} */,
  {32'hbdb6bdee, 32'h3bd44570} /* (5, 24, 28) {real, imag} */,
  {32'h3d819985, 32'hbe03eb5f} /* (5, 24, 27) {real, imag} */,
  {32'h3daebd22, 32'hbd757f84} /* (5, 24, 26) {real, imag} */,
  {32'hbd55349e, 32'h3dcfd253} /* (5, 24, 25) {real, imag} */,
  {32'h3cef22ca, 32'hbcb2d156} /* (5, 24, 24) {real, imag} */,
  {32'h3cfae572, 32'hba827460} /* (5, 24, 23) {real, imag} */,
  {32'h3d30df3c, 32'h3db0b326} /* (5, 24, 22) {real, imag} */,
  {32'hbd6e475a, 32'h3d2574f6} /* (5, 24, 21) {real, imag} */,
  {32'h3a2d7d70, 32'h3d1b85f0} /* (5, 24, 20) {real, imag} */,
  {32'hbd9c148e, 32'h3e106fb2} /* (5, 24, 19) {real, imag} */,
  {32'hbd33c82b, 32'h3d300aee} /* (5, 24, 18) {real, imag} */,
  {32'h3c9ce4c8, 32'h3d4aecce} /* (5, 24, 17) {real, imag} */,
  {32'hbd6bbb43, 32'h00000000} /* (5, 24, 16) {real, imag} */,
  {32'h3c9ce4c8, 32'hbd4aecce} /* (5, 24, 15) {real, imag} */,
  {32'hbd33c82b, 32'hbd300aee} /* (5, 24, 14) {real, imag} */,
  {32'hbd9c148e, 32'hbe106fb2} /* (5, 24, 13) {real, imag} */,
  {32'h3a2d7d70, 32'hbd1b85f0} /* (5, 24, 12) {real, imag} */,
  {32'hbd6e475a, 32'hbd2574f6} /* (5, 24, 11) {real, imag} */,
  {32'h3d30df3c, 32'hbdb0b326} /* (5, 24, 10) {real, imag} */,
  {32'h3cfae572, 32'h3a827460} /* (5, 24, 9) {real, imag} */,
  {32'h3cef22ca, 32'h3cb2d156} /* (5, 24, 8) {real, imag} */,
  {32'hbd55349e, 32'hbdcfd253} /* (5, 24, 7) {real, imag} */,
  {32'h3daebd22, 32'h3d757f84} /* (5, 24, 6) {real, imag} */,
  {32'h3d819985, 32'h3e03eb5f} /* (5, 24, 5) {real, imag} */,
  {32'hbdb6bdee, 32'hbbd44570} /* (5, 24, 4) {real, imag} */,
  {32'h3db89581, 32'h3e0244f8} /* (5, 24, 3) {real, imag} */,
  {32'h3ca46d98, 32'hbe0b0fa6} /* (5, 24, 2) {real, imag} */,
  {32'h3e42172f, 32'h3d95cb1c} /* (5, 24, 1) {real, imag} */,
  {32'h3faf36ff, 32'h00000000} /* (5, 24, 0) {real, imag} */,
  {32'hbd1df27a, 32'hbe618b36} /* (5, 23, 31) {real, imag} */,
  {32'h3d908105, 32'h3d3ad840} /* (5, 23, 30) {real, imag} */,
  {32'hbd1c66f6, 32'hbde9342c} /* (5, 23, 29) {real, imag} */,
  {32'hbcb2375b, 32'hbc2deeca} /* (5, 23, 28) {real, imag} */,
  {32'h3d3a80f0, 32'hbdeb029a} /* (5, 23, 27) {real, imag} */,
  {32'hbd1ee254, 32'hbd996990} /* (5, 23, 26) {real, imag} */,
  {32'hbd050f32, 32'h3c1a8fdc} /* (5, 23, 25) {real, imag} */,
  {32'h3cc67478, 32'h3cd69d1a} /* (5, 23, 24) {real, imag} */,
  {32'h3d6eea66, 32'hbc82bfa2} /* (5, 23, 23) {real, imag} */,
  {32'hbd9f3565, 32'h3c907c17} /* (5, 23, 22) {real, imag} */,
  {32'h3b93d656, 32'h3db089ff} /* (5, 23, 21) {real, imag} */,
  {32'hbc852d9c, 32'h3bd45f80} /* (5, 23, 20) {real, imag} */,
  {32'hbc49537c, 32'h3cbc4f07} /* (5, 23, 19) {real, imag} */,
  {32'hbc1d0e4c, 32'h3d8f97ff} /* (5, 23, 18) {real, imag} */,
  {32'h3d2dc1cd, 32'hbcd73280} /* (5, 23, 17) {real, imag} */,
  {32'h3cbc4300, 32'h00000000} /* (5, 23, 16) {real, imag} */,
  {32'h3d2dc1cd, 32'h3cd73280} /* (5, 23, 15) {real, imag} */,
  {32'hbc1d0e4c, 32'hbd8f97ff} /* (5, 23, 14) {real, imag} */,
  {32'hbc49537c, 32'hbcbc4f07} /* (5, 23, 13) {real, imag} */,
  {32'hbc852d9c, 32'hbbd45f80} /* (5, 23, 12) {real, imag} */,
  {32'h3b93d656, 32'hbdb089ff} /* (5, 23, 11) {real, imag} */,
  {32'hbd9f3565, 32'hbc907c17} /* (5, 23, 10) {real, imag} */,
  {32'h3d6eea66, 32'h3c82bfa2} /* (5, 23, 9) {real, imag} */,
  {32'h3cc67478, 32'hbcd69d1a} /* (5, 23, 8) {real, imag} */,
  {32'hbd050f32, 32'hbc1a8fdc} /* (5, 23, 7) {real, imag} */,
  {32'hbd1ee254, 32'h3d996990} /* (5, 23, 6) {real, imag} */,
  {32'h3d3a80f0, 32'h3deb029a} /* (5, 23, 5) {real, imag} */,
  {32'hbcb2375b, 32'h3c2deeca} /* (5, 23, 4) {real, imag} */,
  {32'hbd1c66f6, 32'h3de9342c} /* (5, 23, 3) {real, imag} */,
  {32'h3d908105, 32'hbd3ad840} /* (5, 23, 2) {real, imag} */,
  {32'hbd1df27a, 32'h3e618b36} /* (5, 23, 1) {real, imag} */,
  {32'h3f9275e4, 32'h00000000} /* (5, 23, 0) {real, imag} */,
  {32'hbe157118, 32'hbe71c773} /* (5, 22, 31) {real, imag} */,
  {32'h3c832f84, 32'h3daa38aa} /* (5, 22, 30) {real, imag} */,
  {32'hbd81430e, 32'hbe3a8b4c} /* (5, 22, 29) {real, imag} */,
  {32'hbdb581d6, 32'h3dacd972} /* (5, 22, 28) {real, imag} */,
  {32'h3ddc38f9, 32'hbd9315aa} /* (5, 22, 27) {real, imag} */,
  {32'h3c67edcf, 32'hbd2c8b1a} /* (5, 22, 26) {real, imag} */,
  {32'h3d775e6e, 32'h3c03d9a6} /* (5, 22, 25) {real, imag} */,
  {32'hbcee2d62, 32'hbd5128e4} /* (5, 22, 24) {real, imag} */,
  {32'hbcd997e7, 32'h3da36408} /* (5, 22, 23) {real, imag} */,
  {32'h3d32b976, 32'h3d3d4d03} /* (5, 22, 22) {real, imag} */,
  {32'hbd72eea5, 32'h3d084db8} /* (5, 22, 21) {real, imag} */,
  {32'hbb2f04c0, 32'hbc2f7f18} /* (5, 22, 20) {real, imag} */,
  {32'hbae0ecb0, 32'h3cc617f6} /* (5, 22, 19) {real, imag} */,
  {32'h3d78778a, 32'hbd328223} /* (5, 22, 18) {real, imag} */,
  {32'hbcc71048, 32'h3cbef18b} /* (5, 22, 17) {real, imag} */,
  {32'hbda99862, 32'h00000000} /* (5, 22, 16) {real, imag} */,
  {32'hbcc71048, 32'hbcbef18b} /* (5, 22, 15) {real, imag} */,
  {32'h3d78778a, 32'h3d328223} /* (5, 22, 14) {real, imag} */,
  {32'hbae0ecb0, 32'hbcc617f6} /* (5, 22, 13) {real, imag} */,
  {32'hbb2f04c0, 32'h3c2f7f18} /* (5, 22, 12) {real, imag} */,
  {32'hbd72eea5, 32'hbd084db8} /* (5, 22, 11) {real, imag} */,
  {32'h3d32b976, 32'hbd3d4d03} /* (5, 22, 10) {real, imag} */,
  {32'hbcd997e7, 32'hbda36408} /* (5, 22, 9) {real, imag} */,
  {32'hbcee2d62, 32'h3d5128e4} /* (5, 22, 8) {real, imag} */,
  {32'h3d775e6e, 32'hbc03d9a6} /* (5, 22, 7) {real, imag} */,
  {32'h3c67edcf, 32'h3d2c8b1a} /* (5, 22, 6) {real, imag} */,
  {32'h3ddc38f9, 32'h3d9315aa} /* (5, 22, 5) {real, imag} */,
  {32'hbdb581d6, 32'hbdacd972} /* (5, 22, 4) {real, imag} */,
  {32'hbd81430e, 32'h3e3a8b4c} /* (5, 22, 3) {real, imag} */,
  {32'h3c832f84, 32'hbdaa38aa} /* (5, 22, 2) {real, imag} */,
  {32'hbe157118, 32'h3e71c773} /* (5, 22, 1) {real, imag} */,
  {32'h3f585d0a, 32'h00000000} /* (5, 22, 0) {real, imag} */,
  {32'hbe054d6b, 32'hbdeef332} /* (5, 21, 31) {real, imag} */,
  {32'hbd905456, 32'h3cc6dc24} /* (5, 21, 30) {real, imag} */,
  {32'h3d1904b2, 32'hbe0d5a76} /* (5, 21, 29) {real, imag} */,
  {32'hbdcdb4a4, 32'h3cf7978c} /* (5, 21, 28) {real, imag} */,
  {32'h3a7de6e0, 32'hbc824c1a} /* (5, 21, 27) {real, imag} */,
  {32'hbdf229d4, 32'hbcfeabc6} /* (5, 21, 26) {real, imag} */,
  {32'h3dc02ea8, 32'h3de3f915} /* (5, 21, 25) {real, imag} */,
  {32'hbd128fd2, 32'hbe01d1b3} /* (5, 21, 24) {real, imag} */,
  {32'h3a443880, 32'h3d1cc1ec} /* (5, 21, 23) {real, imag} */,
  {32'hbbf4c75c, 32'h3cefbd7b} /* (5, 21, 22) {real, imag} */,
  {32'hbc003410, 32'hbdb82dcf} /* (5, 21, 21) {real, imag} */,
  {32'h3ccd4bee, 32'h3c0ff798} /* (5, 21, 20) {real, imag} */,
  {32'h3a2b3440, 32'hbce6d63e} /* (5, 21, 19) {real, imag} */,
  {32'hbcb748b4, 32'h3d64f74d} /* (5, 21, 18) {real, imag} */,
  {32'h3b7eda70, 32'h3d8fc7f0} /* (5, 21, 17) {real, imag} */,
  {32'h3c978d92, 32'h00000000} /* (5, 21, 16) {real, imag} */,
  {32'h3b7eda70, 32'hbd8fc7f0} /* (5, 21, 15) {real, imag} */,
  {32'hbcb748b4, 32'hbd64f74d} /* (5, 21, 14) {real, imag} */,
  {32'h3a2b3440, 32'h3ce6d63e} /* (5, 21, 13) {real, imag} */,
  {32'h3ccd4bee, 32'hbc0ff798} /* (5, 21, 12) {real, imag} */,
  {32'hbc003410, 32'h3db82dcf} /* (5, 21, 11) {real, imag} */,
  {32'hbbf4c75c, 32'hbcefbd7b} /* (5, 21, 10) {real, imag} */,
  {32'h3a443880, 32'hbd1cc1ec} /* (5, 21, 9) {real, imag} */,
  {32'hbd128fd2, 32'h3e01d1b3} /* (5, 21, 8) {real, imag} */,
  {32'h3dc02ea8, 32'hbde3f915} /* (5, 21, 7) {real, imag} */,
  {32'hbdf229d4, 32'h3cfeabc6} /* (5, 21, 6) {real, imag} */,
  {32'h3a7de6e0, 32'h3c824c1a} /* (5, 21, 5) {real, imag} */,
  {32'hbdcdb4a4, 32'hbcf7978c} /* (5, 21, 4) {real, imag} */,
  {32'h3d1904b2, 32'h3e0d5a76} /* (5, 21, 3) {real, imag} */,
  {32'hbd905456, 32'hbcc6dc24} /* (5, 21, 2) {real, imag} */,
  {32'hbe054d6b, 32'h3deef332} /* (5, 21, 1) {real, imag} */,
  {32'h3f403f92, 32'h00000000} /* (5, 21, 0) {real, imag} */,
  {32'hbd5c613c, 32'hbd279a8d} /* (5, 20, 31) {real, imag} */,
  {32'hbdb55a0d, 32'h3c22c6c4} /* (5, 20, 30) {real, imag} */,
  {32'h3d1e9ef8, 32'hbe11a847} /* (5, 20, 29) {real, imag} */,
  {32'hbd703a2c, 32'hbd942f89} /* (5, 20, 28) {real, imag} */,
  {32'hbd918444, 32'hbd729eb2} /* (5, 20, 27) {real, imag} */,
  {32'h3cc7f7b8, 32'hbc878b18} /* (5, 20, 26) {real, imag} */,
  {32'h3cdd9244, 32'h3e4e3271} /* (5, 20, 25) {real, imag} */,
  {32'hbdd5998e, 32'h3cd2825d} /* (5, 20, 24) {real, imag} */,
  {32'hbc8ab74c, 32'hbd1a317b} /* (5, 20, 23) {real, imag} */,
  {32'hbdde1c92, 32'hbd08b17d} /* (5, 20, 22) {real, imag} */,
  {32'hbd339b07, 32'h3dc9d7a0} /* (5, 20, 21) {real, imag} */,
  {32'hbca4e700, 32'hbb50f060} /* (5, 20, 20) {real, imag} */,
  {32'h3de99ede, 32'h3d167a7d} /* (5, 20, 19) {real, imag} */,
  {32'h3c69fcb6, 32'h3d4e108f} /* (5, 20, 18) {real, imag} */,
  {32'hbd0d9d32, 32'hbb594530} /* (5, 20, 17) {real, imag} */,
  {32'hbce89335, 32'h00000000} /* (5, 20, 16) {real, imag} */,
  {32'hbd0d9d32, 32'h3b594530} /* (5, 20, 15) {real, imag} */,
  {32'h3c69fcb6, 32'hbd4e108f} /* (5, 20, 14) {real, imag} */,
  {32'h3de99ede, 32'hbd167a7d} /* (5, 20, 13) {real, imag} */,
  {32'hbca4e700, 32'h3b50f060} /* (5, 20, 12) {real, imag} */,
  {32'hbd339b07, 32'hbdc9d7a0} /* (5, 20, 11) {real, imag} */,
  {32'hbdde1c92, 32'h3d08b17d} /* (5, 20, 10) {real, imag} */,
  {32'hbc8ab74c, 32'h3d1a317b} /* (5, 20, 9) {real, imag} */,
  {32'hbdd5998e, 32'hbcd2825d} /* (5, 20, 8) {real, imag} */,
  {32'h3cdd9244, 32'hbe4e3271} /* (5, 20, 7) {real, imag} */,
  {32'h3cc7f7b8, 32'h3c878b18} /* (5, 20, 6) {real, imag} */,
  {32'hbd918444, 32'h3d729eb2} /* (5, 20, 5) {real, imag} */,
  {32'hbd703a2c, 32'h3d942f89} /* (5, 20, 4) {real, imag} */,
  {32'h3d1e9ef8, 32'h3e11a847} /* (5, 20, 3) {real, imag} */,
  {32'hbdb55a0d, 32'hbc22c6c4} /* (5, 20, 2) {real, imag} */,
  {32'hbd5c613c, 32'h3d279a8d} /* (5, 20, 1) {real, imag} */,
  {32'h3f4612eb, 32'h00000000} /* (5, 20, 0) {real, imag} */,
  {32'hbe3a1410, 32'hbcab89a8} /* (5, 19, 31) {real, imag} */,
  {32'hbdaa292e, 32'hbd36ed44} /* (5, 19, 30) {real, imag} */,
  {32'hbc978d00, 32'hbe1d8f8a} /* (5, 19, 29) {real, imag} */,
  {32'hbdb0cf86, 32'hbd75a038} /* (5, 19, 28) {real, imag} */,
  {32'hbd76ce49, 32'hbd511d7a} /* (5, 19, 27) {real, imag} */,
  {32'h3cec5304, 32'h3d0120a3} /* (5, 19, 26) {real, imag} */,
  {32'h3de45732, 32'h3ccacf12} /* (5, 19, 25) {real, imag} */,
  {32'hbdd11fd0, 32'h3cb4fee0} /* (5, 19, 24) {real, imag} */,
  {32'hbdc0c84c, 32'hbc800e70} /* (5, 19, 23) {real, imag} */,
  {32'hbd2cbd86, 32'hb9f8b800} /* (5, 19, 22) {real, imag} */,
  {32'hbdc7d986, 32'h3d6c02aa} /* (5, 19, 21) {real, imag} */,
  {32'hbdbce2bd, 32'h3c2ea6e8} /* (5, 19, 20) {real, imag} */,
  {32'hbd2b8fa9, 32'hbcd3ee7c} /* (5, 19, 19) {real, imag} */,
  {32'hbac725c0, 32'h3c9c2184} /* (5, 19, 18) {real, imag} */,
  {32'h3c90534a, 32'h3d2792dc} /* (5, 19, 17) {real, imag} */,
  {32'h3b67d948, 32'h00000000} /* (5, 19, 16) {real, imag} */,
  {32'h3c90534a, 32'hbd2792dc} /* (5, 19, 15) {real, imag} */,
  {32'hbac725c0, 32'hbc9c2184} /* (5, 19, 14) {real, imag} */,
  {32'hbd2b8fa9, 32'h3cd3ee7c} /* (5, 19, 13) {real, imag} */,
  {32'hbdbce2bd, 32'hbc2ea6e8} /* (5, 19, 12) {real, imag} */,
  {32'hbdc7d986, 32'hbd6c02aa} /* (5, 19, 11) {real, imag} */,
  {32'hbd2cbd86, 32'h39f8b800} /* (5, 19, 10) {real, imag} */,
  {32'hbdc0c84c, 32'h3c800e70} /* (5, 19, 9) {real, imag} */,
  {32'hbdd11fd0, 32'hbcb4fee0} /* (5, 19, 8) {real, imag} */,
  {32'h3de45732, 32'hbccacf12} /* (5, 19, 7) {real, imag} */,
  {32'h3cec5304, 32'hbd0120a3} /* (5, 19, 6) {real, imag} */,
  {32'hbd76ce49, 32'h3d511d7a} /* (5, 19, 5) {real, imag} */,
  {32'hbdb0cf86, 32'h3d75a038} /* (5, 19, 4) {real, imag} */,
  {32'hbc978d00, 32'h3e1d8f8a} /* (5, 19, 3) {real, imag} */,
  {32'hbdaa292e, 32'h3d36ed44} /* (5, 19, 2) {real, imag} */,
  {32'hbe3a1410, 32'h3cab89a8} /* (5, 19, 1) {real, imag} */,
  {32'h3e921b0c, 32'h00000000} /* (5, 19, 0) {real, imag} */,
  {32'hbe871ec2, 32'h3cad5516} /* (5, 18, 31) {real, imag} */,
  {32'hbccb931c, 32'h3dc65f19} /* (5, 18, 30) {real, imag} */,
  {32'hbd85b697, 32'hbe06b288} /* (5, 18, 29) {real, imag} */,
  {32'hbe093d40, 32'hbdb7884b} /* (5, 18, 28) {real, imag} */,
  {32'h3d88f802, 32'hbc55ef58} /* (5, 18, 27) {real, imag} */,
  {32'h3c816de6, 32'h3c8f2306} /* (5, 18, 26) {real, imag} */,
  {32'h3d2e85f4, 32'h3cb133e4} /* (5, 18, 25) {real, imag} */,
  {32'h3b6002c0, 32'h3d8bc79d} /* (5, 18, 24) {real, imag} */,
  {32'h3d4e0adc, 32'h3d80f9ce} /* (5, 18, 23) {real, imag} */,
  {32'h3b7734ec, 32'hbb80dfd0} /* (5, 18, 22) {real, imag} */,
  {32'h3d008844, 32'hbc7db6fc} /* (5, 18, 21) {real, imag} */,
  {32'hbddc6b40, 32'hbcc439fd} /* (5, 18, 20) {real, imag} */,
  {32'hbccdaf28, 32'h3d942408} /* (5, 18, 19) {real, imag} */,
  {32'hbe0bceed, 32'h3caffbfa} /* (5, 18, 18) {real, imag} */,
  {32'hbceb9f3a, 32'h3d89febc} /* (5, 18, 17) {real, imag} */,
  {32'hbdac5c58, 32'h00000000} /* (5, 18, 16) {real, imag} */,
  {32'hbceb9f3a, 32'hbd89febc} /* (5, 18, 15) {real, imag} */,
  {32'hbe0bceed, 32'hbcaffbfa} /* (5, 18, 14) {real, imag} */,
  {32'hbccdaf28, 32'hbd942408} /* (5, 18, 13) {real, imag} */,
  {32'hbddc6b40, 32'h3cc439fd} /* (5, 18, 12) {real, imag} */,
  {32'h3d008844, 32'h3c7db6fc} /* (5, 18, 11) {real, imag} */,
  {32'h3b7734ec, 32'h3b80dfd0} /* (5, 18, 10) {real, imag} */,
  {32'h3d4e0adc, 32'hbd80f9ce} /* (5, 18, 9) {real, imag} */,
  {32'h3b6002c0, 32'hbd8bc79d} /* (5, 18, 8) {real, imag} */,
  {32'h3d2e85f4, 32'hbcb133e4} /* (5, 18, 7) {real, imag} */,
  {32'h3c816de6, 32'hbc8f2306} /* (5, 18, 6) {real, imag} */,
  {32'h3d88f802, 32'h3c55ef58} /* (5, 18, 5) {real, imag} */,
  {32'hbe093d40, 32'h3db7884b} /* (5, 18, 4) {real, imag} */,
  {32'hbd85b697, 32'h3e06b288} /* (5, 18, 3) {real, imag} */,
  {32'hbccb931c, 32'hbdc65f19} /* (5, 18, 2) {real, imag} */,
  {32'hbe871ec2, 32'hbcad5516} /* (5, 18, 1) {real, imag} */,
  {32'h3d131c80, 32'h00000000} /* (5, 18, 0) {real, imag} */,
  {32'hbed87e0f, 32'h3bd755a0} /* (5, 17, 31) {real, imag} */,
  {32'h3cd7f229, 32'h3e0e05ea} /* (5, 17, 30) {real, imag} */,
  {32'h3cd00589, 32'h3d2c034e} /* (5, 17, 29) {real, imag} */,
  {32'h3d600416, 32'hbc0c7da4} /* (5, 17, 28) {real, imag} */,
  {32'h3c8a2c08, 32'h3dae17ac} /* (5, 17, 27) {real, imag} */,
  {32'h3b5d54e0, 32'hbdb2a34b} /* (5, 17, 26) {real, imag} */,
  {32'hbd82f3d4, 32'h3d14c586} /* (5, 17, 25) {real, imag} */,
  {32'h3bd31f3c, 32'h3cfd69fc} /* (5, 17, 24) {real, imag} */,
  {32'hbd3a368f, 32'h3d07f064} /* (5, 17, 23) {real, imag} */,
  {32'h3cabe4cc, 32'h3cb1a918} /* (5, 17, 22) {real, imag} */,
  {32'hbd10cbde, 32'hbc3a43c8} /* (5, 17, 21) {real, imag} */,
  {32'h3cb13e88, 32'h3d20feee} /* (5, 17, 20) {real, imag} */,
  {32'h3bb47600, 32'h3d3c0ae1} /* (5, 17, 19) {real, imag} */,
  {32'h3c626b1f, 32'hbbd679a8} /* (5, 17, 18) {real, imag} */,
  {32'hbd5f17b9, 32'hbcff65fd} /* (5, 17, 17) {real, imag} */,
  {32'h3d6f0d12, 32'h00000000} /* (5, 17, 16) {real, imag} */,
  {32'hbd5f17b9, 32'h3cff65fd} /* (5, 17, 15) {real, imag} */,
  {32'h3c626b1f, 32'h3bd679a8} /* (5, 17, 14) {real, imag} */,
  {32'h3bb47600, 32'hbd3c0ae1} /* (5, 17, 13) {real, imag} */,
  {32'h3cb13e88, 32'hbd20feee} /* (5, 17, 12) {real, imag} */,
  {32'hbd10cbde, 32'h3c3a43c8} /* (5, 17, 11) {real, imag} */,
  {32'h3cabe4cc, 32'hbcb1a918} /* (5, 17, 10) {real, imag} */,
  {32'hbd3a368f, 32'hbd07f064} /* (5, 17, 9) {real, imag} */,
  {32'h3bd31f3c, 32'hbcfd69fc} /* (5, 17, 8) {real, imag} */,
  {32'hbd82f3d4, 32'hbd14c586} /* (5, 17, 7) {real, imag} */,
  {32'h3b5d54e0, 32'h3db2a34b} /* (5, 17, 6) {real, imag} */,
  {32'h3c8a2c08, 32'hbdae17ac} /* (5, 17, 5) {real, imag} */,
  {32'h3d600416, 32'h3c0c7da4} /* (5, 17, 4) {real, imag} */,
  {32'h3cd00589, 32'hbd2c034e} /* (5, 17, 3) {real, imag} */,
  {32'h3cd7f229, 32'hbe0e05ea} /* (5, 17, 2) {real, imag} */,
  {32'hbed87e0f, 32'hbbd755a0} /* (5, 17, 1) {real, imag} */,
  {32'hbd851e74, 32'h00000000} /* (5, 17, 0) {real, imag} */,
  {32'hbef9e8eb, 32'hbdcc97d6} /* (5, 16, 31) {real, imag} */,
  {32'hbdc35311, 32'h3dcaddd0} /* (5, 16, 30) {real, imag} */,
  {32'h3d7ef099, 32'hbcb1479c} /* (5, 16, 29) {real, imag} */,
  {32'h3bf916c8, 32'hbdc0cd62} /* (5, 16, 28) {real, imag} */,
  {32'h3de3eee3, 32'h3d20a392} /* (5, 16, 27) {real, imag} */,
  {32'hbcf62a0a, 32'hbaaf1058} /* (5, 16, 26) {real, imag} */,
  {32'h3e2eec83, 32'hbc2ac17e} /* (5, 16, 25) {real, imag} */,
  {32'hbd2210d8, 32'h3d4811f0} /* (5, 16, 24) {real, imag} */,
  {32'h3d683723, 32'hbd26b36a} /* (5, 16, 23) {real, imag} */,
  {32'hbd0030c5, 32'h3da54472} /* (5, 16, 22) {real, imag} */,
  {32'hbd58cfad, 32'hbda0bf86} /* (5, 16, 21) {real, imag} */,
  {32'hbd811e3e, 32'hbc3324af} /* (5, 16, 20) {real, imag} */,
  {32'h3c521868, 32'h3d4fb3cb} /* (5, 16, 19) {real, imag} */,
  {32'hbc3ca89a, 32'h3c4b9364} /* (5, 16, 18) {real, imag} */,
  {32'h3d6301e1, 32'hbd286e2a} /* (5, 16, 17) {real, imag} */,
  {32'hbb9111bc, 32'h00000000} /* (5, 16, 16) {real, imag} */,
  {32'h3d6301e1, 32'h3d286e2a} /* (5, 16, 15) {real, imag} */,
  {32'hbc3ca89a, 32'hbc4b9364} /* (5, 16, 14) {real, imag} */,
  {32'h3c521868, 32'hbd4fb3cb} /* (5, 16, 13) {real, imag} */,
  {32'hbd811e3e, 32'h3c3324af} /* (5, 16, 12) {real, imag} */,
  {32'hbd58cfad, 32'h3da0bf86} /* (5, 16, 11) {real, imag} */,
  {32'hbd0030c5, 32'hbda54472} /* (5, 16, 10) {real, imag} */,
  {32'h3d683723, 32'h3d26b36a} /* (5, 16, 9) {real, imag} */,
  {32'hbd2210d8, 32'hbd4811f0} /* (5, 16, 8) {real, imag} */,
  {32'h3e2eec83, 32'h3c2ac17e} /* (5, 16, 7) {real, imag} */,
  {32'hbcf62a0a, 32'h3aaf1058} /* (5, 16, 6) {real, imag} */,
  {32'h3de3eee3, 32'hbd20a392} /* (5, 16, 5) {real, imag} */,
  {32'h3bf916c8, 32'h3dc0cd62} /* (5, 16, 4) {real, imag} */,
  {32'h3d7ef099, 32'h3cb1479c} /* (5, 16, 3) {real, imag} */,
  {32'hbdc35311, 32'hbdcaddd0} /* (5, 16, 2) {real, imag} */,
  {32'hbef9e8eb, 32'h3dcc97d6} /* (5, 16, 1) {real, imag} */,
  {32'hbe0e7064, 32'h00000000} /* (5, 16, 0) {real, imag} */,
  {32'hbeceea47, 32'hbe6888ef} /* (5, 15, 31) {real, imag} */,
  {32'h3b2b42f8, 32'h3de7da21} /* (5, 15, 30) {real, imag} */,
  {32'h3d3f6adc, 32'hbe693328} /* (5, 15, 29) {real, imag} */,
  {32'h3d8d4ec9, 32'hbca6e0e2} /* (5, 15, 28) {real, imag} */,
  {32'hbcac2662, 32'h3c6a07b0} /* (5, 15, 27) {real, imag} */,
  {32'h3da0ae6b, 32'hbd0e6d96} /* (5, 15, 26) {real, imag} */,
  {32'h3db5019c, 32'h3d71c8a2} /* (5, 15, 25) {real, imag} */,
  {32'h3ab47970, 32'h3b849c78} /* (5, 15, 24) {real, imag} */,
  {32'hbd9f2f7a, 32'h3c12412a} /* (5, 15, 23) {real, imag} */,
  {32'hbc178899, 32'h3d9eb7cb} /* (5, 15, 22) {real, imag} */,
  {32'h3d251f94, 32'hbd82afd5} /* (5, 15, 21) {real, imag} */,
  {32'hbd0d9d71, 32'h3db22f71} /* (5, 15, 20) {real, imag} */,
  {32'hbe113a63, 32'hbd96c4af} /* (5, 15, 19) {real, imag} */,
  {32'h3c0688ab, 32'hbcb7c78e} /* (5, 15, 18) {real, imag} */,
  {32'hbdabbb44, 32'h3d666d12} /* (5, 15, 17) {real, imag} */,
  {32'hbd27d99e, 32'h00000000} /* (5, 15, 16) {real, imag} */,
  {32'hbdabbb44, 32'hbd666d12} /* (5, 15, 15) {real, imag} */,
  {32'h3c0688ab, 32'h3cb7c78e} /* (5, 15, 14) {real, imag} */,
  {32'hbe113a63, 32'h3d96c4af} /* (5, 15, 13) {real, imag} */,
  {32'hbd0d9d71, 32'hbdb22f71} /* (5, 15, 12) {real, imag} */,
  {32'h3d251f94, 32'h3d82afd5} /* (5, 15, 11) {real, imag} */,
  {32'hbc178899, 32'hbd9eb7cb} /* (5, 15, 10) {real, imag} */,
  {32'hbd9f2f7a, 32'hbc12412a} /* (5, 15, 9) {real, imag} */,
  {32'h3ab47970, 32'hbb849c78} /* (5, 15, 8) {real, imag} */,
  {32'h3db5019c, 32'hbd71c8a2} /* (5, 15, 7) {real, imag} */,
  {32'h3da0ae6b, 32'h3d0e6d96} /* (5, 15, 6) {real, imag} */,
  {32'hbcac2662, 32'hbc6a07b0} /* (5, 15, 5) {real, imag} */,
  {32'h3d8d4ec9, 32'h3ca6e0e2} /* (5, 15, 4) {real, imag} */,
  {32'h3d3f6adc, 32'h3e693328} /* (5, 15, 3) {real, imag} */,
  {32'h3b2b42f8, 32'hbde7da21} /* (5, 15, 2) {real, imag} */,
  {32'hbeceea47, 32'h3e6888ef} /* (5, 15, 1) {real, imag} */,
  {32'hbee65a8f, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'hbea66182, 32'hbdbd5c0e} /* (5, 14, 31) {real, imag} */,
  {32'h3d27657e, 32'hbdf14d77} /* (5, 14, 30) {real, imag} */,
  {32'h3da8986d, 32'hbe1b2330} /* (5, 14, 29) {real, imag} */,
  {32'h3c513438, 32'hbddf6273} /* (5, 14, 28) {real, imag} */,
  {32'hbd3c8f1a, 32'h3d92f208} /* (5, 14, 27) {real, imag} */,
  {32'h3d34e47c, 32'hbb07a950} /* (5, 14, 26) {real, imag} */,
  {32'h3d61e8cc, 32'hbd71141a} /* (5, 14, 25) {real, imag} */,
  {32'hbb817610, 32'hbd874403} /* (5, 14, 24) {real, imag} */,
  {32'h3abc9e40, 32'h3dcbbaf2} /* (5, 14, 23) {real, imag} */,
  {32'hbb9c63b6, 32'hbd887c4d} /* (5, 14, 22) {real, imag} */,
  {32'h3db5ed72, 32'h3d9b05dc} /* (5, 14, 21) {real, imag} */,
  {32'h3d312329, 32'h3c029a16} /* (5, 14, 20) {real, imag} */,
  {32'hbd29543e, 32'h3c77dfd4} /* (5, 14, 19) {real, imag} */,
  {32'h3d9c9ab8, 32'h3b1468e0} /* (5, 14, 18) {real, imag} */,
  {32'hbd76454b, 32'hbd0f5ba3} /* (5, 14, 17) {real, imag} */,
  {32'h3d8684cc, 32'h00000000} /* (5, 14, 16) {real, imag} */,
  {32'hbd76454b, 32'h3d0f5ba3} /* (5, 14, 15) {real, imag} */,
  {32'h3d9c9ab8, 32'hbb1468e0} /* (5, 14, 14) {real, imag} */,
  {32'hbd29543e, 32'hbc77dfd4} /* (5, 14, 13) {real, imag} */,
  {32'h3d312329, 32'hbc029a16} /* (5, 14, 12) {real, imag} */,
  {32'h3db5ed72, 32'hbd9b05dc} /* (5, 14, 11) {real, imag} */,
  {32'hbb9c63b6, 32'h3d887c4d} /* (5, 14, 10) {real, imag} */,
  {32'h3abc9e40, 32'hbdcbbaf2} /* (5, 14, 9) {real, imag} */,
  {32'hbb817610, 32'h3d874403} /* (5, 14, 8) {real, imag} */,
  {32'h3d61e8cc, 32'h3d71141a} /* (5, 14, 7) {real, imag} */,
  {32'h3d34e47c, 32'h3b07a950} /* (5, 14, 6) {real, imag} */,
  {32'hbd3c8f1a, 32'hbd92f208} /* (5, 14, 5) {real, imag} */,
  {32'h3c513438, 32'h3ddf6273} /* (5, 14, 4) {real, imag} */,
  {32'h3da8986d, 32'h3e1b2330} /* (5, 14, 3) {real, imag} */,
  {32'h3d27657e, 32'h3df14d77} /* (5, 14, 2) {real, imag} */,
  {32'hbea66182, 32'h3dbd5c0e} /* (5, 14, 1) {real, imag} */,
  {32'hbf21ceac, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hbd901a60, 32'hbe5fbf49} /* (5, 13, 31) {real, imag} */,
  {32'hbca0dd72, 32'hbe6c444d} /* (5, 13, 30) {real, imag} */,
  {32'h3dcf1bd8, 32'hbd232b3a} /* (5, 13, 29) {real, imag} */,
  {32'hbd933a6a, 32'hbe1f59ee} /* (5, 13, 28) {real, imag} */,
  {32'hbdb51ca2, 32'h3e475f9e} /* (5, 13, 27) {real, imag} */,
  {32'h3e454778, 32'h3de56574} /* (5, 13, 26) {real, imag} */,
  {32'h3d608ecf, 32'hbd5435dd} /* (5, 13, 25) {real, imag} */,
  {32'hbda7f81e, 32'h3c8ca934} /* (5, 13, 24) {real, imag} */,
  {32'h3d642a71, 32'h3da6ff7e} /* (5, 13, 23) {real, imag} */,
  {32'h3cb16f6c, 32'hbde3da4c} /* (5, 13, 22) {real, imag} */,
  {32'hbd968342, 32'h3a74c8a0} /* (5, 13, 21) {real, imag} */,
  {32'h3d3f306e, 32'hbbebe530} /* (5, 13, 20) {real, imag} */,
  {32'hbd87c768, 32'hbdc6f4bf} /* (5, 13, 19) {real, imag} */,
  {32'hbd3cfc24, 32'h3d83325e} /* (5, 13, 18) {real, imag} */,
  {32'h3d5556ef, 32'hbd0b89fa} /* (5, 13, 17) {real, imag} */,
  {32'hbc573bd6, 32'h00000000} /* (5, 13, 16) {real, imag} */,
  {32'h3d5556ef, 32'h3d0b89fa} /* (5, 13, 15) {real, imag} */,
  {32'hbd3cfc24, 32'hbd83325e} /* (5, 13, 14) {real, imag} */,
  {32'hbd87c768, 32'h3dc6f4bf} /* (5, 13, 13) {real, imag} */,
  {32'h3d3f306e, 32'h3bebe530} /* (5, 13, 12) {real, imag} */,
  {32'hbd968342, 32'hba74c8a0} /* (5, 13, 11) {real, imag} */,
  {32'h3cb16f6c, 32'h3de3da4c} /* (5, 13, 10) {real, imag} */,
  {32'h3d642a71, 32'hbda6ff7e} /* (5, 13, 9) {real, imag} */,
  {32'hbda7f81e, 32'hbc8ca934} /* (5, 13, 8) {real, imag} */,
  {32'h3d608ecf, 32'h3d5435dd} /* (5, 13, 7) {real, imag} */,
  {32'h3e454778, 32'hbde56574} /* (5, 13, 6) {real, imag} */,
  {32'hbdb51ca2, 32'hbe475f9e} /* (5, 13, 5) {real, imag} */,
  {32'hbd933a6a, 32'h3e1f59ee} /* (5, 13, 4) {real, imag} */,
  {32'h3dcf1bd8, 32'h3d232b3a} /* (5, 13, 3) {real, imag} */,
  {32'hbca0dd72, 32'h3e6c444d} /* (5, 13, 2) {real, imag} */,
  {32'hbd901a60, 32'h3e5fbf49} /* (5, 13, 1) {real, imag} */,
  {32'hbef17ebc, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'h3d881c4e, 32'hbdf32dae} /* (5, 12, 31) {real, imag} */,
  {32'h3e1065e0, 32'hbe05f511} /* (5, 12, 30) {real, imag} */,
  {32'h3e0aa958, 32'h3d86d878} /* (5, 12, 29) {real, imag} */,
  {32'hbd9b5092, 32'hbd0c787e} /* (5, 12, 28) {real, imag} */,
  {32'hbe031fa4, 32'h3df1c2df} /* (5, 12, 27) {real, imag} */,
  {32'h3defbd0e, 32'h3e0b108d} /* (5, 12, 26) {real, imag} */,
  {32'hbdab9f7b, 32'hbc1f0d40} /* (5, 12, 25) {real, imag} */,
  {32'h3d3902d7, 32'h3d89cc2d} /* (5, 12, 24) {real, imag} */,
  {32'h3d39087b, 32'hbb832910} /* (5, 12, 23) {real, imag} */,
  {32'hbd4e4b25, 32'hbd7894bf} /* (5, 12, 22) {real, imag} */,
  {32'hbc55b2c4, 32'h3a1b7700} /* (5, 12, 21) {real, imag} */,
  {32'hbcb730d8, 32'hbdb77e05} /* (5, 12, 20) {real, imag} */,
  {32'h3cab4548, 32'h3d98a5d8} /* (5, 12, 19) {real, imag} */,
  {32'h39727280, 32'hbce2ef62} /* (5, 12, 18) {real, imag} */,
  {32'hbc0f014e, 32'hbd9572ba} /* (5, 12, 17) {real, imag} */,
  {32'hbdb11d75, 32'h00000000} /* (5, 12, 16) {real, imag} */,
  {32'hbc0f014e, 32'h3d9572ba} /* (5, 12, 15) {real, imag} */,
  {32'h39727280, 32'h3ce2ef62} /* (5, 12, 14) {real, imag} */,
  {32'h3cab4548, 32'hbd98a5d8} /* (5, 12, 13) {real, imag} */,
  {32'hbcb730d8, 32'h3db77e05} /* (5, 12, 12) {real, imag} */,
  {32'hbc55b2c4, 32'hba1b7700} /* (5, 12, 11) {real, imag} */,
  {32'hbd4e4b25, 32'h3d7894bf} /* (5, 12, 10) {real, imag} */,
  {32'h3d39087b, 32'h3b832910} /* (5, 12, 9) {real, imag} */,
  {32'h3d3902d7, 32'hbd89cc2d} /* (5, 12, 8) {real, imag} */,
  {32'hbdab9f7b, 32'h3c1f0d40} /* (5, 12, 7) {real, imag} */,
  {32'h3defbd0e, 32'hbe0b108d} /* (5, 12, 6) {real, imag} */,
  {32'hbe031fa4, 32'hbdf1c2df} /* (5, 12, 5) {real, imag} */,
  {32'hbd9b5092, 32'h3d0c787e} /* (5, 12, 4) {real, imag} */,
  {32'h3e0aa958, 32'hbd86d878} /* (5, 12, 3) {real, imag} */,
  {32'h3e1065e0, 32'h3e05f511} /* (5, 12, 2) {real, imag} */,
  {32'h3d881c4e, 32'h3df32dae} /* (5, 12, 1) {real, imag} */,
  {32'hbe123ac4, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h3e1e4923, 32'hbe9c77f6} /* (5, 11, 31) {real, imag} */,
  {32'h3d996248, 32'hbd5b77be} /* (5, 11, 30) {real, imag} */,
  {32'h3e49dc36, 32'h3d0599f6} /* (5, 11, 29) {real, imag} */,
  {32'h3d66896b, 32'hbd84e717} /* (5, 11, 28) {real, imag} */,
  {32'hbd06f428, 32'h3dcd19ac} /* (5, 11, 27) {real, imag} */,
  {32'h3e1c1a94, 32'h3bd91450} /* (5, 11, 26) {real, imag} */,
  {32'hbbba8b98, 32'h3d10dc32} /* (5, 11, 25) {real, imag} */,
  {32'h3c42ce88, 32'h3d37888c} /* (5, 11, 24) {real, imag} */,
  {32'h3e04636e, 32'h3db0f99a} /* (5, 11, 23) {real, imag} */,
  {32'hbd664bba, 32'h3d3677e2} /* (5, 11, 22) {real, imag} */,
  {32'hbdb3b7e0, 32'h3daeffb1} /* (5, 11, 21) {real, imag} */,
  {32'hbe00a5a5, 32'h3da3e6d5} /* (5, 11, 20) {real, imag} */,
  {32'h3d0c3067, 32'h3d6af91f} /* (5, 11, 19) {real, imag} */,
  {32'h3d6eef92, 32'hbc94815e} /* (5, 11, 18) {real, imag} */,
  {32'hbdb3a710, 32'h3d22d4de} /* (5, 11, 17) {real, imag} */,
  {32'h3dc901f6, 32'h00000000} /* (5, 11, 16) {real, imag} */,
  {32'hbdb3a710, 32'hbd22d4de} /* (5, 11, 15) {real, imag} */,
  {32'h3d6eef92, 32'h3c94815e} /* (5, 11, 14) {real, imag} */,
  {32'h3d0c3067, 32'hbd6af91f} /* (5, 11, 13) {real, imag} */,
  {32'hbe00a5a5, 32'hbda3e6d5} /* (5, 11, 12) {real, imag} */,
  {32'hbdb3b7e0, 32'hbdaeffb1} /* (5, 11, 11) {real, imag} */,
  {32'hbd664bba, 32'hbd3677e2} /* (5, 11, 10) {real, imag} */,
  {32'h3e04636e, 32'hbdb0f99a} /* (5, 11, 9) {real, imag} */,
  {32'h3c42ce88, 32'hbd37888c} /* (5, 11, 8) {real, imag} */,
  {32'hbbba8b98, 32'hbd10dc32} /* (5, 11, 7) {real, imag} */,
  {32'h3e1c1a94, 32'hbbd91450} /* (5, 11, 6) {real, imag} */,
  {32'hbd06f428, 32'hbdcd19ac} /* (5, 11, 5) {real, imag} */,
  {32'h3d66896b, 32'h3d84e717} /* (5, 11, 4) {real, imag} */,
  {32'h3e49dc36, 32'hbd0599f6} /* (5, 11, 3) {real, imag} */,
  {32'h3d996248, 32'h3d5b77be} /* (5, 11, 2) {real, imag} */,
  {32'h3e1e4923, 32'h3e9c77f6} /* (5, 11, 1) {real, imag} */,
  {32'h3e46d0ba, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'h3dcc1dd5, 32'hbebec316} /* (5, 10, 31) {real, imag} */,
  {32'h3de91543, 32'hbd281a5c} /* (5, 10, 30) {real, imag} */,
  {32'h3d96e0c6, 32'hbc9c2220} /* (5, 10, 29) {real, imag} */,
  {32'h3d433f74, 32'hbdbc8f7a} /* (5, 10, 28) {real, imag} */,
  {32'hbc9c3374, 32'h3ba38f78} /* (5, 10, 27) {real, imag} */,
  {32'hbd30ca1b, 32'hbc6f7cd0} /* (5, 10, 26) {real, imag} */,
  {32'h3c1348c6, 32'hbc323106} /* (5, 10, 25) {real, imag} */,
  {32'h3cb7748e, 32'hbe6bdb65} /* (5, 10, 24) {real, imag} */,
  {32'hbd6b5da0, 32'h3e4d1d0a} /* (5, 10, 23) {real, imag} */,
  {32'h3d97edf5, 32'h3dffbe9e} /* (5, 10, 22) {real, imag} */,
  {32'hbd1b9e13, 32'hbdf5f6d4} /* (5, 10, 21) {real, imag} */,
  {32'h3dac785e, 32'h3d6f292a} /* (5, 10, 20) {real, imag} */,
  {32'h3d54f9d8, 32'h3ca8b8da} /* (5, 10, 19) {real, imag} */,
  {32'hbd16eaec, 32'h3d854518} /* (5, 10, 18) {real, imag} */,
  {32'hbc07432f, 32'h3d349178} /* (5, 10, 17) {real, imag} */,
  {32'hbd7682f4, 32'h00000000} /* (5, 10, 16) {real, imag} */,
  {32'hbc07432f, 32'hbd349178} /* (5, 10, 15) {real, imag} */,
  {32'hbd16eaec, 32'hbd854518} /* (5, 10, 14) {real, imag} */,
  {32'h3d54f9d8, 32'hbca8b8da} /* (5, 10, 13) {real, imag} */,
  {32'h3dac785e, 32'hbd6f292a} /* (5, 10, 12) {real, imag} */,
  {32'hbd1b9e13, 32'h3df5f6d4} /* (5, 10, 11) {real, imag} */,
  {32'h3d97edf5, 32'hbdffbe9e} /* (5, 10, 10) {real, imag} */,
  {32'hbd6b5da0, 32'hbe4d1d0a} /* (5, 10, 9) {real, imag} */,
  {32'h3cb7748e, 32'h3e6bdb65} /* (5, 10, 8) {real, imag} */,
  {32'h3c1348c6, 32'h3c323106} /* (5, 10, 7) {real, imag} */,
  {32'hbd30ca1b, 32'h3c6f7cd0} /* (5, 10, 6) {real, imag} */,
  {32'hbc9c3374, 32'hbba38f78} /* (5, 10, 5) {real, imag} */,
  {32'h3d433f74, 32'h3dbc8f7a} /* (5, 10, 4) {real, imag} */,
  {32'h3d96e0c6, 32'h3c9c2220} /* (5, 10, 3) {real, imag} */,
  {32'h3de91543, 32'h3d281a5c} /* (5, 10, 2) {real, imag} */,
  {32'h3dcc1dd5, 32'h3ebec316} /* (5, 10, 1) {real, imag} */,
  {32'h3ea5b66c, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'h3d9e4805, 32'hbea6c253} /* (5, 9, 31) {real, imag} */,
  {32'h3dbe638d, 32'h3d1b2260} /* (5, 9, 30) {real, imag} */,
  {32'h3d79f48e, 32'h3cafd17e} /* (5, 9, 29) {real, imag} */,
  {32'h3d38a1ec, 32'hbc953085} /* (5, 9, 28) {real, imag} */,
  {32'hbcf382d9, 32'hbd0c950d} /* (5, 9, 27) {real, imag} */,
  {32'h3e02140a, 32'h3d3ed4e4} /* (5, 9, 26) {real, imag} */,
  {32'hbd23472e, 32'h3cf1555a} /* (5, 9, 25) {real, imag} */,
  {32'h3d332f1a, 32'hbda7078a} /* (5, 9, 24) {real, imag} */,
  {32'h3c0de37a, 32'h3d86fa36} /* (5, 9, 23) {real, imag} */,
  {32'h3de71e5d, 32'hbca19a8b} /* (5, 9, 22) {real, imag} */,
  {32'h3cd57e22, 32'h3bc18110} /* (5, 9, 21) {real, imag} */,
  {32'hbdc18fc9, 32'hbce96618} /* (5, 9, 20) {real, imag} */,
  {32'hbd54d48d, 32'h3d697bdc} /* (5, 9, 19) {real, imag} */,
  {32'h3d3c0333, 32'hbd5f5362} /* (5, 9, 18) {real, imag} */,
  {32'h3d0b3909, 32'h3d577b66} /* (5, 9, 17) {real, imag} */,
  {32'hbda3cc98, 32'h00000000} /* (5, 9, 16) {real, imag} */,
  {32'h3d0b3909, 32'hbd577b66} /* (5, 9, 15) {real, imag} */,
  {32'h3d3c0333, 32'h3d5f5362} /* (5, 9, 14) {real, imag} */,
  {32'hbd54d48d, 32'hbd697bdc} /* (5, 9, 13) {real, imag} */,
  {32'hbdc18fc9, 32'h3ce96618} /* (5, 9, 12) {real, imag} */,
  {32'h3cd57e22, 32'hbbc18110} /* (5, 9, 11) {real, imag} */,
  {32'h3de71e5d, 32'h3ca19a8b} /* (5, 9, 10) {real, imag} */,
  {32'h3c0de37a, 32'hbd86fa36} /* (5, 9, 9) {real, imag} */,
  {32'h3d332f1a, 32'h3da7078a} /* (5, 9, 8) {real, imag} */,
  {32'hbd23472e, 32'hbcf1555a} /* (5, 9, 7) {real, imag} */,
  {32'h3e02140a, 32'hbd3ed4e4} /* (5, 9, 6) {real, imag} */,
  {32'hbcf382d9, 32'h3d0c950d} /* (5, 9, 5) {real, imag} */,
  {32'h3d38a1ec, 32'h3c953085} /* (5, 9, 4) {real, imag} */,
  {32'h3d79f48e, 32'hbcafd17e} /* (5, 9, 3) {real, imag} */,
  {32'h3dbe638d, 32'hbd1b2260} /* (5, 9, 2) {real, imag} */,
  {32'h3d9e4805, 32'h3ea6c253} /* (5, 9, 1) {real, imag} */,
  {32'h3f2c0ed7, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'h3e281039, 32'hbeccec91} /* (5, 8, 31) {real, imag} */,
  {32'h3e1e2e54, 32'h3e93dd65} /* (5, 8, 30) {real, imag} */,
  {32'h3e598d04, 32'hbdd0d8be} /* (5, 8, 29) {real, imag} */,
  {32'h3d8f4622, 32'h3d6ef0dc} /* (5, 8, 28) {real, imag} */,
  {32'hbd97f78d, 32'hbc6f8574} /* (5, 8, 27) {real, imag} */,
  {32'h3d323977, 32'h3d15c822} /* (5, 8, 26) {real, imag} */,
  {32'hbd360250, 32'h3d6f3d3e} /* (5, 8, 25) {real, imag} */,
  {32'h3ca9e1ba, 32'hbe0f8c8f} /* (5, 8, 24) {real, imag} */,
  {32'h3d0e2ab9, 32'h3c958d5c} /* (5, 8, 23) {real, imag} */,
  {32'hbdc11280, 32'h3db43374} /* (5, 8, 22) {real, imag} */,
  {32'h3dda8d51, 32'h3baee4bc} /* (5, 8, 21) {real, imag} */,
  {32'h3cb52bf0, 32'hbd46b73c} /* (5, 8, 20) {real, imag} */,
  {32'hbd260b85, 32'hbd05b1f8} /* (5, 8, 19) {real, imag} */,
  {32'hbd9d990a, 32'hbb2925d0} /* (5, 8, 18) {real, imag} */,
  {32'hbc693063, 32'hbc6667f6} /* (5, 8, 17) {real, imag} */,
  {32'hbd8d6063, 32'h00000000} /* (5, 8, 16) {real, imag} */,
  {32'hbc693063, 32'h3c6667f6} /* (5, 8, 15) {real, imag} */,
  {32'hbd9d990a, 32'h3b2925d0} /* (5, 8, 14) {real, imag} */,
  {32'hbd260b85, 32'h3d05b1f8} /* (5, 8, 13) {real, imag} */,
  {32'h3cb52bf0, 32'h3d46b73c} /* (5, 8, 12) {real, imag} */,
  {32'h3dda8d51, 32'hbbaee4bc} /* (5, 8, 11) {real, imag} */,
  {32'hbdc11280, 32'hbdb43374} /* (5, 8, 10) {real, imag} */,
  {32'h3d0e2ab9, 32'hbc958d5c} /* (5, 8, 9) {real, imag} */,
  {32'h3ca9e1ba, 32'h3e0f8c8f} /* (5, 8, 8) {real, imag} */,
  {32'hbd360250, 32'hbd6f3d3e} /* (5, 8, 7) {real, imag} */,
  {32'h3d323977, 32'hbd15c822} /* (5, 8, 6) {real, imag} */,
  {32'hbd97f78d, 32'h3c6f8574} /* (5, 8, 5) {real, imag} */,
  {32'h3d8f4622, 32'hbd6ef0dc} /* (5, 8, 4) {real, imag} */,
  {32'h3e598d04, 32'h3dd0d8be} /* (5, 8, 3) {real, imag} */,
  {32'h3e1e2e54, 32'hbe93dd65} /* (5, 8, 2) {real, imag} */,
  {32'h3e281039, 32'h3eccec91} /* (5, 8, 1) {real, imag} */,
  {32'h3f5a4c22, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'h3ea1046c, 32'hbecfb300} /* (5, 7, 31) {real, imag} */,
  {32'h3e32d838, 32'h3ec46604} /* (5, 7, 30) {real, imag} */,
  {32'h3e71cb39, 32'hbe25ae0a} /* (5, 7, 29) {real, imag} */,
  {32'h3d09d944, 32'h3dd9b7b8} /* (5, 7, 28) {real, imag} */,
  {32'hbdc0b510, 32'h3d099a7e} /* (5, 7, 27) {real, imag} */,
  {32'h3d2b782c, 32'h3e26ae66} /* (5, 7, 26) {real, imag} */,
  {32'hbdfa46b7, 32'hbdee0b30} /* (5, 7, 25) {real, imag} */,
  {32'h3d050f72, 32'hbe43c275} /* (5, 7, 24) {real, imag} */,
  {32'hbe0525f4, 32'h3df47cae} /* (5, 7, 23) {real, imag} */,
  {32'h3a00a1d0, 32'h3d3dc0d6} /* (5, 7, 22) {real, imag} */,
  {32'h3d0cab12, 32'hbe334542} /* (5, 7, 21) {real, imag} */,
  {32'hbdb0baad, 32'hbe0fff2d} /* (5, 7, 20) {real, imag} */,
  {32'h3c9a289e, 32'h3bee46b4} /* (5, 7, 19) {real, imag} */,
  {32'h3ca2f01c, 32'hbd1f7c1e} /* (5, 7, 18) {real, imag} */,
  {32'hbc18f62c, 32'h3d76c855} /* (5, 7, 17) {real, imag} */,
  {32'h3cf4e6e8, 32'h00000000} /* (5, 7, 16) {real, imag} */,
  {32'hbc18f62c, 32'hbd76c855} /* (5, 7, 15) {real, imag} */,
  {32'h3ca2f01c, 32'h3d1f7c1e} /* (5, 7, 14) {real, imag} */,
  {32'h3c9a289e, 32'hbbee46b4} /* (5, 7, 13) {real, imag} */,
  {32'hbdb0baad, 32'h3e0fff2d} /* (5, 7, 12) {real, imag} */,
  {32'h3d0cab12, 32'h3e334542} /* (5, 7, 11) {real, imag} */,
  {32'h3a00a1d0, 32'hbd3dc0d6} /* (5, 7, 10) {real, imag} */,
  {32'hbe0525f4, 32'hbdf47cae} /* (5, 7, 9) {real, imag} */,
  {32'h3d050f72, 32'h3e43c275} /* (5, 7, 8) {real, imag} */,
  {32'hbdfa46b7, 32'h3dee0b30} /* (5, 7, 7) {real, imag} */,
  {32'h3d2b782c, 32'hbe26ae66} /* (5, 7, 6) {real, imag} */,
  {32'hbdc0b510, 32'hbd099a7e} /* (5, 7, 5) {real, imag} */,
  {32'h3d09d944, 32'hbdd9b7b8} /* (5, 7, 4) {real, imag} */,
  {32'h3e71cb39, 32'h3e25ae0a} /* (5, 7, 3) {real, imag} */,
  {32'h3e32d838, 32'hbec46604} /* (5, 7, 2) {real, imag} */,
  {32'h3ea1046c, 32'h3ecfb300} /* (5, 7, 1) {real, imag} */,
  {32'h3f8a2d7f, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'h3ee8ee86, 32'hbeb65ccc} /* (5, 6, 31) {real, imag} */,
  {32'hbd9a4d72, 32'h3e8d7caa} /* (5, 6, 30) {real, imag} */,
  {32'h3e4ea4f6, 32'h3d01ff35} /* (5, 6, 29) {real, imag} */,
  {32'h3d8108cf, 32'hbc189688} /* (5, 6, 28) {real, imag} */,
  {32'hbd078244, 32'hbcce49f8} /* (5, 6, 27) {real, imag} */,
  {32'h3d348035, 32'hbc474846} /* (5, 6, 26) {real, imag} */,
  {32'h3d2e1a76, 32'hbd8fc9a2} /* (5, 6, 25) {real, imag} */,
  {32'hbda613ce, 32'hbc3f71e0} /* (5, 6, 24) {real, imag} */,
  {32'hbd0afbd6, 32'h3c95daa4} /* (5, 6, 23) {real, imag} */,
  {32'hbd689792, 32'hbbd77590} /* (5, 6, 22) {real, imag} */,
  {32'hbd9232aa, 32'hbd86c9f2} /* (5, 6, 21) {real, imag} */,
  {32'h3d31a2f4, 32'h3dd8137c} /* (5, 6, 20) {real, imag} */,
  {32'h3adf67d0, 32'h3d62d0f0} /* (5, 6, 19) {real, imag} */,
  {32'h3dd567ed, 32'hbb46faa8} /* (5, 6, 18) {real, imag} */,
  {32'h3c93ac60, 32'h3c538f5d} /* (5, 6, 17) {real, imag} */,
  {32'h3d4795ae, 32'h00000000} /* (5, 6, 16) {real, imag} */,
  {32'h3c93ac60, 32'hbc538f5d} /* (5, 6, 15) {real, imag} */,
  {32'h3dd567ed, 32'h3b46faa8} /* (5, 6, 14) {real, imag} */,
  {32'h3adf67d0, 32'hbd62d0f0} /* (5, 6, 13) {real, imag} */,
  {32'h3d31a2f4, 32'hbdd8137c} /* (5, 6, 12) {real, imag} */,
  {32'hbd9232aa, 32'h3d86c9f2} /* (5, 6, 11) {real, imag} */,
  {32'hbd689792, 32'h3bd77590} /* (5, 6, 10) {real, imag} */,
  {32'hbd0afbd6, 32'hbc95daa4} /* (5, 6, 9) {real, imag} */,
  {32'hbda613ce, 32'h3c3f71e0} /* (5, 6, 8) {real, imag} */,
  {32'h3d2e1a76, 32'h3d8fc9a2} /* (5, 6, 7) {real, imag} */,
  {32'h3d348035, 32'h3c474846} /* (5, 6, 6) {real, imag} */,
  {32'hbd078244, 32'h3cce49f8} /* (5, 6, 5) {real, imag} */,
  {32'h3d8108cf, 32'h3c189688} /* (5, 6, 4) {real, imag} */,
  {32'h3e4ea4f6, 32'hbd01ff35} /* (5, 6, 3) {real, imag} */,
  {32'hbd9a4d72, 32'hbe8d7caa} /* (5, 6, 2) {real, imag} */,
  {32'h3ee8ee86, 32'h3eb65ccc} /* (5, 6, 1) {real, imag} */,
  {32'h3fb265d8, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'h3f3acd81, 32'hbeb0eedc} /* (5, 5, 31) {real, imag} */,
  {32'hbd85272c, 32'h3e569a33} /* (5, 5, 30) {real, imag} */,
  {32'h3dc2e145, 32'h3dd6434f} /* (5, 5, 29) {real, imag} */,
  {32'h3cadfdf2, 32'hbdeecb6b} /* (5, 5, 28) {real, imag} */,
  {32'hbc44de98, 32'hbd317c31} /* (5, 5, 27) {real, imag} */,
  {32'h3d58f4a7, 32'hbd7a97ba} /* (5, 5, 26) {real, imag} */,
  {32'h3d831162, 32'hbdcd2ba9} /* (5, 5, 25) {real, imag} */,
  {32'hbda240aa, 32'hbd361174} /* (5, 5, 24) {real, imag} */,
  {32'hbccb17c6, 32'h3d89576d} /* (5, 5, 23) {real, imag} */,
  {32'hbda04a15, 32'h3bacec5c} /* (5, 5, 22) {real, imag} */,
  {32'h3ca386cc, 32'h3d922ee0} /* (5, 5, 21) {real, imag} */,
  {32'h3d7a0fba, 32'hbdbcb1a3} /* (5, 5, 20) {real, imag} */,
  {32'h3d17d27b, 32'hbd36b9ec} /* (5, 5, 19) {real, imag} */,
  {32'h3c29a0d7, 32'h3dc783a8} /* (5, 5, 18) {real, imag} */,
  {32'hbde34a46, 32'hbca6f17a} /* (5, 5, 17) {real, imag} */,
  {32'h3ce21306, 32'h00000000} /* (5, 5, 16) {real, imag} */,
  {32'hbde34a46, 32'h3ca6f17a} /* (5, 5, 15) {real, imag} */,
  {32'h3c29a0d7, 32'hbdc783a8} /* (5, 5, 14) {real, imag} */,
  {32'h3d17d27b, 32'h3d36b9ec} /* (5, 5, 13) {real, imag} */,
  {32'h3d7a0fba, 32'h3dbcb1a3} /* (5, 5, 12) {real, imag} */,
  {32'h3ca386cc, 32'hbd922ee0} /* (5, 5, 11) {real, imag} */,
  {32'hbda04a15, 32'hbbacec5c} /* (5, 5, 10) {real, imag} */,
  {32'hbccb17c6, 32'hbd89576d} /* (5, 5, 9) {real, imag} */,
  {32'hbda240aa, 32'h3d361174} /* (5, 5, 8) {real, imag} */,
  {32'h3d831162, 32'h3dcd2ba9} /* (5, 5, 7) {real, imag} */,
  {32'h3d58f4a7, 32'h3d7a97ba} /* (5, 5, 6) {real, imag} */,
  {32'hbc44de98, 32'h3d317c31} /* (5, 5, 5) {real, imag} */,
  {32'h3cadfdf2, 32'h3deecb6b} /* (5, 5, 4) {real, imag} */,
  {32'h3dc2e145, 32'hbdd6434f} /* (5, 5, 3) {real, imag} */,
  {32'hbd85272c, 32'hbe569a33} /* (5, 5, 2) {real, imag} */,
  {32'h3f3acd81, 32'h3eb0eedc} /* (5, 5, 1) {real, imag} */,
  {32'h3fbadec0, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'h3f4de130, 32'hbed070e6} /* (5, 4, 31) {real, imag} */,
  {32'hbdaeb34f, 32'h3e5c89ca} /* (5, 4, 30) {real, imag} */,
  {32'h3dfa4546, 32'h3d0fd9f4} /* (5, 4, 29) {real, imag} */,
  {32'h3d876352, 32'hbd9157c5} /* (5, 4, 28) {real, imag} */,
  {32'h3d5d3d18, 32'hbc290778} /* (5, 4, 27) {real, imag} */,
  {32'h3dd80742, 32'h3d36f9fa} /* (5, 4, 26) {real, imag} */,
  {32'h3d4be568, 32'hbcaa6278} /* (5, 4, 25) {real, imag} */,
  {32'hbc8b9ed6, 32'h3d113e32} /* (5, 4, 24) {real, imag} */,
  {32'hbd85de98, 32'hbcb5bd50} /* (5, 4, 23) {real, imag} */,
  {32'h3d764984, 32'h3d8f489c} /* (5, 4, 22) {real, imag} */,
  {32'h3c8f3fea, 32'hbcd878a4} /* (5, 4, 21) {real, imag} */,
  {32'hbd63a36c, 32'h3d48f64e} /* (5, 4, 20) {real, imag} */,
  {32'h3c5ed97e, 32'hbc58aacc} /* (5, 4, 19) {real, imag} */,
  {32'h3d521bc7, 32'hbc9dd985} /* (5, 4, 18) {real, imag} */,
  {32'hbc4cfb90, 32'hbc46690c} /* (5, 4, 17) {real, imag} */,
  {32'h3d55d5ba, 32'h00000000} /* (5, 4, 16) {real, imag} */,
  {32'hbc4cfb90, 32'h3c46690c} /* (5, 4, 15) {real, imag} */,
  {32'h3d521bc7, 32'h3c9dd985} /* (5, 4, 14) {real, imag} */,
  {32'h3c5ed97e, 32'h3c58aacc} /* (5, 4, 13) {real, imag} */,
  {32'hbd63a36c, 32'hbd48f64e} /* (5, 4, 12) {real, imag} */,
  {32'h3c8f3fea, 32'h3cd878a4} /* (5, 4, 11) {real, imag} */,
  {32'h3d764984, 32'hbd8f489c} /* (5, 4, 10) {real, imag} */,
  {32'hbd85de98, 32'h3cb5bd50} /* (5, 4, 9) {real, imag} */,
  {32'hbc8b9ed6, 32'hbd113e32} /* (5, 4, 8) {real, imag} */,
  {32'h3d4be568, 32'h3caa6278} /* (5, 4, 7) {real, imag} */,
  {32'h3dd80742, 32'hbd36f9fa} /* (5, 4, 6) {real, imag} */,
  {32'h3d5d3d18, 32'h3c290778} /* (5, 4, 5) {real, imag} */,
  {32'h3d876352, 32'h3d9157c5} /* (5, 4, 4) {real, imag} */,
  {32'h3dfa4546, 32'hbd0fd9f4} /* (5, 4, 3) {real, imag} */,
  {32'hbdaeb34f, 32'hbe5c89ca} /* (5, 4, 2) {real, imag} */,
  {32'h3f4de130, 32'h3ed070e6} /* (5, 4, 1) {real, imag} */,
  {32'h3fba11ba, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'h3f3d98f0, 32'hbf0df1a6} /* (5, 3, 31) {real, imag} */,
  {32'hbd760c8e, 32'h3de0c55c} /* (5, 3, 30) {real, imag} */,
  {32'h3e016db9, 32'h3c98a780} /* (5, 3, 29) {real, imag} */,
  {32'h3ccdbb18, 32'h3c11d790} /* (5, 3, 28) {real, imag} */,
  {32'h3def017e, 32'h3b7e9a60} /* (5, 3, 27) {real, imag} */,
  {32'h3d212f0a, 32'hbd9ed2e6} /* (5, 3, 26) {real, imag} */,
  {32'h3cb168b2, 32'hbcc2fc12} /* (5, 3, 25) {real, imag} */,
  {32'h3ca27bb0, 32'h3d657d57} /* (5, 3, 24) {real, imag} */,
  {32'h3dca41cc, 32'h3d633664} /* (5, 3, 23) {real, imag} */,
  {32'h3ce63d28, 32'h3dd5faea} /* (5, 3, 22) {real, imag} */,
  {32'hbc2837a8, 32'h3c6e27a6} /* (5, 3, 21) {real, imag} */,
  {32'hbdaaff99, 32'h3db7c2d6} /* (5, 3, 20) {real, imag} */,
  {32'h3d9d9c62, 32'hbcc1fdaa} /* (5, 3, 19) {real, imag} */,
  {32'h3d254693, 32'hbd41c987} /* (5, 3, 18) {real, imag} */,
  {32'h3d13b1fa, 32'hbca2796e} /* (5, 3, 17) {real, imag} */,
  {32'hbcebcfa5, 32'h00000000} /* (5, 3, 16) {real, imag} */,
  {32'h3d13b1fa, 32'h3ca2796e} /* (5, 3, 15) {real, imag} */,
  {32'h3d254693, 32'h3d41c987} /* (5, 3, 14) {real, imag} */,
  {32'h3d9d9c62, 32'h3cc1fdaa} /* (5, 3, 13) {real, imag} */,
  {32'hbdaaff99, 32'hbdb7c2d6} /* (5, 3, 12) {real, imag} */,
  {32'hbc2837a8, 32'hbc6e27a6} /* (5, 3, 11) {real, imag} */,
  {32'h3ce63d28, 32'hbdd5faea} /* (5, 3, 10) {real, imag} */,
  {32'h3dca41cc, 32'hbd633664} /* (5, 3, 9) {real, imag} */,
  {32'h3ca27bb0, 32'hbd657d57} /* (5, 3, 8) {real, imag} */,
  {32'h3cb168b2, 32'h3cc2fc12} /* (5, 3, 7) {real, imag} */,
  {32'h3d212f0a, 32'h3d9ed2e6} /* (5, 3, 6) {real, imag} */,
  {32'h3def017e, 32'hbb7e9a60} /* (5, 3, 5) {real, imag} */,
  {32'h3ccdbb18, 32'hbc11d790} /* (5, 3, 4) {real, imag} */,
  {32'h3e016db9, 32'hbc98a780} /* (5, 3, 3) {real, imag} */,
  {32'hbd760c8e, 32'hbde0c55c} /* (5, 3, 2) {real, imag} */,
  {32'h3f3d98f0, 32'h3f0df1a6} /* (5, 3, 1) {real, imag} */,
  {32'h3fcae2c5, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'h3f3510cd, 32'hbf03ee29} /* (5, 2, 31) {real, imag} */,
  {32'hbc144cc8, 32'hbcd9fa8e} /* (5, 2, 30) {real, imag} */,
  {32'h3dd9adba, 32'h3d4ae05d} /* (5, 2, 29) {real, imag} */,
  {32'h3d125e2e, 32'hbdb58bb0} /* (5, 2, 28) {real, imag} */,
  {32'h3d77e9f9, 32'h3b1a2360} /* (5, 2, 27) {real, imag} */,
  {32'hbba57e14, 32'hbd2621fa} /* (5, 2, 26) {real, imag} */,
  {32'hbe149383, 32'hbda2afdf} /* (5, 2, 25) {real, imag} */,
  {32'hbd340a56, 32'hbd069033} /* (5, 2, 24) {real, imag} */,
  {32'hbd8e1727, 32'h3d41c4e8} /* (5, 2, 23) {real, imag} */,
  {32'hbd83b5d3, 32'hbd994ff9} /* (5, 2, 22) {real, imag} */,
  {32'h3bbe91f0, 32'h3d96cb9d} /* (5, 2, 21) {real, imag} */,
  {32'h3cadb6c9, 32'hbbc77b54} /* (5, 2, 20) {real, imag} */,
  {32'hbcadb9ec, 32'hbd095f72} /* (5, 2, 19) {real, imag} */,
  {32'hbcc3b983, 32'hbd41b902} /* (5, 2, 18) {real, imag} */,
  {32'h3c23fac3, 32'h3d99dc32} /* (5, 2, 17) {real, imag} */,
  {32'hbcc7ac14, 32'h00000000} /* (5, 2, 16) {real, imag} */,
  {32'h3c23fac3, 32'hbd99dc32} /* (5, 2, 15) {real, imag} */,
  {32'hbcc3b983, 32'h3d41b902} /* (5, 2, 14) {real, imag} */,
  {32'hbcadb9ec, 32'h3d095f72} /* (5, 2, 13) {real, imag} */,
  {32'h3cadb6c9, 32'h3bc77b54} /* (5, 2, 12) {real, imag} */,
  {32'h3bbe91f0, 32'hbd96cb9d} /* (5, 2, 11) {real, imag} */,
  {32'hbd83b5d3, 32'h3d994ff9} /* (5, 2, 10) {real, imag} */,
  {32'hbd8e1727, 32'hbd41c4e8} /* (5, 2, 9) {real, imag} */,
  {32'hbd340a56, 32'h3d069033} /* (5, 2, 8) {real, imag} */,
  {32'hbe149383, 32'h3da2afdf} /* (5, 2, 7) {real, imag} */,
  {32'hbba57e14, 32'h3d2621fa} /* (5, 2, 6) {real, imag} */,
  {32'h3d77e9f9, 32'hbb1a2360} /* (5, 2, 5) {real, imag} */,
  {32'h3d125e2e, 32'h3db58bb0} /* (5, 2, 4) {real, imag} */,
  {32'h3dd9adba, 32'hbd4ae05d} /* (5, 2, 3) {real, imag} */,
  {32'hbc144cc8, 32'h3cd9fa8e} /* (5, 2, 2) {real, imag} */,
  {32'h3f3510cd, 32'h3f03ee29} /* (5, 2, 1) {real, imag} */,
  {32'h3fe66f2d, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'h3f47ae08, 32'hbecff9b3} /* (5, 1, 31) {real, imag} */,
  {32'hbd2687e8, 32'hbe2823a8} /* (5, 1, 30) {real, imag} */,
  {32'h3de3e257, 32'hbc3059b8} /* (5, 1, 29) {real, imag} */,
  {32'h3db95bb3, 32'hbe0098bb} /* (5, 1, 28) {real, imag} */,
  {32'hbdc577b0, 32'h3d12f376} /* (5, 1, 27) {real, imag} */,
  {32'hbd4932c2, 32'hbc80c422} /* (5, 1, 26) {real, imag} */,
  {32'hbd4dee94, 32'h3e324262} /* (5, 1, 25) {real, imag} */,
  {32'h3de23ebe, 32'hbdddcae6} /* (5, 1, 24) {real, imag} */,
  {32'hbcc486f9, 32'hbcf03f2a} /* (5, 1, 23) {real, imag} */,
  {32'hbc0db809, 32'h3d14cb33} /* (5, 1, 22) {real, imag} */,
  {32'hbca2ff4a, 32'h3c1d2e88} /* (5, 1, 21) {real, imag} */,
  {32'h3d40ed93, 32'h3cba28e3} /* (5, 1, 20) {real, imag} */,
  {32'hbdbf42ec, 32'hbd2760bc} /* (5, 1, 19) {real, imag} */,
  {32'h3cd94afa, 32'hbc322920} /* (5, 1, 18) {real, imag} */,
  {32'h39cf1e80, 32'hbd298f90} /* (5, 1, 17) {real, imag} */,
  {32'hba1db480, 32'h00000000} /* (5, 1, 16) {real, imag} */,
  {32'h39cf1e80, 32'h3d298f90} /* (5, 1, 15) {real, imag} */,
  {32'h3cd94afa, 32'h3c322920} /* (5, 1, 14) {real, imag} */,
  {32'hbdbf42ec, 32'h3d2760bc} /* (5, 1, 13) {real, imag} */,
  {32'h3d40ed93, 32'hbcba28e3} /* (5, 1, 12) {real, imag} */,
  {32'hbca2ff4a, 32'hbc1d2e88} /* (5, 1, 11) {real, imag} */,
  {32'hbc0db809, 32'hbd14cb33} /* (5, 1, 10) {real, imag} */,
  {32'hbcc486f9, 32'h3cf03f2a} /* (5, 1, 9) {real, imag} */,
  {32'h3de23ebe, 32'h3dddcae6} /* (5, 1, 8) {real, imag} */,
  {32'hbd4dee94, 32'hbe324262} /* (5, 1, 7) {real, imag} */,
  {32'hbd4932c2, 32'h3c80c422} /* (5, 1, 6) {real, imag} */,
  {32'hbdc577b0, 32'hbd12f376} /* (5, 1, 5) {real, imag} */,
  {32'h3db95bb3, 32'h3e0098bb} /* (5, 1, 4) {real, imag} */,
  {32'h3de3e257, 32'h3c3059b8} /* (5, 1, 3) {real, imag} */,
  {32'hbd2687e8, 32'h3e2823a8} /* (5, 1, 2) {real, imag} */,
  {32'h3f47ae08, 32'h3ecff9b3} /* (5, 1, 1) {real, imag} */,
  {32'h3ff4a426, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'h3f588a52, 32'hbf15dae1} /* (5, 0, 31) {real, imag} */,
  {32'h3d47967e, 32'hbddee23e} /* (5, 0, 30) {real, imag} */,
  {32'h3ddbe5ac, 32'h3d54ffaa} /* (5, 0, 29) {real, imag} */,
  {32'hbc829b56, 32'hbd71b0d3} /* (5, 0, 28) {real, imag} */,
  {32'hbd5c5a1a, 32'hbc4b4642} /* (5, 0, 27) {real, imag} */,
  {32'hbd808254, 32'h3cc186e0} /* (5, 0, 26) {real, imag} */,
  {32'hbd3a297c, 32'h3d176e5c} /* (5, 0, 25) {real, imag} */,
  {32'h3d4f1056, 32'hbbdab984} /* (5, 0, 24) {real, imag} */,
  {32'hbcb7f0aa, 32'hbd2024ca} /* (5, 0, 23) {real, imag} */,
  {32'hbcf10ab8, 32'h3c16f3a0} /* (5, 0, 22) {real, imag} */,
  {32'hbbef6838, 32'hbce02a70} /* (5, 0, 21) {real, imag} */,
  {32'h3cf3265e, 32'h3d05f818} /* (5, 0, 20) {real, imag} */,
  {32'h3ce67428, 32'hbc7cbddc} /* (5, 0, 19) {real, imag} */,
  {32'hbcb83a43, 32'h3d9c8bae} /* (5, 0, 18) {real, imag} */,
  {32'hbd10932f, 32'hbc7796f4} /* (5, 0, 17) {real, imag} */,
  {32'h3d24425a, 32'h00000000} /* (5, 0, 16) {real, imag} */,
  {32'hbd10932f, 32'h3c7796f4} /* (5, 0, 15) {real, imag} */,
  {32'hbcb83a43, 32'hbd9c8bae} /* (5, 0, 14) {real, imag} */,
  {32'h3ce67428, 32'h3c7cbddc} /* (5, 0, 13) {real, imag} */,
  {32'h3cf3265e, 32'hbd05f818} /* (5, 0, 12) {real, imag} */,
  {32'hbbef6838, 32'h3ce02a70} /* (5, 0, 11) {real, imag} */,
  {32'hbcf10ab8, 32'hbc16f3a0} /* (5, 0, 10) {real, imag} */,
  {32'hbcb7f0aa, 32'h3d2024ca} /* (5, 0, 9) {real, imag} */,
  {32'h3d4f1056, 32'h3bdab984} /* (5, 0, 8) {real, imag} */,
  {32'hbd3a297c, 32'hbd176e5c} /* (5, 0, 7) {real, imag} */,
  {32'hbd808254, 32'hbcc186e0} /* (5, 0, 6) {real, imag} */,
  {32'hbd5c5a1a, 32'h3c4b4642} /* (5, 0, 5) {real, imag} */,
  {32'hbc829b56, 32'h3d71b0d3} /* (5, 0, 4) {real, imag} */,
  {32'h3ddbe5ac, 32'hbd54ffaa} /* (5, 0, 3) {real, imag} */,
  {32'h3d47967e, 32'h3ddee23e} /* (5, 0, 2) {real, imag} */,
  {32'h3f588a52, 32'h3f15dae1} /* (5, 0, 1) {real, imag} */,
  {32'h400283e6, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hbe462a88, 32'h3d6d6720} /* (4, 31, 31) {real, imag} */,
  {32'h3ed0de82, 32'hbdf61456} /* (4, 31, 30) {real, imag} */,
  {32'h3e36da98, 32'hbd59bc15} /* (4, 31, 29) {real, imag} */,
  {32'hbdf4ef42, 32'hbdab94b8} /* (4, 31, 28) {real, imag} */,
  {32'h3d57e92e, 32'hbc5c5690} /* (4, 31, 27) {real, imag} */,
  {32'hbd8e6c5e, 32'h3d9d11ed} /* (4, 31, 26) {real, imag} */,
  {32'hbbda0330, 32'hbcf10099} /* (4, 31, 25) {real, imag} */,
  {32'h3d52be99, 32'h3c89823a} /* (4, 31, 24) {real, imag} */,
  {32'hbd0eb817, 32'h3d49b103} /* (4, 31, 23) {real, imag} */,
  {32'h3d142641, 32'h3d076d31} /* (4, 31, 22) {real, imag} */,
  {32'hbd0e0c79, 32'hbd2d8768} /* (4, 31, 21) {real, imag} */,
  {32'hbd026823, 32'h3b372724} /* (4, 31, 20) {real, imag} */,
  {32'h3cbcfbba, 32'h3d01d45a} /* (4, 31, 19) {real, imag} */,
  {32'h3bf70dac, 32'hbd05e93a} /* (4, 31, 18) {real, imag} */,
  {32'h3d22f756, 32'hbcafa3a4} /* (4, 31, 17) {real, imag} */,
  {32'hbdb0f278, 32'h00000000} /* (4, 31, 16) {real, imag} */,
  {32'h3d22f756, 32'h3cafa3a4} /* (4, 31, 15) {real, imag} */,
  {32'h3bf70dac, 32'h3d05e93a} /* (4, 31, 14) {real, imag} */,
  {32'h3cbcfbba, 32'hbd01d45a} /* (4, 31, 13) {real, imag} */,
  {32'hbd026823, 32'hbb372724} /* (4, 31, 12) {real, imag} */,
  {32'hbd0e0c79, 32'h3d2d8768} /* (4, 31, 11) {real, imag} */,
  {32'h3d142641, 32'hbd076d31} /* (4, 31, 10) {real, imag} */,
  {32'hbd0eb817, 32'hbd49b103} /* (4, 31, 9) {real, imag} */,
  {32'h3d52be99, 32'hbc89823a} /* (4, 31, 8) {real, imag} */,
  {32'hbbda0330, 32'h3cf10099} /* (4, 31, 7) {real, imag} */,
  {32'hbd8e6c5e, 32'hbd9d11ed} /* (4, 31, 6) {real, imag} */,
  {32'h3d57e92e, 32'h3c5c5690} /* (4, 31, 5) {real, imag} */,
  {32'hbdf4ef42, 32'h3dab94b8} /* (4, 31, 4) {real, imag} */,
  {32'h3e36da98, 32'h3d59bc15} /* (4, 31, 3) {real, imag} */,
  {32'h3ed0de82, 32'h3df61456} /* (4, 31, 2) {real, imag} */,
  {32'hbe462a88, 32'hbd6d6720} /* (4, 31, 1) {real, imag} */,
  {32'h3f604fbc, 32'h00000000} /* (4, 31, 0) {real, imag} */,
  {32'hbf08da75, 32'h3d0f6070} /* (4, 30, 31) {real, imag} */,
  {32'h3f20cc7e, 32'hbe09d191} /* (4, 30, 30) {real, imag} */,
  {32'h3e3e44fe, 32'hbd00241b} /* (4, 30, 29) {real, imag} */,
  {32'hbe1e7236, 32'h3c099b60} /* (4, 30, 28) {real, imag} */,
  {32'h3d64081c, 32'hbcf3c99c} /* (4, 30, 27) {real, imag} */,
  {32'hbd6bc67e, 32'h3d9b5ad9} /* (4, 30, 26) {real, imag} */,
  {32'hbc4b14dc, 32'h3b827d78} /* (4, 30, 25) {real, imag} */,
  {32'h3da8abf4, 32'hbcc0572a} /* (4, 30, 24) {real, imag} */,
  {32'h3cacdc7a, 32'h3c87b744} /* (4, 30, 23) {real, imag} */,
  {32'h3b666990, 32'hbd45cfd5} /* (4, 30, 22) {real, imag} */,
  {32'h3bfa0d9c, 32'hbd283ea4} /* (4, 30, 21) {real, imag} */,
  {32'h3d0b5665, 32'hbbc355c2} /* (4, 30, 20) {real, imag} */,
  {32'h3cd78d36, 32'hbc01ea58} /* (4, 30, 19) {real, imag} */,
  {32'hbced353e, 32'hbd9ef0de} /* (4, 30, 18) {real, imag} */,
  {32'h3d3ee5f5, 32'hbd0ba779} /* (4, 30, 17) {real, imag} */,
  {32'hbd6e71d4, 32'h00000000} /* (4, 30, 16) {real, imag} */,
  {32'h3d3ee5f5, 32'h3d0ba779} /* (4, 30, 15) {real, imag} */,
  {32'hbced353e, 32'h3d9ef0de} /* (4, 30, 14) {real, imag} */,
  {32'h3cd78d36, 32'h3c01ea58} /* (4, 30, 13) {real, imag} */,
  {32'h3d0b5665, 32'h3bc355c2} /* (4, 30, 12) {real, imag} */,
  {32'h3bfa0d9c, 32'h3d283ea4} /* (4, 30, 11) {real, imag} */,
  {32'h3b666990, 32'h3d45cfd5} /* (4, 30, 10) {real, imag} */,
  {32'h3cacdc7a, 32'hbc87b744} /* (4, 30, 9) {real, imag} */,
  {32'h3da8abf4, 32'h3cc0572a} /* (4, 30, 8) {real, imag} */,
  {32'hbc4b14dc, 32'hbb827d78} /* (4, 30, 7) {real, imag} */,
  {32'hbd6bc67e, 32'hbd9b5ad9} /* (4, 30, 6) {real, imag} */,
  {32'h3d64081c, 32'h3cf3c99c} /* (4, 30, 5) {real, imag} */,
  {32'hbe1e7236, 32'hbc099b60} /* (4, 30, 4) {real, imag} */,
  {32'h3e3e44fe, 32'h3d00241b} /* (4, 30, 3) {real, imag} */,
  {32'h3f20cc7e, 32'h3e09d191} /* (4, 30, 2) {real, imag} */,
  {32'hbf08da75, 32'hbd0f6070} /* (4, 30, 1) {real, imag} */,
  {32'h3f2b6bb4, 32'h00000000} /* (4, 30, 0) {real, imag} */,
  {32'hbf2d4510, 32'hbc0d4000} /* (4, 29, 31) {real, imag} */,
  {32'h3f3ec81d, 32'hbd56a988} /* (4, 29, 30) {real, imag} */,
  {32'hbb021490, 32'hbcfe2773} /* (4, 29, 29) {real, imag} */,
  {32'hbe0f596a, 32'h3dc1da0c} /* (4, 29, 28) {real, imag} */,
  {32'h3d81ba64, 32'h3b821e50} /* (4, 29, 27) {real, imag} */,
  {32'h3d8e12f7, 32'h3db5d56d} /* (4, 29, 26) {real, imag} */,
  {32'hbe0abc5b, 32'hbc0e8728} /* (4, 29, 25) {real, imag} */,
  {32'h3df33dab, 32'hbdcb9e28} /* (4, 29, 24) {real, imag} */,
  {32'hbd8d6100, 32'hbd1c4afc} /* (4, 29, 23) {real, imag} */,
  {32'hbd1512df, 32'hbdcdff92} /* (4, 29, 22) {real, imag} */,
  {32'h3cf592e9, 32'hbdc15568} /* (4, 29, 21) {real, imag} */,
  {32'h3d299c19, 32'h3dbeb600} /* (4, 29, 20) {real, imag} */,
  {32'hbc92d030, 32'hbd576a9b} /* (4, 29, 19) {real, imag} */,
  {32'hbd25e483, 32'hbce62835} /* (4, 29, 18) {real, imag} */,
  {32'h3cccf21a, 32'hbba1d1b0} /* (4, 29, 17) {real, imag} */,
  {32'hbd49a9ae, 32'h00000000} /* (4, 29, 16) {real, imag} */,
  {32'h3cccf21a, 32'h3ba1d1b0} /* (4, 29, 15) {real, imag} */,
  {32'hbd25e483, 32'h3ce62835} /* (4, 29, 14) {real, imag} */,
  {32'hbc92d030, 32'h3d576a9b} /* (4, 29, 13) {real, imag} */,
  {32'h3d299c19, 32'hbdbeb600} /* (4, 29, 12) {real, imag} */,
  {32'h3cf592e9, 32'h3dc15568} /* (4, 29, 11) {real, imag} */,
  {32'hbd1512df, 32'h3dcdff92} /* (4, 29, 10) {real, imag} */,
  {32'hbd8d6100, 32'h3d1c4afc} /* (4, 29, 9) {real, imag} */,
  {32'h3df33dab, 32'h3dcb9e28} /* (4, 29, 8) {real, imag} */,
  {32'hbe0abc5b, 32'h3c0e8728} /* (4, 29, 7) {real, imag} */,
  {32'h3d8e12f7, 32'hbdb5d56d} /* (4, 29, 6) {real, imag} */,
  {32'h3d81ba64, 32'hbb821e50} /* (4, 29, 5) {real, imag} */,
  {32'hbe0f596a, 32'hbdc1da0c} /* (4, 29, 4) {real, imag} */,
  {32'hbb021490, 32'h3cfe2773} /* (4, 29, 3) {real, imag} */,
  {32'h3f3ec81d, 32'h3d56a988} /* (4, 29, 2) {real, imag} */,
  {32'hbf2d4510, 32'h3c0d4000} /* (4, 29, 1) {real, imag} */,
  {32'h3f14e045, 32'h00000000} /* (4, 29, 0) {real, imag} */,
  {32'hbf392fd3, 32'hbc4bcda0} /* (4, 28, 31) {real, imag} */,
  {32'h3f195331, 32'hbbb7d420} /* (4, 28, 30) {real, imag} */,
  {32'h3e5c82e5, 32'hbdb4552e} /* (4, 28, 29) {real, imag} */,
  {32'hbe64ab64, 32'h3c977520} /* (4, 28, 28) {real, imag} */,
  {32'h3e3492a4, 32'hbd8f18fe} /* (4, 28, 27) {real, imag} */,
  {32'h3e45f3d7, 32'h3c6e8312} /* (4, 28, 26) {real, imag} */,
  {32'hbdd9fdb0, 32'h3d09a34a} /* (4, 28, 25) {real, imag} */,
  {32'h3d3ada98, 32'hbdaa3d09} /* (4, 28, 24) {real, imag} */,
  {32'h3c7c0fd4, 32'hbdbe40ee} /* (4, 28, 23) {real, imag} */,
  {32'hbce44111, 32'h3d086372} /* (4, 28, 22) {real, imag} */,
  {32'hbdda4696, 32'hbd534596} /* (4, 28, 21) {real, imag} */,
  {32'hbab8f768, 32'hbc74b74a} /* (4, 28, 20) {real, imag} */,
  {32'hbcd5939d, 32'h3d2f1f40} /* (4, 28, 19) {real, imag} */,
  {32'h3cd7f64c, 32'h3cc0a91b} /* (4, 28, 18) {real, imag} */,
  {32'h3d179692, 32'h3cd50e6f} /* (4, 28, 17) {real, imag} */,
  {32'hbd37cac8, 32'h00000000} /* (4, 28, 16) {real, imag} */,
  {32'h3d179692, 32'hbcd50e6f} /* (4, 28, 15) {real, imag} */,
  {32'h3cd7f64c, 32'hbcc0a91b} /* (4, 28, 14) {real, imag} */,
  {32'hbcd5939d, 32'hbd2f1f40} /* (4, 28, 13) {real, imag} */,
  {32'hbab8f768, 32'h3c74b74a} /* (4, 28, 12) {real, imag} */,
  {32'hbdda4696, 32'h3d534596} /* (4, 28, 11) {real, imag} */,
  {32'hbce44111, 32'hbd086372} /* (4, 28, 10) {real, imag} */,
  {32'h3c7c0fd4, 32'h3dbe40ee} /* (4, 28, 9) {real, imag} */,
  {32'h3d3ada98, 32'h3daa3d09} /* (4, 28, 8) {real, imag} */,
  {32'hbdd9fdb0, 32'hbd09a34a} /* (4, 28, 7) {real, imag} */,
  {32'h3e45f3d7, 32'hbc6e8312} /* (4, 28, 6) {real, imag} */,
  {32'h3e3492a4, 32'h3d8f18fe} /* (4, 28, 5) {real, imag} */,
  {32'hbe64ab64, 32'hbc977520} /* (4, 28, 4) {real, imag} */,
  {32'h3e5c82e5, 32'h3db4552e} /* (4, 28, 3) {real, imag} */,
  {32'h3f195331, 32'h3bb7d420} /* (4, 28, 2) {real, imag} */,
  {32'hbf392fd3, 32'h3c4bcda0} /* (4, 28, 1) {real, imag} */,
  {32'h3f15f723, 32'h00000000} /* (4, 28, 0) {real, imag} */,
  {32'hbf65b10a, 32'h3df4f6bc} /* (4, 27, 31) {real, imag} */,
  {32'h3f2ce203, 32'hbbdc9e98} /* (4, 27, 30) {real, imag} */,
  {32'h3dd116a1, 32'hbe00afc9} /* (4, 27, 29) {real, imag} */,
  {32'hbe8944b9, 32'h3ce6429c} /* (4, 27, 28) {real, imag} */,
  {32'h3e1eb158, 32'hbddaf0db} /* (4, 27, 27) {real, imag} */,
  {32'h3c1d0288, 32'hbd2cce7c} /* (4, 27, 26) {real, imag} */,
  {32'hbd84a832, 32'h3cecd8e5} /* (4, 27, 25) {real, imag} */,
  {32'h3d4f8078, 32'hbe18b16e} /* (4, 27, 24) {real, imag} */,
  {32'h3c936bba, 32'h3e05d34e} /* (4, 27, 23) {real, imag} */,
  {32'hbd7df722, 32'h3d1a51c8} /* (4, 27, 22) {real, imag} */,
  {32'h3dd43f5a, 32'hbd2b54b6} /* (4, 27, 21) {real, imag} */,
  {32'hbdf4ae96, 32'hbdf2202e} /* (4, 27, 20) {real, imag} */,
  {32'h3c8151ca, 32'h3c8d0061} /* (4, 27, 19) {real, imag} */,
  {32'h3c9abde8, 32'hbe01a751} /* (4, 27, 18) {real, imag} */,
  {32'hbbe01b09, 32'h3cc16c3f} /* (4, 27, 17) {real, imag} */,
  {32'hbdb94ad5, 32'h00000000} /* (4, 27, 16) {real, imag} */,
  {32'hbbe01b09, 32'hbcc16c3f} /* (4, 27, 15) {real, imag} */,
  {32'h3c9abde8, 32'h3e01a751} /* (4, 27, 14) {real, imag} */,
  {32'h3c8151ca, 32'hbc8d0061} /* (4, 27, 13) {real, imag} */,
  {32'hbdf4ae96, 32'h3df2202e} /* (4, 27, 12) {real, imag} */,
  {32'h3dd43f5a, 32'h3d2b54b6} /* (4, 27, 11) {real, imag} */,
  {32'hbd7df722, 32'hbd1a51c8} /* (4, 27, 10) {real, imag} */,
  {32'h3c936bba, 32'hbe05d34e} /* (4, 27, 9) {real, imag} */,
  {32'h3d4f8078, 32'h3e18b16e} /* (4, 27, 8) {real, imag} */,
  {32'hbd84a832, 32'hbcecd8e5} /* (4, 27, 7) {real, imag} */,
  {32'h3c1d0288, 32'h3d2cce7c} /* (4, 27, 6) {real, imag} */,
  {32'h3e1eb158, 32'h3ddaf0db} /* (4, 27, 5) {real, imag} */,
  {32'hbe8944b9, 32'hbce6429c} /* (4, 27, 4) {real, imag} */,
  {32'h3dd116a1, 32'h3e00afc9} /* (4, 27, 3) {real, imag} */,
  {32'h3f2ce203, 32'h3bdc9e98} /* (4, 27, 2) {real, imag} */,
  {32'hbf65b10a, 32'hbdf4f6bc} /* (4, 27, 1) {real, imag} */,
  {32'h3f1c03cc, 32'h00000000} /* (4, 27, 0) {real, imag} */,
  {32'hbf62ec6f, 32'h3e6ec5dc} /* (4, 26, 31) {real, imag} */,
  {32'h3f3bf48b, 32'hbd2d2816} /* (4, 26, 30) {real, imag} */,
  {32'hbc4a50d0, 32'hbdf9923c} /* (4, 26, 29) {real, imag} */,
  {32'hbe3783dc, 32'hbcf1be06} /* (4, 26, 28) {real, imag} */,
  {32'h3e29ee63, 32'h3d065bd1} /* (4, 26, 27) {real, imag} */,
  {32'h3d685516, 32'h3be2870c} /* (4, 26, 26) {real, imag} */,
  {32'hbc5fcfbc, 32'hbd05b5d0} /* (4, 26, 25) {real, imag} */,
  {32'h3be9d858, 32'hbd8cac05} /* (4, 26, 24) {real, imag} */,
  {32'h3d99c794, 32'hbabb3500} /* (4, 26, 23) {real, imag} */,
  {32'hbcc5fe6e, 32'hbd4284bb} /* (4, 26, 22) {real, imag} */,
  {32'h3d301782, 32'hbce49f20} /* (4, 26, 21) {real, imag} */,
  {32'hbcc83206, 32'h3d6ead7c} /* (4, 26, 20) {real, imag} */,
  {32'h3da31692, 32'hbc7beacc} /* (4, 26, 19) {real, imag} */,
  {32'hbc3a6a10, 32'h3cb2126e} /* (4, 26, 18) {real, imag} */,
  {32'hbd0e634c, 32'hbd12ab48} /* (4, 26, 17) {real, imag} */,
  {32'hbd03d2b2, 32'h00000000} /* (4, 26, 16) {real, imag} */,
  {32'hbd0e634c, 32'h3d12ab48} /* (4, 26, 15) {real, imag} */,
  {32'hbc3a6a10, 32'hbcb2126e} /* (4, 26, 14) {real, imag} */,
  {32'h3da31692, 32'h3c7beacc} /* (4, 26, 13) {real, imag} */,
  {32'hbcc83206, 32'hbd6ead7c} /* (4, 26, 12) {real, imag} */,
  {32'h3d301782, 32'h3ce49f20} /* (4, 26, 11) {real, imag} */,
  {32'hbcc5fe6e, 32'h3d4284bb} /* (4, 26, 10) {real, imag} */,
  {32'h3d99c794, 32'h3abb3500} /* (4, 26, 9) {real, imag} */,
  {32'h3be9d858, 32'h3d8cac05} /* (4, 26, 8) {real, imag} */,
  {32'hbc5fcfbc, 32'h3d05b5d0} /* (4, 26, 7) {real, imag} */,
  {32'h3d685516, 32'hbbe2870c} /* (4, 26, 6) {real, imag} */,
  {32'h3e29ee63, 32'hbd065bd1} /* (4, 26, 5) {real, imag} */,
  {32'hbe3783dc, 32'h3cf1be06} /* (4, 26, 4) {real, imag} */,
  {32'hbc4a50d0, 32'h3df9923c} /* (4, 26, 3) {real, imag} */,
  {32'h3f3bf48b, 32'h3d2d2816} /* (4, 26, 2) {real, imag} */,
  {32'hbf62ec6f, 32'hbe6ec5dc} /* (4, 26, 1) {real, imag} */,
  {32'h3f04ff53, 32'h00000000} /* (4, 26, 0) {real, imag} */,
  {32'hbf886cd2, 32'h3e291975} /* (4, 25, 31) {real, imag} */,
  {32'h3f3f5c10, 32'hbccc2802} /* (4, 25, 30) {real, imag} */,
  {32'h3dc74ce9, 32'hbe29170c} /* (4, 25, 29) {real, imag} */,
  {32'hbe3182b2, 32'h3d878efb} /* (4, 25, 28) {real, imag} */,
  {32'h3e329900, 32'hbd1677ad} /* (4, 25, 27) {real, imag} */,
  {32'h3c9b335a, 32'hbc9cbfda} /* (4, 25, 26) {real, imag} */,
  {32'hbd5cba1d, 32'h3df696da} /* (4, 25, 25) {real, imag} */,
  {32'h3d54f288, 32'hbdeb1740} /* (4, 25, 24) {real, imag} */,
  {32'hbc327bbe, 32'hbdb9ef54} /* (4, 25, 23) {real, imag} */,
  {32'h3dca71ef, 32'h3d97929c} /* (4, 25, 22) {real, imag} */,
  {32'h3da98b9e, 32'h3d06abfe} /* (4, 25, 21) {real, imag} */,
  {32'hbbf68fc8, 32'h3d49bc93} /* (4, 25, 20) {real, imag} */,
  {32'hbd6105da, 32'h3c82c408} /* (4, 25, 19) {real, imag} */,
  {32'hbd425f03, 32'hbdc3e443} /* (4, 25, 18) {real, imag} */,
  {32'h3cfbd412, 32'h3de9507e} /* (4, 25, 17) {real, imag} */,
  {32'hbd428e09, 32'h00000000} /* (4, 25, 16) {real, imag} */,
  {32'h3cfbd412, 32'hbde9507e} /* (4, 25, 15) {real, imag} */,
  {32'hbd425f03, 32'h3dc3e443} /* (4, 25, 14) {real, imag} */,
  {32'hbd6105da, 32'hbc82c408} /* (4, 25, 13) {real, imag} */,
  {32'hbbf68fc8, 32'hbd49bc93} /* (4, 25, 12) {real, imag} */,
  {32'h3da98b9e, 32'hbd06abfe} /* (4, 25, 11) {real, imag} */,
  {32'h3dca71ef, 32'hbd97929c} /* (4, 25, 10) {real, imag} */,
  {32'hbc327bbe, 32'h3db9ef54} /* (4, 25, 9) {real, imag} */,
  {32'h3d54f288, 32'h3deb1740} /* (4, 25, 8) {real, imag} */,
  {32'hbd5cba1d, 32'hbdf696da} /* (4, 25, 7) {real, imag} */,
  {32'h3c9b335a, 32'h3c9cbfda} /* (4, 25, 6) {real, imag} */,
  {32'h3e329900, 32'h3d1677ad} /* (4, 25, 5) {real, imag} */,
  {32'hbe3182b2, 32'hbd878efb} /* (4, 25, 4) {real, imag} */,
  {32'h3dc74ce9, 32'h3e29170c} /* (4, 25, 3) {real, imag} */,
  {32'h3f3f5c10, 32'h3ccc2802} /* (4, 25, 2) {real, imag} */,
  {32'hbf886cd2, 32'hbe291975} /* (4, 25, 1) {real, imag} */,
  {32'h3dc7aa7c, 32'h00000000} /* (4, 25, 0) {real, imag} */,
  {32'hbfa3aaa8, 32'h3db010a2} /* (4, 24, 31) {real, imag} */,
  {32'h3f294120, 32'h3e04c7b0} /* (4, 24, 30) {real, imag} */,
  {32'hbd239084, 32'hbdb9b1aa} /* (4, 24, 29) {real, imag} */,
  {32'hbe324164, 32'hbc98199f} /* (4, 24, 28) {real, imag} */,
  {32'h3e144038, 32'hbdeda0a9} /* (4, 24, 27) {real, imag} */,
  {32'hbcadd771, 32'hbdefaa1c} /* (4, 24, 26) {real, imag} */,
  {32'hbbd1be08, 32'h3c0f6804} /* (4, 24, 25) {real, imag} */,
  {32'h3db4890d, 32'hbe5da5fa} /* (4, 24, 24) {real, imag} */,
  {32'h3c6b19fc, 32'hbd130f11} /* (4, 24, 23) {real, imag} */,
  {32'hbbacc850, 32'hbcf96dbb} /* (4, 24, 22) {real, imag} */,
  {32'h3c66322a, 32'h3b50cce0} /* (4, 24, 21) {real, imag} */,
  {32'hbc687d58, 32'h3ccb7940} /* (4, 24, 20) {real, imag} */,
  {32'h3ce51a39, 32'h3d108554} /* (4, 24, 19) {real, imag} */,
  {32'h3cf2d7e8, 32'hbd9e4d73} /* (4, 24, 18) {real, imag} */,
  {32'hbce0c3b4, 32'h3d9c2f1a} /* (4, 24, 17) {real, imag} */,
  {32'hbd595b63, 32'h00000000} /* (4, 24, 16) {real, imag} */,
  {32'hbce0c3b4, 32'hbd9c2f1a} /* (4, 24, 15) {real, imag} */,
  {32'h3cf2d7e8, 32'h3d9e4d73} /* (4, 24, 14) {real, imag} */,
  {32'h3ce51a39, 32'hbd108554} /* (4, 24, 13) {real, imag} */,
  {32'hbc687d58, 32'hbccb7940} /* (4, 24, 12) {real, imag} */,
  {32'h3c66322a, 32'hbb50cce0} /* (4, 24, 11) {real, imag} */,
  {32'hbbacc850, 32'h3cf96dbb} /* (4, 24, 10) {real, imag} */,
  {32'h3c6b19fc, 32'h3d130f11} /* (4, 24, 9) {real, imag} */,
  {32'h3db4890d, 32'h3e5da5fa} /* (4, 24, 8) {real, imag} */,
  {32'hbbd1be08, 32'hbc0f6804} /* (4, 24, 7) {real, imag} */,
  {32'hbcadd771, 32'h3defaa1c} /* (4, 24, 6) {real, imag} */,
  {32'h3e144038, 32'h3deda0a9} /* (4, 24, 5) {real, imag} */,
  {32'hbe324164, 32'h3c98199f} /* (4, 24, 4) {real, imag} */,
  {32'hbd239084, 32'h3db9b1aa} /* (4, 24, 3) {real, imag} */,
  {32'h3f294120, 32'hbe04c7b0} /* (4, 24, 2) {real, imag} */,
  {32'hbfa3aaa8, 32'hbdb010a2} /* (4, 24, 1) {real, imag} */,
  {32'h3e6934f6, 32'h00000000} /* (4, 24, 0) {real, imag} */,
  {32'hbfa0d6b7, 32'hbd0453f8} /* (4, 23, 31) {real, imag} */,
  {32'h3f236956, 32'h3e493776} /* (4, 23, 30) {real, imag} */,
  {32'hbd40485c, 32'hbcd9cc42} /* (4, 23, 29) {real, imag} */,
  {32'hbe5375f6, 32'h3cedcf7b} /* (4, 23, 28) {real, imag} */,
  {32'h3e02321b, 32'hbe1fda2e} /* (4, 23, 27) {real, imag} */,
  {32'h3d53c9b8, 32'hbd0e9856} /* (4, 23, 26) {real, imag} */,
  {32'hbd0846c7, 32'h3d48741c} /* (4, 23, 25) {real, imag} */,
  {32'hbd71446e, 32'hbcd72cfc} /* (4, 23, 24) {real, imag} */,
  {32'h3d8fd996, 32'hbc803fc8} /* (4, 23, 23) {real, imag} */,
  {32'hbcda7f05, 32'h3da43c4f} /* (4, 23, 22) {real, imag} */,
  {32'h3d3f72cf, 32'hbdec552a} /* (4, 23, 21) {real, imag} */,
  {32'hbcbb463f, 32'hbd3e4e10} /* (4, 23, 20) {real, imag} */,
  {32'hbcafcc7e, 32'hbc99d660} /* (4, 23, 19) {real, imag} */,
  {32'h3d19d198, 32'hbd99a902} /* (4, 23, 18) {real, imag} */,
  {32'h3cd44a62, 32'h3c5d7646} /* (4, 23, 17) {real, imag} */,
  {32'h3d11a6cf, 32'h00000000} /* (4, 23, 16) {real, imag} */,
  {32'h3cd44a62, 32'hbc5d7646} /* (4, 23, 15) {real, imag} */,
  {32'h3d19d198, 32'h3d99a902} /* (4, 23, 14) {real, imag} */,
  {32'hbcafcc7e, 32'h3c99d660} /* (4, 23, 13) {real, imag} */,
  {32'hbcbb463f, 32'h3d3e4e10} /* (4, 23, 12) {real, imag} */,
  {32'h3d3f72cf, 32'h3dec552a} /* (4, 23, 11) {real, imag} */,
  {32'hbcda7f05, 32'hbda43c4f} /* (4, 23, 10) {real, imag} */,
  {32'h3d8fd996, 32'h3c803fc8} /* (4, 23, 9) {real, imag} */,
  {32'hbd71446e, 32'h3cd72cfc} /* (4, 23, 8) {real, imag} */,
  {32'hbd0846c7, 32'hbd48741c} /* (4, 23, 7) {real, imag} */,
  {32'h3d53c9b8, 32'h3d0e9856} /* (4, 23, 6) {real, imag} */,
  {32'h3e02321b, 32'h3e1fda2e} /* (4, 23, 5) {real, imag} */,
  {32'hbe5375f6, 32'hbcedcf7b} /* (4, 23, 4) {real, imag} */,
  {32'hbd40485c, 32'h3cd9cc42} /* (4, 23, 3) {real, imag} */,
  {32'h3f236956, 32'hbe493776} /* (4, 23, 2) {real, imag} */,
  {32'hbfa0d6b7, 32'h3d0453f8} /* (4, 23, 1) {real, imag} */,
  {32'h3e160522, 32'h00000000} /* (4, 23, 0) {real, imag} */,
  {32'hbf810f06, 32'hbdc08a34} /* (4, 22, 31) {real, imag} */,
  {32'h3f038c9a, 32'h3e013128} /* (4, 22, 30) {real, imag} */,
  {32'hbd2db437, 32'hbdb724e2} /* (4, 22, 29) {real, imag} */,
  {32'hbe45778b, 32'h3d7e03b1} /* (4, 22, 28) {real, imag} */,
  {32'h3e4f2057, 32'hbcbcc592} /* (4, 22, 27) {real, imag} */,
  {32'hbcc86c02, 32'hbb46d2c8} /* (4, 22, 26) {real, imag} */,
  {32'hbd0b9b64, 32'hbd2aa0e4} /* (4, 22, 25) {real, imag} */,
  {32'hbc7b9514, 32'hbda00803} /* (4, 22, 24) {real, imag} */,
  {32'h3d9cdb3d, 32'hbca90ac6} /* (4, 22, 23) {real, imag} */,
  {32'hbcb6459a, 32'h3c94b2ef} /* (4, 22, 22) {real, imag} */,
  {32'h3d3410e3, 32'hbe249f22} /* (4, 22, 21) {real, imag} */,
  {32'hbd348ad4, 32'hbd0c745c} /* (4, 22, 20) {real, imag} */,
  {32'h3d292254, 32'hbde807ae} /* (4, 22, 19) {real, imag} */,
  {32'hbd326352, 32'hbd8453ce} /* (4, 22, 18) {real, imag} */,
  {32'hbb229378, 32'h3d9443a2} /* (4, 22, 17) {real, imag} */,
  {32'h3d1d565f, 32'h00000000} /* (4, 22, 16) {real, imag} */,
  {32'hbb229378, 32'hbd9443a2} /* (4, 22, 15) {real, imag} */,
  {32'hbd326352, 32'h3d8453ce} /* (4, 22, 14) {real, imag} */,
  {32'h3d292254, 32'h3de807ae} /* (4, 22, 13) {real, imag} */,
  {32'hbd348ad4, 32'h3d0c745c} /* (4, 22, 12) {real, imag} */,
  {32'h3d3410e3, 32'h3e249f22} /* (4, 22, 11) {real, imag} */,
  {32'hbcb6459a, 32'hbc94b2ef} /* (4, 22, 10) {real, imag} */,
  {32'h3d9cdb3d, 32'h3ca90ac6} /* (4, 22, 9) {real, imag} */,
  {32'hbc7b9514, 32'h3da00803} /* (4, 22, 8) {real, imag} */,
  {32'hbd0b9b64, 32'h3d2aa0e4} /* (4, 22, 7) {real, imag} */,
  {32'hbcc86c02, 32'h3b46d2c8} /* (4, 22, 6) {real, imag} */,
  {32'h3e4f2057, 32'h3cbcc592} /* (4, 22, 5) {real, imag} */,
  {32'hbe45778b, 32'hbd7e03b1} /* (4, 22, 4) {real, imag} */,
  {32'hbd2db437, 32'h3db724e2} /* (4, 22, 3) {real, imag} */,
  {32'h3f038c9a, 32'hbe013128} /* (4, 22, 2) {real, imag} */,
  {32'hbf810f06, 32'h3dc08a34} /* (4, 22, 1) {real, imag} */,
  {32'h3d87e7b5, 32'h00000000} /* (4, 22, 0) {real, imag} */,
  {32'hbee42cf0, 32'hbddd603e} /* (4, 21, 31) {real, imag} */,
  {32'h3de4abca, 32'h3ca75d12} /* (4, 21, 30) {real, imag} */,
  {32'h3d033b60, 32'hbd5d2bdb} /* (4, 21, 29) {real, imag} */,
  {32'hbd2dbad0, 32'h3be827e0} /* (4, 21, 28) {real, imag} */,
  {32'h3d89c4d3, 32'hbd7a191b} /* (4, 21, 27) {real, imag} */,
  {32'hbdb336bd, 32'hbd783c22} /* (4, 21, 26) {real, imag} */,
  {32'h3d870a23, 32'h3d35f51c} /* (4, 21, 25) {real, imag} */,
  {32'hbcbae8b9, 32'h3cbc3790} /* (4, 21, 24) {real, imag} */,
  {32'h3c824b9c, 32'hbd7f701f} /* (4, 21, 23) {real, imag} */,
  {32'hbe19c4e3, 32'hbcbed5d5} /* (4, 21, 22) {real, imag} */,
  {32'hbe1a5ce0, 32'hbd2942c9} /* (4, 21, 21) {real, imag} */,
  {32'h3c23725c, 32'h3dbdc4fa} /* (4, 21, 20) {real, imag} */,
  {32'h3dd3ce5e, 32'hbc80c90f} /* (4, 21, 19) {real, imag} */,
  {32'h3d40fa48, 32'hbd37afb5} /* (4, 21, 18) {real, imag} */,
  {32'h3d47dff4, 32'hbd84602a} /* (4, 21, 17) {real, imag} */,
  {32'hbd214716, 32'h00000000} /* (4, 21, 16) {real, imag} */,
  {32'h3d47dff4, 32'h3d84602a} /* (4, 21, 15) {real, imag} */,
  {32'h3d40fa48, 32'h3d37afb5} /* (4, 21, 14) {real, imag} */,
  {32'h3dd3ce5e, 32'h3c80c90f} /* (4, 21, 13) {real, imag} */,
  {32'h3c23725c, 32'hbdbdc4fa} /* (4, 21, 12) {real, imag} */,
  {32'hbe1a5ce0, 32'h3d2942c9} /* (4, 21, 11) {real, imag} */,
  {32'hbe19c4e3, 32'h3cbed5d5} /* (4, 21, 10) {real, imag} */,
  {32'h3c824b9c, 32'h3d7f701f} /* (4, 21, 9) {real, imag} */,
  {32'hbcbae8b9, 32'hbcbc3790} /* (4, 21, 8) {real, imag} */,
  {32'h3d870a23, 32'hbd35f51c} /* (4, 21, 7) {real, imag} */,
  {32'hbdb336bd, 32'h3d783c22} /* (4, 21, 6) {real, imag} */,
  {32'h3d89c4d3, 32'h3d7a191b} /* (4, 21, 5) {real, imag} */,
  {32'hbd2dbad0, 32'hbbe827e0} /* (4, 21, 4) {real, imag} */,
  {32'h3d033b60, 32'h3d5d2bdb} /* (4, 21, 3) {real, imag} */,
  {32'h3de4abca, 32'hbca75d12} /* (4, 21, 2) {real, imag} */,
  {32'hbee42cf0, 32'h3ddd603e} /* (4, 21, 1) {real, imag} */,
  {32'h3eef6b8a, 32'h00000000} /* (4, 21, 0) {real, imag} */,
  {32'h3efe0a34, 32'hbe9c9f6a} /* (4, 20, 31) {real, imag} */,
  {32'hbed4a6a2, 32'hbda5be6a} /* (4, 20, 30) {real, imag} */,
  {32'hbd12cbfe, 32'hbdbdd6c6} /* (4, 20, 29) {real, imag} */,
  {32'h3d942773, 32'hbd8668b2} /* (4, 20, 28) {real, imag} */,
  {32'hbe081c99, 32'hbdf25f0c} /* (4, 20, 27) {real, imag} */,
  {32'hbd230af2, 32'hbd329528} /* (4, 20, 26) {real, imag} */,
  {32'h3d64f21d, 32'h3e1f4c9c} /* (4, 20, 25) {real, imag} */,
  {32'hbdd8a8aa, 32'hbb8f8ca0} /* (4, 20, 24) {real, imag} */,
  {32'hbd84b616, 32'hbd3107fb} /* (4, 20, 23) {real, imag} */,
  {32'hbdd05062, 32'hbcbe846c} /* (4, 20, 22) {real, imag} */,
  {32'hbdd5fe6c, 32'hbc99630e} /* (4, 20, 21) {real, imag} */,
  {32'hbd1790c6, 32'hbd00d9b1} /* (4, 20, 20) {real, imag} */,
  {32'hbd7ebfe6, 32'h3d8a209b} /* (4, 20, 19) {real, imag} */,
  {32'h3cc3b8fc, 32'h3d45dac8} /* (4, 20, 18) {real, imag} */,
  {32'h3d51a810, 32'hbda3ee98} /* (4, 20, 17) {real, imag} */,
  {32'hbd1415b8, 32'h00000000} /* (4, 20, 16) {real, imag} */,
  {32'h3d51a810, 32'h3da3ee98} /* (4, 20, 15) {real, imag} */,
  {32'h3cc3b8fc, 32'hbd45dac8} /* (4, 20, 14) {real, imag} */,
  {32'hbd7ebfe6, 32'hbd8a209b} /* (4, 20, 13) {real, imag} */,
  {32'hbd1790c6, 32'h3d00d9b1} /* (4, 20, 12) {real, imag} */,
  {32'hbdd5fe6c, 32'h3c99630e} /* (4, 20, 11) {real, imag} */,
  {32'hbdd05062, 32'h3cbe846c} /* (4, 20, 10) {real, imag} */,
  {32'hbd84b616, 32'h3d3107fb} /* (4, 20, 9) {real, imag} */,
  {32'hbdd8a8aa, 32'h3b8f8ca0} /* (4, 20, 8) {real, imag} */,
  {32'h3d64f21d, 32'hbe1f4c9c} /* (4, 20, 7) {real, imag} */,
  {32'hbd230af2, 32'h3d329528} /* (4, 20, 6) {real, imag} */,
  {32'hbe081c99, 32'h3df25f0c} /* (4, 20, 5) {real, imag} */,
  {32'h3d942773, 32'h3d8668b2} /* (4, 20, 4) {real, imag} */,
  {32'hbd12cbfe, 32'h3dbdd6c6} /* (4, 20, 3) {real, imag} */,
  {32'hbed4a6a2, 32'h3da5be6a} /* (4, 20, 2) {real, imag} */,
  {32'h3efe0a34, 32'h3e9c9f6a} /* (4, 20, 1) {real, imag} */,
  {32'h3f8a0758, 32'h00000000} /* (4, 20, 0) {real, imag} */,
  {32'h3f51b273, 32'hbe2fb1b4} /* (4, 19, 31) {real, imag} */,
  {32'hbf0d3c5f, 32'h3c7b44e8} /* (4, 19, 30) {real, imag} */,
  {32'hbd97ad2a, 32'hbc6155e6} /* (4, 19, 29) {real, imag} */,
  {32'h3d30f0a0, 32'hbe298242} /* (4, 19, 28) {real, imag} */,
  {32'hbddeee80, 32'hbd0eb7d0} /* (4, 19, 27) {real, imag} */,
  {32'hbd022b06, 32'hbdc7e0b0} /* (4, 19, 26) {real, imag} */,
  {32'h3d602714, 32'h38a33800} /* (4, 19, 25) {real, imag} */,
  {32'hbc0a9d2c, 32'h3c9aa724} /* (4, 19, 24) {real, imag} */,
  {32'h3d81477b, 32'h3c12d9c6} /* (4, 19, 23) {real, imag} */,
  {32'h3d004a48, 32'hbc0e65e0} /* (4, 19, 22) {real, imag} */,
  {32'hbd675cb8, 32'h3ddd0b4d} /* (4, 19, 21) {real, imag} */,
  {32'h3c817fa4, 32'h3beaa6b0} /* (4, 19, 20) {real, imag} */,
  {32'h3b9dd17c, 32'h3d990436} /* (4, 19, 19) {real, imag} */,
  {32'h3dab7870, 32'h3d89e9f6} /* (4, 19, 18) {real, imag} */,
  {32'hbcca6c8a, 32'h3dae2fc5} /* (4, 19, 17) {real, imag} */,
  {32'h3d9a3dcd, 32'h00000000} /* (4, 19, 16) {real, imag} */,
  {32'hbcca6c8a, 32'hbdae2fc5} /* (4, 19, 15) {real, imag} */,
  {32'h3dab7870, 32'hbd89e9f6} /* (4, 19, 14) {real, imag} */,
  {32'h3b9dd17c, 32'hbd990436} /* (4, 19, 13) {real, imag} */,
  {32'h3c817fa4, 32'hbbeaa6b0} /* (4, 19, 12) {real, imag} */,
  {32'hbd675cb8, 32'hbddd0b4d} /* (4, 19, 11) {real, imag} */,
  {32'h3d004a48, 32'h3c0e65e0} /* (4, 19, 10) {real, imag} */,
  {32'h3d81477b, 32'hbc12d9c6} /* (4, 19, 9) {real, imag} */,
  {32'hbc0a9d2c, 32'hbc9aa724} /* (4, 19, 8) {real, imag} */,
  {32'h3d602714, 32'hb8a33800} /* (4, 19, 7) {real, imag} */,
  {32'hbd022b06, 32'h3dc7e0b0} /* (4, 19, 6) {real, imag} */,
  {32'hbddeee80, 32'h3d0eb7d0} /* (4, 19, 5) {real, imag} */,
  {32'h3d30f0a0, 32'h3e298242} /* (4, 19, 4) {real, imag} */,
  {32'hbd97ad2a, 32'h3c6155e6} /* (4, 19, 3) {real, imag} */,
  {32'hbf0d3c5f, 32'hbc7b44e8} /* (4, 19, 2) {real, imag} */,
  {32'h3f51b273, 32'h3e2fb1b4} /* (4, 19, 1) {real, imag} */,
  {32'h3f563718, 32'h00000000} /* (4, 19, 0) {real, imag} */,
  {32'h3f6056fc, 32'hbde8e2c8} /* (4, 18, 31) {real, imag} */,
  {32'hbf08b655, 32'h3e5f29c7} /* (4, 18, 30) {real, imag} */,
  {32'hbdb1adb1, 32'hbdb44668} /* (4, 18, 29) {real, imag} */,
  {32'h3db09169, 32'hbe1bdc24} /* (4, 18, 28) {real, imag} */,
  {32'hbe1911f4, 32'hbd205754} /* (4, 18, 27) {real, imag} */,
  {32'h3d00455c, 32'hbab82700} /* (4, 18, 26) {real, imag} */,
  {32'h3d7e2b9c, 32'hbc7af444} /* (4, 18, 25) {real, imag} */,
  {32'hbced06f6, 32'h3e009c72} /* (4, 18, 24) {real, imag} */,
  {32'hbb937ed0, 32'hbb59cb98} /* (4, 18, 23) {real, imag} */,
  {32'hbd646a1a, 32'hbd814d42} /* (4, 18, 22) {real, imag} */,
  {32'h3c61ded8, 32'h3e032cce} /* (4, 18, 21) {real, imag} */,
  {32'hbd4fc546, 32'h3cade3fa} /* (4, 18, 20) {real, imag} */,
  {32'hbd749f61, 32'hbcde2356} /* (4, 18, 19) {real, imag} */,
  {32'h3d22f122, 32'h3d096e1e} /* (4, 18, 18) {real, imag} */,
  {32'hbc9b4a9e, 32'hbd387abb} /* (4, 18, 17) {real, imag} */,
  {32'h3d433779, 32'h00000000} /* (4, 18, 16) {real, imag} */,
  {32'hbc9b4a9e, 32'h3d387abb} /* (4, 18, 15) {real, imag} */,
  {32'h3d22f122, 32'hbd096e1e} /* (4, 18, 14) {real, imag} */,
  {32'hbd749f61, 32'h3cde2356} /* (4, 18, 13) {real, imag} */,
  {32'hbd4fc546, 32'hbcade3fa} /* (4, 18, 12) {real, imag} */,
  {32'h3c61ded8, 32'hbe032cce} /* (4, 18, 11) {real, imag} */,
  {32'hbd646a1a, 32'h3d814d42} /* (4, 18, 10) {real, imag} */,
  {32'hbb937ed0, 32'h3b59cb98} /* (4, 18, 9) {real, imag} */,
  {32'hbced06f6, 32'hbe009c72} /* (4, 18, 8) {real, imag} */,
  {32'h3d7e2b9c, 32'h3c7af444} /* (4, 18, 7) {real, imag} */,
  {32'h3d00455c, 32'h3ab82700} /* (4, 18, 6) {real, imag} */,
  {32'hbe1911f4, 32'h3d205754} /* (4, 18, 5) {real, imag} */,
  {32'h3db09169, 32'h3e1bdc24} /* (4, 18, 4) {real, imag} */,
  {32'hbdb1adb1, 32'h3db44668} /* (4, 18, 3) {real, imag} */,
  {32'hbf08b655, 32'hbe5f29c7} /* (4, 18, 2) {real, imag} */,
  {32'h3f6056fc, 32'h3de8e2c8} /* (4, 18, 1) {real, imag} */,
  {32'h3f5664eb, 32'h00000000} /* (4, 18, 0) {real, imag} */,
  {32'h3f80949d, 32'hbdb42c08} /* (4, 17, 31) {real, imag} */,
  {32'hbf1023fa, 32'h3e6842d1} /* (4, 17, 30) {real, imag} */,
  {32'hbdbb9ae4, 32'h3b047aa0} /* (4, 17, 29) {real, imag} */,
  {32'h3c320538, 32'hbd6793ac} /* (4, 17, 28) {real, imag} */,
  {32'hbe304680, 32'hbb43a980} /* (4, 17, 27) {real, imag} */,
  {32'hbb2bf558, 32'hbd0cdb24} /* (4, 17, 26) {real, imag} */,
  {32'h3de63e9a, 32'hbd7e87ee} /* (4, 17, 25) {real, imag} */,
  {32'hbe2a3d83, 32'h3dc8e8b8} /* (4, 17, 24) {real, imag} */,
  {32'hbd41ce10, 32'hbd05dace} /* (4, 17, 23) {real, imag} */,
  {32'hbd74b834, 32'h3cc0dc08} /* (4, 17, 22) {real, imag} */,
  {32'hbce0a273, 32'h3d02b2dd} /* (4, 17, 21) {real, imag} */,
  {32'hbcdd34c6, 32'hbdb36450} /* (4, 17, 20) {real, imag} */,
  {32'h3d3823e4, 32'h3cb935ad} /* (4, 17, 19) {real, imag} */,
  {32'h3a2e22e0, 32'h3db8e817} /* (4, 17, 18) {real, imag} */,
  {32'hbd64f0a0, 32'h3b3a0240} /* (4, 17, 17) {real, imag} */,
  {32'h3c6ae786, 32'h00000000} /* (4, 17, 16) {real, imag} */,
  {32'hbd64f0a0, 32'hbb3a0240} /* (4, 17, 15) {real, imag} */,
  {32'h3a2e22e0, 32'hbdb8e817} /* (4, 17, 14) {real, imag} */,
  {32'h3d3823e4, 32'hbcb935ad} /* (4, 17, 13) {real, imag} */,
  {32'hbcdd34c6, 32'h3db36450} /* (4, 17, 12) {real, imag} */,
  {32'hbce0a273, 32'hbd02b2dd} /* (4, 17, 11) {real, imag} */,
  {32'hbd74b834, 32'hbcc0dc08} /* (4, 17, 10) {real, imag} */,
  {32'hbd41ce10, 32'h3d05dace} /* (4, 17, 9) {real, imag} */,
  {32'hbe2a3d83, 32'hbdc8e8b8} /* (4, 17, 8) {real, imag} */,
  {32'h3de63e9a, 32'h3d7e87ee} /* (4, 17, 7) {real, imag} */,
  {32'hbb2bf558, 32'h3d0cdb24} /* (4, 17, 6) {real, imag} */,
  {32'hbe304680, 32'h3b43a980} /* (4, 17, 5) {real, imag} */,
  {32'h3c320538, 32'h3d6793ac} /* (4, 17, 4) {real, imag} */,
  {32'hbdbb9ae4, 32'hbb047aa0} /* (4, 17, 3) {real, imag} */,
  {32'hbf1023fa, 32'hbe6842d1} /* (4, 17, 2) {real, imag} */,
  {32'h3f80949d, 32'h3db42c08} /* (4, 17, 1) {real, imag} */,
  {32'h3f4c2e3f, 32'h00000000} /* (4, 17, 0) {real, imag} */,
  {32'h3f83c284, 32'hbe576417} /* (4, 16, 31) {real, imag} */,
  {32'hbf1ea174, 32'h3e4d3afc} /* (4, 16, 30) {real, imag} */,
  {32'hbc9f5451, 32'hbb8539b0} /* (4, 16, 29) {real, imag} */,
  {32'h3e081b22, 32'hbdf07758} /* (4, 16, 28) {real, imag} */,
  {32'hbda640fc, 32'h3e205a7c} /* (4, 16, 27) {real, imag} */,
  {32'hbd232c34, 32'hbce6898b} /* (4, 16, 26) {real, imag} */,
  {32'h3cb84d3a, 32'hbe0a104e} /* (4, 16, 25) {real, imag} */,
  {32'hbdb5f66c, 32'h3df4851f} /* (4, 16, 24) {real, imag} */,
  {32'h3d66a1ad, 32'hbc2be414} /* (4, 16, 23) {real, imag} */,
  {32'h3c925283, 32'h3da6bb10} /* (4, 16, 22) {real, imag} */,
  {32'h3d258732, 32'hbd45a170} /* (4, 16, 21) {real, imag} */,
  {32'h3d247930, 32'hbd70af54} /* (4, 16, 20) {real, imag} */,
  {32'h3d6f8f8c, 32'hbc984ee6} /* (4, 16, 19) {real, imag} */,
  {32'h3d3eb334, 32'h3bbe6564} /* (4, 16, 18) {real, imag} */,
  {32'hbc5c44c1, 32'hbd2b5a75} /* (4, 16, 17) {real, imag} */,
  {32'hbcdb9c98, 32'h00000000} /* (4, 16, 16) {real, imag} */,
  {32'hbc5c44c1, 32'h3d2b5a75} /* (4, 16, 15) {real, imag} */,
  {32'h3d3eb334, 32'hbbbe6564} /* (4, 16, 14) {real, imag} */,
  {32'h3d6f8f8c, 32'h3c984ee6} /* (4, 16, 13) {real, imag} */,
  {32'h3d247930, 32'h3d70af54} /* (4, 16, 12) {real, imag} */,
  {32'h3d258732, 32'h3d45a170} /* (4, 16, 11) {real, imag} */,
  {32'h3c925283, 32'hbda6bb10} /* (4, 16, 10) {real, imag} */,
  {32'h3d66a1ad, 32'h3c2be414} /* (4, 16, 9) {real, imag} */,
  {32'hbdb5f66c, 32'hbdf4851f} /* (4, 16, 8) {real, imag} */,
  {32'h3cb84d3a, 32'h3e0a104e} /* (4, 16, 7) {real, imag} */,
  {32'hbd232c34, 32'h3ce6898b} /* (4, 16, 6) {real, imag} */,
  {32'hbda640fc, 32'hbe205a7c} /* (4, 16, 5) {real, imag} */,
  {32'h3e081b22, 32'h3df07758} /* (4, 16, 4) {real, imag} */,
  {32'hbc9f5451, 32'h3b8539b0} /* (4, 16, 3) {real, imag} */,
  {32'hbf1ea174, 32'hbe4d3afc} /* (4, 16, 2) {real, imag} */,
  {32'h3f83c284, 32'h3e576417} /* (4, 16, 1) {real, imag} */,
  {32'h3f2344fe, 32'h00000000} /* (4, 16, 0) {real, imag} */,
  {32'h3f7f9516, 32'hbecee3e4} /* (4, 15, 31) {real, imag} */,
  {32'hbf17e74a, 32'h3da12162} /* (4, 15, 30) {real, imag} */,
  {32'h3dc58430, 32'hbe065016} /* (4, 15, 29) {real, imag} */,
  {32'h3e4ddcec, 32'hbd51f126} /* (4, 15, 28) {real, imag} */,
  {32'hbe8b6c10, 32'h3e01b739} /* (4, 15, 27) {real, imag} */,
  {32'h3d27467a, 32'h3d646a08} /* (4, 15, 26) {real, imag} */,
  {32'h3ceab590, 32'h3c0bfb2e} /* (4, 15, 25) {real, imag} */,
  {32'hbd670dfc, 32'h3d490f99} /* (4, 15, 24) {real, imag} */,
  {32'h3d38d08c, 32'h3dad368a} /* (4, 15, 23) {real, imag} */,
  {32'h3ca1c524, 32'h3d1fe158} /* (4, 15, 22) {real, imag} */,
  {32'h3af6aff0, 32'h3d5b812d} /* (4, 15, 21) {real, imag} */,
  {32'h3bf26288, 32'h3d816acc} /* (4, 15, 20) {real, imag} */,
  {32'hbc40d5a6, 32'h3bef33a4} /* (4, 15, 19) {real, imag} */,
  {32'h3d5de5cc, 32'h3db84365} /* (4, 15, 18) {real, imag} */,
  {32'h3955d080, 32'hbdc031b9} /* (4, 15, 17) {real, imag} */,
  {32'h3d541b7e, 32'h00000000} /* (4, 15, 16) {real, imag} */,
  {32'h3955d080, 32'h3dc031b9} /* (4, 15, 15) {real, imag} */,
  {32'h3d5de5cc, 32'hbdb84365} /* (4, 15, 14) {real, imag} */,
  {32'hbc40d5a6, 32'hbbef33a4} /* (4, 15, 13) {real, imag} */,
  {32'h3bf26288, 32'hbd816acc} /* (4, 15, 12) {real, imag} */,
  {32'h3af6aff0, 32'hbd5b812d} /* (4, 15, 11) {real, imag} */,
  {32'h3ca1c524, 32'hbd1fe158} /* (4, 15, 10) {real, imag} */,
  {32'h3d38d08c, 32'hbdad368a} /* (4, 15, 9) {real, imag} */,
  {32'hbd670dfc, 32'hbd490f99} /* (4, 15, 8) {real, imag} */,
  {32'h3ceab590, 32'hbc0bfb2e} /* (4, 15, 7) {real, imag} */,
  {32'h3d27467a, 32'hbd646a08} /* (4, 15, 6) {real, imag} */,
  {32'hbe8b6c10, 32'hbe01b739} /* (4, 15, 5) {real, imag} */,
  {32'h3e4ddcec, 32'h3d51f126} /* (4, 15, 4) {real, imag} */,
  {32'h3dc58430, 32'h3e065016} /* (4, 15, 3) {real, imag} */,
  {32'hbf17e74a, 32'hbda12162} /* (4, 15, 2) {real, imag} */,
  {32'h3f7f9516, 32'h3ecee3e4} /* (4, 15, 1) {real, imag} */,
  {32'h3f2a43e5, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'h3f808084, 32'hbe8715ac} /* (4, 14, 31) {real, imag} */,
  {32'hbf0cbedf, 32'hbca1ba48} /* (4, 14, 30) {real, imag} */,
  {32'h3df6e325, 32'hbe523594} /* (4, 14, 29) {real, imag} */,
  {32'h3de313ab, 32'hbdee9fdf} /* (4, 14, 28) {real, imag} */,
  {32'hbd86aa61, 32'h3e05b187} /* (4, 14, 27) {real, imag} */,
  {32'h3da34e74, 32'h3dbd3420} /* (4, 14, 26) {real, imag} */,
  {32'h3dc51ae2, 32'hbc2a49ec} /* (4, 14, 25) {real, imag} */,
  {32'hbc296a4d, 32'h3ccbdf5c} /* (4, 14, 24) {real, imag} */,
  {32'h3d9237bb, 32'h3d1a3ed6} /* (4, 14, 23) {real, imag} */,
  {32'h3d2c3874, 32'hbc873a5e} /* (4, 14, 22) {real, imag} */,
  {32'hbe0c2d8e, 32'h3c79663c} /* (4, 14, 21) {real, imag} */,
  {32'hbd3c1714, 32'h3c923054} /* (4, 14, 20) {real, imag} */,
  {32'hbdd0bace, 32'hbadc05c0} /* (4, 14, 19) {real, imag} */,
  {32'h3bb0409c, 32'h3d647810} /* (4, 14, 18) {real, imag} */,
  {32'hbdb30ca0, 32'h3d4f187d} /* (4, 14, 17) {real, imag} */,
  {32'hbd2c5a5f, 32'h00000000} /* (4, 14, 16) {real, imag} */,
  {32'hbdb30ca0, 32'hbd4f187d} /* (4, 14, 15) {real, imag} */,
  {32'h3bb0409c, 32'hbd647810} /* (4, 14, 14) {real, imag} */,
  {32'hbdd0bace, 32'h3adc05c0} /* (4, 14, 13) {real, imag} */,
  {32'hbd3c1714, 32'hbc923054} /* (4, 14, 12) {real, imag} */,
  {32'hbe0c2d8e, 32'hbc79663c} /* (4, 14, 11) {real, imag} */,
  {32'h3d2c3874, 32'h3c873a5e} /* (4, 14, 10) {real, imag} */,
  {32'h3d9237bb, 32'hbd1a3ed6} /* (4, 14, 9) {real, imag} */,
  {32'hbc296a4d, 32'hbccbdf5c} /* (4, 14, 8) {real, imag} */,
  {32'h3dc51ae2, 32'h3c2a49ec} /* (4, 14, 7) {real, imag} */,
  {32'h3da34e74, 32'hbdbd3420} /* (4, 14, 6) {real, imag} */,
  {32'hbd86aa61, 32'hbe05b187} /* (4, 14, 5) {real, imag} */,
  {32'h3de313ab, 32'h3dee9fdf} /* (4, 14, 4) {real, imag} */,
  {32'h3df6e325, 32'h3e523594} /* (4, 14, 3) {real, imag} */,
  {32'hbf0cbedf, 32'h3ca1ba48} /* (4, 14, 2) {real, imag} */,
  {32'h3f808084, 32'h3e8715ac} /* (4, 14, 1) {real, imag} */,
  {32'h3f34b3a1, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'h3f83c8b6, 32'hbe7c5a98} /* (4, 13, 31) {real, imag} */,
  {32'hbedff9f6, 32'hbd8dd99d} /* (4, 13, 30) {real, imag} */,
  {32'h3e24f51c, 32'h3d37fd1a} /* (4, 13, 29) {real, imag} */,
  {32'h3dc9ff3a, 32'hbd91b028} /* (4, 13, 28) {real, imag} */,
  {32'hbdec4474, 32'h3e7e86e4} /* (4, 13, 27) {real, imag} */,
  {32'h3e490994, 32'h3dbf517c} /* (4, 13, 26) {real, imag} */,
  {32'hbba9a4fc, 32'hbcae6c6f} /* (4, 13, 25) {real, imag} */,
  {32'hbdae2e22, 32'h3d16785a} /* (4, 13, 24) {real, imag} */,
  {32'h3d7658d4, 32'h3c3c7b22} /* (4, 13, 23) {real, imag} */,
  {32'hbcdd2a3d, 32'hbd803444} /* (4, 13, 22) {real, imag} */,
  {32'h3ca20cf0, 32'h3de4c13b} /* (4, 13, 21) {real, imag} */,
  {32'h3d9cbe62, 32'hbd725ff2} /* (4, 13, 20) {real, imag} */,
  {32'h3cc81197, 32'hbd593cd3} /* (4, 13, 19) {real, imag} */,
  {32'h3cf2a07c, 32'h3c11364e} /* (4, 13, 18) {real, imag} */,
  {32'hbbcfee8e, 32'hbcd0e23c} /* (4, 13, 17) {real, imag} */,
  {32'h3d22c33a, 32'h00000000} /* (4, 13, 16) {real, imag} */,
  {32'hbbcfee8e, 32'h3cd0e23c} /* (4, 13, 15) {real, imag} */,
  {32'h3cf2a07c, 32'hbc11364e} /* (4, 13, 14) {real, imag} */,
  {32'h3cc81197, 32'h3d593cd3} /* (4, 13, 13) {real, imag} */,
  {32'h3d9cbe62, 32'h3d725ff2} /* (4, 13, 12) {real, imag} */,
  {32'h3ca20cf0, 32'hbde4c13b} /* (4, 13, 11) {real, imag} */,
  {32'hbcdd2a3d, 32'h3d803444} /* (4, 13, 10) {real, imag} */,
  {32'h3d7658d4, 32'hbc3c7b22} /* (4, 13, 9) {real, imag} */,
  {32'hbdae2e22, 32'hbd16785a} /* (4, 13, 8) {real, imag} */,
  {32'hbba9a4fc, 32'h3cae6c6f} /* (4, 13, 7) {real, imag} */,
  {32'h3e490994, 32'hbdbf517c} /* (4, 13, 6) {real, imag} */,
  {32'hbdec4474, 32'hbe7e86e4} /* (4, 13, 5) {real, imag} */,
  {32'h3dc9ff3a, 32'h3d91b028} /* (4, 13, 4) {real, imag} */,
  {32'h3e24f51c, 32'hbd37fd1a} /* (4, 13, 3) {real, imag} */,
  {32'hbedff9f6, 32'h3d8dd99d} /* (4, 13, 2) {real, imag} */,
  {32'h3f83c8b6, 32'h3e7c5a98} /* (4, 13, 1) {real, imag} */,
  {32'h3f1dd89a, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'h3f626e9e, 32'hbe629d19} /* (4, 12, 31) {real, imag} */,
  {32'hbee1ef8a, 32'hbd0a021b} /* (4, 12, 30) {real, imag} */,
  {32'h3e297e28, 32'h3daac09c} /* (4, 12, 29) {real, imag} */,
  {32'h3da3cf69, 32'hbd7b949c} /* (4, 12, 28) {real, imag} */,
  {32'hbe7601f9, 32'h3da79694} /* (4, 12, 27) {real, imag} */,
  {32'h3dbc5f19, 32'h3db7f0ce} /* (4, 12, 26) {real, imag} */,
  {32'h3cbeabb6, 32'h3ce3c684} /* (4, 12, 25) {real, imag} */,
  {32'hbd7ca46d, 32'h3d86356c} /* (4, 12, 24) {real, imag} */,
  {32'h3d86e81a, 32'hb8511000} /* (4, 12, 23) {real, imag} */,
  {32'h3b2fbcb0, 32'h3c793bc4} /* (4, 12, 22) {real, imag} */,
  {32'hbcf71938, 32'h3dd80e8a} /* (4, 12, 21) {real, imag} */,
  {32'h3b0584b8, 32'hbd25280b} /* (4, 12, 20) {real, imag} */,
  {32'h3cabe06b, 32'hbd2b9f62} /* (4, 12, 19) {real, imag} */,
  {32'h3c2ead40, 32'hbd852ab8} /* (4, 12, 18) {real, imag} */,
  {32'h3c0371ea, 32'h3cc69922} /* (4, 12, 17) {real, imag} */,
  {32'h3dded54c, 32'h00000000} /* (4, 12, 16) {real, imag} */,
  {32'h3c0371ea, 32'hbcc69922} /* (4, 12, 15) {real, imag} */,
  {32'h3c2ead40, 32'h3d852ab8} /* (4, 12, 14) {real, imag} */,
  {32'h3cabe06b, 32'h3d2b9f62} /* (4, 12, 13) {real, imag} */,
  {32'h3b0584b8, 32'h3d25280b} /* (4, 12, 12) {real, imag} */,
  {32'hbcf71938, 32'hbdd80e8a} /* (4, 12, 11) {real, imag} */,
  {32'h3b2fbcb0, 32'hbc793bc4} /* (4, 12, 10) {real, imag} */,
  {32'h3d86e81a, 32'h38511000} /* (4, 12, 9) {real, imag} */,
  {32'hbd7ca46d, 32'hbd86356c} /* (4, 12, 8) {real, imag} */,
  {32'h3cbeabb6, 32'hbce3c684} /* (4, 12, 7) {real, imag} */,
  {32'h3dbc5f19, 32'hbdb7f0ce} /* (4, 12, 6) {real, imag} */,
  {32'hbe7601f9, 32'hbda79694} /* (4, 12, 5) {real, imag} */,
  {32'h3da3cf69, 32'h3d7b949c} /* (4, 12, 4) {real, imag} */,
  {32'h3e297e28, 32'hbdaac09c} /* (4, 12, 3) {real, imag} */,
  {32'hbee1ef8a, 32'h3d0a021b} /* (4, 12, 2) {real, imag} */,
  {32'h3f626e9e, 32'h3e629d19} /* (4, 12, 1) {real, imag} */,
  {32'h3f335a46, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'h3f3380d2, 32'hbe62c373} /* (4, 11, 31) {real, imag} */,
  {32'hbeb58202, 32'hbcae7276} /* (4, 11, 30) {real, imag} */,
  {32'h3e23f03d, 32'hbcc1df66} /* (4, 11, 29) {real, imag} */,
  {32'h3d447898, 32'hbd31b898} /* (4, 11, 28) {real, imag} */,
  {32'hbe50f924, 32'h3da33230} /* (4, 11, 27) {real, imag} */,
  {32'h3e32660a, 32'h3d5fe128} /* (4, 11, 26) {real, imag} */,
  {32'h3d2a5b9a, 32'h3d74f5e8} /* (4, 11, 25) {real, imag} */,
  {32'hbd3a7174, 32'h3cfb1908} /* (4, 11, 24) {real, imag} */,
  {32'hbd2db3ba, 32'hbd19b641} /* (4, 11, 23) {real, imag} */,
  {32'h3e01169f, 32'h3cd33d6b} /* (4, 11, 22) {real, imag} */,
  {32'hbd9241ad, 32'h3ce77fbe} /* (4, 11, 21) {real, imag} */,
  {32'hbd344435, 32'h3bdf90a0} /* (4, 11, 20) {real, imag} */,
  {32'h3c62efcc, 32'h3d7585ce} /* (4, 11, 19) {real, imag} */,
  {32'h3bf094a4, 32'h3df11a9a} /* (4, 11, 18) {real, imag} */,
  {32'hbcdfb640, 32'hbc43d8a2} /* (4, 11, 17) {real, imag} */,
  {32'h3d0379b0, 32'h00000000} /* (4, 11, 16) {real, imag} */,
  {32'hbcdfb640, 32'h3c43d8a2} /* (4, 11, 15) {real, imag} */,
  {32'h3bf094a4, 32'hbdf11a9a} /* (4, 11, 14) {real, imag} */,
  {32'h3c62efcc, 32'hbd7585ce} /* (4, 11, 13) {real, imag} */,
  {32'hbd344435, 32'hbbdf90a0} /* (4, 11, 12) {real, imag} */,
  {32'hbd9241ad, 32'hbce77fbe} /* (4, 11, 11) {real, imag} */,
  {32'h3e01169f, 32'hbcd33d6b} /* (4, 11, 10) {real, imag} */,
  {32'hbd2db3ba, 32'h3d19b641} /* (4, 11, 9) {real, imag} */,
  {32'hbd3a7174, 32'hbcfb1908} /* (4, 11, 8) {real, imag} */,
  {32'h3d2a5b9a, 32'hbd74f5e8} /* (4, 11, 7) {real, imag} */,
  {32'h3e32660a, 32'hbd5fe128} /* (4, 11, 6) {real, imag} */,
  {32'hbe50f924, 32'hbda33230} /* (4, 11, 5) {real, imag} */,
  {32'h3d447898, 32'h3d31b898} /* (4, 11, 4) {real, imag} */,
  {32'h3e23f03d, 32'h3cc1df66} /* (4, 11, 3) {real, imag} */,
  {32'hbeb58202, 32'h3cae7276} /* (4, 11, 2) {real, imag} */,
  {32'h3f3380d2, 32'h3e62c373} /* (4, 11, 1) {real, imag} */,
  {32'h3f1a2f81, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'hbdc5ce50, 32'hbe01ce7f} /* (4, 10, 31) {real, imag} */,
  {32'h3e5598de, 32'hbdb753a7} /* (4, 10, 30) {real, imag} */,
  {32'h3e169152, 32'hbc863946} /* (4, 10, 29) {real, imag} */,
  {32'hbd8e3d8a, 32'hbcd54892} /* (4, 10, 28) {real, imag} */,
  {32'h3d466534, 32'hbdb59702} /* (4, 10, 27) {real, imag} */,
  {32'h3dea221c, 32'hbd09f3d8} /* (4, 10, 26) {real, imag} */,
  {32'hbdeb29b4, 32'h3dfbbc20} /* (4, 10, 25) {real, imag} */,
  {32'h3d4ca7c9, 32'hbd4615a6} /* (4, 10, 24) {real, imag} */,
  {32'hbdcdf8f5, 32'h3dbdf1d4} /* (4, 10, 23) {real, imag} */,
  {32'hbba5e1e6, 32'hbcbb63ed} /* (4, 10, 22) {real, imag} */,
  {32'hbcf94b2b, 32'hbd9f7a5d} /* (4, 10, 21) {real, imag} */,
  {32'h3cf8bb98, 32'h3dccfe5a} /* (4, 10, 20) {real, imag} */,
  {32'hbbe5a9b8, 32'hbd5a66d5} /* (4, 10, 19) {real, imag} */,
  {32'hbd99f92f, 32'h3be89978} /* (4, 10, 18) {real, imag} */,
  {32'h3d08f0d8, 32'h3d4e09d0} /* (4, 10, 17) {real, imag} */,
  {32'hbc9861fe, 32'h00000000} /* (4, 10, 16) {real, imag} */,
  {32'h3d08f0d8, 32'hbd4e09d0} /* (4, 10, 15) {real, imag} */,
  {32'hbd99f92f, 32'hbbe89978} /* (4, 10, 14) {real, imag} */,
  {32'hbbe5a9b8, 32'h3d5a66d5} /* (4, 10, 13) {real, imag} */,
  {32'h3cf8bb98, 32'hbdccfe5a} /* (4, 10, 12) {real, imag} */,
  {32'hbcf94b2b, 32'h3d9f7a5d} /* (4, 10, 11) {real, imag} */,
  {32'hbba5e1e6, 32'h3cbb63ed} /* (4, 10, 10) {real, imag} */,
  {32'hbdcdf8f5, 32'hbdbdf1d4} /* (4, 10, 9) {real, imag} */,
  {32'h3d4ca7c9, 32'h3d4615a6} /* (4, 10, 8) {real, imag} */,
  {32'hbdeb29b4, 32'hbdfbbc20} /* (4, 10, 7) {real, imag} */,
  {32'h3dea221c, 32'h3d09f3d8} /* (4, 10, 6) {real, imag} */,
  {32'h3d466534, 32'h3db59702} /* (4, 10, 5) {real, imag} */,
  {32'hbd8e3d8a, 32'h3cd54892} /* (4, 10, 4) {real, imag} */,
  {32'h3e169152, 32'h3c863946} /* (4, 10, 3) {real, imag} */,
  {32'h3e5598de, 32'h3db753a7} /* (4, 10, 2) {real, imag} */,
  {32'hbdc5ce50, 32'h3e01ce7f} /* (4, 10, 1) {real, imag} */,
  {32'hbd5b9da2, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'hbf1daf98, 32'hbda39b8e} /* (4, 9, 31) {real, imag} */,
  {32'h3edd0fd5, 32'hbb901ff0} /* (4, 9, 30) {real, imag} */,
  {32'h3da36cc4, 32'hbd1286e9} /* (4, 9, 29) {real, imag} */,
  {32'hbddd836f, 32'h3d2a0302} /* (4, 9, 28) {real, imag} */,
  {32'h3e4c6487, 32'hbe294f4e} /* (4, 9, 27) {real, imag} */,
  {32'h3de97880, 32'hbd08d3b4} /* (4, 9, 26) {real, imag} */,
  {32'hbd83c132, 32'h3d4de248} /* (4, 9, 25) {real, imag} */,
  {32'h3d6858bc, 32'hbdb31c6e} /* (4, 9, 24) {real, imag} */,
  {32'h3d013860, 32'h3c5ed4b8} /* (4, 9, 23) {real, imag} */,
  {32'h3c87e13d, 32'h3ce0d6e4} /* (4, 9, 22) {real, imag} */,
  {32'hb9001f00, 32'hbc4f6140} /* (4, 9, 21) {real, imag} */,
  {32'hbcc67e53, 32'h3d9bfc1d} /* (4, 9, 20) {real, imag} */,
  {32'h3d18058f, 32'h3d94eab8} /* (4, 9, 19) {real, imag} */,
  {32'hbd629840, 32'hbd5c6d4f} /* (4, 9, 18) {real, imag} */,
  {32'hbdc54ed2, 32'h3d1e5b8e} /* (4, 9, 17) {real, imag} */,
  {32'h3d89d0fa, 32'h00000000} /* (4, 9, 16) {real, imag} */,
  {32'hbdc54ed2, 32'hbd1e5b8e} /* (4, 9, 15) {real, imag} */,
  {32'hbd629840, 32'h3d5c6d4f} /* (4, 9, 14) {real, imag} */,
  {32'h3d18058f, 32'hbd94eab8} /* (4, 9, 13) {real, imag} */,
  {32'hbcc67e53, 32'hbd9bfc1d} /* (4, 9, 12) {real, imag} */,
  {32'hb9001f00, 32'h3c4f6140} /* (4, 9, 11) {real, imag} */,
  {32'h3c87e13d, 32'hbce0d6e4} /* (4, 9, 10) {real, imag} */,
  {32'h3d013860, 32'hbc5ed4b8} /* (4, 9, 9) {real, imag} */,
  {32'h3d6858bc, 32'h3db31c6e} /* (4, 9, 8) {real, imag} */,
  {32'hbd83c132, 32'hbd4de248} /* (4, 9, 7) {real, imag} */,
  {32'h3de97880, 32'h3d08d3b4} /* (4, 9, 6) {real, imag} */,
  {32'h3e4c6487, 32'h3e294f4e} /* (4, 9, 5) {real, imag} */,
  {32'hbddd836f, 32'hbd2a0302} /* (4, 9, 4) {real, imag} */,
  {32'h3da36cc4, 32'h3d1286e9} /* (4, 9, 3) {real, imag} */,
  {32'h3edd0fd5, 32'h3b901ff0} /* (4, 9, 2) {real, imag} */,
  {32'hbf1daf98, 32'h3da39b8e} /* (4, 9, 1) {real, imag} */,
  {32'hbdf1793c, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'hbf4c0b48, 32'hbdddaa3a} /* (4, 8, 31) {real, imag} */,
  {32'h3f0843b4, 32'h3dbafe97} /* (4, 8, 30) {real, imag} */,
  {32'h3e181eb1, 32'hbd94ea3a} /* (4, 8, 29) {real, imag} */,
  {32'h3b9028c0, 32'h3c0a057e} /* (4, 8, 28) {real, imag} */,
  {32'h3de5fea1, 32'hbdebd2ff} /* (4, 8, 27) {real, imag} */,
  {32'h3d0d9c72, 32'h3d797924} /* (4, 8, 26) {real, imag} */,
  {32'hbdd4fa74, 32'h3d0e8730} /* (4, 8, 25) {real, imag} */,
  {32'h3d3d286e, 32'hbe0e981a} /* (4, 8, 24) {real, imag} */,
  {32'hbd4246f3, 32'hbc599cc4} /* (4, 8, 23) {real, imag} */,
  {32'h39fdb700, 32'hbd96cc38} /* (4, 8, 22) {real, imag} */,
  {32'h3d1a7542, 32'h3dc15ff5} /* (4, 8, 21) {real, imag} */,
  {32'hbd806722, 32'hbdabf0a2} /* (4, 8, 20) {real, imag} */,
  {32'h3d92bcef, 32'hbc8edf48} /* (4, 8, 19) {real, imag} */,
  {32'h3d10208c, 32'h3af615c0} /* (4, 8, 18) {real, imag} */,
  {32'hbb3d8934, 32'h3c8f6b7b} /* (4, 8, 17) {real, imag} */,
  {32'hbce29906, 32'h00000000} /* (4, 8, 16) {real, imag} */,
  {32'hbb3d8934, 32'hbc8f6b7b} /* (4, 8, 15) {real, imag} */,
  {32'h3d10208c, 32'hbaf615c0} /* (4, 8, 14) {real, imag} */,
  {32'h3d92bcef, 32'h3c8edf48} /* (4, 8, 13) {real, imag} */,
  {32'hbd806722, 32'h3dabf0a2} /* (4, 8, 12) {real, imag} */,
  {32'h3d1a7542, 32'hbdc15ff5} /* (4, 8, 11) {real, imag} */,
  {32'h39fdb700, 32'h3d96cc38} /* (4, 8, 10) {real, imag} */,
  {32'hbd4246f3, 32'h3c599cc4} /* (4, 8, 9) {real, imag} */,
  {32'h3d3d286e, 32'h3e0e981a} /* (4, 8, 8) {real, imag} */,
  {32'hbdd4fa74, 32'hbd0e8730} /* (4, 8, 7) {real, imag} */,
  {32'h3d0d9c72, 32'hbd797924} /* (4, 8, 6) {real, imag} */,
  {32'h3de5fea1, 32'h3debd2ff} /* (4, 8, 5) {real, imag} */,
  {32'h3b9028c0, 32'hbc0a057e} /* (4, 8, 4) {real, imag} */,
  {32'h3e181eb1, 32'h3d94ea3a} /* (4, 8, 3) {real, imag} */,
  {32'h3f0843b4, 32'hbdbafe97} /* (4, 8, 2) {real, imag} */,
  {32'hbf4c0b48, 32'h3dddaa3a} /* (4, 8, 1) {real, imag} */,
  {32'hbd08d678, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'hbf55fa23, 32'h3da3454c} /* (4, 7, 31) {real, imag} */,
  {32'h3f206f50, 32'h3d068963} /* (4, 7, 30) {real, imag} */,
  {32'h3e7f0584, 32'hbe008de4} /* (4, 7, 29) {real, imag} */,
  {32'h3d84f14d, 32'hbd4a2d1e} /* (4, 7, 28) {real, imag} */,
  {32'h3b0513a0, 32'h3c7aeb14} /* (4, 7, 27) {real, imag} */,
  {32'hbc6bab6c, 32'h3dbdf560} /* (4, 7, 26) {real, imag} */,
  {32'hbd0e89ef, 32'h3d730b28} /* (4, 7, 25) {real, imag} */,
  {32'h3c13aaa8, 32'hbd2fef51} /* (4, 7, 24) {real, imag} */,
  {32'h3d1079ac, 32'h3ba9fb28} /* (4, 7, 23) {real, imag} */,
  {32'hbd6ab5ea, 32'hbd1d4120} /* (4, 7, 22) {real, imag} */,
  {32'h3db69396, 32'hbd39c4ce} /* (4, 7, 21) {real, imag} */,
  {32'hbd58682e, 32'h3d9bf482} /* (4, 7, 20) {real, imag} */,
  {32'hbb037d00, 32'hbc4873a8} /* (4, 7, 19) {real, imag} */,
  {32'h3d695f75, 32'h39a6b900} /* (4, 7, 18) {real, imag} */,
  {32'hbc9dd4e4, 32'h3ccf9870} /* (4, 7, 17) {real, imag} */,
  {32'hbe28ab3f, 32'h00000000} /* (4, 7, 16) {real, imag} */,
  {32'hbc9dd4e4, 32'hbccf9870} /* (4, 7, 15) {real, imag} */,
  {32'h3d695f75, 32'hb9a6b900} /* (4, 7, 14) {real, imag} */,
  {32'hbb037d00, 32'h3c4873a8} /* (4, 7, 13) {real, imag} */,
  {32'hbd58682e, 32'hbd9bf482} /* (4, 7, 12) {real, imag} */,
  {32'h3db69396, 32'h3d39c4ce} /* (4, 7, 11) {real, imag} */,
  {32'hbd6ab5ea, 32'h3d1d4120} /* (4, 7, 10) {real, imag} */,
  {32'h3d1079ac, 32'hbba9fb28} /* (4, 7, 9) {real, imag} */,
  {32'h3c13aaa8, 32'h3d2fef51} /* (4, 7, 8) {real, imag} */,
  {32'hbd0e89ef, 32'hbd730b28} /* (4, 7, 7) {real, imag} */,
  {32'hbc6bab6c, 32'hbdbdf560} /* (4, 7, 6) {real, imag} */,
  {32'h3b0513a0, 32'hbc7aeb14} /* (4, 7, 5) {real, imag} */,
  {32'h3d84f14d, 32'h3d4a2d1e} /* (4, 7, 4) {real, imag} */,
  {32'h3e7f0584, 32'h3e008de4} /* (4, 7, 3) {real, imag} */,
  {32'h3f206f50, 32'hbd068963} /* (4, 7, 2) {real, imag} */,
  {32'hbf55fa23, 32'hbda3454c} /* (4, 7, 1) {real, imag} */,
  {32'h3e91810f, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'hbf2b9e87, 32'h3df07c51} /* (4, 6, 31) {real, imag} */,
  {32'h3ed93cbe, 32'h3bb870d0} /* (4, 6, 30) {real, imag} */,
  {32'h3e3a60f7, 32'h3d604f80} /* (4, 6, 29) {real, imag} */,
  {32'h3d956467, 32'hbd30639d} /* (4, 6, 28) {real, imag} */,
  {32'h3c8d4508, 32'hbd7e6443} /* (4, 6, 27) {real, imag} */,
  {32'h3d811cbe, 32'h3d4023c8} /* (4, 6, 26) {real, imag} */,
  {32'h3dcfff9a, 32'hbe01abf3} /* (4, 6, 25) {real, imag} */,
  {32'hbd29b4db, 32'hbcdd882b} /* (4, 6, 24) {real, imag} */,
  {32'hbd9c6cb2, 32'hbd167c36} /* (4, 6, 23) {real, imag} */,
  {32'hbda7edb0, 32'h3d4fba97} /* (4, 6, 22) {real, imag} */,
  {32'hbdaff515, 32'hbc3a42d0} /* (4, 6, 21) {real, imag} */,
  {32'hbcf6356e, 32'h3ce72d79} /* (4, 6, 20) {real, imag} */,
  {32'h3d8bfd1e, 32'h3d6a07ef} /* (4, 6, 19) {real, imag} */,
  {32'h3d93e0f4, 32'h3db2bf3a} /* (4, 6, 18) {real, imag} */,
  {32'h3cbca5d0, 32'h3c9d114f} /* (4, 6, 17) {real, imag} */,
  {32'hbcde661f, 32'h00000000} /* (4, 6, 16) {real, imag} */,
  {32'h3cbca5d0, 32'hbc9d114f} /* (4, 6, 15) {real, imag} */,
  {32'h3d93e0f4, 32'hbdb2bf3a} /* (4, 6, 14) {real, imag} */,
  {32'h3d8bfd1e, 32'hbd6a07ef} /* (4, 6, 13) {real, imag} */,
  {32'hbcf6356e, 32'hbce72d79} /* (4, 6, 12) {real, imag} */,
  {32'hbdaff515, 32'h3c3a42d0} /* (4, 6, 11) {real, imag} */,
  {32'hbda7edb0, 32'hbd4fba97} /* (4, 6, 10) {real, imag} */,
  {32'hbd9c6cb2, 32'h3d167c36} /* (4, 6, 9) {real, imag} */,
  {32'hbd29b4db, 32'h3cdd882b} /* (4, 6, 8) {real, imag} */,
  {32'h3dcfff9a, 32'h3e01abf3} /* (4, 6, 7) {real, imag} */,
  {32'h3d811cbe, 32'hbd4023c8} /* (4, 6, 6) {real, imag} */,
  {32'h3c8d4508, 32'h3d7e6443} /* (4, 6, 5) {real, imag} */,
  {32'h3d956467, 32'h3d30639d} /* (4, 6, 4) {real, imag} */,
  {32'h3e3a60f7, 32'hbd604f80} /* (4, 6, 3) {real, imag} */,
  {32'h3ed93cbe, 32'hbbb870d0} /* (4, 6, 2) {real, imag} */,
  {32'hbf2b9e87, 32'hbdf07c51} /* (4, 6, 1) {real, imag} */,
  {32'h3e95be7e, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'hbea0ee50, 32'h3f30aa7a} /* (4, 5, 31) {real, imag} */,
  {32'h3e0cc474, 32'hbc57c73c} /* (4, 5, 30) {real, imag} */,
  {32'h3e77bf44, 32'hbd7cbe94} /* (4, 5, 29) {real, imag} */,
  {32'h3cb9ae80, 32'hbe7abb40} /* (4, 5, 28) {real, imag} */,
  {32'h3dd43f90, 32'hbc994714} /* (4, 5, 27) {real, imag} */,
  {32'hbd19b006, 32'h3e0197cf} /* (4, 5, 26) {real, imag} */,
  {32'h3d2aa86c, 32'hbd3b3646} /* (4, 5, 25) {real, imag} */,
  {32'hbd081ebc, 32'hbdbbc6c3} /* (4, 5, 24) {real, imag} */,
  {32'h3caa0a36, 32'hbca8785c} /* (4, 5, 23) {real, imag} */,
  {32'hbcd49294, 32'hbdca2b98} /* (4, 5, 22) {real, imag} */,
  {32'hbd2ba03d, 32'h3d2db562} /* (4, 5, 21) {real, imag} */,
  {32'hbdaed27a, 32'h3b4842c0} /* (4, 5, 20) {real, imag} */,
  {32'hbcd603de, 32'hbd39a88a} /* (4, 5, 19) {real, imag} */,
  {32'h3db5fb9e, 32'h3d574b2b} /* (4, 5, 18) {real, imag} */,
  {32'hbbdd7b89, 32'h3d2d7dfc} /* (4, 5, 17) {real, imag} */,
  {32'h3dc39893, 32'h00000000} /* (4, 5, 16) {real, imag} */,
  {32'hbbdd7b89, 32'hbd2d7dfc} /* (4, 5, 15) {real, imag} */,
  {32'h3db5fb9e, 32'hbd574b2b} /* (4, 5, 14) {real, imag} */,
  {32'hbcd603de, 32'h3d39a88a} /* (4, 5, 13) {real, imag} */,
  {32'hbdaed27a, 32'hbb4842c0} /* (4, 5, 12) {real, imag} */,
  {32'hbd2ba03d, 32'hbd2db562} /* (4, 5, 11) {real, imag} */,
  {32'hbcd49294, 32'h3dca2b98} /* (4, 5, 10) {real, imag} */,
  {32'h3caa0a36, 32'h3ca8785c} /* (4, 5, 9) {real, imag} */,
  {32'hbd081ebc, 32'h3dbbc6c3} /* (4, 5, 8) {real, imag} */,
  {32'h3d2aa86c, 32'h3d3b3646} /* (4, 5, 7) {real, imag} */,
  {32'hbd19b006, 32'hbe0197cf} /* (4, 5, 6) {real, imag} */,
  {32'h3dd43f90, 32'h3c994714} /* (4, 5, 5) {real, imag} */,
  {32'h3cb9ae80, 32'h3e7abb40} /* (4, 5, 4) {real, imag} */,
  {32'h3e77bf44, 32'h3d7cbe94} /* (4, 5, 3) {real, imag} */,
  {32'h3e0cc474, 32'h3c57c73c} /* (4, 5, 2) {real, imag} */,
  {32'hbea0ee50, 32'hbf30aa7a} /* (4, 5, 1) {real, imag} */,
  {32'h3e41d8dd, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'hbe7cbde3, 32'h3f5903e8} /* (4, 4, 31) {real, imag} */,
  {32'hbe026e7f, 32'hbe4f05e7} /* (4, 4, 30) {real, imag} */,
  {32'h3e2fedab, 32'hbd2583e8} /* (4, 4, 29) {real, imag} */,
  {32'h3d7d4370, 32'hbe8b6a0b} /* (4, 4, 28) {real, imag} */,
  {32'h3e8bfed5, 32'h3d3d09bb} /* (4, 4, 27) {real, imag} */,
  {32'h3db0f4fa, 32'hbd8f3344} /* (4, 4, 26) {real, imag} */,
  {32'hbcf168d6, 32'hbdf403d3} /* (4, 4, 25) {real, imag} */,
  {32'hbe452a7e, 32'hbceae17c} /* (4, 4, 24) {real, imag} */,
  {32'hbd359465, 32'h3d5c68b0} /* (4, 4, 23) {real, imag} */,
  {32'hbcaa6a23, 32'hbd14dc7e} /* (4, 4, 22) {real, imag} */,
  {32'h3bea9568, 32'hbda1ca23} /* (4, 4, 21) {real, imag} */,
  {32'h3d0538c0, 32'h3d21951c} /* (4, 4, 20) {real, imag} */,
  {32'h3d64a8ea, 32'h3d4e3f94} /* (4, 4, 19) {real, imag} */,
  {32'hbd9536eb, 32'hbd9e2977} /* (4, 4, 18) {real, imag} */,
  {32'hbb8d76c4, 32'h3c0ec06a} /* (4, 4, 17) {real, imag} */,
  {32'hbc0b4f5e, 32'h00000000} /* (4, 4, 16) {real, imag} */,
  {32'hbb8d76c4, 32'hbc0ec06a} /* (4, 4, 15) {real, imag} */,
  {32'hbd9536eb, 32'h3d9e2977} /* (4, 4, 14) {real, imag} */,
  {32'h3d64a8ea, 32'hbd4e3f94} /* (4, 4, 13) {real, imag} */,
  {32'h3d0538c0, 32'hbd21951c} /* (4, 4, 12) {real, imag} */,
  {32'h3bea9568, 32'h3da1ca23} /* (4, 4, 11) {real, imag} */,
  {32'hbcaa6a23, 32'h3d14dc7e} /* (4, 4, 10) {real, imag} */,
  {32'hbd359465, 32'hbd5c68b0} /* (4, 4, 9) {real, imag} */,
  {32'hbe452a7e, 32'h3ceae17c} /* (4, 4, 8) {real, imag} */,
  {32'hbcf168d6, 32'h3df403d3} /* (4, 4, 7) {real, imag} */,
  {32'h3db0f4fa, 32'h3d8f3344} /* (4, 4, 6) {real, imag} */,
  {32'h3e8bfed5, 32'hbd3d09bb} /* (4, 4, 5) {real, imag} */,
  {32'h3d7d4370, 32'h3e8b6a0b} /* (4, 4, 4) {real, imag} */,
  {32'h3e2fedab, 32'h3d2583e8} /* (4, 4, 3) {real, imag} */,
  {32'hbe026e7f, 32'h3e4f05e7} /* (4, 4, 2) {real, imag} */,
  {32'hbe7cbde3, 32'hbf5903e8} /* (4, 4, 1) {real, imag} */,
  {32'h3e5bbf7b, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'hbdd33e40, 32'h3f49c635} /* (4, 3, 31) {real, imag} */,
  {32'hbeb0a2ee, 32'hbea09109} /* (4, 3, 30) {real, imag} */,
  {32'h3de7886a, 32'h3d9d8ba1} /* (4, 3, 29) {real, imag} */,
  {32'h3d51a26e, 32'hbe9c01ae} /* (4, 3, 28) {real, imag} */,
  {32'h3e9f1eea, 32'h3da19293} /* (4, 3, 27) {real, imag} */,
  {32'h3e0e2cd4, 32'hbe0a3358} /* (4, 3, 26) {real, imag} */,
  {32'h3da4bb50, 32'h3d35faa8} /* (4, 3, 25) {real, imag} */,
  {32'hbe02b846, 32'h3d6309f5} /* (4, 3, 24) {real, imag} */,
  {32'hbd21af9a, 32'hbd53b53e} /* (4, 3, 23) {real, imag} */,
  {32'hbc7057bf, 32'h3da73662} /* (4, 3, 22) {real, imag} */,
  {32'h3c18db7e, 32'hbb197d00} /* (4, 3, 21) {real, imag} */,
  {32'h3d258621, 32'hbd23314d} /* (4, 3, 20) {real, imag} */,
  {32'h3cbf94f8, 32'h3ba1a298} /* (4, 3, 19) {real, imag} */,
  {32'h3c5b2c64, 32'hbd058a46} /* (4, 3, 18) {real, imag} */,
  {32'h3d1d7f33, 32'hbd22af3e} /* (4, 3, 17) {real, imag} */,
  {32'hbc4f0c4a, 32'h00000000} /* (4, 3, 16) {real, imag} */,
  {32'h3d1d7f33, 32'h3d22af3e} /* (4, 3, 15) {real, imag} */,
  {32'h3c5b2c64, 32'h3d058a46} /* (4, 3, 14) {real, imag} */,
  {32'h3cbf94f8, 32'hbba1a298} /* (4, 3, 13) {real, imag} */,
  {32'h3d258621, 32'h3d23314d} /* (4, 3, 12) {real, imag} */,
  {32'h3c18db7e, 32'h3b197d00} /* (4, 3, 11) {real, imag} */,
  {32'hbc7057bf, 32'hbda73662} /* (4, 3, 10) {real, imag} */,
  {32'hbd21af9a, 32'h3d53b53e} /* (4, 3, 9) {real, imag} */,
  {32'hbe02b846, 32'hbd6309f5} /* (4, 3, 8) {real, imag} */,
  {32'h3da4bb50, 32'hbd35faa8} /* (4, 3, 7) {real, imag} */,
  {32'h3e0e2cd4, 32'h3e0a3358} /* (4, 3, 6) {real, imag} */,
  {32'h3e9f1eea, 32'hbda19293} /* (4, 3, 5) {real, imag} */,
  {32'h3d51a26e, 32'h3e9c01ae} /* (4, 3, 4) {real, imag} */,
  {32'h3de7886a, 32'hbd9d8ba1} /* (4, 3, 3) {real, imag} */,
  {32'hbeb0a2ee, 32'h3ea09109} /* (4, 3, 2) {real, imag} */,
  {32'hbdd33e40, 32'hbf49c635} /* (4, 3, 1) {real, imag} */,
  {32'h3ee68661, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'hbdc54276, 32'h3f3d54ac} /* (4, 2, 31) {real, imag} */,
  {32'hbeaebfe1, 32'hbec56f14} /* (4, 2, 30) {real, imag} */,
  {32'h3ddd65d3, 32'h3d94792e} /* (4, 2, 29) {real, imag} */,
  {32'h3e46066a, 32'hbeac8e89} /* (4, 2, 28) {real, imag} */,
  {32'h3dad787a, 32'hbd59e396} /* (4, 2, 27) {real, imag} */,
  {32'h3d03f3fa, 32'h3d84bf2d} /* (4, 2, 26) {real, imag} */,
  {32'hbb796950, 32'h3d4ac0f7} /* (4, 2, 25) {real, imag} */,
  {32'h3cf51c06, 32'hbc2abd24} /* (4, 2, 24) {real, imag} */,
  {32'h3c4796ec, 32'h3da2fdbb} /* (4, 2, 23) {real, imag} */,
  {32'hbd8f49d6, 32'hbe0f8986} /* (4, 2, 22) {real, imag} */,
  {32'h3d6ff39c, 32'h3d5dc4ae} /* (4, 2, 21) {real, imag} */,
  {32'hbc1cac04, 32'hbc900992} /* (4, 2, 20) {real, imag} */,
  {32'h3e06c5b4, 32'hbda6a6b3} /* (4, 2, 19) {real, imag} */,
  {32'hbd19ddf1, 32'hbb6f42d0} /* (4, 2, 18) {real, imag} */,
  {32'hbc880eea, 32'hbd8639f0} /* (4, 2, 17) {real, imag} */,
  {32'h3cbec5c0, 32'h00000000} /* (4, 2, 16) {real, imag} */,
  {32'hbc880eea, 32'h3d8639f0} /* (4, 2, 15) {real, imag} */,
  {32'hbd19ddf1, 32'h3b6f42d0} /* (4, 2, 14) {real, imag} */,
  {32'h3e06c5b4, 32'h3da6a6b3} /* (4, 2, 13) {real, imag} */,
  {32'hbc1cac04, 32'h3c900992} /* (4, 2, 12) {real, imag} */,
  {32'h3d6ff39c, 32'hbd5dc4ae} /* (4, 2, 11) {real, imag} */,
  {32'hbd8f49d6, 32'h3e0f8986} /* (4, 2, 10) {real, imag} */,
  {32'h3c4796ec, 32'hbda2fdbb} /* (4, 2, 9) {real, imag} */,
  {32'h3cf51c06, 32'h3c2abd24} /* (4, 2, 8) {real, imag} */,
  {32'hbb796950, 32'hbd4ac0f7} /* (4, 2, 7) {real, imag} */,
  {32'h3d03f3fa, 32'hbd84bf2d} /* (4, 2, 6) {real, imag} */,
  {32'h3dad787a, 32'h3d59e396} /* (4, 2, 5) {real, imag} */,
  {32'h3e46066a, 32'h3eac8e89} /* (4, 2, 4) {real, imag} */,
  {32'h3ddd65d3, 32'hbd94792e} /* (4, 2, 3) {real, imag} */,
  {32'hbeaebfe1, 32'h3ec56f14} /* (4, 2, 2) {real, imag} */,
  {32'hbdc54276, 32'hbf3d54ac} /* (4, 2, 1) {real, imag} */,
  {32'h3f176c58, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'hbd3221c0, 32'h3f2a75e5} /* (4, 1, 31) {real, imag} */,
  {32'hbe483878, 32'hbee12f36} /* (4, 1, 30) {real, imag} */,
  {32'h3e06deac, 32'hbcab8082} /* (4, 1, 29) {real, imag} */,
  {32'h3e5236bf, 32'hbe4951ce} /* (4, 1, 28) {real, imag} */,
  {32'h3e5d437c, 32'h3e07b2c0} /* (4, 1, 27) {real, imag} */,
  {32'hbcc2d56e, 32'h3c43c248} /* (4, 1, 26) {real, imag} */,
  {32'hbca0201a, 32'h3d55830a} /* (4, 1, 25) {real, imag} */,
  {32'hbe0c8314, 32'h3c7f8b0c} /* (4, 1, 24) {real, imag} */,
  {32'hbd6a2d9d, 32'hbe03f6df} /* (4, 1, 23) {real, imag} */,
  {32'h3ddba704, 32'hbd934bb4} /* (4, 1, 22) {real, imag} */,
  {32'hbd0aabc5, 32'h3c8937c4} /* (4, 1, 21) {real, imag} */,
  {32'hbcac2866, 32'h3cc9bf20} /* (4, 1, 20) {real, imag} */,
  {32'h3b00a584, 32'hbcf0dfd5} /* (4, 1, 19) {real, imag} */,
  {32'hbd4aef48, 32'hbbe7b374} /* (4, 1, 18) {real, imag} */,
  {32'h3d3061c2, 32'h3d60fdec} /* (4, 1, 17) {real, imag} */,
  {32'h3d2221d8, 32'h00000000} /* (4, 1, 16) {real, imag} */,
  {32'h3d3061c2, 32'hbd60fdec} /* (4, 1, 15) {real, imag} */,
  {32'hbd4aef48, 32'h3be7b374} /* (4, 1, 14) {real, imag} */,
  {32'h3b00a584, 32'h3cf0dfd5} /* (4, 1, 13) {real, imag} */,
  {32'hbcac2866, 32'hbcc9bf20} /* (4, 1, 12) {real, imag} */,
  {32'hbd0aabc5, 32'hbc8937c4} /* (4, 1, 11) {real, imag} */,
  {32'h3ddba704, 32'h3d934bb4} /* (4, 1, 10) {real, imag} */,
  {32'hbd6a2d9d, 32'h3e03f6df} /* (4, 1, 9) {real, imag} */,
  {32'hbe0c8314, 32'hbc7f8b0c} /* (4, 1, 8) {real, imag} */,
  {32'hbca0201a, 32'hbd55830a} /* (4, 1, 7) {real, imag} */,
  {32'hbcc2d56e, 32'hbc43c248} /* (4, 1, 6) {real, imag} */,
  {32'h3e5d437c, 32'hbe07b2c0} /* (4, 1, 5) {real, imag} */,
  {32'h3e5236bf, 32'h3e4951ce} /* (4, 1, 4) {real, imag} */,
  {32'h3e06deac, 32'h3cab8082} /* (4, 1, 3) {real, imag} */,
  {32'hbe483878, 32'h3ee12f36} /* (4, 1, 2) {real, imag} */,
  {32'hbd3221c0, 32'hbf2a75e5} /* (4, 1, 1) {real, imag} */,
  {32'h3f444fac, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'hbd7bf8b8, 32'h3eba1aa6} /* (4, 0, 31) {real, imag} */,
  {32'h3c9bc570, 32'hbea8660a} /* (4, 0, 30) {real, imag} */,
  {32'h3d4a2e52, 32'hbd22c478} /* (4, 0, 29) {real, imag} */,
  {32'h3d8129c8, 32'hbe1bb62e} /* (4, 0, 28) {real, imag} */,
  {32'h3e55c92e, 32'h3da5c08d} /* (4, 0, 27) {real, imag} */,
  {32'hbb5acb08, 32'h39624680} /* (4, 0, 26) {real, imag} */,
  {32'hbd29663b, 32'hbc6b1e80} /* (4, 0, 25) {real, imag} */,
  {32'hbdcd60dc, 32'hbc8ffd64} /* (4, 0, 24) {real, imag} */,
  {32'hbd2d4d1b, 32'hbe057d21} /* (4, 0, 23) {real, imag} */,
  {32'hbbd0494c, 32'hbd53f12f} /* (4, 0, 22) {real, imag} */,
  {32'hbd6fe052, 32'h3daa142c} /* (4, 0, 21) {real, imag} */,
  {32'h3d06ac6a, 32'h3cbbbe14} /* (4, 0, 20) {real, imag} */,
  {32'hbd24dffc, 32'h3b516cc4} /* (4, 0, 19) {real, imag} */,
  {32'h3ab9c900, 32'hbd02ed28} /* (4, 0, 18) {real, imag} */,
  {32'h3c8ede9a, 32'h3d1df923} /* (4, 0, 17) {real, imag} */,
  {32'h3cc5448c, 32'h00000000} /* (4, 0, 16) {real, imag} */,
  {32'h3c8ede9a, 32'hbd1df923} /* (4, 0, 15) {real, imag} */,
  {32'h3ab9c900, 32'h3d02ed28} /* (4, 0, 14) {real, imag} */,
  {32'hbd24dffc, 32'hbb516cc4} /* (4, 0, 13) {real, imag} */,
  {32'h3d06ac6a, 32'hbcbbbe14} /* (4, 0, 12) {real, imag} */,
  {32'hbd6fe052, 32'hbdaa142c} /* (4, 0, 11) {real, imag} */,
  {32'hbbd0494c, 32'h3d53f12f} /* (4, 0, 10) {real, imag} */,
  {32'hbd2d4d1b, 32'h3e057d21} /* (4, 0, 9) {real, imag} */,
  {32'hbdcd60dc, 32'h3c8ffd64} /* (4, 0, 8) {real, imag} */,
  {32'hbd29663b, 32'h3c6b1e80} /* (4, 0, 7) {real, imag} */,
  {32'hbb5acb08, 32'hb9624680} /* (4, 0, 6) {real, imag} */,
  {32'h3e55c92e, 32'hbda5c08d} /* (4, 0, 5) {real, imag} */,
  {32'h3d8129c8, 32'h3e1bb62e} /* (4, 0, 4) {real, imag} */,
  {32'h3d4a2e52, 32'h3d22c478} /* (4, 0, 3) {real, imag} */,
  {32'h3c9bc570, 32'h3ea8660a} /* (4, 0, 2) {real, imag} */,
  {32'hbd7bf8b8, 32'hbeba1aa6} /* (4, 0, 1) {real, imag} */,
  {32'h3f67531c, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hbf64e8e5, 32'h3ed8b39f} /* (3, 31, 31) {real, imag} */,
  {32'h3eeaa161, 32'hbe8238fd} /* (3, 31, 30) {real, imag} */,
  {32'h3dd16516, 32'hbc8f752c} /* (3, 31, 29) {real, imag} */,
  {32'hbe0246a0, 32'hbe0d597e} /* (3, 31, 28) {real, imag} */,
  {32'h3e2dcc56, 32'hbdd3e0e9} /* (3, 31, 27) {real, imag} */,
  {32'hbcb2a054, 32'hbda723ae} /* (3, 31, 26) {real, imag} */,
  {32'h3ba64d80, 32'h3c2a9c0c} /* (3, 31, 25) {real, imag} */,
  {32'hbd77a12a, 32'hbd09419c} /* (3, 31, 24) {real, imag} */,
  {32'h3d7a42f8, 32'hbcb30842} /* (3, 31, 23) {real, imag} */,
  {32'hbb0365a0, 32'h3d638480} /* (3, 31, 22) {real, imag} */,
  {32'hbce3daff, 32'hbd190182} /* (3, 31, 21) {real, imag} */,
  {32'h3ca1346f, 32'h3cd5e72d} /* (3, 31, 20) {real, imag} */,
  {32'hbdadc98e, 32'hbd7d84f2} /* (3, 31, 19) {real, imag} */,
  {32'h3cb91514, 32'h3d0c226b} /* (3, 31, 18) {real, imag} */,
  {32'h3bf26278, 32'h3cea1c53} /* (3, 31, 17) {real, imag} */,
  {32'h3b926c48, 32'h00000000} /* (3, 31, 16) {real, imag} */,
  {32'h3bf26278, 32'hbcea1c53} /* (3, 31, 15) {real, imag} */,
  {32'h3cb91514, 32'hbd0c226b} /* (3, 31, 14) {real, imag} */,
  {32'hbdadc98e, 32'h3d7d84f2} /* (3, 31, 13) {real, imag} */,
  {32'h3ca1346f, 32'hbcd5e72d} /* (3, 31, 12) {real, imag} */,
  {32'hbce3daff, 32'h3d190182} /* (3, 31, 11) {real, imag} */,
  {32'hbb0365a0, 32'hbd638480} /* (3, 31, 10) {real, imag} */,
  {32'h3d7a42f8, 32'h3cb30842} /* (3, 31, 9) {real, imag} */,
  {32'hbd77a12a, 32'h3d09419c} /* (3, 31, 8) {real, imag} */,
  {32'h3ba64d80, 32'hbc2a9c0c} /* (3, 31, 7) {real, imag} */,
  {32'hbcb2a054, 32'h3da723ae} /* (3, 31, 6) {real, imag} */,
  {32'h3e2dcc56, 32'h3dd3e0e9} /* (3, 31, 5) {real, imag} */,
  {32'hbe0246a0, 32'h3e0d597e} /* (3, 31, 4) {real, imag} */,
  {32'h3dd16516, 32'h3c8f752c} /* (3, 31, 3) {real, imag} */,
  {32'h3eeaa161, 32'h3e8238fd} /* (3, 31, 2) {real, imag} */,
  {32'hbf64e8e5, 32'hbed8b39f} /* (3, 31, 1) {real, imag} */,
  {32'h3cd7d49e, 32'h00000000} /* (3, 31, 0) {real, imag} */,
  {32'hbf983df4, 32'h3e86d55a} /* (3, 30, 31) {real, imag} */,
  {32'h3f57da4c, 32'hbe53431e} /* (3, 30, 30) {real, imag} */,
  {32'h3e463afb, 32'hbcb69f1c} /* (3, 30, 29) {real, imag} */,
  {32'hbe1baa64, 32'hbd848804} /* (3, 30, 28) {real, imag} */,
  {32'h3e7563da, 32'hbe59921c} /* (3, 30, 27) {real, imag} */,
  {32'h3be25a40, 32'h3c09adc0} /* (3, 30, 26) {real, imag} */,
  {32'hbc9cbeb6, 32'h3d8632f2} /* (3, 30, 25) {real, imag} */,
  {32'h3dc11a11, 32'hbc8f0f85} /* (3, 30, 24) {real, imag} */,
  {32'h3d5f6dc4, 32'h3e17cb78} /* (3, 30, 23) {real, imag} */,
  {32'hbb70a2a8, 32'h3b2d6140} /* (3, 30, 22) {real, imag} */,
  {32'hbccd7c04, 32'hbd9b9352} /* (3, 30, 21) {real, imag} */,
  {32'h3d778514, 32'h3c7b58f6} /* (3, 30, 20) {real, imag} */,
  {32'h3d8c57e9, 32'h3d51aafc} /* (3, 30, 19) {real, imag} */,
  {32'h3ce8059c, 32'h3c521cfc} /* (3, 30, 18) {real, imag} */,
  {32'hbb9f8030, 32'h3d212b86} /* (3, 30, 17) {real, imag} */,
  {32'hbcf60225, 32'h00000000} /* (3, 30, 16) {real, imag} */,
  {32'hbb9f8030, 32'hbd212b86} /* (3, 30, 15) {real, imag} */,
  {32'h3ce8059c, 32'hbc521cfc} /* (3, 30, 14) {real, imag} */,
  {32'h3d8c57e9, 32'hbd51aafc} /* (3, 30, 13) {real, imag} */,
  {32'h3d778514, 32'hbc7b58f6} /* (3, 30, 12) {real, imag} */,
  {32'hbccd7c04, 32'h3d9b9352} /* (3, 30, 11) {real, imag} */,
  {32'hbb70a2a8, 32'hbb2d6140} /* (3, 30, 10) {real, imag} */,
  {32'h3d5f6dc4, 32'hbe17cb78} /* (3, 30, 9) {real, imag} */,
  {32'h3dc11a11, 32'h3c8f0f85} /* (3, 30, 8) {real, imag} */,
  {32'hbc9cbeb6, 32'hbd8632f2} /* (3, 30, 7) {real, imag} */,
  {32'h3be25a40, 32'hbc09adc0} /* (3, 30, 6) {real, imag} */,
  {32'h3e7563da, 32'h3e59921c} /* (3, 30, 5) {real, imag} */,
  {32'hbe1baa64, 32'h3d848804} /* (3, 30, 4) {real, imag} */,
  {32'h3e463afb, 32'h3cb69f1c} /* (3, 30, 3) {real, imag} */,
  {32'h3f57da4c, 32'h3e53431e} /* (3, 30, 2) {real, imag} */,
  {32'hbf983df4, 32'hbe86d55a} /* (3, 30, 1) {real, imag} */,
  {32'hbe0eb332, 32'h00000000} /* (3, 30, 0) {real, imag} */,
  {32'hbfbd00cc, 32'h3e5842d4} /* (3, 29, 31) {real, imag} */,
  {32'h3f72b250, 32'hbd3b4328} /* (3, 29, 30) {real, imag} */,
  {32'h3e62d306, 32'hbe0d97c6} /* (3, 29, 29) {real, imag} */,
  {32'hbe5d244b, 32'h3dffad80} /* (3, 29, 28) {real, imag} */,
  {32'h3e8449e0, 32'hbe2054c2} /* (3, 29, 27) {real, imag} */,
  {32'h3d9b8a0d, 32'h3e33170f} /* (3, 29, 26) {real, imag} */,
  {32'hbdbdf93e, 32'h3dd9092a} /* (3, 29, 25) {real, imag} */,
  {32'h3ddb7598, 32'hbdb5def2} /* (3, 29, 24) {real, imag} */,
  {32'hbdac9462, 32'h3e28aa4d} /* (3, 29, 23) {real, imag} */,
  {32'hbc7a43e6, 32'hbd972daf} /* (3, 29, 22) {real, imag} */,
  {32'h3ddf393c, 32'hbde00074} /* (3, 29, 21) {real, imag} */,
  {32'h3cfa2d05, 32'hbcb4b24b} /* (3, 29, 20) {real, imag} */,
  {32'h3cbaf6b6, 32'hbdaa9ae8} /* (3, 29, 19) {real, imag} */,
  {32'hbd0af8d4, 32'h3d939178} /* (3, 29, 18) {real, imag} */,
  {32'h3d085812, 32'hbc3a4b5c} /* (3, 29, 17) {real, imag} */,
  {32'h3d3092ee, 32'h00000000} /* (3, 29, 16) {real, imag} */,
  {32'h3d085812, 32'h3c3a4b5c} /* (3, 29, 15) {real, imag} */,
  {32'hbd0af8d4, 32'hbd939178} /* (3, 29, 14) {real, imag} */,
  {32'h3cbaf6b6, 32'h3daa9ae8} /* (3, 29, 13) {real, imag} */,
  {32'h3cfa2d05, 32'h3cb4b24b} /* (3, 29, 12) {real, imag} */,
  {32'h3ddf393c, 32'h3de00074} /* (3, 29, 11) {real, imag} */,
  {32'hbc7a43e6, 32'h3d972daf} /* (3, 29, 10) {real, imag} */,
  {32'hbdac9462, 32'hbe28aa4d} /* (3, 29, 9) {real, imag} */,
  {32'h3ddb7598, 32'h3db5def2} /* (3, 29, 8) {real, imag} */,
  {32'hbdbdf93e, 32'hbdd9092a} /* (3, 29, 7) {real, imag} */,
  {32'h3d9b8a0d, 32'hbe33170f} /* (3, 29, 6) {real, imag} */,
  {32'h3e8449e0, 32'h3e2054c2} /* (3, 29, 5) {real, imag} */,
  {32'hbe5d244b, 32'hbdffad80} /* (3, 29, 4) {real, imag} */,
  {32'h3e62d306, 32'h3e0d97c6} /* (3, 29, 3) {real, imag} */,
  {32'h3f72b250, 32'h3d3b4328} /* (3, 29, 2) {real, imag} */,
  {32'hbfbd00cc, 32'hbe5842d4} /* (3, 29, 1) {real, imag} */,
  {32'hbd5f7230, 32'h00000000} /* (3, 29, 0) {real, imag} */,
  {32'hbfc60a33, 32'h3e5154b4} /* (3, 28, 31) {real, imag} */,
  {32'h3f6e40ac, 32'hbd4e5490} /* (3, 28, 30) {real, imag} */,
  {32'h3e07166b, 32'hbda4d3f2} /* (3, 28, 29) {real, imag} */,
  {32'hbdc47b8a, 32'h3d43be18} /* (3, 28, 28) {real, imag} */,
  {32'h3e78983f, 32'hbe40c61a} /* (3, 28, 27) {real, imag} */,
  {32'h3d2ab758, 32'hbd1c5139} /* (3, 28, 26) {real, imag} */,
  {32'hbe0c9add, 32'h3db233f3} /* (3, 28, 25) {real, imag} */,
  {32'h3da0e498, 32'hbcbe1a17} /* (3, 28, 24) {real, imag} */,
  {32'hbdb898f0, 32'h3d7ed28d} /* (3, 28, 23) {real, imag} */,
  {32'h3d9eb91b, 32'h3c274fbc} /* (3, 28, 22) {real, imag} */,
  {32'h3d9f8baa, 32'hbda8f441} /* (3, 28, 21) {real, imag} */,
  {32'hbd9852e0, 32'h3c561e40} /* (3, 28, 20) {real, imag} */,
  {32'hbda02b6a, 32'hbd7f8bd8} /* (3, 28, 19) {real, imag} */,
  {32'hbcca87a2, 32'h3d7e4d03} /* (3, 28, 18) {real, imag} */,
  {32'hbc9752c4, 32'hbd580c38} /* (3, 28, 17) {real, imag} */,
  {32'h3d99997a, 32'h00000000} /* (3, 28, 16) {real, imag} */,
  {32'hbc9752c4, 32'h3d580c38} /* (3, 28, 15) {real, imag} */,
  {32'hbcca87a2, 32'hbd7e4d03} /* (3, 28, 14) {real, imag} */,
  {32'hbda02b6a, 32'h3d7f8bd8} /* (3, 28, 13) {real, imag} */,
  {32'hbd9852e0, 32'hbc561e40} /* (3, 28, 12) {real, imag} */,
  {32'h3d9f8baa, 32'h3da8f441} /* (3, 28, 11) {real, imag} */,
  {32'h3d9eb91b, 32'hbc274fbc} /* (3, 28, 10) {real, imag} */,
  {32'hbdb898f0, 32'hbd7ed28d} /* (3, 28, 9) {real, imag} */,
  {32'h3da0e498, 32'h3cbe1a17} /* (3, 28, 8) {real, imag} */,
  {32'hbe0c9add, 32'hbdb233f3} /* (3, 28, 7) {real, imag} */,
  {32'h3d2ab758, 32'h3d1c5139} /* (3, 28, 6) {real, imag} */,
  {32'h3e78983f, 32'h3e40c61a} /* (3, 28, 5) {real, imag} */,
  {32'hbdc47b8a, 32'hbd43be18} /* (3, 28, 4) {real, imag} */,
  {32'h3e07166b, 32'h3da4d3f2} /* (3, 28, 3) {real, imag} */,
  {32'h3f6e40ac, 32'h3d4e5490} /* (3, 28, 2) {real, imag} */,
  {32'hbfc60a33, 32'hbe5154b4} /* (3, 28, 1) {real, imag} */,
  {32'hbe0a229e, 32'h00000000} /* (3, 28, 0) {real, imag} */,
  {32'hbfc9d310, 32'h3e5365fc} /* (3, 27, 31) {real, imag} */,
  {32'h3f6699d0, 32'hbe0c634a} /* (3, 27, 30) {real, imag} */,
  {32'h3de74080, 32'hbe38f329} /* (3, 27, 29) {real, imag} */,
  {32'hbe709a96, 32'h3cb0a880} /* (3, 27, 28) {real, imag} */,
  {32'h3e9e1683, 32'hbdb9de13} /* (3, 27, 27) {real, imag} */,
  {32'hbda52ffb, 32'h3b9d7162} /* (3, 27, 26) {real, imag} */,
  {32'hbd00996a, 32'hbc529380} /* (3, 27, 25) {real, imag} */,
  {32'h3df3aa50, 32'hbccb8dba} /* (3, 27, 24) {real, imag} */,
  {32'h3be57340, 32'hbc5b1bba} /* (3, 27, 23) {real, imag} */,
  {32'hbd5be0ca, 32'hbd6601e4} /* (3, 27, 22) {real, imag} */,
  {32'h3b748b90, 32'hbca6d175} /* (3, 27, 21) {real, imag} */,
  {32'h3d99027f, 32'h3bd178ac} /* (3, 27, 20) {real, imag} */,
  {32'h3cc357c6, 32'hbd423ca3} /* (3, 27, 19) {real, imag} */,
  {32'h3d47b34c, 32'hbc8fec66} /* (3, 27, 18) {real, imag} */,
  {32'h3e0658ff, 32'h3d377bb4} /* (3, 27, 17) {real, imag} */,
  {32'hbd4cd1be, 32'h00000000} /* (3, 27, 16) {real, imag} */,
  {32'h3e0658ff, 32'hbd377bb4} /* (3, 27, 15) {real, imag} */,
  {32'h3d47b34c, 32'h3c8fec66} /* (3, 27, 14) {real, imag} */,
  {32'h3cc357c6, 32'h3d423ca3} /* (3, 27, 13) {real, imag} */,
  {32'h3d99027f, 32'hbbd178ac} /* (3, 27, 12) {real, imag} */,
  {32'h3b748b90, 32'h3ca6d175} /* (3, 27, 11) {real, imag} */,
  {32'hbd5be0ca, 32'h3d6601e4} /* (3, 27, 10) {real, imag} */,
  {32'h3be57340, 32'h3c5b1bba} /* (3, 27, 9) {real, imag} */,
  {32'h3df3aa50, 32'h3ccb8dba} /* (3, 27, 8) {real, imag} */,
  {32'hbd00996a, 32'h3c529380} /* (3, 27, 7) {real, imag} */,
  {32'hbda52ffb, 32'hbb9d7162} /* (3, 27, 6) {real, imag} */,
  {32'h3e9e1683, 32'h3db9de13} /* (3, 27, 5) {real, imag} */,
  {32'hbe709a96, 32'hbcb0a880} /* (3, 27, 4) {real, imag} */,
  {32'h3de74080, 32'h3e38f329} /* (3, 27, 3) {real, imag} */,
  {32'h3f6699d0, 32'h3e0c634a} /* (3, 27, 2) {real, imag} */,
  {32'hbfc9d310, 32'hbe5365fc} /* (3, 27, 1) {real, imag} */,
  {32'hbe642319, 32'h00000000} /* (3, 27, 0) {real, imag} */,
  {32'hbfd83ec4, 32'h3e5de436} /* (3, 26, 31) {real, imag} */,
  {32'h3f78e066, 32'hbd66a843} /* (3, 26, 30) {real, imag} */,
  {32'h3dbfee93, 32'hbe47d18a} /* (3, 26, 29) {real, imag} */,
  {32'hbe9c720a, 32'h3d3e5144} /* (3, 26, 28) {real, imag} */,
  {32'h3e492139, 32'hbc5ad504} /* (3, 26, 27) {real, imag} */,
  {32'h3d617054, 32'hbdc52d30} /* (3, 26, 26) {real, imag} */,
  {32'hbd613278, 32'h3c096d74} /* (3, 26, 25) {real, imag} */,
  {32'h3d28939b, 32'hbdc6f64a} /* (3, 26, 24) {real, imag} */,
  {32'h3da881f0, 32'hbd86f9f6} /* (3, 26, 23) {real, imag} */,
  {32'h3c192288, 32'h3c487a1c} /* (3, 26, 22) {real, imag} */,
  {32'h3d732255, 32'h3d4a39f3} /* (3, 26, 21) {real, imag} */,
  {32'hbdfcb133, 32'h3cfef283} /* (3, 26, 20) {real, imag} */,
  {32'h3c0e4e88, 32'h3d85a1e1} /* (3, 26, 19) {real, imag} */,
  {32'hbd5cca30, 32'hb94c1c80} /* (3, 26, 18) {real, imag} */,
  {32'h3d03b766, 32'h3c8f1328} /* (3, 26, 17) {real, imag} */,
  {32'h3ccff680, 32'h00000000} /* (3, 26, 16) {real, imag} */,
  {32'h3d03b766, 32'hbc8f1328} /* (3, 26, 15) {real, imag} */,
  {32'hbd5cca30, 32'h394c1c80} /* (3, 26, 14) {real, imag} */,
  {32'h3c0e4e88, 32'hbd85a1e1} /* (3, 26, 13) {real, imag} */,
  {32'hbdfcb133, 32'hbcfef283} /* (3, 26, 12) {real, imag} */,
  {32'h3d732255, 32'hbd4a39f3} /* (3, 26, 11) {real, imag} */,
  {32'h3c192288, 32'hbc487a1c} /* (3, 26, 10) {real, imag} */,
  {32'h3da881f0, 32'h3d86f9f6} /* (3, 26, 9) {real, imag} */,
  {32'h3d28939b, 32'h3dc6f64a} /* (3, 26, 8) {real, imag} */,
  {32'hbd613278, 32'hbc096d74} /* (3, 26, 7) {real, imag} */,
  {32'h3d617054, 32'h3dc52d30} /* (3, 26, 6) {real, imag} */,
  {32'h3e492139, 32'h3c5ad504} /* (3, 26, 5) {real, imag} */,
  {32'hbe9c720a, 32'hbd3e5144} /* (3, 26, 4) {real, imag} */,
  {32'h3dbfee93, 32'h3e47d18a} /* (3, 26, 3) {real, imag} */,
  {32'h3f78e066, 32'h3d66a843} /* (3, 26, 2) {real, imag} */,
  {32'hbfd83ec4, 32'hbe5de436} /* (3, 26, 1) {real, imag} */,
  {32'hbe236832, 32'h00000000} /* (3, 26, 0) {real, imag} */,
  {32'hbfede8f4, 32'h3e3fbcd6} /* (3, 25, 31) {real, imag} */,
  {32'h3f812c05, 32'h3cbb38a0} /* (3, 25, 30) {real, imag} */,
  {32'h3dd32e56, 32'hbe07a146} /* (3, 25, 29) {real, imag} */,
  {32'hbe47106c, 32'h3cf149f4} /* (3, 25, 28) {real, imag} */,
  {32'h3e1e3a0e, 32'hbe2c0cad} /* (3, 25, 27) {real, imag} */,
  {32'h3ac1e6a0, 32'hbdc32ee0} /* (3, 25, 26) {real, imag} */,
  {32'hbde919e4, 32'h3d4a8a59} /* (3, 25, 25) {real, imag} */,
  {32'h3d0b5d14, 32'hbdafcd1f} /* (3, 25, 24) {real, imag} */,
  {32'h3d95f0de, 32'hbcca3ede} /* (3, 25, 23) {real, imag} */,
  {32'hbc8d4860, 32'hbcbb3a96} /* (3, 25, 22) {real, imag} */,
  {32'h3d886f5e, 32'hbc2f97d8} /* (3, 25, 21) {real, imag} */,
  {32'hbd23cc10, 32'h3d2221d9} /* (3, 25, 20) {real, imag} */,
  {32'h3d81c768, 32'h3d3881c7} /* (3, 25, 19) {real, imag} */,
  {32'h3c165097, 32'h3d52cedd} /* (3, 25, 18) {real, imag} */,
  {32'hbd1646fc, 32'hbd9c29c6} /* (3, 25, 17) {real, imag} */,
  {32'hbc1dfd8a, 32'h00000000} /* (3, 25, 16) {real, imag} */,
  {32'hbd1646fc, 32'h3d9c29c6} /* (3, 25, 15) {real, imag} */,
  {32'h3c165097, 32'hbd52cedd} /* (3, 25, 14) {real, imag} */,
  {32'h3d81c768, 32'hbd3881c7} /* (3, 25, 13) {real, imag} */,
  {32'hbd23cc10, 32'hbd2221d9} /* (3, 25, 12) {real, imag} */,
  {32'h3d886f5e, 32'h3c2f97d8} /* (3, 25, 11) {real, imag} */,
  {32'hbc8d4860, 32'h3cbb3a96} /* (3, 25, 10) {real, imag} */,
  {32'h3d95f0de, 32'h3cca3ede} /* (3, 25, 9) {real, imag} */,
  {32'h3d0b5d14, 32'h3dafcd1f} /* (3, 25, 8) {real, imag} */,
  {32'hbde919e4, 32'hbd4a8a59} /* (3, 25, 7) {real, imag} */,
  {32'h3ac1e6a0, 32'h3dc32ee0} /* (3, 25, 6) {real, imag} */,
  {32'h3e1e3a0e, 32'h3e2c0cad} /* (3, 25, 5) {real, imag} */,
  {32'hbe47106c, 32'hbcf149f4} /* (3, 25, 4) {real, imag} */,
  {32'h3dd32e56, 32'h3e07a146} /* (3, 25, 3) {real, imag} */,
  {32'h3f812c05, 32'hbcbb38a0} /* (3, 25, 2) {real, imag} */,
  {32'hbfede8f4, 32'hbe3fbcd6} /* (3, 25, 1) {real, imag} */,
  {32'hbe9b0aa2, 32'h00000000} /* (3, 25, 0) {real, imag} */,
  {32'hbfedb06b, 32'h3e511e32} /* (3, 24, 31) {real, imag} */,
  {32'h3f66a370, 32'h3cb6199e} /* (3, 24, 30) {real, imag} */,
  {32'h3d0b2e12, 32'hbccb1bfc} /* (3, 24, 29) {real, imag} */,
  {32'hbe7cba0e, 32'h3c2e56cc} /* (3, 24, 28) {real, imag} */,
  {32'h3e44bbfb, 32'hbdd0d414} /* (3, 24, 27) {real, imag} */,
  {32'h3d8be9ac, 32'hbd523243} /* (3, 24, 26) {real, imag} */,
  {32'hbd31a31e, 32'hbc651a56} /* (3, 24, 25) {real, imag} */,
  {32'hbbdc4d2c, 32'hbdb60d2c} /* (3, 24, 24) {real, imag} */,
  {32'h3d43f84c, 32'h3c977534} /* (3, 24, 23) {real, imag} */,
  {32'hbdbbcd6c, 32'h3dae5dc5} /* (3, 24, 22) {real, imag} */,
  {32'h3dd7fe55, 32'h3c737994} /* (3, 24, 21) {real, imag} */,
  {32'h3c736e20, 32'hbce90599} /* (3, 24, 20) {real, imag} */,
  {32'hbba1056c, 32'hbe5541de} /* (3, 24, 19) {real, imag} */,
  {32'hbd21a9ed, 32'hbc536e5a} /* (3, 24, 18) {real, imag} */,
  {32'hbe06af85, 32'hbbc66b97} /* (3, 24, 17) {real, imag} */,
  {32'h3b45d0ac, 32'h00000000} /* (3, 24, 16) {real, imag} */,
  {32'hbe06af85, 32'h3bc66b97} /* (3, 24, 15) {real, imag} */,
  {32'hbd21a9ed, 32'h3c536e5a} /* (3, 24, 14) {real, imag} */,
  {32'hbba1056c, 32'h3e5541de} /* (3, 24, 13) {real, imag} */,
  {32'h3c736e20, 32'h3ce90599} /* (3, 24, 12) {real, imag} */,
  {32'h3dd7fe55, 32'hbc737994} /* (3, 24, 11) {real, imag} */,
  {32'hbdbbcd6c, 32'hbdae5dc5} /* (3, 24, 10) {real, imag} */,
  {32'h3d43f84c, 32'hbc977534} /* (3, 24, 9) {real, imag} */,
  {32'hbbdc4d2c, 32'h3db60d2c} /* (3, 24, 8) {real, imag} */,
  {32'hbd31a31e, 32'h3c651a56} /* (3, 24, 7) {real, imag} */,
  {32'h3d8be9ac, 32'h3d523243} /* (3, 24, 6) {real, imag} */,
  {32'h3e44bbfb, 32'h3dd0d414} /* (3, 24, 5) {real, imag} */,
  {32'hbe7cba0e, 32'hbc2e56cc} /* (3, 24, 4) {real, imag} */,
  {32'h3d0b2e12, 32'h3ccb1bfc} /* (3, 24, 3) {real, imag} */,
  {32'h3f66a370, 32'hbcb6199e} /* (3, 24, 2) {real, imag} */,
  {32'hbfedb06b, 32'hbe511e32} /* (3, 24, 1) {real, imag} */,
  {32'hbed3bd76, 32'h00000000} /* (3, 24, 0) {real, imag} */,
  {32'hbfd769aa, 32'h3e06e386} /* (3, 23, 31) {real, imag} */,
  {32'h3f2debbf, 32'hbd2ab350} /* (3, 23, 30) {real, imag} */,
  {32'h3dd8bca6, 32'h3c4571d6} /* (3, 23, 29) {real, imag} */,
  {32'hbe3b26d9, 32'hbd9f1b27} /* (3, 23, 28) {real, imag} */,
  {32'h3e79f7a6, 32'hbe202de2} /* (3, 23, 27) {real, imag} */,
  {32'h3aac2760, 32'hbb411760} /* (3, 23, 26) {real, imag} */,
  {32'hbb00e140, 32'h3d66b118} /* (3, 23, 25) {real, imag} */,
  {32'h3d950894, 32'h3c8b97b2} /* (3, 23, 24) {real, imag} */,
  {32'h3c2b8ce0, 32'h3d6792ae} /* (3, 23, 23) {real, imag} */,
  {32'hbd34cc56, 32'h3dded8f5} /* (3, 23, 22) {real, imag} */,
  {32'h3d23ae14, 32'hbcb461e2} /* (3, 23, 21) {real, imag} */,
  {32'hbd91f9d5, 32'hbc1e07e4} /* (3, 23, 20) {real, imag} */,
  {32'hbde87109, 32'hbc923980} /* (3, 23, 19) {real, imag} */,
  {32'h3d50d4e0, 32'hbd3d2233} /* (3, 23, 18) {real, imag} */,
  {32'h3d3d9566, 32'hbd07efa2} /* (3, 23, 17) {real, imag} */,
  {32'h3d046944, 32'h00000000} /* (3, 23, 16) {real, imag} */,
  {32'h3d3d9566, 32'h3d07efa2} /* (3, 23, 15) {real, imag} */,
  {32'h3d50d4e0, 32'h3d3d2233} /* (3, 23, 14) {real, imag} */,
  {32'hbde87109, 32'h3c923980} /* (3, 23, 13) {real, imag} */,
  {32'hbd91f9d5, 32'h3c1e07e4} /* (3, 23, 12) {real, imag} */,
  {32'h3d23ae14, 32'h3cb461e2} /* (3, 23, 11) {real, imag} */,
  {32'hbd34cc56, 32'hbdded8f5} /* (3, 23, 10) {real, imag} */,
  {32'h3c2b8ce0, 32'hbd6792ae} /* (3, 23, 9) {real, imag} */,
  {32'h3d950894, 32'hbc8b97b2} /* (3, 23, 8) {real, imag} */,
  {32'hbb00e140, 32'hbd66b118} /* (3, 23, 7) {real, imag} */,
  {32'h3aac2760, 32'h3b411760} /* (3, 23, 6) {real, imag} */,
  {32'h3e79f7a6, 32'h3e202de2} /* (3, 23, 5) {real, imag} */,
  {32'hbe3b26d9, 32'h3d9f1b27} /* (3, 23, 4) {real, imag} */,
  {32'h3dd8bca6, 32'hbc4571d6} /* (3, 23, 3) {real, imag} */,
  {32'h3f2debbf, 32'h3d2ab350} /* (3, 23, 2) {real, imag} */,
  {32'hbfd769aa, 32'hbe06e386} /* (3, 23, 1) {real, imag} */,
  {32'hbec0857e, 32'h00000000} /* (3, 23, 0) {real, imag} */,
  {32'hbfaa1683, 32'h3bcad910} /* (3, 22, 31) {real, imag} */,
  {32'h3ef2f46e, 32'h3d51b955} /* (3, 22, 30) {real, imag} */,
  {32'h3dfd9ae9, 32'h3dcaa426} /* (3, 22, 29) {real, imag} */,
  {32'hbdb35828, 32'hbd8e3f91} /* (3, 22, 28) {real, imag} */,
  {32'h3e27262e, 32'hbe0455d6} /* (3, 22, 27) {real, imag} */,
  {32'hbcab80d0, 32'hbc4ff440} /* (3, 22, 26) {real, imag} */,
  {32'h3d5dd04c, 32'hbd8a31fc} /* (3, 22, 25) {real, imag} */,
  {32'h3d3e8e48, 32'h3d586b4d} /* (3, 22, 24) {real, imag} */,
  {32'h3de7374e, 32'hbde43646} /* (3, 22, 23) {real, imag} */,
  {32'h3d68c785, 32'hbc12499f} /* (3, 22, 22) {real, imag} */,
  {32'hbbd73928, 32'hbd99e9e0} /* (3, 22, 21) {real, imag} */,
  {32'h3ac1e1c0, 32'h3d9a1f6c} /* (3, 22, 20) {real, imag} */,
  {32'hbb5f4b60, 32'h3d9d80d9} /* (3, 22, 19) {real, imag} */,
  {32'hbd8edf87, 32'hbd1f8c50} /* (3, 22, 18) {real, imag} */,
  {32'h3cb077c0, 32'hbda3c962} /* (3, 22, 17) {real, imag} */,
  {32'h3cb3e946, 32'h00000000} /* (3, 22, 16) {real, imag} */,
  {32'h3cb077c0, 32'h3da3c962} /* (3, 22, 15) {real, imag} */,
  {32'hbd8edf87, 32'h3d1f8c50} /* (3, 22, 14) {real, imag} */,
  {32'hbb5f4b60, 32'hbd9d80d9} /* (3, 22, 13) {real, imag} */,
  {32'h3ac1e1c0, 32'hbd9a1f6c} /* (3, 22, 12) {real, imag} */,
  {32'hbbd73928, 32'h3d99e9e0} /* (3, 22, 11) {real, imag} */,
  {32'h3d68c785, 32'h3c12499f} /* (3, 22, 10) {real, imag} */,
  {32'h3de7374e, 32'h3de43646} /* (3, 22, 9) {real, imag} */,
  {32'h3d3e8e48, 32'hbd586b4d} /* (3, 22, 8) {real, imag} */,
  {32'h3d5dd04c, 32'h3d8a31fc} /* (3, 22, 7) {real, imag} */,
  {32'hbcab80d0, 32'h3c4ff440} /* (3, 22, 6) {real, imag} */,
  {32'h3e27262e, 32'h3e0455d6} /* (3, 22, 5) {real, imag} */,
  {32'hbdb35828, 32'h3d8e3f91} /* (3, 22, 4) {real, imag} */,
  {32'h3dfd9ae9, 32'hbdcaa426} /* (3, 22, 3) {real, imag} */,
  {32'h3ef2f46e, 32'hbd51b955} /* (3, 22, 2) {real, imag} */,
  {32'hbfaa1683, 32'hbbcad910} /* (3, 22, 1) {real, imag} */,
  {32'hbeb6df4d, 32'h00000000} /* (3, 22, 0) {real, imag} */,
  {32'hbedbf8a2, 32'hbe2e74f4} /* (3, 21, 31) {real, imag} */,
  {32'h3e202238, 32'hbd064858} /* (3, 21, 30) {real, imag} */,
  {32'hbd81a59e, 32'hbd47b68f} /* (3, 21, 29) {real, imag} */,
  {32'h3d63dc2e, 32'hbdd23f48} /* (3, 21, 28) {real, imag} */,
  {32'h3d95ad7c, 32'hbe003f30} /* (3, 21, 27) {real, imag} */,
  {32'hbd0e735f, 32'h3d8790fd} /* (3, 21, 26) {real, imag} */,
  {32'hbdc17232, 32'h3d8f5583} /* (3, 21, 25) {real, imag} */,
  {32'h3aa72650, 32'h3d939d9a} /* (3, 21, 24) {real, imag} */,
  {32'h3dcb74d7, 32'hbcb344a4} /* (3, 21, 23) {real, imag} */,
  {32'h3d6ae4d5, 32'h3d15a894} /* (3, 21, 22) {real, imag} */,
  {32'hbdb92c74, 32'hbb071d10} /* (3, 21, 21) {real, imag} */,
  {32'h3d0ddc2a, 32'hbcc51581} /* (3, 21, 20) {real, imag} */,
  {32'hbc99ab76, 32'hbd76a5ca} /* (3, 21, 19) {real, imag} */,
  {32'hbc2c2db9, 32'hbc67f92d} /* (3, 21, 18) {real, imag} */,
  {32'hbcf38768, 32'h3c742a9b} /* (3, 21, 17) {real, imag} */,
  {32'h3cb813c4, 32'h00000000} /* (3, 21, 16) {real, imag} */,
  {32'hbcf38768, 32'hbc742a9b} /* (3, 21, 15) {real, imag} */,
  {32'hbc2c2db9, 32'h3c67f92d} /* (3, 21, 14) {real, imag} */,
  {32'hbc99ab76, 32'h3d76a5ca} /* (3, 21, 13) {real, imag} */,
  {32'h3d0ddc2a, 32'h3cc51581} /* (3, 21, 12) {real, imag} */,
  {32'hbdb92c74, 32'h3b071d10} /* (3, 21, 11) {real, imag} */,
  {32'h3d6ae4d5, 32'hbd15a894} /* (3, 21, 10) {real, imag} */,
  {32'h3dcb74d7, 32'h3cb344a4} /* (3, 21, 9) {real, imag} */,
  {32'h3aa72650, 32'hbd939d9a} /* (3, 21, 8) {real, imag} */,
  {32'hbdc17232, 32'hbd8f5583} /* (3, 21, 7) {real, imag} */,
  {32'hbd0e735f, 32'hbd8790fd} /* (3, 21, 6) {real, imag} */,
  {32'h3d95ad7c, 32'h3e003f30} /* (3, 21, 5) {real, imag} */,
  {32'h3d63dc2e, 32'h3dd23f48} /* (3, 21, 4) {real, imag} */,
  {32'hbd81a59e, 32'h3d47b68f} /* (3, 21, 3) {real, imag} */,
  {32'h3e202238, 32'h3d064858} /* (3, 21, 2) {real, imag} */,
  {32'hbedbf8a2, 32'h3e2e74f4} /* (3, 21, 1) {real, imag} */,
  {32'h3e6a76db, 32'h00000000} /* (3, 21, 0) {real, imag} */,
  {32'h3f25aeb0, 32'hbeaa32a8} /* (3, 20, 31) {real, imag} */,
  {32'hbef4ea57, 32'hbc90c25e} /* (3, 20, 30) {real, imag} */,
  {32'hbe720404, 32'h3c5bb653} /* (3, 20, 29) {real, imag} */,
  {32'h3e28ef94, 32'hbd911b54} /* (3, 20, 28) {real, imag} */,
  {32'hbdeceb42, 32'hbe19b204} /* (3, 20, 27) {real, imag} */,
  {32'hbb83b4d4, 32'h3c81253c} /* (3, 20, 26) {real, imag} */,
  {32'hbc1ea0fa, 32'h3df45bcf} /* (3, 20, 25) {real, imag} */,
  {32'hbdb90d18, 32'h3ca36a8f} /* (3, 20, 24) {real, imag} */,
  {32'h3d98c029, 32'hbd8f4550} /* (3, 20, 23) {real, imag} */,
  {32'h3b9f35aa, 32'h3d0c2f6b} /* (3, 20, 22) {real, imag} */,
  {32'hbe21b0e4, 32'hb92c1000} /* (3, 20, 21) {real, imag} */,
  {32'h3c815652, 32'hbdad4d62} /* (3, 20, 20) {real, imag} */,
  {32'h3cf4c2db, 32'hbd1bf312} /* (3, 20, 19) {real, imag} */,
  {32'h3d527eaf, 32'h3c7a876a} /* (3, 20, 18) {real, imag} */,
  {32'h3b5b1db8, 32'hbbd526d6} /* (3, 20, 17) {real, imag} */,
  {32'hbe25bce8, 32'h00000000} /* (3, 20, 16) {real, imag} */,
  {32'h3b5b1db8, 32'h3bd526d6} /* (3, 20, 15) {real, imag} */,
  {32'h3d527eaf, 32'hbc7a876a} /* (3, 20, 14) {real, imag} */,
  {32'h3cf4c2db, 32'h3d1bf312} /* (3, 20, 13) {real, imag} */,
  {32'h3c815652, 32'h3dad4d62} /* (3, 20, 12) {real, imag} */,
  {32'hbe21b0e4, 32'h392c1000} /* (3, 20, 11) {real, imag} */,
  {32'h3b9f35aa, 32'hbd0c2f6b} /* (3, 20, 10) {real, imag} */,
  {32'h3d98c029, 32'h3d8f4550} /* (3, 20, 9) {real, imag} */,
  {32'hbdb90d18, 32'hbca36a8f} /* (3, 20, 8) {real, imag} */,
  {32'hbc1ea0fa, 32'hbdf45bcf} /* (3, 20, 7) {real, imag} */,
  {32'hbb83b4d4, 32'hbc81253c} /* (3, 20, 6) {real, imag} */,
  {32'hbdeceb42, 32'h3e19b204} /* (3, 20, 5) {real, imag} */,
  {32'h3e28ef94, 32'h3d911b54} /* (3, 20, 4) {real, imag} */,
  {32'hbe720404, 32'hbc5bb653} /* (3, 20, 3) {real, imag} */,
  {32'hbef4ea57, 32'h3c90c25e} /* (3, 20, 2) {real, imag} */,
  {32'h3f25aeb0, 32'h3eaa32a8} /* (3, 20, 1) {real, imag} */,
  {32'h3f730034, 32'h00000000} /* (3, 20, 0) {real, imag} */,
  {32'h3f9b8ef3, 32'hbe98abfe} /* (3, 19, 31) {real, imag} */,
  {32'hbf3aaa48, 32'h3cc4d5d8} /* (3, 19, 30) {real, imag} */,
  {32'hbe461148, 32'h3d058e1a} /* (3, 19, 29) {real, imag} */,
  {32'h3e8a32f5, 32'hbc9f8964} /* (3, 19, 28) {real, imag} */,
  {32'hbe1b8d9a, 32'h3bf3d030} /* (3, 19, 27) {real, imag} */,
  {32'hbd6c5ad8, 32'hbd682b13} /* (3, 19, 26) {real, imag} */,
  {32'h3df4c060, 32'h3d0c2202} /* (3, 19, 25) {real, imag} */,
  {32'hbcfaa434, 32'h3d9a3efb} /* (3, 19, 24) {real, imag} */,
  {32'h3dbe1cd8, 32'hbc1c547c} /* (3, 19, 23) {real, imag} */,
  {32'h3cf817cc, 32'h3c5d98e0} /* (3, 19, 22) {real, imag} */,
  {32'hbe5a0f76, 32'h3d86f3fd} /* (3, 19, 21) {real, imag} */,
  {32'h3bc339f8, 32'h3b152ed0} /* (3, 19, 20) {real, imag} */,
  {32'h3d3242b5, 32'hbc46fd80} /* (3, 19, 19) {real, imag} */,
  {32'h3d0da5f6, 32'h3cae7550} /* (3, 19, 18) {real, imag} */,
  {32'hbd436270, 32'hbcc0a79e} /* (3, 19, 17) {real, imag} */,
  {32'hbd9b95a6, 32'h00000000} /* (3, 19, 16) {real, imag} */,
  {32'hbd436270, 32'h3cc0a79e} /* (3, 19, 15) {real, imag} */,
  {32'h3d0da5f6, 32'hbcae7550} /* (3, 19, 14) {real, imag} */,
  {32'h3d3242b5, 32'h3c46fd80} /* (3, 19, 13) {real, imag} */,
  {32'h3bc339f8, 32'hbb152ed0} /* (3, 19, 12) {real, imag} */,
  {32'hbe5a0f76, 32'hbd86f3fd} /* (3, 19, 11) {real, imag} */,
  {32'h3cf817cc, 32'hbc5d98e0} /* (3, 19, 10) {real, imag} */,
  {32'h3dbe1cd8, 32'h3c1c547c} /* (3, 19, 9) {real, imag} */,
  {32'hbcfaa434, 32'hbd9a3efb} /* (3, 19, 8) {real, imag} */,
  {32'h3df4c060, 32'hbd0c2202} /* (3, 19, 7) {real, imag} */,
  {32'hbd6c5ad8, 32'h3d682b13} /* (3, 19, 6) {real, imag} */,
  {32'hbe1b8d9a, 32'hbbf3d030} /* (3, 19, 5) {real, imag} */,
  {32'h3e8a32f5, 32'h3c9f8964} /* (3, 19, 4) {real, imag} */,
  {32'hbe461148, 32'hbd058e1a} /* (3, 19, 3) {real, imag} */,
  {32'hbf3aaa48, 32'hbcc4d5d8} /* (3, 19, 2) {real, imag} */,
  {32'h3f9b8ef3, 32'h3e98abfe} /* (3, 19, 1) {real, imag} */,
  {32'h3f855cd5, 32'h00000000} /* (3, 19, 0) {real, imag} */,
  {32'h3fc4da00, 32'hbea64579} /* (3, 18, 31) {real, imag} */,
  {32'hbf69b140, 32'h3e4edc60} /* (3, 18, 30) {real, imag} */,
  {32'hbe43c27a, 32'hbce91c1f} /* (3, 18, 29) {real, imag} */,
  {32'h3e96c238, 32'hbdc6906c} /* (3, 18, 28) {real, imag} */,
  {32'hbe3b046c, 32'h3e14bbaf} /* (3, 18, 27) {real, imag} */,
  {32'hbdd827be, 32'hbd4662e8} /* (3, 18, 26) {real, imag} */,
  {32'h3cf6cd20, 32'hbc8ccfa8} /* (3, 18, 25) {real, imag} */,
  {32'h3d11e10a, 32'h3d1e859e} /* (3, 18, 24) {real, imag} */,
  {32'hbc2085e2, 32'h3d66fda2} /* (3, 18, 23) {real, imag} */,
  {32'h3d81cd50, 32'hbd6f1cee} /* (3, 18, 22) {real, imag} */,
  {32'hbdfbbd84, 32'h3d6fb701} /* (3, 18, 21) {real, imag} */,
  {32'h3e297311, 32'hbd99a3c7} /* (3, 18, 20) {real, imag} */,
  {32'hbe1186b2, 32'hbd7ad386} /* (3, 18, 19) {real, imag} */,
  {32'hbd0285e7, 32'h3e365e78} /* (3, 18, 18) {real, imag} */,
  {32'h3c937f6b, 32'h3cfa8c93} /* (3, 18, 17) {real, imag} */,
  {32'h3d9dcc5f, 32'h00000000} /* (3, 18, 16) {real, imag} */,
  {32'h3c937f6b, 32'hbcfa8c93} /* (3, 18, 15) {real, imag} */,
  {32'hbd0285e7, 32'hbe365e78} /* (3, 18, 14) {real, imag} */,
  {32'hbe1186b2, 32'h3d7ad386} /* (3, 18, 13) {real, imag} */,
  {32'h3e297311, 32'h3d99a3c7} /* (3, 18, 12) {real, imag} */,
  {32'hbdfbbd84, 32'hbd6fb701} /* (3, 18, 11) {real, imag} */,
  {32'h3d81cd50, 32'h3d6f1cee} /* (3, 18, 10) {real, imag} */,
  {32'hbc2085e2, 32'hbd66fda2} /* (3, 18, 9) {real, imag} */,
  {32'h3d11e10a, 32'hbd1e859e} /* (3, 18, 8) {real, imag} */,
  {32'h3cf6cd20, 32'h3c8ccfa8} /* (3, 18, 7) {real, imag} */,
  {32'hbdd827be, 32'h3d4662e8} /* (3, 18, 6) {real, imag} */,
  {32'hbe3b046c, 32'hbe14bbaf} /* (3, 18, 5) {real, imag} */,
  {32'h3e96c238, 32'h3dc6906c} /* (3, 18, 4) {real, imag} */,
  {32'hbe43c27a, 32'h3ce91c1f} /* (3, 18, 3) {real, imag} */,
  {32'hbf69b140, 32'hbe4edc60} /* (3, 18, 2) {real, imag} */,
  {32'h3fc4da00, 32'h3ea64579} /* (3, 18, 1) {real, imag} */,
  {32'h3f7a603a, 32'h00000000} /* (3, 18, 0) {real, imag} */,
  {32'h3fd0ecee, 32'hbe895918} /* (3, 17, 31) {real, imag} */,
  {32'hbf62778e, 32'h3db5f8ee} /* (3, 17, 30) {real, imag} */,
  {32'hbdd6ba25, 32'h3cf7f168} /* (3, 17, 29) {real, imag} */,
  {32'h3dbf8b10, 32'hbdc74668} /* (3, 17, 28) {real, imag} */,
  {32'hbdebf0f0, 32'h3b7a4200} /* (3, 17, 27) {real, imag} */,
  {32'hbb574770, 32'hbd354137} /* (3, 17, 26) {real, imag} */,
  {32'h3dc7569f, 32'hbe066c8a} /* (3, 17, 25) {real, imag} */,
  {32'hbd34dd06, 32'h3cf5fe40} /* (3, 17, 24) {real, imag} */,
  {32'h3c4c1714, 32'h3d518e04} /* (3, 17, 23) {real, imag} */,
  {32'h3d90b0b5, 32'hbcf48df5} /* (3, 17, 22) {real, imag} */,
  {32'hbcc3f7f4, 32'h3d776145} /* (3, 17, 21) {real, imag} */,
  {32'hbd6c4dee, 32'hbccc4a9f} /* (3, 17, 20) {real, imag} */,
  {32'hbc5476b0, 32'hbd650bbd} /* (3, 17, 19) {real, imag} */,
  {32'hbccfe782, 32'h3d73f2c9} /* (3, 17, 18) {real, imag} */,
  {32'h3d59836d, 32'hbd180e0f} /* (3, 17, 17) {real, imag} */,
  {32'h3cb4dd16, 32'h00000000} /* (3, 17, 16) {real, imag} */,
  {32'h3d59836d, 32'h3d180e0f} /* (3, 17, 15) {real, imag} */,
  {32'hbccfe782, 32'hbd73f2c9} /* (3, 17, 14) {real, imag} */,
  {32'hbc5476b0, 32'h3d650bbd} /* (3, 17, 13) {real, imag} */,
  {32'hbd6c4dee, 32'h3ccc4a9f} /* (3, 17, 12) {real, imag} */,
  {32'hbcc3f7f4, 32'hbd776145} /* (3, 17, 11) {real, imag} */,
  {32'h3d90b0b5, 32'h3cf48df5} /* (3, 17, 10) {real, imag} */,
  {32'h3c4c1714, 32'hbd518e04} /* (3, 17, 9) {real, imag} */,
  {32'hbd34dd06, 32'hbcf5fe40} /* (3, 17, 8) {real, imag} */,
  {32'h3dc7569f, 32'h3e066c8a} /* (3, 17, 7) {real, imag} */,
  {32'hbb574770, 32'h3d354137} /* (3, 17, 6) {real, imag} */,
  {32'hbdebf0f0, 32'hbb7a4200} /* (3, 17, 5) {real, imag} */,
  {32'h3dbf8b10, 32'h3dc74668} /* (3, 17, 4) {real, imag} */,
  {32'hbdd6ba25, 32'hbcf7f168} /* (3, 17, 3) {real, imag} */,
  {32'hbf62778e, 32'hbdb5f8ee} /* (3, 17, 2) {real, imag} */,
  {32'h3fd0ecee, 32'h3e895918} /* (3, 17, 1) {real, imag} */,
  {32'h3f84b9a4, 32'h00000000} /* (3, 17, 0) {real, imag} */,
  {32'h3fea1bb9, 32'hbe59d10e} /* (3, 16, 31) {real, imag} */,
  {32'hbf55d647, 32'h3e1bf9a8} /* (3, 16, 30) {real, imag} */,
  {32'h3dfe41b8, 32'hbc2884de} /* (3, 16, 29) {real, imag} */,
  {32'h3e42840c, 32'hbdab550b} /* (3, 16, 28) {real, imag} */,
  {32'hbe20dd64, 32'h3d952e7d} /* (3, 16, 27) {real, imag} */,
  {32'hbd99ed7c, 32'hbd490adc} /* (3, 16, 26) {real, imag} */,
  {32'h3cf24610, 32'hbd2e9a62} /* (3, 16, 25) {real, imag} */,
  {32'hbdd7f3e6, 32'h3da9507a} /* (3, 16, 24) {real, imag} */,
  {32'h3d6be222, 32'h3cf44ba4} /* (3, 16, 23) {real, imag} */,
  {32'hbd2ed07c, 32'hbc930a55} /* (3, 16, 22) {real, imag} */,
  {32'h3c15383c, 32'h3d8cf89c} /* (3, 16, 21) {real, imag} */,
  {32'hbc877651, 32'h3daf3aba} /* (3, 16, 20) {real, imag} */,
  {32'h3cb37304, 32'hbd3e408c} /* (3, 16, 19) {real, imag} */,
  {32'h3dd2a777, 32'h3da37ac5} /* (3, 16, 18) {real, imag} */,
  {32'hbc77b108, 32'hbcaa5be3} /* (3, 16, 17) {real, imag} */,
  {32'h3cfaec94, 32'h00000000} /* (3, 16, 16) {real, imag} */,
  {32'hbc77b108, 32'h3caa5be3} /* (3, 16, 15) {real, imag} */,
  {32'h3dd2a777, 32'hbda37ac5} /* (3, 16, 14) {real, imag} */,
  {32'h3cb37304, 32'h3d3e408c} /* (3, 16, 13) {real, imag} */,
  {32'hbc877651, 32'hbdaf3aba} /* (3, 16, 12) {real, imag} */,
  {32'h3c15383c, 32'hbd8cf89c} /* (3, 16, 11) {real, imag} */,
  {32'hbd2ed07c, 32'h3c930a55} /* (3, 16, 10) {real, imag} */,
  {32'h3d6be222, 32'hbcf44ba4} /* (3, 16, 9) {real, imag} */,
  {32'hbdd7f3e6, 32'hbda9507a} /* (3, 16, 8) {real, imag} */,
  {32'h3cf24610, 32'h3d2e9a62} /* (3, 16, 7) {real, imag} */,
  {32'hbd99ed7c, 32'h3d490adc} /* (3, 16, 6) {real, imag} */,
  {32'hbe20dd64, 32'hbd952e7d} /* (3, 16, 5) {real, imag} */,
  {32'h3e42840c, 32'h3dab550b} /* (3, 16, 4) {real, imag} */,
  {32'h3dfe41b8, 32'h3c2884de} /* (3, 16, 3) {real, imag} */,
  {32'hbf55d647, 32'hbe1bf9a8} /* (3, 16, 2) {real, imag} */,
  {32'h3fea1bb9, 32'h3e59d10e} /* (3, 16, 1) {real, imag} */,
  {32'h3f7db468, 32'h00000000} /* (3, 16, 0) {real, imag} */,
  {32'h3fd42f2a, 32'hbea494aa} /* (3, 15, 31) {real, imag} */,
  {32'hbf4e0c26, 32'h3e5942d3} /* (3, 15, 30) {real, imag} */,
  {32'h3dad9605, 32'h3c9a2252} /* (3, 15, 29) {real, imag} */,
  {32'h3e58386c, 32'hbdaf05ee} /* (3, 15, 28) {real, imag} */,
  {32'hbe4d9958, 32'h3dbfa458} /* (3, 15, 27) {real, imag} */,
  {32'h3d220c93, 32'hba2d1d80} /* (3, 15, 26) {real, imag} */,
  {32'h3d6af63a, 32'hbd880f37} /* (3, 15, 25) {real, imag} */,
  {32'hbe0f5e62, 32'h3c910880} /* (3, 15, 24) {real, imag} */,
  {32'hbd181902, 32'hbb6dd988} /* (3, 15, 23) {real, imag} */,
  {32'h3cf4bfcc, 32'hbcd8019b} /* (3, 15, 22) {real, imag} */,
  {32'hbd756eea, 32'h3cf24a76} /* (3, 15, 21) {real, imag} */,
  {32'h3d927075, 32'hbccc8e77} /* (3, 15, 20) {real, imag} */,
  {32'h3d8a14da, 32'hbc65e3bc} /* (3, 15, 19) {real, imag} */,
  {32'h3dab91c6, 32'h39f7e900} /* (3, 15, 18) {real, imag} */,
  {32'hbbf318f8, 32'h3d6ac249} /* (3, 15, 17) {real, imag} */,
  {32'hbd958154, 32'h00000000} /* (3, 15, 16) {real, imag} */,
  {32'hbbf318f8, 32'hbd6ac249} /* (3, 15, 15) {real, imag} */,
  {32'h3dab91c6, 32'hb9f7e900} /* (3, 15, 14) {real, imag} */,
  {32'h3d8a14da, 32'h3c65e3bc} /* (3, 15, 13) {real, imag} */,
  {32'h3d927075, 32'h3ccc8e77} /* (3, 15, 12) {real, imag} */,
  {32'hbd756eea, 32'hbcf24a76} /* (3, 15, 11) {real, imag} */,
  {32'h3cf4bfcc, 32'h3cd8019b} /* (3, 15, 10) {real, imag} */,
  {32'hbd181902, 32'h3b6dd988} /* (3, 15, 9) {real, imag} */,
  {32'hbe0f5e62, 32'hbc910880} /* (3, 15, 8) {real, imag} */,
  {32'h3d6af63a, 32'h3d880f37} /* (3, 15, 7) {real, imag} */,
  {32'h3d220c93, 32'h3a2d1d80} /* (3, 15, 6) {real, imag} */,
  {32'hbe4d9958, 32'hbdbfa458} /* (3, 15, 5) {real, imag} */,
  {32'h3e58386c, 32'h3daf05ee} /* (3, 15, 4) {real, imag} */,
  {32'h3dad9605, 32'hbc9a2252} /* (3, 15, 3) {real, imag} */,
  {32'hbf4e0c26, 32'hbe5942d3} /* (3, 15, 2) {real, imag} */,
  {32'h3fd42f2a, 32'h3ea494aa} /* (3, 15, 1) {real, imag} */,
  {32'h3f9c167a, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'h3fd006fc, 32'hbe905243} /* (3, 14, 31) {real, imag} */,
  {32'hbf53e808, 32'h3dee1bfb} /* (3, 14, 30) {real, imag} */,
  {32'h3e41ff80, 32'h3cc53c15} /* (3, 14, 29) {real, imag} */,
  {32'h3e04389d, 32'hbe2fdf5a} /* (3, 14, 28) {real, imag} */,
  {32'hbe4fa836, 32'h3e8152a2} /* (3, 14, 27) {real, imag} */,
  {32'h3dac3332, 32'h3d61967c} /* (3, 14, 26) {real, imag} */,
  {32'h3df367c8, 32'hbdda4bb3} /* (3, 14, 25) {real, imag} */,
  {32'hbde2f24b, 32'h3da0a491} /* (3, 14, 24) {real, imag} */,
  {32'h3cc102b5, 32'hbbe08e80} /* (3, 14, 23) {real, imag} */,
  {32'hbd64065f, 32'h3ca34800} /* (3, 14, 22) {real, imag} */,
  {32'h3d31212c, 32'hbc48081c} /* (3, 14, 21) {real, imag} */,
  {32'h3d77b16c, 32'h3d90994d} /* (3, 14, 20) {real, imag} */,
  {32'h3c0e5c50, 32'hbd3c081a} /* (3, 14, 19) {real, imag} */,
  {32'hbd13faf1, 32'h3daaf9e0} /* (3, 14, 18) {real, imag} */,
  {32'h3d8194d3, 32'hbd22694a} /* (3, 14, 17) {real, imag} */,
  {32'h3c982ffd, 32'h00000000} /* (3, 14, 16) {real, imag} */,
  {32'h3d8194d3, 32'h3d22694a} /* (3, 14, 15) {real, imag} */,
  {32'hbd13faf1, 32'hbdaaf9e0} /* (3, 14, 14) {real, imag} */,
  {32'h3c0e5c50, 32'h3d3c081a} /* (3, 14, 13) {real, imag} */,
  {32'h3d77b16c, 32'hbd90994d} /* (3, 14, 12) {real, imag} */,
  {32'h3d31212c, 32'h3c48081c} /* (3, 14, 11) {real, imag} */,
  {32'hbd64065f, 32'hbca34800} /* (3, 14, 10) {real, imag} */,
  {32'h3cc102b5, 32'h3be08e80} /* (3, 14, 9) {real, imag} */,
  {32'hbde2f24b, 32'hbda0a491} /* (3, 14, 8) {real, imag} */,
  {32'h3df367c8, 32'h3dda4bb3} /* (3, 14, 7) {real, imag} */,
  {32'h3dac3332, 32'hbd61967c} /* (3, 14, 6) {real, imag} */,
  {32'hbe4fa836, 32'hbe8152a2} /* (3, 14, 5) {real, imag} */,
  {32'h3e04389d, 32'h3e2fdf5a} /* (3, 14, 4) {real, imag} */,
  {32'h3e41ff80, 32'hbcc53c15} /* (3, 14, 3) {real, imag} */,
  {32'hbf53e808, 32'hbdee1bfb} /* (3, 14, 2) {real, imag} */,
  {32'h3fd006fc, 32'h3e905243} /* (3, 14, 1) {real, imag} */,
  {32'h3fa171b3, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'h3fd33c3d, 32'hbeb15a3a} /* (3, 13, 31) {real, imag} */,
  {32'hbf2fb5c0, 32'h3d0ad1ac} /* (3, 13, 30) {real, imag} */,
  {32'h3e333b44, 32'h3c21b558} /* (3, 13, 29) {real, imag} */,
  {32'h3e36cd33, 32'hbe1c777e} /* (3, 13, 28) {real, imag} */,
  {32'hbe2cd4e4, 32'h3e2a7028} /* (3, 13, 27) {real, imag} */,
  {32'hbd1d22fc, 32'h3df0f0c6} /* (3, 13, 26) {real, imag} */,
  {32'h3c442830, 32'h3d8cd941} /* (3, 13, 25) {real, imag} */,
  {32'hbddef0fb, 32'h3de9c5fd} /* (3, 13, 24) {real, imag} */,
  {32'h3dc82ac8, 32'h3dcdd59e} /* (3, 13, 23) {real, imag} */,
  {32'hbd158f00, 32'hbd30a39e} /* (3, 13, 22) {real, imag} */,
  {32'hbd106e82, 32'h3d719352} /* (3, 13, 21) {real, imag} */,
  {32'hbdc7a176, 32'hbdd92b12} /* (3, 13, 20) {real, imag} */,
  {32'hbd01362d, 32'h3dfad6cc} /* (3, 13, 19) {real, imag} */,
  {32'h3c569817, 32'h3d02ed96} /* (3, 13, 18) {real, imag} */,
  {32'hbd45b0c0, 32'h3d96afce} /* (3, 13, 17) {real, imag} */,
  {32'hb9a52c80, 32'h00000000} /* (3, 13, 16) {real, imag} */,
  {32'hbd45b0c0, 32'hbd96afce} /* (3, 13, 15) {real, imag} */,
  {32'h3c569817, 32'hbd02ed96} /* (3, 13, 14) {real, imag} */,
  {32'hbd01362d, 32'hbdfad6cc} /* (3, 13, 13) {real, imag} */,
  {32'hbdc7a176, 32'h3dd92b12} /* (3, 13, 12) {real, imag} */,
  {32'hbd106e82, 32'hbd719352} /* (3, 13, 11) {real, imag} */,
  {32'hbd158f00, 32'h3d30a39e} /* (3, 13, 10) {real, imag} */,
  {32'h3dc82ac8, 32'hbdcdd59e} /* (3, 13, 9) {real, imag} */,
  {32'hbddef0fb, 32'hbde9c5fd} /* (3, 13, 8) {real, imag} */,
  {32'h3c442830, 32'hbd8cd941} /* (3, 13, 7) {real, imag} */,
  {32'hbd1d22fc, 32'hbdf0f0c6} /* (3, 13, 6) {real, imag} */,
  {32'hbe2cd4e4, 32'hbe2a7028} /* (3, 13, 5) {real, imag} */,
  {32'h3e36cd33, 32'h3e1c777e} /* (3, 13, 4) {real, imag} */,
  {32'h3e333b44, 32'hbc21b558} /* (3, 13, 3) {real, imag} */,
  {32'hbf2fb5c0, 32'hbd0ad1ac} /* (3, 13, 2) {real, imag} */,
  {32'h3fd33c3d, 32'h3eb15a3a} /* (3, 13, 1) {real, imag} */,
  {32'h3f971ed1, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'h3fb4d41c, 32'hbe8021e4} /* (3, 12, 31) {real, imag} */,
  {32'hbf155e1a, 32'h3cd75b1e} /* (3, 12, 30) {real, imag} */,
  {32'h3e199eb6, 32'hbc8bdcdf} /* (3, 12, 29) {real, imag} */,
  {32'h3e12dea8, 32'hbdabaa9c} /* (3, 12, 28) {real, imag} */,
  {32'hbd90b9ba, 32'h3d7215d2} /* (3, 12, 27) {real, imag} */,
  {32'hbd37f14c, 32'h3e425cae} /* (3, 12, 26) {real, imag} */,
  {32'hba8e03b0, 32'h3e023dd3} /* (3, 12, 25) {real, imag} */,
  {32'hbcac1602, 32'h3d8c3670} /* (3, 12, 24) {real, imag} */,
  {32'h3d65cbbe, 32'h3d7a8ddd} /* (3, 12, 23) {real, imag} */,
  {32'h3d05439f, 32'hbbbaaf52} /* (3, 12, 22) {real, imag} */,
  {32'hbd015ad0, 32'h3e0fd3be} /* (3, 12, 21) {real, imag} */,
  {32'hbc062771, 32'h3e06326a} /* (3, 12, 20) {real, imag} */,
  {32'h3c91c487, 32'hbc8b802a} /* (3, 12, 19) {real, imag} */,
  {32'hbddb0f2a, 32'h3d8edd26} /* (3, 12, 18) {real, imag} */,
  {32'hbcef1a75, 32'h3c3659bb} /* (3, 12, 17) {real, imag} */,
  {32'hbd6feb98, 32'h00000000} /* (3, 12, 16) {real, imag} */,
  {32'hbcef1a75, 32'hbc3659bb} /* (3, 12, 15) {real, imag} */,
  {32'hbddb0f2a, 32'hbd8edd26} /* (3, 12, 14) {real, imag} */,
  {32'h3c91c487, 32'h3c8b802a} /* (3, 12, 13) {real, imag} */,
  {32'hbc062771, 32'hbe06326a} /* (3, 12, 12) {real, imag} */,
  {32'hbd015ad0, 32'hbe0fd3be} /* (3, 12, 11) {real, imag} */,
  {32'h3d05439f, 32'h3bbaaf52} /* (3, 12, 10) {real, imag} */,
  {32'h3d65cbbe, 32'hbd7a8ddd} /* (3, 12, 9) {real, imag} */,
  {32'hbcac1602, 32'hbd8c3670} /* (3, 12, 8) {real, imag} */,
  {32'hba8e03b0, 32'hbe023dd3} /* (3, 12, 7) {real, imag} */,
  {32'hbd37f14c, 32'hbe425cae} /* (3, 12, 6) {real, imag} */,
  {32'hbd90b9ba, 32'hbd7215d2} /* (3, 12, 5) {real, imag} */,
  {32'h3e12dea8, 32'h3dabaa9c} /* (3, 12, 4) {real, imag} */,
  {32'h3e199eb6, 32'h3c8bdcdf} /* (3, 12, 3) {real, imag} */,
  {32'hbf155e1a, 32'hbcd75b1e} /* (3, 12, 2) {real, imag} */,
  {32'h3fb4d41c, 32'h3e8021e4} /* (3, 12, 1) {real, imag} */,
  {32'h3f83458f, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'h3f70b997, 32'hbd20fb30} /* (3, 11, 31) {real, imag} */,
  {32'hbeebb9be, 32'hbd1db798} /* (3, 11, 30) {real, imag} */,
  {32'h3d5f7ead, 32'hbd7f2aa7} /* (3, 11, 29) {real, imag} */,
  {32'h3ded4f3b, 32'hbdd07b2e} /* (3, 11, 28) {real, imag} */,
  {32'hbe50046e, 32'h3dd6b182} /* (3, 11, 27) {real, imag} */,
  {32'hbbc28b98, 32'h3c0967e8} /* (3, 11, 26) {real, imag} */,
  {32'h3b8482b8, 32'hbda15d91} /* (3, 11, 25) {real, imag} */,
  {32'hbc8ae4e3, 32'h3dbe47ac} /* (3, 11, 24) {real, imag} */,
  {32'h3bcfc940, 32'hbddc3447} /* (3, 11, 23) {real, imag} */,
  {32'hbd3316e1, 32'h3d97b37c} /* (3, 11, 22) {real, imag} */,
  {32'h3d4f7d31, 32'h3dc81478} /* (3, 11, 21) {real, imag} */,
  {32'h3cd5d553, 32'h3c39285e} /* (3, 11, 20) {real, imag} */,
  {32'h3ca2e35e, 32'hbd1f1530} /* (3, 11, 19) {real, imag} */,
  {32'h3bc1788e, 32'hbc01e2ed} /* (3, 11, 18) {real, imag} */,
  {32'hbc57a630, 32'h3c81a5f8} /* (3, 11, 17) {real, imag} */,
  {32'h3baea346, 32'h00000000} /* (3, 11, 16) {real, imag} */,
  {32'hbc57a630, 32'hbc81a5f8} /* (3, 11, 15) {real, imag} */,
  {32'h3bc1788e, 32'h3c01e2ed} /* (3, 11, 14) {real, imag} */,
  {32'h3ca2e35e, 32'h3d1f1530} /* (3, 11, 13) {real, imag} */,
  {32'h3cd5d553, 32'hbc39285e} /* (3, 11, 12) {real, imag} */,
  {32'h3d4f7d31, 32'hbdc81478} /* (3, 11, 11) {real, imag} */,
  {32'hbd3316e1, 32'hbd97b37c} /* (3, 11, 10) {real, imag} */,
  {32'h3bcfc940, 32'h3ddc3447} /* (3, 11, 9) {real, imag} */,
  {32'hbc8ae4e3, 32'hbdbe47ac} /* (3, 11, 8) {real, imag} */,
  {32'h3b8482b8, 32'h3da15d91} /* (3, 11, 7) {real, imag} */,
  {32'hbbc28b98, 32'hbc0967e8} /* (3, 11, 6) {real, imag} */,
  {32'hbe50046e, 32'hbdd6b182} /* (3, 11, 5) {real, imag} */,
  {32'h3ded4f3b, 32'h3dd07b2e} /* (3, 11, 4) {real, imag} */,
  {32'h3d5f7ead, 32'h3d7f2aa7} /* (3, 11, 3) {real, imag} */,
  {32'hbeebb9be, 32'h3d1db798} /* (3, 11, 2) {real, imag} */,
  {32'h3f70b997, 32'h3d20fb30} /* (3, 11, 1) {real, imag} */,
  {32'h3f1f28c5, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'hbe2fba58, 32'h3d94f587} /* (3, 10, 31) {real, imag} */,
  {32'h3dc2f5c0, 32'hbdec1e7a} /* (3, 10, 30) {real, imag} */,
  {32'h3d032eee, 32'hbe335521} /* (3, 10, 29) {real, imag} */,
  {32'hbc7e7d54, 32'h3d296a96} /* (3, 10, 28) {real, imag} */,
  {32'hbcfae384, 32'hbd19e607} /* (3, 10, 27) {real, imag} */,
  {32'h3dab4608, 32'h3d0cca80} /* (3, 10, 26) {real, imag} */,
  {32'hbd3ecb82, 32'h3cf58c8e} /* (3, 10, 25) {real, imag} */,
  {32'h3c6f1c56, 32'h3cda35d6} /* (3, 10, 24) {real, imag} */,
  {32'h3cd57a02, 32'h3a25fc00} /* (3, 10, 23) {real, imag} */,
  {32'h3ab93d80, 32'h3ca57f18} /* (3, 10, 22) {real, imag} */,
  {32'hbd91aa80, 32'hbceaf942} /* (3, 10, 21) {real, imag} */,
  {32'hbd76135e, 32'h3bdc31c0} /* (3, 10, 20) {real, imag} */,
  {32'hbd83e88c, 32'h3d254c40} /* (3, 10, 19) {real, imag} */,
  {32'h3dda4813, 32'hbd5eee68} /* (3, 10, 18) {real, imag} */,
  {32'hbdbfc774, 32'hbd5a6675} /* (3, 10, 17) {real, imag} */,
  {32'hbd38b40d, 32'h00000000} /* (3, 10, 16) {real, imag} */,
  {32'hbdbfc774, 32'h3d5a6675} /* (3, 10, 15) {real, imag} */,
  {32'h3dda4813, 32'h3d5eee68} /* (3, 10, 14) {real, imag} */,
  {32'hbd83e88c, 32'hbd254c40} /* (3, 10, 13) {real, imag} */,
  {32'hbd76135e, 32'hbbdc31c0} /* (3, 10, 12) {real, imag} */,
  {32'hbd91aa80, 32'h3ceaf942} /* (3, 10, 11) {real, imag} */,
  {32'h3ab93d80, 32'hbca57f18} /* (3, 10, 10) {real, imag} */,
  {32'h3cd57a02, 32'hba25fc00} /* (3, 10, 9) {real, imag} */,
  {32'h3c6f1c56, 32'hbcda35d6} /* (3, 10, 8) {real, imag} */,
  {32'hbd3ecb82, 32'hbcf58c8e} /* (3, 10, 7) {real, imag} */,
  {32'h3dab4608, 32'hbd0cca80} /* (3, 10, 6) {real, imag} */,
  {32'hbcfae384, 32'h3d19e607} /* (3, 10, 5) {real, imag} */,
  {32'hbc7e7d54, 32'hbd296a96} /* (3, 10, 4) {real, imag} */,
  {32'h3d032eee, 32'h3e335521} /* (3, 10, 3) {real, imag} */,
  {32'h3dc2f5c0, 32'h3dec1e7a} /* (3, 10, 2) {real, imag} */,
  {32'hbe2fba58, 32'hbd94f587} /* (3, 10, 1) {real, imag} */,
  {32'hbdc69c54, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'hbf75d5df, 32'h3dc76e2d} /* (3, 9, 31) {real, imag} */,
  {32'h3ee5e7b2, 32'hbe5d8e1c} /* (3, 9, 30) {real, imag} */,
  {32'h3cf7f520, 32'hbd245e08} /* (3, 9, 29) {real, imag} */,
  {32'hbd58a7e4, 32'h3dc3e883} /* (3, 9, 28) {real, imag} */,
  {32'h3e421ec0, 32'hbe204236} /* (3, 9, 27) {real, imag} */,
  {32'h3d5aefe3, 32'h3dd06ba9} /* (3, 9, 26) {real, imag} */,
  {32'hbdd45b86, 32'h3d214f88} /* (3, 9, 25) {real, imag} */,
  {32'h3e08bc84, 32'hbd2ef991} /* (3, 9, 24) {real, imag} */,
  {32'h3d522a24, 32'h3c9ab55f} /* (3, 9, 23) {real, imag} */,
  {32'hbd4a82c4, 32'hbd0f996e} /* (3, 9, 22) {real, imag} */,
  {32'h3cb86ae1, 32'hbd2f38a9} /* (3, 9, 21) {real, imag} */,
  {32'hbcd0f1ed, 32'hbc68878c} /* (3, 9, 20) {real, imag} */,
  {32'h3d5ea9d6, 32'hbe28a150} /* (3, 9, 19) {real, imag} */,
  {32'h3d7e6312, 32'h3d852a1e} /* (3, 9, 18) {real, imag} */,
  {32'hbd1a74b2, 32'hbd5e79ca} /* (3, 9, 17) {real, imag} */,
  {32'hbc86f04b, 32'h00000000} /* (3, 9, 16) {real, imag} */,
  {32'hbd1a74b2, 32'h3d5e79ca} /* (3, 9, 15) {real, imag} */,
  {32'h3d7e6312, 32'hbd852a1e} /* (3, 9, 14) {real, imag} */,
  {32'h3d5ea9d6, 32'h3e28a150} /* (3, 9, 13) {real, imag} */,
  {32'hbcd0f1ed, 32'h3c68878c} /* (3, 9, 12) {real, imag} */,
  {32'h3cb86ae1, 32'h3d2f38a9} /* (3, 9, 11) {real, imag} */,
  {32'hbd4a82c4, 32'h3d0f996e} /* (3, 9, 10) {real, imag} */,
  {32'h3d522a24, 32'hbc9ab55f} /* (3, 9, 9) {real, imag} */,
  {32'h3e08bc84, 32'h3d2ef991} /* (3, 9, 8) {real, imag} */,
  {32'hbdd45b86, 32'hbd214f88} /* (3, 9, 7) {real, imag} */,
  {32'h3d5aefe3, 32'hbdd06ba9} /* (3, 9, 6) {real, imag} */,
  {32'h3e421ec0, 32'h3e204236} /* (3, 9, 5) {real, imag} */,
  {32'hbd58a7e4, 32'hbdc3e883} /* (3, 9, 4) {real, imag} */,
  {32'h3cf7f520, 32'h3d245e08} /* (3, 9, 3) {real, imag} */,
  {32'h3ee5e7b2, 32'h3e5d8e1c} /* (3, 9, 2) {real, imag} */,
  {32'hbf75d5df, 32'hbdc76e2d} /* (3, 9, 1) {real, imag} */,
  {32'hbed6a2ac, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'hbf995621, 32'h3cca1510} /* (3, 8, 31) {real, imag} */,
  {32'h3f31c39e, 32'hbc10d4c4} /* (3, 8, 30) {real, imag} */,
  {32'h3dcc96c7, 32'hbd206622} /* (3, 8, 29) {real, imag} */,
  {32'hbe0d4696, 32'hbd9f0de0} /* (3, 8, 28) {real, imag} */,
  {32'h3e60835d, 32'hbe1d1722} /* (3, 8, 27) {real, imag} */,
  {32'hbc9e44e5, 32'h3d8d1c3c} /* (3, 8, 26) {real, imag} */,
  {32'hbd9a713a, 32'h3d0cd578} /* (3, 8, 25) {real, imag} */,
  {32'h3d533db4, 32'hbdb5540c} /* (3, 8, 24) {real, imag} */,
  {32'h3d5b1c4c, 32'h3df78c47} /* (3, 8, 23) {real, imag} */,
  {32'hbdc3308c, 32'hbe17ec0a} /* (3, 8, 22) {real, imag} */,
  {32'h3d14e5aa, 32'h3d42c243} /* (3, 8, 21) {real, imag} */,
  {32'hbda82682, 32'hbc94ea9d} /* (3, 8, 20) {real, imag} */,
  {32'h3d0871ca, 32'hbdb912fd} /* (3, 8, 19) {real, imag} */,
  {32'h3d3ec7dd, 32'hbcc18933} /* (3, 8, 18) {real, imag} */,
  {32'h3cb5fe58, 32'h3c8b3c50} /* (3, 8, 17) {real, imag} */,
  {32'hbc672c67, 32'h00000000} /* (3, 8, 16) {real, imag} */,
  {32'h3cb5fe58, 32'hbc8b3c50} /* (3, 8, 15) {real, imag} */,
  {32'h3d3ec7dd, 32'h3cc18933} /* (3, 8, 14) {real, imag} */,
  {32'h3d0871ca, 32'h3db912fd} /* (3, 8, 13) {real, imag} */,
  {32'hbda82682, 32'h3c94ea9d} /* (3, 8, 12) {real, imag} */,
  {32'h3d14e5aa, 32'hbd42c243} /* (3, 8, 11) {real, imag} */,
  {32'hbdc3308c, 32'h3e17ec0a} /* (3, 8, 10) {real, imag} */,
  {32'h3d5b1c4c, 32'hbdf78c47} /* (3, 8, 9) {real, imag} */,
  {32'h3d533db4, 32'h3db5540c} /* (3, 8, 8) {real, imag} */,
  {32'hbd9a713a, 32'hbd0cd578} /* (3, 8, 7) {real, imag} */,
  {32'hbc9e44e5, 32'hbd8d1c3c} /* (3, 8, 6) {real, imag} */,
  {32'h3e60835d, 32'h3e1d1722} /* (3, 8, 5) {real, imag} */,
  {32'hbe0d4696, 32'h3d9f0de0} /* (3, 8, 4) {real, imag} */,
  {32'h3dcc96c7, 32'h3d206622} /* (3, 8, 3) {real, imag} */,
  {32'h3f31c39e, 32'h3c10d4c4} /* (3, 8, 2) {real, imag} */,
  {32'hbf995621, 32'hbcca1510} /* (3, 8, 1) {real, imag} */,
  {32'hbf2f3e6f, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'hbfaeb2e6, 32'h3e7c74f6} /* (3, 7, 31) {real, imag} */,
  {32'h3f410b06, 32'h3d927bc8} /* (3, 7, 30) {real, imag} */,
  {32'h3e2836b1, 32'hbd9dff4f} /* (3, 7, 29) {real, imag} */,
  {32'h3d426298, 32'hbe133b96} /* (3, 7, 28) {real, imag} */,
  {32'h3e5081d4, 32'hbe282ec3} /* (3, 7, 27) {real, imag} */,
  {32'h3c834a6a, 32'h3dc49e7c} /* (3, 7, 26) {real, imag} */,
  {32'hbdd7bfc0, 32'h3ccd160e} /* (3, 7, 25) {real, imag} */,
  {32'h3d1317ac, 32'h3d256ca2} /* (3, 7, 24) {real, imag} */,
  {32'hbd021d21, 32'h3c17b11f} /* (3, 7, 23) {real, imag} */,
  {32'hbdc08a51, 32'h3d8db4b6} /* (3, 7, 22) {real, imag} */,
  {32'hbc92ffd8, 32'hbd8bafb4} /* (3, 7, 21) {real, imag} */,
  {32'h3b8cbbc4, 32'h3e0cfa75} /* (3, 7, 20) {real, imag} */,
  {32'h3d74f530, 32'hbd4228c7} /* (3, 7, 19) {real, imag} */,
  {32'h3bdab9c2, 32'hbd9dfd2a} /* (3, 7, 18) {real, imag} */,
  {32'hbaf2f600, 32'hbdfd5354} /* (3, 7, 17) {real, imag} */,
  {32'h3d89b344, 32'h00000000} /* (3, 7, 16) {real, imag} */,
  {32'hbaf2f600, 32'h3dfd5354} /* (3, 7, 15) {real, imag} */,
  {32'h3bdab9c2, 32'h3d9dfd2a} /* (3, 7, 14) {real, imag} */,
  {32'h3d74f530, 32'h3d4228c7} /* (3, 7, 13) {real, imag} */,
  {32'h3b8cbbc4, 32'hbe0cfa75} /* (3, 7, 12) {real, imag} */,
  {32'hbc92ffd8, 32'h3d8bafb4} /* (3, 7, 11) {real, imag} */,
  {32'hbdc08a51, 32'hbd8db4b6} /* (3, 7, 10) {real, imag} */,
  {32'hbd021d21, 32'hbc17b11f} /* (3, 7, 9) {real, imag} */,
  {32'h3d1317ac, 32'hbd256ca2} /* (3, 7, 8) {real, imag} */,
  {32'hbdd7bfc0, 32'hbccd160e} /* (3, 7, 7) {real, imag} */,
  {32'h3c834a6a, 32'hbdc49e7c} /* (3, 7, 6) {real, imag} */,
  {32'h3e5081d4, 32'h3e282ec3} /* (3, 7, 5) {real, imag} */,
  {32'h3d426298, 32'h3e133b96} /* (3, 7, 4) {real, imag} */,
  {32'h3e2836b1, 32'h3d9dff4f} /* (3, 7, 3) {real, imag} */,
  {32'h3f410b06, 32'hbd927bc8} /* (3, 7, 2) {real, imag} */,
  {32'hbfaeb2e6, 32'hbe7c74f6} /* (3, 7, 1) {real, imag} */,
  {32'hbf3a6d5d, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'hbfa15e22, 32'h3f0520fa} /* (3, 6, 31) {real, imag} */,
  {32'h3f05a61e, 32'hbd83072e} /* (3, 6, 30) {real, imag} */,
  {32'h3e36d7d4, 32'hbd4769ea} /* (3, 6, 29) {real, imag} */,
  {32'hbd110544, 32'hbe226951} /* (3, 6, 28) {real, imag} */,
  {32'h3d937296, 32'hbd5b8e63} /* (3, 6, 27) {real, imag} */,
  {32'h3b008430, 32'hbd9ef5e4} /* (3, 6, 26) {real, imag} */,
  {32'hbc1d9e38, 32'hbd7e31ff} /* (3, 6, 25) {real, imag} */,
  {32'h3ddb9e08, 32'hbdd3e76a} /* (3, 6, 24) {real, imag} */,
  {32'h3de2f856, 32'h3d26aaf4} /* (3, 6, 23) {real, imag} */,
  {32'hbd413639, 32'h3d69ec25} /* (3, 6, 22) {real, imag} */,
  {32'h3ce1ffbe, 32'hbdb87a0c} /* (3, 6, 21) {real, imag} */,
  {32'h3aa4a0c0, 32'h3cb8fead} /* (3, 6, 20) {real, imag} */,
  {32'hbd7dc770, 32'hbcf35578} /* (3, 6, 19) {real, imag} */,
  {32'hbbabc25c, 32'hbb7e72f8} /* (3, 6, 18) {real, imag} */,
  {32'h3c0499dc, 32'h3d80a599} /* (3, 6, 17) {real, imag} */,
  {32'hbd6d5ffc, 32'h00000000} /* (3, 6, 16) {real, imag} */,
  {32'h3c0499dc, 32'hbd80a599} /* (3, 6, 15) {real, imag} */,
  {32'hbbabc25c, 32'h3b7e72f8} /* (3, 6, 14) {real, imag} */,
  {32'hbd7dc770, 32'h3cf35578} /* (3, 6, 13) {real, imag} */,
  {32'h3aa4a0c0, 32'hbcb8fead} /* (3, 6, 12) {real, imag} */,
  {32'h3ce1ffbe, 32'h3db87a0c} /* (3, 6, 11) {real, imag} */,
  {32'hbd413639, 32'hbd69ec25} /* (3, 6, 10) {real, imag} */,
  {32'h3de2f856, 32'hbd26aaf4} /* (3, 6, 9) {real, imag} */,
  {32'h3ddb9e08, 32'h3dd3e76a} /* (3, 6, 8) {real, imag} */,
  {32'hbc1d9e38, 32'h3d7e31ff} /* (3, 6, 7) {real, imag} */,
  {32'h3b008430, 32'h3d9ef5e4} /* (3, 6, 6) {real, imag} */,
  {32'h3d937296, 32'h3d5b8e63} /* (3, 6, 5) {real, imag} */,
  {32'hbd110544, 32'h3e226951} /* (3, 6, 4) {real, imag} */,
  {32'h3e36d7d4, 32'h3d4769ea} /* (3, 6, 3) {real, imag} */,
  {32'h3f05a61e, 32'h3d83072e} /* (3, 6, 2) {real, imag} */,
  {32'hbfa15e22, 32'hbf0520fa} /* (3, 6, 1) {real, imag} */,
  {32'hbf2a6f7a, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hbf7734e0, 32'h3f8125c0} /* (3, 5, 31) {real, imag} */,
  {32'h3e1f3532, 32'hbe4fba76} /* (3, 5, 30) {real, imag} */,
  {32'h3e96c1cb, 32'hbcc28af8} /* (3, 5, 29) {real, imag} */,
  {32'hbdb4db3b, 32'hbe1e978b} /* (3, 5, 28) {real, imag} */,
  {32'h3d800f75, 32'h3c3b97b8} /* (3, 5, 27) {real, imag} */,
  {32'h3d9f156f, 32'h3ca0b5b8} /* (3, 5, 26) {real, imag} */,
  {32'h3d59213a, 32'hbd1549ea} /* (3, 5, 25) {real, imag} */,
  {32'hbd9ec2d6, 32'hbd84983c} /* (3, 5, 24) {real, imag} */,
  {32'h3d2c074e, 32'h3cc9d869} /* (3, 5, 23) {real, imag} */,
  {32'h3d808f5a, 32'h388a0200} /* (3, 5, 22) {real, imag} */,
  {32'hbda3fe6c, 32'h3c9b48a7} /* (3, 5, 21) {real, imag} */,
  {32'hbbf1ab70, 32'hbd6dff78} /* (3, 5, 20) {real, imag} */,
  {32'h3cc589ba, 32'h3cc84fa2} /* (3, 5, 19) {real, imag} */,
  {32'h3c14be8a, 32'h3d9ca830} /* (3, 5, 18) {real, imag} */,
  {32'hbd3a89e4, 32'hbd81ed82} /* (3, 5, 17) {real, imag} */,
  {32'hbc22d85a, 32'h00000000} /* (3, 5, 16) {real, imag} */,
  {32'hbd3a89e4, 32'h3d81ed82} /* (3, 5, 15) {real, imag} */,
  {32'h3c14be8a, 32'hbd9ca830} /* (3, 5, 14) {real, imag} */,
  {32'h3cc589ba, 32'hbcc84fa2} /* (3, 5, 13) {real, imag} */,
  {32'hbbf1ab70, 32'h3d6dff78} /* (3, 5, 12) {real, imag} */,
  {32'hbda3fe6c, 32'hbc9b48a7} /* (3, 5, 11) {real, imag} */,
  {32'h3d808f5a, 32'hb88a0200} /* (3, 5, 10) {real, imag} */,
  {32'h3d2c074e, 32'hbcc9d869} /* (3, 5, 9) {real, imag} */,
  {32'hbd9ec2d6, 32'h3d84983c} /* (3, 5, 8) {real, imag} */,
  {32'h3d59213a, 32'h3d1549ea} /* (3, 5, 7) {real, imag} */,
  {32'h3d9f156f, 32'hbca0b5b8} /* (3, 5, 6) {real, imag} */,
  {32'h3d800f75, 32'hbc3b97b8} /* (3, 5, 5) {real, imag} */,
  {32'hbdb4db3b, 32'h3e1e978b} /* (3, 5, 4) {real, imag} */,
  {32'h3e96c1cb, 32'h3cc28af8} /* (3, 5, 3) {real, imag} */,
  {32'h3e1f3532, 32'h3e4fba76} /* (3, 5, 2) {real, imag} */,
  {32'hbf7734e0, 32'hbf8125c0} /* (3, 5, 1) {real, imag} */,
  {32'hbf05f6b8, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hbf523ef2, 32'h3fbaa9e8} /* (3, 4, 31) {real, imag} */,
  {32'hbe22463e, 32'hbe7e736c} /* (3, 4, 30) {real, imag} */,
  {32'h3e6255ad, 32'h3da4e42c} /* (3, 4, 29) {real, imag} */,
  {32'h3d80c424, 32'hbe6c638a} /* (3, 4, 28) {real, imag} */,
  {32'h3e17c1f3, 32'h3d6e53d2} /* (3, 4, 27) {real, imag} */,
  {32'h3d718f9c, 32'hbccb57c6} /* (3, 4, 26) {real, imag} */,
  {32'hbd276aa4, 32'h3cbd74e8} /* (3, 4, 25) {real, imag} */,
  {32'h3c50aa34, 32'h3d66762c} /* (3, 4, 24) {real, imag} */,
  {32'h3d47bd53, 32'hbd4ccbb5} /* (3, 4, 23) {real, imag} */,
  {32'h3bf1cf50, 32'hbd7cea61} /* (3, 4, 22) {real, imag} */,
  {32'h3cac0dd4, 32'h3d907a73} /* (3, 4, 21) {real, imag} */,
  {32'h3d23f8fb, 32'hbd4236fc} /* (3, 4, 20) {real, imag} */,
  {32'h3cb4b4e7, 32'h3d4905f0} /* (3, 4, 19) {real, imag} */,
  {32'hbc4e43f4, 32'hbca85a62} /* (3, 4, 18) {real, imag} */,
  {32'h3c4617e0, 32'hbcec38a4} /* (3, 4, 17) {real, imag} */,
  {32'h3d965d82, 32'h00000000} /* (3, 4, 16) {real, imag} */,
  {32'h3c4617e0, 32'h3cec38a4} /* (3, 4, 15) {real, imag} */,
  {32'hbc4e43f4, 32'h3ca85a62} /* (3, 4, 14) {real, imag} */,
  {32'h3cb4b4e7, 32'hbd4905f0} /* (3, 4, 13) {real, imag} */,
  {32'h3d23f8fb, 32'h3d4236fc} /* (3, 4, 12) {real, imag} */,
  {32'h3cac0dd4, 32'hbd907a73} /* (3, 4, 11) {real, imag} */,
  {32'h3bf1cf50, 32'h3d7cea61} /* (3, 4, 10) {real, imag} */,
  {32'h3d47bd53, 32'h3d4ccbb5} /* (3, 4, 9) {real, imag} */,
  {32'h3c50aa34, 32'hbd66762c} /* (3, 4, 8) {real, imag} */,
  {32'hbd276aa4, 32'hbcbd74e8} /* (3, 4, 7) {real, imag} */,
  {32'h3d718f9c, 32'h3ccb57c6} /* (3, 4, 6) {real, imag} */,
  {32'h3e17c1f3, 32'hbd6e53d2} /* (3, 4, 5) {real, imag} */,
  {32'h3d80c424, 32'h3e6c638a} /* (3, 4, 4) {real, imag} */,
  {32'h3e6255ad, 32'hbda4e42c} /* (3, 4, 3) {real, imag} */,
  {32'hbe22463e, 32'h3e7e736c} /* (3, 4, 2) {real, imag} */,
  {32'hbf523ef2, 32'hbfbaa9e8} /* (3, 4, 1) {real, imag} */,
  {32'hbeb805ed, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hbf36cc18, 32'h3fc10ebc} /* (3, 3, 31) {real, imag} */,
  {32'hbeae1108, 32'hbeeda99b} /* (3, 3, 30) {real, imag} */,
  {32'h3e6b30aa, 32'h3d9ed403} /* (3, 3, 29) {real, imag} */,
  {32'h3d1af264, 32'hbe5cb320} /* (3, 3, 28) {real, imag} */,
  {32'h3e5cd293, 32'h3d21f893} /* (3, 3, 27) {real, imag} */,
  {32'h3da3cd7d, 32'hbc5e6610} /* (3, 3, 26) {real, imag} */,
  {32'h3d8d7a84, 32'hbce70430} /* (3, 3, 25) {real, imag} */,
  {32'hbcde8c02, 32'hbd70b10c} /* (3, 3, 24) {real, imag} */,
  {32'h3c070e1c, 32'hbd8ddd42} /* (3, 3, 23) {real, imag} */,
  {32'hbb9bef9c, 32'hbd96b52d} /* (3, 3, 22) {real, imag} */,
  {32'h39709b00, 32'hbd27c3bc} /* (3, 3, 21) {real, imag} */,
  {32'hbd391efc, 32'hbd21955c} /* (3, 3, 20) {real, imag} */,
  {32'h3d172b29, 32'h3c6c6c10} /* (3, 3, 19) {real, imag} */,
  {32'hbd85cbc8, 32'h3c9f947c} /* (3, 3, 18) {real, imag} */,
  {32'h3dc20db1, 32'hbd980ee2} /* (3, 3, 17) {real, imag} */,
  {32'h3d410bf4, 32'h00000000} /* (3, 3, 16) {real, imag} */,
  {32'h3dc20db1, 32'h3d980ee2} /* (3, 3, 15) {real, imag} */,
  {32'hbd85cbc8, 32'hbc9f947c} /* (3, 3, 14) {real, imag} */,
  {32'h3d172b29, 32'hbc6c6c10} /* (3, 3, 13) {real, imag} */,
  {32'hbd391efc, 32'h3d21955c} /* (3, 3, 12) {real, imag} */,
  {32'h39709b00, 32'h3d27c3bc} /* (3, 3, 11) {real, imag} */,
  {32'hbb9bef9c, 32'h3d96b52d} /* (3, 3, 10) {real, imag} */,
  {32'h3c070e1c, 32'h3d8ddd42} /* (3, 3, 9) {real, imag} */,
  {32'hbcde8c02, 32'h3d70b10c} /* (3, 3, 8) {real, imag} */,
  {32'h3d8d7a84, 32'h3ce70430} /* (3, 3, 7) {real, imag} */,
  {32'h3da3cd7d, 32'h3c5e6610} /* (3, 3, 6) {real, imag} */,
  {32'h3e5cd293, 32'hbd21f893} /* (3, 3, 5) {real, imag} */,
  {32'h3d1af264, 32'h3e5cb320} /* (3, 3, 4) {real, imag} */,
  {32'h3e6b30aa, 32'hbd9ed403} /* (3, 3, 3) {real, imag} */,
  {32'hbeae1108, 32'h3eeda99b} /* (3, 3, 2) {real, imag} */,
  {32'hbf36cc18, 32'hbfc10ebc} /* (3, 3, 1) {real, imag} */,
  {32'hbef6eb4c, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hbf16e6cf, 32'h3fb2dbca} /* (3, 2, 31) {real, imag} */,
  {32'hbeb87d18, 32'hbf086084} /* (3, 2, 30) {real, imag} */,
  {32'h3e24d781, 32'h3dec0f21} /* (3, 2, 29) {real, imag} */,
  {32'h3e2894c0, 32'hbe628f22} /* (3, 2, 28) {real, imag} */,
  {32'h3da9adb9, 32'h3d92e8c4} /* (3, 2, 27) {real, imag} */,
  {32'h3dcb4088, 32'h3c90210e} /* (3, 2, 26) {real, imag} */,
  {32'h3d976e7e, 32'h3d9dae5a} /* (3, 2, 25) {real, imag} */,
  {32'hbde8b24f, 32'hbd946677} /* (3, 2, 24) {real, imag} */,
  {32'h3d008ea2, 32'hbd9caff0} /* (3, 2, 23) {real, imag} */,
  {32'h3cfa6feb, 32'hbd490322} /* (3, 2, 22) {real, imag} */,
  {32'h3db5e5a5, 32'h3d1b70b1} /* (3, 2, 21) {real, imag} */,
  {32'h3b5b23e8, 32'h3d58a1ae} /* (3, 2, 20) {real, imag} */,
  {32'hbdb8c8f9, 32'hbcee55af} /* (3, 2, 19) {real, imag} */,
  {32'h3b740774, 32'h3d7b6ac5} /* (3, 2, 18) {real, imag} */,
  {32'hbc8b2626, 32'h3cd1ab0c} /* (3, 2, 17) {real, imag} */,
  {32'hb97dd180, 32'h00000000} /* (3, 2, 16) {real, imag} */,
  {32'hbc8b2626, 32'hbcd1ab0c} /* (3, 2, 15) {real, imag} */,
  {32'h3b740774, 32'hbd7b6ac5} /* (3, 2, 14) {real, imag} */,
  {32'hbdb8c8f9, 32'h3cee55af} /* (3, 2, 13) {real, imag} */,
  {32'h3b5b23e8, 32'hbd58a1ae} /* (3, 2, 12) {real, imag} */,
  {32'h3db5e5a5, 32'hbd1b70b1} /* (3, 2, 11) {real, imag} */,
  {32'h3cfa6feb, 32'h3d490322} /* (3, 2, 10) {real, imag} */,
  {32'h3d008ea2, 32'h3d9caff0} /* (3, 2, 9) {real, imag} */,
  {32'hbde8b24f, 32'h3d946677} /* (3, 2, 8) {real, imag} */,
  {32'h3d976e7e, 32'hbd9dae5a} /* (3, 2, 7) {real, imag} */,
  {32'h3dcb4088, 32'hbc90210e} /* (3, 2, 6) {real, imag} */,
  {32'h3da9adb9, 32'hbd92e8c4} /* (3, 2, 5) {real, imag} */,
  {32'h3e2894c0, 32'h3e628f22} /* (3, 2, 4) {real, imag} */,
  {32'h3e24d781, 32'hbdec0f21} /* (3, 2, 3) {real, imag} */,
  {32'hbeb87d18, 32'h3f086084} /* (3, 2, 2) {real, imag} */,
  {32'hbf16e6cf, 32'hbfb2dbca} /* (3, 2, 1) {real, imag} */,
  {32'hbe7883b6, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hbf1281ab, 32'h3fa143f0} /* (3, 1, 31) {real, imag} */,
  {32'hbeb2aa4d, 32'hbefd2d6b} /* (3, 1, 30) {real, imag} */,
  {32'h3d9dfe6a, 32'hbd05c217} /* (3, 1, 29) {real, imag} */,
  {32'h3dec2c6b, 32'hbe8620c7} /* (3, 1, 28) {real, imag} */,
  {32'h3e019672, 32'hbd9fca6f} /* (3, 1, 27) {real, imag} */,
  {32'h3ccae78c, 32'h3da5c8b8} /* (3, 1, 26) {real, imag} */,
  {32'h3cac97fc, 32'h3d89026a} /* (3, 1, 25) {real, imag} */,
  {32'hbd9d4c87, 32'hbe118d27} /* (3, 1, 24) {real, imag} */,
  {32'h3d00fe80, 32'hbdd32d16} /* (3, 1, 23) {real, imag} */,
  {32'h3d9e5cff, 32'hbcd4dd10} /* (3, 1, 22) {real, imag} */,
  {32'h3c6275d2, 32'hbcca126e} /* (3, 1, 21) {real, imag} */,
  {32'hbd4ca7c8, 32'hbd36d2aa} /* (3, 1, 20) {real, imag} */,
  {32'h3d3e5143, 32'h3c389732} /* (3, 1, 19) {real, imag} */,
  {32'hbccf5cf6, 32'hbc7e4bb8} /* (3, 1, 18) {real, imag} */,
  {32'h3d276aeb, 32'h3bbba264} /* (3, 1, 17) {real, imag} */,
  {32'h3d5ff871, 32'h00000000} /* (3, 1, 16) {real, imag} */,
  {32'h3d276aeb, 32'hbbbba264} /* (3, 1, 15) {real, imag} */,
  {32'hbccf5cf6, 32'h3c7e4bb8} /* (3, 1, 14) {real, imag} */,
  {32'h3d3e5143, 32'hbc389732} /* (3, 1, 13) {real, imag} */,
  {32'hbd4ca7c8, 32'h3d36d2aa} /* (3, 1, 12) {real, imag} */,
  {32'h3c6275d2, 32'h3cca126e} /* (3, 1, 11) {real, imag} */,
  {32'h3d9e5cff, 32'h3cd4dd10} /* (3, 1, 10) {real, imag} */,
  {32'h3d00fe80, 32'h3dd32d16} /* (3, 1, 9) {real, imag} */,
  {32'hbd9d4c87, 32'h3e118d27} /* (3, 1, 8) {real, imag} */,
  {32'h3cac97fc, 32'hbd89026a} /* (3, 1, 7) {real, imag} */,
  {32'h3ccae78c, 32'hbda5c8b8} /* (3, 1, 6) {real, imag} */,
  {32'h3e019672, 32'h3d9fca6f} /* (3, 1, 5) {real, imag} */,
  {32'h3dec2c6b, 32'h3e8620c7} /* (3, 1, 4) {real, imag} */,
  {32'h3d9dfe6a, 32'h3d05c217} /* (3, 1, 3) {real, imag} */,
  {32'hbeb2aa4d, 32'h3efd2d6b} /* (3, 1, 2) {real, imag} */,
  {32'hbf1281ab, 32'hbfa143f0} /* (3, 1, 1) {real, imag} */,
  {32'h3c089ec4, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'hbf124592, 32'h3f561210} /* (3, 0, 31) {real, imag} */,
  {32'hbe047fcc, 32'hbebd8ba0} /* (3, 0, 30) {real, imag} */,
  {32'h3d866d08, 32'hbd05acd8} /* (3, 0, 29) {real, imag} */,
  {32'h3d72ce60, 32'hbe52e882} /* (3, 0, 28) {real, imag} */,
  {32'h3e2c58cc, 32'h3d503e36} /* (3, 0, 27) {real, imag} */,
  {32'h3d20aa6e, 32'h3cf47164} /* (3, 0, 26) {real, imag} */,
  {32'h3d4bb656, 32'h3ac5f450} /* (3, 0, 25) {real, imag} */,
  {32'hbc85ba4a, 32'hba9b1bc0} /* (3, 0, 24) {real, imag} */,
  {32'hbd9f20c7, 32'hbcad5c84} /* (3, 0, 23) {real, imag} */,
  {32'hbac81440, 32'hbc0232f2} /* (3, 0, 22) {real, imag} */,
  {32'hbcaba97e, 32'h3cc3ecf9} /* (3, 0, 21) {real, imag} */,
  {32'hbcd5cfb5, 32'h3d004ff0} /* (3, 0, 20) {real, imag} */,
  {32'hbcb1ac5c, 32'h3b51a3c8} /* (3, 0, 19) {real, imag} */,
  {32'h3b7b15a0, 32'hbd9bfc57} /* (3, 0, 18) {real, imag} */,
  {32'h3d4b082e, 32'hbca168cb} /* (3, 0, 17) {real, imag} */,
  {32'hbc188870, 32'h00000000} /* (3, 0, 16) {real, imag} */,
  {32'h3d4b082e, 32'h3ca168cb} /* (3, 0, 15) {real, imag} */,
  {32'h3b7b15a0, 32'h3d9bfc57} /* (3, 0, 14) {real, imag} */,
  {32'hbcb1ac5c, 32'hbb51a3c8} /* (3, 0, 13) {real, imag} */,
  {32'hbcd5cfb5, 32'hbd004ff0} /* (3, 0, 12) {real, imag} */,
  {32'hbcaba97e, 32'hbcc3ecf9} /* (3, 0, 11) {real, imag} */,
  {32'hbac81440, 32'h3c0232f2} /* (3, 0, 10) {real, imag} */,
  {32'hbd9f20c7, 32'h3cad5c84} /* (3, 0, 9) {real, imag} */,
  {32'hbc85ba4a, 32'h3a9b1bc0} /* (3, 0, 8) {real, imag} */,
  {32'h3d4bb656, 32'hbac5f450} /* (3, 0, 7) {real, imag} */,
  {32'h3d20aa6e, 32'hbcf47164} /* (3, 0, 6) {real, imag} */,
  {32'h3e2c58cc, 32'hbd503e36} /* (3, 0, 5) {real, imag} */,
  {32'h3d72ce60, 32'h3e52e882} /* (3, 0, 4) {real, imag} */,
  {32'h3d866d08, 32'h3d05acd8} /* (3, 0, 3) {real, imag} */,
  {32'hbe047fcc, 32'h3ebd8ba0} /* (3, 0, 2) {real, imag} */,
  {32'hbf124592, 32'hbf561210} /* (3, 0, 1) {real, imag} */,
  {32'h3e4dfa9a, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hbf8b5903, 32'h3ec995f0} /* (2, 31, 31) {real, imag} */,
  {32'h3ee34841, 32'hbe9d9d6e} /* (2, 31, 30) {real, imag} */,
  {32'h3d728d0d, 32'h3d39d3b0} /* (2, 31, 29) {real, imag} */,
  {32'hbd8538c4, 32'hbdd1403e} /* (2, 31, 28) {real, imag} */,
  {32'h3dc98b1c, 32'hbd9f64b4} /* (2, 31, 27) {real, imag} */,
  {32'hbd10e51c, 32'hbded4b70} /* (2, 31, 26) {real, imag} */,
  {32'h3ce9744a, 32'h3ac3ace0} /* (2, 31, 25) {real, imag} */,
  {32'h3daa4a55, 32'hbd743a42} /* (2, 31, 24) {real, imag} */,
  {32'h3d4f9148, 32'h3cfef4de} /* (2, 31, 23) {real, imag} */,
  {32'h3d550dfa, 32'h3d0bcfa1} /* (2, 31, 22) {real, imag} */,
  {32'hbc7bd9d4, 32'hbde783e9} /* (2, 31, 21) {real, imag} */,
  {32'h3c0b74a8, 32'hbbd7cda0} /* (2, 31, 20) {real, imag} */,
  {32'h3d552d4f, 32'h3d031178} /* (2, 31, 19) {real, imag} */,
  {32'hbce895b5, 32'hbd067566} /* (2, 31, 18) {real, imag} */,
  {32'h3d3426be, 32'h3c4850c8} /* (2, 31, 17) {real, imag} */,
  {32'h3d64088f, 32'h00000000} /* (2, 31, 16) {real, imag} */,
  {32'h3d3426be, 32'hbc4850c8} /* (2, 31, 15) {real, imag} */,
  {32'hbce895b5, 32'h3d067566} /* (2, 31, 14) {real, imag} */,
  {32'h3d552d4f, 32'hbd031178} /* (2, 31, 13) {real, imag} */,
  {32'h3c0b74a8, 32'h3bd7cda0} /* (2, 31, 12) {real, imag} */,
  {32'hbc7bd9d4, 32'h3de783e9} /* (2, 31, 11) {real, imag} */,
  {32'h3d550dfa, 32'hbd0bcfa1} /* (2, 31, 10) {real, imag} */,
  {32'h3d4f9148, 32'hbcfef4de} /* (2, 31, 9) {real, imag} */,
  {32'h3daa4a55, 32'h3d743a42} /* (2, 31, 8) {real, imag} */,
  {32'h3ce9744a, 32'hbac3ace0} /* (2, 31, 7) {real, imag} */,
  {32'hbd10e51c, 32'h3ded4b70} /* (2, 31, 6) {real, imag} */,
  {32'h3dc98b1c, 32'h3d9f64b4} /* (2, 31, 5) {real, imag} */,
  {32'hbd8538c4, 32'h3dd1403e} /* (2, 31, 4) {real, imag} */,
  {32'h3d728d0d, 32'hbd39d3b0} /* (2, 31, 3) {real, imag} */,
  {32'h3ee34841, 32'h3e9d9d6e} /* (2, 31, 2) {real, imag} */,
  {32'hbf8b5903, 32'hbec995f0} /* (2, 31, 1) {real, imag} */,
  {32'hbed50de2, 32'h00000000} /* (2, 31, 0) {real, imag} */,
  {32'hbfba18fc, 32'h3e6fc7d8} /* (2, 30, 31) {real, imag} */,
  {32'h3f408630, 32'hbe54ef78} /* (2, 30, 30) {real, imag} */,
  {32'h3dc09fd8, 32'hbcd81e3e} /* (2, 30, 29) {real, imag} */,
  {32'hbd8e0f71, 32'hbd4b3d9c} /* (2, 30, 28) {real, imag} */,
  {32'h3e6dcb20, 32'hbdbe23c7} /* (2, 30, 27) {real, imag} */,
  {32'hbd23b794, 32'hbdb72c3c} /* (2, 30, 26) {real, imag} */,
  {32'hbb6aaef8, 32'h3d6fb155} /* (2, 30, 25) {real, imag} */,
  {32'h3e1a9a38, 32'hbdb02cd4} /* (2, 30, 24) {real, imag} */,
  {32'hbc978379, 32'h3c5624d3} /* (2, 30, 23) {real, imag} */,
  {32'h3d817ada, 32'h3dd3133c} /* (2, 30, 22) {real, imag} */,
  {32'h3e22901a, 32'hbd4e5121} /* (2, 30, 21) {real, imag} */,
  {32'h3db67872, 32'h3d8a0b86} /* (2, 30, 20) {real, imag} */,
  {32'hbab4f6e0, 32'h3c289e56} /* (2, 30, 19) {real, imag} */,
  {32'hbdb51a30, 32'h3d62a1ae} /* (2, 30, 18) {real, imag} */,
  {32'hbd8a5c14, 32'h3baff3d4} /* (2, 30, 17) {real, imag} */,
  {32'hbe0ec0fc, 32'h00000000} /* (2, 30, 16) {real, imag} */,
  {32'hbd8a5c14, 32'hbbaff3d4} /* (2, 30, 15) {real, imag} */,
  {32'hbdb51a30, 32'hbd62a1ae} /* (2, 30, 14) {real, imag} */,
  {32'hbab4f6e0, 32'hbc289e56} /* (2, 30, 13) {real, imag} */,
  {32'h3db67872, 32'hbd8a0b86} /* (2, 30, 12) {real, imag} */,
  {32'h3e22901a, 32'h3d4e5121} /* (2, 30, 11) {real, imag} */,
  {32'h3d817ada, 32'hbdd3133c} /* (2, 30, 10) {real, imag} */,
  {32'hbc978379, 32'hbc5624d3} /* (2, 30, 9) {real, imag} */,
  {32'h3e1a9a38, 32'h3db02cd4} /* (2, 30, 8) {real, imag} */,
  {32'hbb6aaef8, 32'hbd6fb155} /* (2, 30, 7) {real, imag} */,
  {32'hbd23b794, 32'h3db72c3c} /* (2, 30, 6) {real, imag} */,
  {32'h3e6dcb20, 32'h3dbe23c7} /* (2, 30, 5) {real, imag} */,
  {32'hbd8e0f71, 32'h3d4b3d9c} /* (2, 30, 4) {real, imag} */,
  {32'h3dc09fd8, 32'h3cd81e3e} /* (2, 30, 3) {real, imag} */,
  {32'h3f408630, 32'h3e54ef78} /* (2, 30, 2) {real, imag} */,
  {32'hbfba18fc, 32'hbe6fc7d8} /* (2, 30, 1) {real, imag} */,
  {32'hbf00a990, 32'h00000000} /* (2, 30, 0) {real, imag} */,
  {32'hbfd64dc6, 32'h3e7b2d58} /* (2, 29, 31) {real, imag} */,
  {32'h3f75c000, 32'hbbf21ec0} /* (2, 29, 30) {real, imag} */,
  {32'h3df5f60e, 32'hbe718a87} /* (2, 29, 29) {real, imag} */,
  {32'hbdd1846a, 32'h3cc5d9f4} /* (2, 29, 28) {real, imag} */,
  {32'h3e93a75b, 32'hbdd71922} /* (2, 29, 27) {real, imag} */,
  {32'hbc6c67e0, 32'h3c50abe4} /* (2, 29, 26) {real, imag} */,
  {32'h3d14e1d8, 32'h3cd2013a} /* (2, 29, 25) {real, imag} */,
  {32'h3e07c660, 32'hbda8209e} /* (2, 29, 24) {real, imag} */,
  {32'hbce9359c, 32'h3db9f0eb} /* (2, 29, 23) {real, imag} */,
  {32'h3d1e03e0, 32'h3c9a60b3} /* (2, 29, 22) {real, imag} */,
  {32'hbcf13add, 32'hbd30a678} /* (2, 29, 21) {real, imag} */,
  {32'h3b14d7a0, 32'h3cf698c0} /* (2, 29, 20) {real, imag} */,
  {32'hbcc693ad, 32'h3e0853ce} /* (2, 29, 19) {real, imag} */,
  {32'h3dbccd05, 32'h3cf437fe} /* (2, 29, 18) {real, imag} */,
  {32'hbd0be510, 32'hbc2f35bf} /* (2, 29, 17) {real, imag} */,
  {32'hbdcc1c6b, 32'h00000000} /* (2, 29, 16) {real, imag} */,
  {32'hbd0be510, 32'h3c2f35bf} /* (2, 29, 15) {real, imag} */,
  {32'h3dbccd05, 32'hbcf437fe} /* (2, 29, 14) {real, imag} */,
  {32'hbcc693ad, 32'hbe0853ce} /* (2, 29, 13) {real, imag} */,
  {32'h3b14d7a0, 32'hbcf698c0} /* (2, 29, 12) {real, imag} */,
  {32'hbcf13add, 32'h3d30a678} /* (2, 29, 11) {real, imag} */,
  {32'h3d1e03e0, 32'hbc9a60b3} /* (2, 29, 10) {real, imag} */,
  {32'hbce9359c, 32'hbdb9f0eb} /* (2, 29, 9) {real, imag} */,
  {32'h3e07c660, 32'h3da8209e} /* (2, 29, 8) {real, imag} */,
  {32'h3d14e1d8, 32'hbcd2013a} /* (2, 29, 7) {real, imag} */,
  {32'hbc6c67e0, 32'hbc50abe4} /* (2, 29, 6) {real, imag} */,
  {32'h3e93a75b, 32'h3dd71922} /* (2, 29, 5) {real, imag} */,
  {32'hbdd1846a, 32'hbcc5d9f4} /* (2, 29, 4) {real, imag} */,
  {32'h3df5f60e, 32'h3e718a87} /* (2, 29, 3) {real, imag} */,
  {32'h3f75c000, 32'h3bf21ec0} /* (2, 29, 2) {real, imag} */,
  {32'hbfd64dc6, 32'hbe7b2d58} /* (2, 29, 1) {real, imag} */,
  {32'hbf1325e4, 32'h00000000} /* (2, 29, 0) {real, imag} */,
  {32'hbfecfb29, 32'h3df6a888} /* (2, 28, 31) {real, imag} */,
  {32'h3f8d2378, 32'h3d1d8a2a} /* (2, 28, 30) {real, imag} */,
  {32'h3d8291f3, 32'hbe05f861} /* (2, 28, 29) {real, imag} */,
  {32'hbe05b184, 32'h3e0cb0d8} /* (2, 28, 28) {real, imag} */,
  {32'h3ea8f5a4, 32'hbe3655b4} /* (2, 28, 27) {real, imag} */,
  {32'h3c61e0a6, 32'hbc0c04f0} /* (2, 28, 26) {real, imag} */,
  {32'hbd9d1894, 32'h3e3c7d9d} /* (2, 28, 25) {real, imag} */,
  {32'h3d96c092, 32'h3d291555} /* (2, 28, 24) {real, imag} */,
  {32'hbd9f0158, 32'hbd8f8a09} /* (2, 28, 23) {real, imag} */,
  {32'hbc2f0429, 32'h3bcd5e90} /* (2, 28, 22) {real, imag} */,
  {32'h3d736f61, 32'hbd303064} /* (2, 28, 21) {real, imag} */,
  {32'h3da4ac29, 32'h3cbf34e8} /* (2, 28, 20) {real, imag} */,
  {32'h3c20e8e0, 32'h3d55339a} /* (2, 28, 19) {real, imag} */,
  {32'h3cedee1d, 32'h3be627fe} /* (2, 28, 18) {real, imag} */,
  {32'hbd5ad449, 32'hbd8b8da4} /* (2, 28, 17) {real, imag} */,
  {32'h3d648277, 32'h00000000} /* (2, 28, 16) {real, imag} */,
  {32'hbd5ad449, 32'h3d8b8da4} /* (2, 28, 15) {real, imag} */,
  {32'h3cedee1d, 32'hbbe627fe} /* (2, 28, 14) {real, imag} */,
  {32'h3c20e8e0, 32'hbd55339a} /* (2, 28, 13) {real, imag} */,
  {32'h3da4ac29, 32'hbcbf34e8} /* (2, 28, 12) {real, imag} */,
  {32'h3d736f61, 32'h3d303064} /* (2, 28, 11) {real, imag} */,
  {32'hbc2f0429, 32'hbbcd5e90} /* (2, 28, 10) {real, imag} */,
  {32'hbd9f0158, 32'h3d8f8a09} /* (2, 28, 9) {real, imag} */,
  {32'h3d96c092, 32'hbd291555} /* (2, 28, 8) {real, imag} */,
  {32'hbd9d1894, 32'hbe3c7d9d} /* (2, 28, 7) {real, imag} */,
  {32'h3c61e0a6, 32'h3c0c04f0} /* (2, 28, 6) {real, imag} */,
  {32'h3ea8f5a4, 32'h3e3655b4} /* (2, 28, 5) {real, imag} */,
  {32'hbe05b184, 32'hbe0cb0d8} /* (2, 28, 4) {real, imag} */,
  {32'h3d8291f3, 32'h3e05f861} /* (2, 28, 3) {real, imag} */,
  {32'h3f8d2378, 32'hbd1d8a2a} /* (2, 28, 2) {real, imag} */,
  {32'hbfecfb29, 32'hbdf6a888} /* (2, 28, 1) {real, imag} */,
  {32'hbf2b9c34, 32'h00000000} /* (2, 28, 0) {real, imag} */,
  {32'hbff64b7e, 32'h3dfa6c90} /* (2, 27, 31) {real, imag} */,
  {32'h3f797d96, 32'hbdcd985f} /* (2, 27, 30) {real, imag} */,
  {32'h3e0425b8, 32'hbe2d09e8} /* (2, 27, 29) {real, imag} */,
  {32'hbe345c40, 32'h3d1a704d} /* (2, 27, 28) {real, imag} */,
  {32'h3e5f5e1a, 32'hbe30c00c} /* (2, 27, 27) {real, imag} */,
  {32'hbcdc4b69, 32'hbcb48a16} /* (2, 27, 26) {real, imag} */,
  {32'h3c8d30aa, 32'h3d14d1ea} /* (2, 27, 25) {real, imag} */,
  {32'h3e44bd1e, 32'hbcb298dd} /* (2, 27, 24) {real, imag} */,
  {32'h3cf453c8, 32'h3d2e4d2a} /* (2, 27, 23) {real, imag} */,
  {32'h3d93ced9, 32'h3cbd261f} /* (2, 27, 22) {real, imag} */,
  {32'h3b002820, 32'hbd15e6e4} /* (2, 27, 21) {real, imag} */,
  {32'h3c648678, 32'h3dbcced9} /* (2, 27, 20) {real, imag} */,
  {32'hbdd9f0ff, 32'h3d28aba6} /* (2, 27, 19) {real, imag} */,
  {32'hbdc4975f, 32'hbce52c58} /* (2, 27, 18) {real, imag} */,
  {32'hbbabd578, 32'h3bc9fefc} /* (2, 27, 17) {real, imag} */,
  {32'hbdbb3816, 32'h00000000} /* (2, 27, 16) {real, imag} */,
  {32'hbbabd578, 32'hbbc9fefc} /* (2, 27, 15) {real, imag} */,
  {32'hbdc4975f, 32'h3ce52c58} /* (2, 27, 14) {real, imag} */,
  {32'hbdd9f0ff, 32'hbd28aba6} /* (2, 27, 13) {real, imag} */,
  {32'h3c648678, 32'hbdbcced9} /* (2, 27, 12) {real, imag} */,
  {32'h3b002820, 32'h3d15e6e4} /* (2, 27, 11) {real, imag} */,
  {32'h3d93ced9, 32'hbcbd261f} /* (2, 27, 10) {real, imag} */,
  {32'h3cf453c8, 32'hbd2e4d2a} /* (2, 27, 9) {real, imag} */,
  {32'h3e44bd1e, 32'h3cb298dd} /* (2, 27, 8) {real, imag} */,
  {32'h3c8d30aa, 32'hbd14d1ea} /* (2, 27, 7) {real, imag} */,
  {32'hbcdc4b69, 32'h3cb48a16} /* (2, 27, 6) {real, imag} */,
  {32'h3e5f5e1a, 32'h3e30c00c} /* (2, 27, 5) {real, imag} */,
  {32'hbe345c40, 32'hbd1a704d} /* (2, 27, 4) {real, imag} */,
  {32'h3e0425b8, 32'h3e2d09e8} /* (2, 27, 3) {real, imag} */,
  {32'h3f797d96, 32'h3dcd985f} /* (2, 27, 2) {real, imag} */,
  {32'hbff64b7e, 32'hbdfa6c90} /* (2, 27, 1) {real, imag} */,
  {32'hbf1a3520, 32'h00000000} /* (2, 27, 0) {real, imag} */,
  {32'hbff90fbb, 32'h3e592860} /* (2, 26, 31) {real, imag} */,
  {32'h3f550220, 32'hbd5d00f4} /* (2, 26, 30) {real, imag} */,
  {32'h3df31d94, 32'hbdc24364} /* (2, 26, 29) {real, imag} */,
  {32'hbe89fc3c, 32'h3d261cf2} /* (2, 26, 28) {real, imag} */,
  {32'h3e66c6ec, 32'hbde7c840} /* (2, 26, 27) {real, imag} */,
  {32'h3cfd18ce, 32'hbdc366a9} /* (2, 26, 26) {real, imag} */,
  {32'hbd520d71, 32'hbd77a026} /* (2, 26, 25) {real, imag} */,
  {32'h3e0a2718, 32'h3cceb9a5} /* (2, 26, 24) {real, imag} */,
  {32'hbc42eb8a, 32'h3d0beadd} /* (2, 26, 23) {real, imag} */,
  {32'h3d00d20c, 32'h3df8bed8} /* (2, 26, 22) {real, imag} */,
  {32'h3d706023, 32'hbd6cf621} /* (2, 26, 21) {real, imag} */,
  {32'hba4dc6c0, 32'hbc0b6d10} /* (2, 26, 20) {real, imag} */,
  {32'h3db5a7bd, 32'hbde5ebec} /* (2, 26, 19) {real, imag} */,
  {32'hbcaa705f, 32'h3d103a86} /* (2, 26, 18) {real, imag} */,
  {32'hbd6c005f, 32'h3accc590} /* (2, 26, 17) {real, imag} */,
  {32'h3da87456, 32'h00000000} /* (2, 26, 16) {real, imag} */,
  {32'hbd6c005f, 32'hbaccc590} /* (2, 26, 15) {real, imag} */,
  {32'hbcaa705f, 32'hbd103a86} /* (2, 26, 14) {real, imag} */,
  {32'h3db5a7bd, 32'h3de5ebec} /* (2, 26, 13) {real, imag} */,
  {32'hba4dc6c0, 32'h3c0b6d10} /* (2, 26, 12) {real, imag} */,
  {32'h3d706023, 32'h3d6cf621} /* (2, 26, 11) {real, imag} */,
  {32'h3d00d20c, 32'hbdf8bed8} /* (2, 26, 10) {real, imag} */,
  {32'hbc42eb8a, 32'hbd0beadd} /* (2, 26, 9) {real, imag} */,
  {32'h3e0a2718, 32'hbcceb9a5} /* (2, 26, 8) {real, imag} */,
  {32'hbd520d71, 32'h3d77a026} /* (2, 26, 7) {real, imag} */,
  {32'h3cfd18ce, 32'h3dc366a9} /* (2, 26, 6) {real, imag} */,
  {32'h3e66c6ec, 32'h3de7c840} /* (2, 26, 5) {real, imag} */,
  {32'hbe89fc3c, 32'hbd261cf2} /* (2, 26, 4) {real, imag} */,
  {32'h3df31d94, 32'h3dc24364} /* (2, 26, 3) {real, imag} */,
  {32'h3f550220, 32'h3d5d00f4} /* (2, 26, 2) {real, imag} */,
  {32'hbff90fbb, 32'hbe592860} /* (2, 26, 1) {real, imag} */,
  {32'hbee7416e, 32'h00000000} /* (2, 26, 0) {real, imag} */,
  {32'hc0003bbd, 32'h3e2f920c} /* (2, 25, 31) {real, imag} */,
  {32'h3f634fac, 32'hbd7a4a7a} /* (2, 25, 30) {real, imag} */,
  {32'h3db65f2c, 32'hbde28299} /* (2, 25, 29) {real, imag} */,
  {32'hbea9c8e6, 32'h3dad6016} /* (2, 25, 28) {real, imag} */,
  {32'h3dce57d4, 32'hbd807738} /* (2, 25, 27) {real, imag} */,
  {32'h3d37a780, 32'hbdaca2a5} /* (2, 25, 26) {real, imag} */,
  {32'hbcd99f08, 32'h3d9cb5ce} /* (2, 25, 25) {real, imag} */,
  {32'h3cc1e119, 32'hbdd477f2} /* (2, 25, 24) {real, imag} */,
  {32'h3dd73bcc, 32'h3c655a18} /* (2, 25, 23) {real, imag} */,
  {32'hbd89c7d3, 32'h3de7cd40} /* (2, 25, 22) {real, imag} */,
  {32'h3d545d51, 32'hbd928e7c} /* (2, 25, 21) {real, imag} */,
  {32'hbd8c3086, 32'hbd50e904} /* (2, 25, 20) {real, imag} */,
  {32'hbdda92c1, 32'h39f0c700} /* (2, 25, 19) {real, imag} */,
  {32'hbc8d441a, 32'hbc907e7a} /* (2, 25, 18) {real, imag} */,
  {32'hbd588ec4, 32'h3c6c9c50} /* (2, 25, 17) {real, imag} */,
  {32'hbd48845d, 32'h00000000} /* (2, 25, 16) {real, imag} */,
  {32'hbd588ec4, 32'hbc6c9c50} /* (2, 25, 15) {real, imag} */,
  {32'hbc8d441a, 32'h3c907e7a} /* (2, 25, 14) {real, imag} */,
  {32'hbdda92c1, 32'hb9f0c700} /* (2, 25, 13) {real, imag} */,
  {32'hbd8c3086, 32'h3d50e904} /* (2, 25, 12) {real, imag} */,
  {32'h3d545d51, 32'h3d928e7c} /* (2, 25, 11) {real, imag} */,
  {32'hbd89c7d3, 32'hbde7cd40} /* (2, 25, 10) {real, imag} */,
  {32'h3dd73bcc, 32'hbc655a18} /* (2, 25, 9) {real, imag} */,
  {32'h3cc1e119, 32'h3dd477f2} /* (2, 25, 8) {real, imag} */,
  {32'hbcd99f08, 32'hbd9cb5ce} /* (2, 25, 7) {real, imag} */,
  {32'h3d37a780, 32'h3daca2a5} /* (2, 25, 6) {real, imag} */,
  {32'h3dce57d4, 32'h3d807738} /* (2, 25, 5) {real, imag} */,
  {32'hbea9c8e6, 32'hbdad6016} /* (2, 25, 4) {real, imag} */,
  {32'h3db65f2c, 32'h3de28299} /* (2, 25, 3) {real, imag} */,
  {32'h3f634fac, 32'h3d7a4a7a} /* (2, 25, 2) {real, imag} */,
  {32'hc0003bbd, 32'hbe2f920c} /* (2, 25, 1) {real, imag} */,
  {32'hbf18c7d9, 32'h00000000} /* (2, 25, 0) {real, imag} */,
  {32'hbff82a5d, 32'h3d2f9b14} /* (2, 24, 31) {real, imag} */,
  {32'h3f4fba2c, 32'h3d256cd0} /* (2, 24, 30) {real, imag} */,
  {32'h3c80a906, 32'hbe35876c} /* (2, 24, 29) {real, imag} */,
  {32'hbe7c12c2, 32'hbba6b2e0} /* (2, 24, 28) {real, imag} */,
  {32'h3defa661, 32'hbdec054e} /* (2, 24, 27) {real, imag} */,
  {32'hbd639d5e, 32'h3d6f44d5} /* (2, 24, 26) {real, imag} */,
  {32'hbd6ccab8, 32'hbc97a788} /* (2, 24, 25) {real, imag} */,
  {32'h3e4343e3, 32'hbd45f767} /* (2, 24, 24) {real, imag} */,
  {32'h3ce82cbe, 32'h3ce84ca1} /* (2, 24, 23) {real, imag} */,
  {32'hbdbfc672, 32'hbccf30b4} /* (2, 24, 22) {real, imag} */,
  {32'h3d9dd1d0, 32'hbd02281c} /* (2, 24, 21) {real, imag} */,
  {32'h3d3ba2eb, 32'hbd18c0c5} /* (2, 24, 20) {real, imag} */,
  {32'hbd55bd40, 32'h3d86e9ea} /* (2, 24, 19) {real, imag} */,
  {32'h3a801360, 32'hbd875463} /* (2, 24, 18) {real, imag} */,
  {32'h3d3ecd66, 32'hbd696c0b} /* (2, 24, 17) {real, imag} */,
  {32'h3cf2eb33, 32'h00000000} /* (2, 24, 16) {real, imag} */,
  {32'h3d3ecd66, 32'h3d696c0b} /* (2, 24, 15) {real, imag} */,
  {32'h3a801360, 32'h3d875463} /* (2, 24, 14) {real, imag} */,
  {32'hbd55bd40, 32'hbd86e9ea} /* (2, 24, 13) {real, imag} */,
  {32'h3d3ba2eb, 32'h3d18c0c5} /* (2, 24, 12) {real, imag} */,
  {32'h3d9dd1d0, 32'h3d02281c} /* (2, 24, 11) {real, imag} */,
  {32'hbdbfc672, 32'h3ccf30b4} /* (2, 24, 10) {real, imag} */,
  {32'h3ce82cbe, 32'hbce84ca1} /* (2, 24, 9) {real, imag} */,
  {32'h3e4343e3, 32'h3d45f767} /* (2, 24, 8) {real, imag} */,
  {32'hbd6ccab8, 32'h3c97a788} /* (2, 24, 7) {real, imag} */,
  {32'hbd639d5e, 32'hbd6f44d5} /* (2, 24, 6) {real, imag} */,
  {32'h3defa661, 32'h3dec054e} /* (2, 24, 5) {real, imag} */,
  {32'hbe7c12c2, 32'h3ba6b2e0} /* (2, 24, 4) {real, imag} */,
  {32'h3c80a906, 32'h3e35876c} /* (2, 24, 3) {real, imag} */,
  {32'h3f4fba2c, 32'hbd256cd0} /* (2, 24, 2) {real, imag} */,
  {32'hbff82a5d, 32'hbd2f9b14} /* (2, 24, 1) {real, imag} */,
  {32'hbf414f50, 32'h00000000} /* (2, 24, 0) {real, imag} */,
  {32'hbfde55de, 32'h3d2d4ea4} /* (2, 23, 31) {real, imag} */,
  {32'h3f23fb19, 32'h3d74597e} /* (2, 23, 30) {real, imag} */,
  {32'hbd5bdbd0, 32'hbdd1b60e} /* (2, 23, 29) {real, imag} */,
  {32'hbe57c014, 32'h3c8afe38} /* (2, 23, 28) {real, imag} */,
  {32'h3dfe002e, 32'hbe6d3ff2} /* (2, 23, 27) {real, imag} */,
  {32'hbc662854, 32'hbbfd5a34} /* (2, 23, 26) {real, imag} */,
  {32'hbce5ef49, 32'hbd162d58} /* (2, 23, 25) {real, imag} */,
  {32'h3d758a50, 32'hbdf138b4} /* (2, 23, 24) {real, imag} */,
  {32'h3d376254, 32'hbe2020e0} /* (2, 23, 23) {real, imag} */,
  {32'hbd1b872f, 32'h3d25cdc0} /* (2, 23, 22) {real, imag} */,
  {32'h3d57bf8d, 32'hbe12e28c} /* (2, 23, 21) {real, imag} */,
  {32'h3d725586, 32'h3d2d13da} /* (2, 23, 20) {real, imag} */,
  {32'h3d5adbb2, 32'h3d254c22} /* (2, 23, 19) {real, imag} */,
  {32'hbc83a022, 32'h3d0be862} /* (2, 23, 18) {real, imag} */,
  {32'h3de85dae, 32'h3b587a00} /* (2, 23, 17) {real, imag} */,
  {32'h3d60bb50, 32'h00000000} /* (2, 23, 16) {real, imag} */,
  {32'h3de85dae, 32'hbb587a00} /* (2, 23, 15) {real, imag} */,
  {32'hbc83a022, 32'hbd0be862} /* (2, 23, 14) {real, imag} */,
  {32'h3d5adbb2, 32'hbd254c22} /* (2, 23, 13) {real, imag} */,
  {32'h3d725586, 32'hbd2d13da} /* (2, 23, 12) {real, imag} */,
  {32'h3d57bf8d, 32'h3e12e28c} /* (2, 23, 11) {real, imag} */,
  {32'hbd1b872f, 32'hbd25cdc0} /* (2, 23, 10) {real, imag} */,
  {32'h3d376254, 32'h3e2020e0} /* (2, 23, 9) {real, imag} */,
  {32'h3d758a50, 32'h3df138b4} /* (2, 23, 8) {real, imag} */,
  {32'hbce5ef49, 32'h3d162d58} /* (2, 23, 7) {real, imag} */,
  {32'hbc662854, 32'h3bfd5a34} /* (2, 23, 6) {real, imag} */,
  {32'h3dfe002e, 32'h3e6d3ff2} /* (2, 23, 5) {real, imag} */,
  {32'hbe57c014, 32'hbc8afe38} /* (2, 23, 4) {real, imag} */,
  {32'hbd5bdbd0, 32'h3dd1b60e} /* (2, 23, 3) {real, imag} */,
  {32'h3f23fb19, 32'hbd74597e} /* (2, 23, 2) {real, imag} */,
  {32'hbfde55de, 32'hbd2d4ea4} /* (2, 23, 1) {real, imag} */,
  {32'hbf0cacc7, 32'h00000000} /* (2, 23, 0) {real, imag} */,
  {32'hbfa9d95a, 32'hbc26a7d0} /* (2, 22, 31) {real, imag} */,
  {32'h3f0dae01, 32'hbcec6178} /* (2, 22, 30) {real, imag} */,
  {32'hbd94a4e4, 32'h3e0f4463} /* (2, 22, 29) {real, imag} */,
  {32'hbe499d8b, 32'hbce4f424} /* (2, 22, 28) {real, imag} */,
  {32'h3e478f3a, 32'hbe2881af} /* (2, 22, 27) {real, imag} */,
  {32'hbd99fe32, 32'h3cb08350} /* (2, 22, 26) {real, imag} */,
  {32'h3d4c0a8c, 32'h3d1b7832} /* (2, 22, 25) {real, imag} */,
  {32'hbd618dfc, 32'hbd9fd098} /* (2, 22, 24) {real, imag} */,
  {32'hbc9cc198, 32'h3d2fb4ab} /* (2, 22, 23) {real, imag} */,
  {32'h3db613cc, 32'h3a5d8400} /* (2, 22, 22) {real, imag} */,
  {32'hbdb8d642, 32'hbd6df531} /* (2, 22, 21) {real, imag} */,
  {32'hbe091f16, 32'h3dbfb556} /* (2, 22, 20) {real, imag} */,
  {32'hbd85f37a, 32'hbcc5cbbe} /* (2, 22, 19) {real, imag} */,
  {32'h3cebbd55, 32'hbcb53b0e} /* (2, 22, 18) {real, imag} */,
  {32'hbd265c22, 32'h3d7c463e} /* (2, 22, 17) {real, imag} */,
  {32'h3cd01c10, 32'h00000000} /* (2, 22, 16) {real, imag} */,
  {32'hbd265c22, 32'hbd7c463e} /* (2, 22, 15) {real, imag} */,
  {32'h3cebbd55, 32'h3cb53b0e} /* (2, 22, 14) {real, imag} */,
  {32'hbd85f37a, 32'h3cc5cbbe} /* (2, 22, 13) {real, imag} */,
  {32'hbe091f16, 32'hbdbfb556} /* (2, 22, 12) {real, imag} */,
  {32'hbdb8d642, 32'h3d6df531} /* (2, 22, 11) {real, imag} */,
  {32'h3db613cc, 32'hba5d8400} /* (2, 22, 10) {real, imag} */,
  {32'hbc9cc198, 32'hbd2fb4ab} /* (2, 22, 9) {real, imag} */,
  {32'hbd618dfc, 32'h3d9fd098} /* (2, 22, 8) {real, imag} */,
  {32'h3d4c0a8c, 32'hbd1b7832} /* (2, 22, 7) {real, imag} */,
  {32'hbd99fe32, 32'hbcb08350} /* (2, 22, 6) {real, imag} */,
  {32'h3e478f3a, 32'h3e2881af} /* (2, 22, 5) {real, imag} */,
  {32'hbe499d8b, 32'h3ce4f424} /* (2, 22, 4) {real, imag} */,
  {32'hbd94a4e4, 32'hbe0f4463} /* (2, 22, 3) {real, imag} */,
  {32'h3f0dae01, 32'h3cec6178} /* (2, 22, 2) {real, imag} */,
  {32'hbfa9d95a, 32'h3c26a7d0} /* (2, 22, 1) {real, imag} */,
  {32'hbec501ea, 32'h00000000} /* (2, 22, 0) {real, imag} */,
  {32'hbf138ae5, 32'hbdceda50} /* (2, 21, 31) {real, imag} */,
  {32'h3db914b0, 32'hbd00009b} /* (2, 21, 30) {real, imag} */,
  {32'hbdc49330, 32'h3c902fe4} /* (2, 21, 29) {real, imag} */,
  {32'hbc7dac50, 32'h3cd8e346} /* (2, 21, 28) {real, imag} */,
  {32'h3cca807c, 32'hbe48f586} /* (2, 21, 27) {real, imag} */,
  {32'h3ad44060, 32'h3b9168e0} /* (2, 21, 26) {real, imag} */,
  {32'hbcfc0446, 32'h3dc4ad44} /* (2, 21, 25) {real, imag} */,
  {32'hbc9d4da0, 32'h3c87d93e} /* (2, 21, 24) {real, imag} */,
  {32'hbd244bf1, 32'hbcc208c1} /* (2, 21, 23) {real, imag} */,
  {32'h3df9c4f4, 32'h3d90ba86} /* (2, 21, 22) {real, imag} */,
  {32'h3c02fe90, 32'hbdecdbd6} /* (2, 21, 21) {real, imag} */,
  {32'h3d108346, 32'h3c584106} /* (2, 21, 20) {real, imag} */,
  {32'hbd240b6e, 32'h3cf8619e} /* (2, 21, 19) {real, imag} */,
  {32'h3d326026, 32'hbd05bb6d} /* (2, 21, 18) {real, imag} */,
  {32'hbcc1b7ef, 32'h3c87e687} /* (2, 21, 17) {real, imag} */,
  {32'h3ce5a811, 32'h00000000} /* (2, 21, 16) {real, imag} */,
  {32'hbcc1b7ef, 32'hbc87e687} /* (2, 21, 15) {real, imag} */,
  {32'h3d326026, 32'h3d05bb6d} /* (2, 21, 14) {real, imag} */,
  {32'hbd240b6e, 32'hbcf8619e} /* (2, 21, 13) {real, imag} */,
  {32'h3d108346, 32'hbc584106} /* (2, 21, 12) {real, imag} */,
  {32'h3c02fe90, 32'h3decdbd6} /* (2, 21, 11) {real, imag} */,
  {32'h3df9c4f4, 32'hbd90ba86} /* (2, 21, 10) {real, imag} */,
  {32'hbd244bf1, 32'h3cc208c1} /* (2, 21, 9) {real, imag} */,
  {32'hbc9d4da0, 32'hbc87d93e} /* (2, 21, 8) {real, imag} */,
  {32'hbcfc0446, 32'hbdc4ad44} /* (2, 21, 7) {real, imag} */,
  {32'h3ad44060, 32'hbb9168e0} /* (2, 21, 6) {real, imag} */,
  {32'h3cca807c, 32'h3e48f586} /* (2, 21, 5) {real, imag} */,
  {32'hbc7dac50, 32'hbcd8e346} /* (2, 21, 4) {real, imag} */,
  {32'hbdc49330, 32'hbc902fe4} /* (2, 21, 3) {real, imag} */,
  {32'h3db914b0, 32'h3d00009b} /* (2, 21, 2) {real, imag} */,
  {32'hbf138ae5, 32'h3dceda50} /* (2, 21, 1) {real, imag} */,
  {32'h3d8ab888, 32'h00000000} /* (2, 21, 0) {real, imag} */,
  {32'h3f2dec8d, 32'hbea943e1} /* (2, 20, 31) {real, imag} */,
  {32'hbf02f12b, 32'h3d97af58} /* (2, 20, 30) {real, imag} */,
  {32'hbe4603ba, 32'hbc14f602} /* (2, 20, 29) {real, imag} */,
  {32'h3d37cb54, 32'hbcdff3c6} /* (2, 20, 28) {real, imag} */,
  {32'hbe0b0db2, 32'hbd911e8f} /* (2, 20, 27) {real, imag} */,
  {32'h3b50d0a0, 32'h3d922b8c} /* (2, 20, 26) {real, imag} */,
  {32'hba5da420, 32'h3dacdefa} /* (2, 20, 25) {real, imag} */,
  {32'h3b906bea, 32'h3dd9c80e} /* (2, 20, 24) {real, imag} */,
  {32'hbce5c19d, 32'h3be7b954} /* (2, 20, 23) {real, imag} */,
  {32'h3b001118, 32'hbe3f1014} /* (2, 20, 22) {real, imag} */,
  {32'hbd4f4f2e, 32'h3dbb78b6} /* (2, 20, 21) {real, imag} */,
  {32'hbc5a5924, 32'h3d232210} /* (2, 20, 20) {real, imag} */,
  {32'h3d05ad32, 32'h3d897ea8} /* (2, 20, 19) {real, imag} */,
  {32'h3d8046da, 32'hbd5a9960} /* (2, 20, 18) {real, imag} */,
  {32'h3d176a84, 32'h3bafeab2} /* (2, 20, 17) {real, imag} */,
  {32'h3b9bcda0, 32'h00000000} /* (2, 20, 16) {real, imag} */,
  {32'h3d176a84, 32'hbbafeab2} /* (2, 20, 15) {real, imag} */,
  {32'h3d8046da, 32'h3d5a9960} /* (2, 20, 14) {real, imag} */,
  {32'h3d05ad32, 32'hbd897ea8} /* (2, 20, 13) {real, imag} */,
  {32'hbc5a5924, 32'hbd232210} /* (2, 20, 12) {real, imag} */,
  {32'hbd4f4f2e, 32'hbdbb78b6} /* (2, 20, 11) {real, imag} */,
  {32'h3b001118, 32'h3e3f1014} /* (2, 20, 10) {real, imag} */,
  {32'hbce5c19d, 32'hbbe7b954} /* (2, 20, 9) {real, imag} */,
  {32'h3b906bea, 32'hbdd9c80e} /* (2, 20, 8) {real, imag} */,
  {32'hba5da420, 32'hbdacdefa} /* (2, 20, 7) {real, imag} */,
  {32'h3b50d0a0, 32'hbd922b8c} /* (2, 20, 6) {real, imag} */,
  {32'hbe0b0db2, 32'h3d911e8f} /* (2, 20, 5) {real, imag} */,
  {32'h3d37cb54, 32'h3cdff3c6} /* (2, 20, 4) {real, imag} */,
  {32'hbe4603ba, 32'h3c14f602} /* (2, 20, 3) {real, imag} */,
  {32'hbf02f12b, 32'hbd97af58} /* (2, 20, 2) {real, imag} */,
  {32'h3f2dec8d, 32'h3ea943e1} /* (2, 20, 1) {real, imag} */,
  {32'h3f466964, 32'h00000000} /* (2, 20, 0) {real, imag} */,
  {32'h3fa1774f, 32'hbebe1754} /* (2, 19, 31) {real, imag} */,
  {32'hbf48bd10, 32'h3c15ab98} /* (2, 19, 30) {real, imag} */,
  {32'hbdc6135e, 32'h3e046cb4} /* (2, 19, 29) {real, imag} */,
  {32'h3e2cf01f, 32'hbd8b41b1} /* (2, 19, 28) {real, imag} */,
  {32'hbe44f50d, 32'h3d8a1d5f} /* (2, 19, 27) {real, imag} */,
  {32'hbd0e5d02, 32'h3d3fab80} /* (2, 19, 26) {real, imag} */,
  {32'h3c8c47a8, 32'h3d4c9d52} /* (2, 19, 25) {real, imag} */,
  {32'hbb9e3400, 32'hbc5c6720} /* (2, 19, 24) {real, imag} */,
  {32'hbcde8e8c, 32'hbe006ce9} /* (2, 19, 23) {real, imag} */,
  {32'hbce89904, 32'hbd4e1807} /* (2, 19, 22) {real, imag} */,
  {32'hbe1f15bc, 32'h3c1a74e0} /* (2, 19, 21) {real, imag} */,
  {32'h3c8e1640, 32'h3cf281ad} /* (2, 19, 20) {real, imag} */,
  {32'h3c2d1986, 32'hbdaf036c} /* (2, 19, 19) {real, imag} */,
  {32'hbd51beb4, 32'h3d9ffac8} /* (2, 19, 18) {real, imag} */,
  {32'hbc3fefa8, 32'h3c98077e} /* (2, 19, 17) {real, imag} */,
  {32'h3d462c37, 32'h00000000} /* (2, 19, 16) {real, imag} */,
  {32'hbc3fefa8, 32'hbc98077e} /* (2, 19, 15) {real, imag} */,
  {32'hbd51beb4, 32'hbd9ffac8} /* (2, 19, 14) {real, imag} */,
  {32'h3c2d1986, 32'h3daf036c} /* (2, 19, 13) {real, imag} */,
  {32'h3c8e1640, 32'hbcf281ad} /* (2, 19, 12) {real, imag} */,
  {32'hbe1f15bc, 32'hbc1a74e0} /* (2, 19, 11) {real, imag} */,
  {32'hbce89904, 32'h3d4e1807} /* (2, 19, 10) {real, imag} */,
  {32'hbcde8e8c, 32'h3e006ce9} /* (2, 19, 9) {real, imag} */,
  {32'hbb9e3400, 32'h3c5c6720} /* (2, 19, 8) {real, imag} */,
  {32'h3c8c47a8, 32'hbd4c9d52} /* (2, 19, 7) {real, imag} */,
  {32'hbd0e5d02, 32'hbd3fab80} /* (2, 19, 6) {real, imag} */,
  {32'hbe44f50d, 32'hbd8a1d5f} /* (2, 19, 5) {real, imag} */,
  {32'h3e2cf01f, 32'h3d8b41b1} /* (2, 19, 4) {real, imag} */,
  {32'hbdc6135e, 32'hbe046cb4} /* (2, 19, 3) {real, imag} */,
  {32'hbf48bd10, 32'hbc15ab98} /* (2, 19, 2) {real, imag} */,
  {32'h3fa1774f, 32'h3ebe1754} /* (2, 19, 1) {real, imag} */,
  {32'h3f909813, 32'h00000000} /* (2, 19, 0) {real, imag} */,
  {32'h3fc78701, 32'hbe996ed0} /* (2, 18, 31) {real, imag} */,
  {32'hbf5ab0ea, 32'hbca80910} /* (2, 18, 30) {real, imag} */,
  {32'hbe27faca, 32'h3d81ac5c} /* (2, 18, 29) {real, imag} */,
  {32'h3e69408c, 32'hbda3f7e0} /* (2, 18, 28) {real, imag} */,
  {32'hbe0aa292, 32'h3e3c3ff1} /* (2, 18, 27) {real, imag} */,
  {32'hbd300c28, 32'hbcfb95c3} /* (2, 18, 26) {real, imag} */,
  {32'h38ad5300, 32'hbd337d34} /* (2, 18, 25) {real, imag} */,
  {32'hbd7e0d3a, 32'h3db3cc8d} /* (2, 18, 24) {real, imag} */,
  {32'hbb60d766, 32'h3be71797} /* (2, 18, 23) {real, imag} */,
  {32'h3b2df800, 32'h3d34a267} /* (2, 18, 22) {real, imag} */,
  {32'hbe18a243, 32'h3bde4122} /* (2, 18, 21) {real, imag} */,
  {32'hbd7ade6e, 32'hbd164d91} /* (2, 18, 20) {real, imag} */,
  {32'h3d2af93f, 32'hbd04d9ac} /* (2, 18, 19) {real, imag} */,
  {32'h3d114321, 32'h3d7d0192} /* (2, 18, 18) {real, imag} */,
  {32'h3d1734e2, 32'hbcc047ad} /* (2, 18, 17) {real, imag} */,
  {32'hbb249440, 32'h00000000} /* (2, 18, 16) {real, imag} */,
  {32'h3d1734e2, 32'h3cc047ad} /* (2, 18, 15) {real, imag} */,
  {32'h3d114321, 32'hbd7d0192} /* (2, 18, 14) {real, imag} */,
  {32'h3d2af93f, 32'h3d04d9ac} /* (2, 18, 13) {real, imag} */,
  {32'hbd7ade6e, 32'h3d164d91} /* (2, 18, 12) {real, imag} */,
  {32'hbe18a243, 32'hbbde4122} /* (2, 18, 11) {real, imag} */,
  {32'h3b2df800, 32'hbd34a267} /* (2, 18, 10) {real, imag} */,
  {32'hbb60d766, 32'hbbe71797} /* (2, 18, 9) {real, imag} */,
  {32'hbd7e0d3a, 32'hbdb3cc8d} /* (2, 18, 8) {real, imag} */,
  {32'h38ad5300, 32'h3d337d34} /* (2, 18, 7) {real, imag} */,
  {32'hbd300c28, 32'h3cfb95c3} /* (2, 18, 6) {real, imag} */,
  {32'hbe0aa292, 32'hbe3c3ff1} /* (2, 18, 5) {real, imag} */,
  {32'h3e69408c, 32'h3da3f7e0} /* (2, 18, 4) {real, imag} */,
  {32'hbe27faca, 32'hbd81ac5c} /* (2, 18, 3) {real, imag} */,
  {32'hbf5ab0ea, 32'h3ca80910} /* (2, 18, 2) {real, imag} */,
  {32'h3fc78701, 32'h3e996ed0} /* (2, 18, 1) {real, imag} */,
  {32'h3f8f053e, 32'h00000000} /* (2, 18, 0) {real, imag} */,
  {32'h3fd86287, 32'hbe6e8093} /* (2, 17, 31) {real, imag} */,
  {32'hbf75082a, 32'h3de49f38} /* (2, 17, 30) {real, imag} */,
  {32'h3b2ae4b0, 32'hbca247af} /* (2, 17, 29) {real, imag} */,
  {32'h3dc255b7, 32'hbe657edd} /* (2, 17, 28) {real, imag} */,
  {32'hbd859522, 32'h3e10f6aa} /* (2, 17, 27) {real, imag} */,
  {32'h3c9b74dc, 32'h398895e0} /* (2, 17, 26) {real, imag} */,
  {32'h3c46e49e, 32'h3d731701} /* (2, 17, 25) {real, imag} */,
  {32'hbd8b888e, 32'hbd7791ef} /* (2, 17, 24) {real, imag} */,
  {32'hbc96f035, 32'h3dd0f829} /* (2, 17, 23) {real, imag} */,
  {32'h3db7b442, 32'hbdbc7b87} /* (2, 17, 22) {real, imag} */,
  {32'h3dbcefe4, 32'h3d99e201} /* (2, 17, 21) {real, imag} */,
  {32'h3bd79440, 32'h3c3f5c98} /* (2, 17, 20) {real, imag} */,
  {32'hb996c280, 32'h3bd51116} /* (2, 17, 19) {real, imag} */,
  {32'h3d3fb16d, 32'hbdbb9e40} /* (2, 17, 18) {real, imag} */,
  {32'hbd034ac2, 32'hbcac7a10} /* (2, 17, 17) {real, imag} */,
  {32'h3c497d40, 32'h00000000} /* (2, 17, 16) {real, imag} */,
  {32'hbd034ac2, 32'h3cac7a10} /* (2, 17, 15) {real, imag} */,
  {32'h3d3fb16d, 32'h3dbb9e40} /* (2, 17, 14) {real, imag} */,
  {32'hb996c280, 32'hbbd51116} /* (2, 17, 13) {real, imag} */,
  {32'h3bd79440, 32'hbc3f5c98} /* (2, 17, 12) {real, imag} */,
  {32'h3dbcefe4, 32'hbd99e201} /* (2, 17, 11) {real, imag} */,
  {32'h3db7b442, 32'h3dbc7b87} /* (2, 17, 10) {real, imag} */,
  {32'hbc96f035, 32'hbdd0f829} /* (2, 17, 9) {real, imag} */,
  {32'hbd8b888e, 32'h3d7791ef} /* (2, 17, 8) {real, imag} */,
  {32'h3c46e49e, 32'hbd731701} /* (2, 17, 7) {real, imag} */,
  {32'h3c9b74dc, 32'hb98895e0} /* (2, 17, 6) {real, imag} */,
  {32'hbd859522, 32'hbe10f6aa} /* (2, 17, 5) {real, imag} */,
  {32'h3dc255b7, 32'h3e657edd} /* (2, 17, 4) {real, imag} */,
  {32'h3b2ae4b0, 32'h3ca247af} /* (2, 17, 3) {real, imag} */,
  {32'hbf75082a, 32'hbde49f38} /* (2, 17, 2) {real, imag} */,
  {32'h3fd86287, 32'h3e6e8093} /* (2, 17, 1) {real, imag} */,
  {32'h3f8ea7b3, 32'h00000000} /* (2, 17, 0) {real, imag} */,
  {32'h3fe14996, 32'hbe587a34} /* (2, 16, 31) {real, imag} */,
  {32'hbf61adae, 32'h3e240e60} /* (2, 16, 30) {real, imag} */,
  {32'h3db08626, 32'h3d7bb436} /* (2, 16, 29) {real, imag} */,
  {32'h3e5b42b1, 32'hbe0d230d} /* (2, 16, 28) {real, imag} */,
  {32'hbe1a1e2e, 32'h3da7d12f} /* (2, 16, 27) {real, imag} */,
  {32'hbc25d8d2, 32'h3d3b030b} /* (2, 16, 26) {real, imag} */,
  {32'h3bd2e618, 32'hbdec8a38} /* (2, 16, 25) {real, imag} */,
  {32'hbe258804, 32'h3c93f2c0} /* (2, 16, 24) {real, imag} */,
  {32'h3c11f9ea, 32'hbdbdc523} /* (2, 16, 23) {real, imag} */,
  {32'h3d3d19c0, 32'hbd9def97} /* (2, 16, 22) {real, imag} */,
  {32'h3b459c80, 32'hbcd9cf30} /* (2, 16, 21) {real, imag} */,
  {32'h3d81a096, 32'hbd39cba9} /* (2, 16, 20) {real, imag} */,
  {32'h3c93596b, 32'h3d0f449c} /* (2, 16, 19) {real, imag} */,
  {32'hbc883dd4, 32'h3dcb642e} /* (2, 16, 18) {real, imag} */,
  {32'h3c860f3e, 32'h3b0b9370} /* (2, 16, 17) {real, imag} */,
  {32'h3d01d1a0, 32'h00000000} /* (2, 16, 16) {real, imag} */,
  {32'h3c860f3e, 32'hbb0b9370} /* (2, 16, 15) {real, imag} */,
  {32'hbc883dd4, 32'hbdcb642e} /* (2, 16, 14) {real, imag} */,
  {32'h3c93596b, 32'hbd0f449c} /* (2, 16, 13) {real, imag} */,
  {32'h3d81a096, 32'h3d39cba9} /* (2, 16, 12) {real, imag} */,
  {32'h3b459c80, 32'h3cd9cf30} /* (2, 16, 11) {real, imag} */,
  {32'h3d3d19c0, 32'h3d9def97} /* (2, 16, 10) {real, imag} */,
  {32'h3c11f9ea, 32'h3dbdc523} /* (2, 16, 9) {real, imag} */,
  {32'hbe258804, 32'hbc93f2c0} /* (2, 16, 8) {real, imag} */,
  {32'h3bd2e618, 32'h3dec8a38} /* (2, 16, 7) {real, imag} */,
  {32'hbc25d8d2, 32'hbd3b030b} /* (2, 16, 6) {real, imag} */,
  {32'hbe1a1e2e, 32'hbda7d12f} /* (2, 16, 5) {real, imag} */,
  {32'h3e5b42b1, 32'h3e0d230d} /* (2, 16, 4) {real, imag} */,
  {32'h3db08626, 32'hbd7bb436} /* (2, 16, 3) {real, imag} */,
  {32'hbf61adae, 32'hbe240e60} /* (2, 16, 2) {real, imag} */,
  {32'h3fe14996, 32'h3e587a34} /* (2, 16, 1) {real, imag} */,
  {32'h3fa2e624, 32'h00000000} /* (2, 16, 0) {real, imag} */,
  {32'h3fe1a4cd, 32'hbe8458c8} /* (2, 15, 31) {real, imag} */,
  {32'hbf4a9112, 32'h3e0a2c30} /* (2, 15, 30) {real, imag} */,
  {32'h3d82965e, 32'hbd126220} /* (2, 15, 29) {real, imag} */,
  {32'h3e2e0488, 32'hbddeb526} /* (2, 15, 28) {real, imag} */,
  {32'hbe2d48c2, 32'h3e20cea0} /* (2, 15, 27) {real, imag} */,
  {32'hbdd08703, 32'h3bc71d7e} /* (2, 15, 26) {real, imag} */,
  {32'h3b93831c, 32'hbd8b0f0e} /* (2, 15, 25) {real, imag} */,
  {32'hbc44769c, 32'hbd09e0c9} /* (2, 15, 24) {real, imag} */,
  {32'h3d4a5bee, 32'h3c8374e8} /* (2, 15, 23) {real, imag} */,
  {32'hbd2efcac, 32'hbd19e48e} /* (2, 15, 22) {real, imag} */,
  {32'hbe097bc2, 32'h3d37794c} /* (2, 15, 21) {real, imag} */,
  {32'hbcd05494, 32'hbdaa7308} /* (2, 15, 20) {real, imag} */,
  {32'hbd0bbaec, 32'hbc7a1027} /* (2, 15, 19) {real, imag} */,
  {32'hbce50aee, 32'h3cf44122} /* (2, 15, 18) {real, imag} */,
  {32'h3b33fd20, 32'h3d2331a8} /* (2, 15, 17) {real, imag} */,
  {32'h3d3d945a, 32'h00000000} /* (2, 15, 16) {real, imag} */,
  {32'h3b33fd20, 32'hbd2331a8} /* (2, 15, 15) {real, imag} */,
  {32'hbce50aee, 32'hbcf44122} /* (2, 15, 14) {real, imag} */,
  {32'hbd0bbaec, 32'h3c7a1027} /* (2, 15, 13) {real, imag} */,
  {32'hbcd05494, 32'h3daa7308} /* (2, 15, 12) {real, imag} */,
  {32'hbe097bc2, 32'hbd37794c} /* (2, 15, 11) {real, imag} */,
  {32'hbd2efcac, 32'h3d19e48e} /* (2, 15, 10) {real, imag} */,
  {32'h3d4a5bee, 32'hbc8374e8} /* (2, 15, 9) {real, imag} */,
  {32'hbc44769c, 32'h3d09e0c9} /* (2, 15, 8) {real, imag} */,
  {32'h3b93831c, 32'h3d8b0f0e} /* (2, 15, 7) {real, imag} */,
  {32'hbdd08703, 32'hbbc71d7e} /* (2, 15, 6) {real, imag} */,
  {32'hbe2d48c2, 32'hbe20cea0} /* (2, 15, 5) {real, imag} */,
  {32'h3e2e0488, 32'h3ddeb526} /* (2, 15, 4) {real, imag} */,
  {32'h3d82965e, 32'h3d126220} /* (2, 15, 3) {real, imag} */,
  {32'hbf4a9112, 32'hbe0a2c30} /* (2, 15, 2) {real, imag} */,
  {32'h3fe1a4cd, 32'h3e8458c8} /* (2, 15, 1) {real, imag} */,
  {32'h3fa1d59d, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'h3ff2d2b1, 32'hbe5e6264} /* (2, 14, 31) {real, imag} */,
  {32'hbf512bce, 32'h3df9f698} /* (2, 14, 30) {real, imag} */,
  {32'h3deb75fd, 32'hbd8a9628} /* (2, 14, 29) {real, imag} */,
  {32'h3e1d2fe8, 32'hbc497b84} /* (2, 14, 28) {real, imag} */,
  {32'hbe7986d4, 32'h3e5d0f53} /* (2, 14, 27) {real, imag} */,
  {32'hbd78cf16, 32'h3af7b2d0} /* (2, 14, 26) {real, imag} */,
  {32'hbd248442, 32'hbd457a22} /* (2, 14, 25) {real, imag} */,
  {32'hbdd9637d, 32'h3ca7d9c4} /* (2, 14, 24) {real, imag} */,
  {32'hbc98b1b3, 32'h3ba3ff5b} /* (2, 14, 23) {real, imag} */,
  {32'hbd1b83e7, 32'hbda8ca14} /* (2, 14, 22) {real, imag} */,
  {32'h3cd6e04a, 32'h3cb8b9de} /* (2, 14, 21) {real, imag} */,
  {32'hbd35e926, 32'hbdec8aac} /* (2, 14, 20) {real, imag} */,
  {32'h3d8c85be, 32'h3d0fc854} /* (2, 14, 19) {real, imag} */,
  {32'hbd77e7c3, 32'hb8f7e100} /* (2, 14, 18) {real, imag} */,
  {32'hbc9670a7, 32'hbcd961ad} /* (2, 14, 17) {real, imag} */,
  {32'hbd0cd594, 32'h00000000} /* (2, 14, 16) {real, imag} */,
  {32'hbc9670a7, 32'h3cd961ad} /* (2, 14, 15) {real, imag} */,
  {32'hbd77e7c3, 32'h38f7e100} /* (2, 14, 14) {real, imag} */,
  {32'h3d8c85be, 32'hbd0fc854} /* (2, 14, 13) {real, imag} */,
  {32'hbd35e926, 32'h3dec8aac} /* (2, 14, 12) {real, imag} */,
  {32'h3cd6e04a, 32'hbcb8b9de} /* (2, 14, 11) {real, imag} */,
  {32'hbd1b83e7, 32'h3da8ca14} /* (2, 14, 10) {real, imag} */,
  {32'hbc98b1b3, 32'hbba3ff5b} /* (2, 14, 9) {real, imag} */,
  {32'hbdd9637d, 32'hbca7d9c4} /* (2, 14, 8) {real, imag} */,
  {32'hbd248442, 32'h3d457a22} /* (2, 14, 7) {real, imag} */,
  {32'hbd78cf16, 32'hbaf7b2d0} /* (2, 14, 6) {real, imag} */,
  {32'hbe7986d4, 32'hbe5d0f53} /* (2, 14, 5) {real, imag} */,
  {32'h3e1d2fe8, 32'h3c497b84} /* (2, 14, 4) {real, imag} */,
  {32'h3deb75fd, 32'h3d8a9628} /* (2, 14, 3) {real, imag} */,
  {32'hbf512bce, 32'hbdf9f698} /* (2, 14, 2) {real, imag} */,
  {32'h3ff2d2b1, 32'h3e5e6264} /* (2, 14, 1) {real, imag} */,
  {32'h3fae4e76, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h3fe99c5f, 32'hbeda7c8a} /* (2, 13, 31) {real, imag} */,
  {32'hbf531050, 32'hbcc0e28c} /* (2, 13, 30) {real, imag} */,
  {32'h3d81a766, 32'hbdceb8db} /* (2, 13, 29) {real, imag} */,
  {32'h3dee80c2, 32'hbe16498a} /* (2, 13, 28) {real, imag} */,
  {32'hbe6e6127, 32'h3d3e2a50} /* (2, 13, 27) {real, imag} */,
  {32'hbc812afc, 32'h3ddf92d8} /* (2, 13, 26) {real, imag} */,
  {32'h3d00e178, 32'h3d403058} /* (2, 13, 25) {real, imag} */,
  {32'hbdb0e4ae, 32'h3d964a28} /* (2, 13, 24) {real, imag} */,
  {32'h3c1c4c28, 32'h3dd2c533} /* (2, 13, 23) {real, imag} */,
  {32'h3d92024f, 32'hbd4c72e1} /* (2, 13, 22) {real, imag} */,
  {32'h3c7a79e0, 32'h3cb82e2c} /* (2, 13, 21) {real, imag} */,
  {32'hbcda4d64, 32'hbcde1671} /* (2, 13, 20) {real, imag} */,
  {32'h3d5bd464, 32'hbb30b6c0} /* (2, 13, 19) {real, imag} */,
  {32'hbdb7e8c8, 32'h3dc69adc} /* (2, 13, 18) {real, imag} */,
  {32'h3ccb9f7e, 32'h3cb3a178} /* (2, 13, 17) {real, imag} */,
  {32'h3d768361, 32'h00000000} /* (2, 13, 16) {real, imag} */,
  {32'h3ccb9f7e, 32'hbcb3a178} /* (2, 13, 15) {real, imag} */,
  {32'hbdb7e8c8, 32'hbdc69adc} /* (2, 13, 14) {real, imag} */,
  {32'h3d5bd464, 32'h3b30b6c0} /* (2, 13, 13) {real, imag} */,
  {32'hbcda4d64, 32'h3cde1671} /* (2, 13, 12) {real, imag} */,
  {32'h3c7a79e0, 32'hbcb82e2c} /* (2, 13, 11) {real, imag} */,
  {32'h3d92024f, 32'h3d4c72e1} /* (2, 13, 10) {real, imag} */,
  {32'h3c1c4c28, 32'hbdd2c533} /* (2, 13, 9) {real, imag} */,
  {32'hbdb0e4ae, 32'hbd964a28} /* (2, 13, 8) {real, imag} */,
  {32'h3d00e178, 32'hbd403058} /* (2, 13, 7) {real, imag} */,
  {32'hbc812afc, 32'hbddf92d8} /* (2, 13, 6) {real, imag} */,
  {32'hbe6e6127, 32'hbd3e2a50} /* (2, 13, 5) {real, imag} */,
  {32'h3dee80c2, 32'h3e16498a} /* (2, 13, 4) {real, imag} */,
  {32'h3d81a766, 32'h3dceb8db} /* (2, 13, 3) {real, imag} */,
  {32'hbf531050, 32'h3cc0e28c} /* (2, 13, 2) {real, imag} */,
  {32'h3fe99c5f, 32'h3eda7c8a} /* (2, 13, 1) {real, imag} */,
  {32'h3facf92f, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'h3fcdae8a, 32'hbea7eb6d} /* (2, 12, 31) {real, imag} */,
  {32'hbf2b54e9, 32'h3db83836} /* (2, 12, 30) {real, imag} */,
  {32'hbbf23490, 32'h3d5b8602} /* (2, 12, 29) {real, imag} */,
  {32'h3e1bfa46, 32'hbdb8d382} /* (2, 12, 28) {real, imag} */,
  {32'hbe283882, 32'h3dae4a65} /* (2, 12, 27) {real, imag} */,
  {32'hbe036fe6, 32'h3e2a967a} /* (2, 12, 26) {real, imag} */,
  {32'h3d0e86f6, 32'h3d853138} /* (2, 12, 25) {real, imag} */,
  {32'h3af78be8, 32'h3d7575dc} /* (2, 12, 24) {real, imag} */,
  {32'h3a76b6e0, 32'hbd5ba55c} /* (2, 12, 23) {real, imag} */,
  {32'h3d0ca32a, 32'hbbaa6ad0} /* (2, 12, 22) {real, imag} */,
  {32'hbda7d089, 32'hbc6fc8b0} /* (2, 12, 21) {real, imag} */,
  {32'h3d5eeca1, 32'hbb0595e8} /* (2, 12, 20) {real, imag} */,
  {32'h3b6eec24, 32'h3da10c64} /* (2, 12, 19) {real, imag} */,
  {32'h3d082289, 32'hbcac26a8} /* (2, 12, 18) {real, imag} */,
  {32'h3cb095c4, 32'hbb9b1552} /* (2, 12, 17) {real, imag} */,
  {32'hbd36878b, 32'h00000000} /* (2, 12, 16) {real, imag} */,
  {32'h3cb095c4, 32'h3b9b1552} /* (2, 12, 15) {real, imag} */,
  {32'h3d082289, 32'h3cac26a8} /* (2, 12, 14) {real, imag} */,
  {32'h3b6eec24, 32'hbda10c64} /* (2, 12, 13) {real, imag} */,
  {32'h3d5eeca1, 32'h3b0595e8} /* (2, 12, 12) {real, imag} */,
  {32'hbda7d089, 32'h3c6fc8b0} /* (2, 12, 11) {real, imag} */,
  {32'h3d0ca32a, 32'h3baa6ad0} /* (2, 12, 10) {real, imag} */,
  {32'h3a76b6e0, 32'h3d5ba55c} /* (2, 12, 9) {real, imag} */,
  {32'h3af78be8, 32'hbd7575dc} /* (2, 12, 8) {real, imag} */,
  {32'h3d0e86f6, 32'hbd853138} /* (2, 12, 7) {real, imag} */,
  {32'hbe036fe6, 32'hbe2a967a} /* (2, 12, 6) {real, imag} */,
  {32'hbe283882, 32'hbdae4a65} /* (2, 12, 5) {real, imag} */,
  {32'h3e1bfa46, 32'h3db8d382} /* (2, 12, 4) {real, imag} */,
  {32'hbbf23490, 32'hbd5b8602} /* (2, 12, 3) {real, imag} */,
  {32'hbf2b54e9, 32'hbdb83836} /* (2, 12, 2) {real, imag} */,
  {32'h3fcdae8a, 32'h3ea7eb6d} /* (2, 12, 1) {real, imag} */,
  {32'h3f886524, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h3f8dec80, 32'hbdadd5b8} /* (2, 11, 31) {real, imag} */,
  {32'hbf015805, 32'h3e1ee94e} /* (2, 11, 30) {real, imag} */,
  {32'hbd5317cf, 32'hbe3708c4} /* (2, 11, 29) {real, imag} */,
  {32'h3e29a35a, 32'hbe019700} /* (2, 11, 28) {real, imag} */,
  {32'hbdd36051, 32'h3daf42f4} /* (2, 11, 27) {real, imag} */,
  {32'hbdd48cfc, 32'h3b7b3a40} /* (2, 11, 26) {real, imag} */,
  {32'h3d659f47, 32'hbd36665b} /* (2, 11, 25) {real, imag} */,
  {32'h3d830c02, 32'h3db76cee} /* (2, 11, 24) {real, imag} */,
  {32'h3db1dd5c, 32'hbc936ceb} /* (2, 11, 23) {real, imag} */,
  {32'h3d8adb62, 32'hbcafdf81} /* (2, 11, 22) {real, imag} */,
  {32'hba475040, 32'h3dc18fbe} /* (2, 11, 21) {real, imag} */,
  {32'hbd9840dd, 32'h3d7dc546} /* (2, 11, 20) {real, imag} */,
  {32'hbc3a8a22, 32'h39b256c0} /* (2, 11, 19) {real, imag} */,
  {32'hbd025356, 32'h3cef0696} /* (2, 11, 18) {real, imag} */,
  {32'h3c28b9a6, 32'hbd319636} /* (2, 11, 17) {real, imag} */,
  {32'hbb6a77b8, 32'h00000000} /* (2, 11, 16) {real, imag} */,
  {32'h3c28b9a6, 32'h3d319636} /* (2, 11, 15) {real, imag} */,
  {32'hbd025356, 32'hbcef0696} /* (2, 11, 14) {real, imag} */,
  {32'hbc3a8a22, 32'hb9b256c0} /* (2, 11, 13) {real, imag} */,
  {32'hbd9840dd, 32'hbd7dc546} /* (2, 11, 12) {real, imag} */,
  {32'hba475040, 32'hbdc18fbe} /* (2, 11, 11) {real, imag} */,
  {32'h3d8adb62, 32'h3cafdf81} /* (2, 11, 10) {real, imag} */,
  {32'h3db1dd5c, 32'h3c936ceb} /* (2, 11, 9) {real, imag} */,
  {32'h3d830c02, 32'hbdb76cee} /* (2, 11, 8) {real, imag} */,
  {32'h3d659f47, 32'h3d36665b} /* (2, 11, 7) {real, imag} */,
  {32'hbdd48cfc, 32'hbb7b3a40} /* (2, 11, 6) {real, imag} */,
  {32'hbdd36051, 32'hbdaf42f4} /* (2, 11, 5) {real, imag} */,
  {32'h3e29a35a, 32'h3e019700} /* (2, 11, 4) {real, imag} */,
  {32'hbd5317cf, 32'h3e3708c4} /* (2, 11, 3) {real, imag} */,
  {32'hbf015805, 32'hbe1ee94e} /* (2, 11, 2) {real, imag} */,
  {32'h3f8dec80, 32'h3dadd5b8} /* (2, 11, 1) {real, imag} */,
  {32'h3f168693, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'hbe95e368, 32'h3c5f29b0} /* (2, 10, 31) {real, imag} */,
  {32'h3c18a5c0, 32'hbdff7c46} /* (2, 10, 30) {real, imag} */,
  {32'hbd70ca44, 32'hbe53a7bd} /* (2, 10, 29) {real, imag} */,
  {32'hbdc8b18a, 32'hbe18d050} /* (2, 10, 28) {real, imag} */,
  {32'hbd805a2f, 32'hbdee5a47} /* (2, 10, 27) {real, imag} */,
  {32'h3be279a8, 32'hbc4d2174} /* (2, 10, 26) {real, imag} */,
  {32'h3d016bae, 32'hbb4d8400} /* (2, 10, 25) {real, imag} */,
  {32'h3c27c400, 32'hbccfae62} /* (2, 10, 24) {real, imag} */,
  {32'hb8f52880, 32'hbe07a7f4} /* (2, 10, 23) {real, imag} */,
  {32'hbd7f6d34, 32'hbb1695e0} /* (2, 10, 22) {real, imag} */,
  {32'h3d196003, 32'h3bb62618} /* (2, 10, 21) {real, imag} */,
  {32'h3b68e380, 32'hbba70800} /* (2, 10, 20) {real, imag} */,
  {32'h3dd20cea, 32'hbd814a7c} /* (2, 10, 19) {real, imag} */,
  {32'h3d2ccaca, 32'hbdd5d1f0} /* (2, 10, 18) {real, imag} */,
  {32'h3d3bc89e, 32'h3b050888} /* (2, 10, 17) {real, imag} */,
  {32'hbd680d88, 32'h00000000} /* (2, 10, 16) {real, imag} */,
  {32'h3d3bc89e, 32'hbb050888} /* (2, 10, 15) {real, imag} */,
  {32'h3d2ccaca, 32'h3dd5d1f0} /* (2, 10, 14) {real, imag} */,
  {32'h3dd20cea, 32'h3d814a7c} /* (2, 10, 13) {real, imag} */,
  {32'h3b68e380, 32'h3ba70800} /* (2, 10, 12) {real, imag} */,
  {32'h3d196003, 32'hbbb62618} /* (2, 10, 11) {real, imag} */,
  {32'hbd7f6d34, 32'h3b1695e0} /* (2, 10, 10) {real, imag} */,
  {32'hb8f52880, 32'h3e07a7f4} /* (2, 10, 9) {real, imag} */,
  {32'h3c27c400, 32'h3ccfae62} /* (2, 10, 8) {real, imag} */,
  {32'h3d016bae, 32'h3b4d8400} /* (2, 10, 7) {real, imag} */,
  {32'h3be279a8, 32'h3c4d2174} /* (2, 10, 6) {real, imag} */,
  {32'hbd805a2f, 32'h3dee5a47} /* (2, 10, 5) {real, imag} */,
  {32'hbdc8b18a, 32'h3e18d050} /* (2, 10, 4) {real, imag} */,
  {32'hbd70ca44, 32'h3e53a7bd} /* (2, 10, 3) {real, imag} */,
  {32'h3c18a5c0, 32'h3dff7c46} /* (2, 10, 2) {real, imag} */,
  {32'hbe95e368, 32'hbc5f29b0} /* (2, 10, 1) {real, imag} */,
  {32'hbe4ff884, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'hbf82dc4e, 32'h3e58bc01} /* (2, 9, 31) {real, imag} */,
  {32'h3eb98166, 32'hbe84c700} /* (2, 9, 30) {real, imag} */,
  {32'h3cd64db4, 32'hbe45f5dd} /* (2, 9, 29) {real, imag} */,
  {32'hbdb5d0f1, 32'hbd61e420} /* (2, 9, 28) {real, imag} */,
  {32'h3ddf47ea, 32'hbce0d7c0} /* (2, 9, 27) {real, imag} */,
  {32'h3c7b74ec, 32'h3d57740e} /* (2, 9, 26) {real, imag} */,
  {32'h3d0c0d7c, 32'h3e1e9eb6} /* (2, 9, 25) {real, imag} */,
  {32'h3e0eaa2f, 32'hbd9f5462} /* (2, 9, 24) {real, imag} */,
  {32'hbd29bc8a, 32'h3dc61285} /* (2, 9, 23) {real, imag} */,
  {32'h3d0dde69, 32'h3d4a39e8} /* (2, 9, 22) {real, imag} */,
  {32'h3d33ad69, 32'h3d1c7ea7} /* (2, 9, 21) {real, imag} */,
  {32'h3bd4b780, 32'hbc958e1f} /* (2, 9, 20) {real, imag} */,
  {32'h3c36e948, 32'h3c3a30e6} /* (2, 9, 19) {real, imag} */,
  {32'h3c4abb2b, 32'hbd4bc524} /* (2, 9, 18) {real, imag} */,
  {32'h3d6e468c, 32'h3c09a49e} /* (2, 9, 17) {real, imag} */,
  {32'hbdea8262, 32'h00000000} /* (2, 9, 16) {real, imag} */,
  {32'h3d6e468c, 32'hbc09a49e} /* (2, 9, 15) {real, imag} */,
  {32'h3c4abb2b, 32'h3d4bc524} /* (2, 9, 14) {real, imag} */,
  {32'h3c36e948, 32'hbc3a30e6} /* (2, 9, 13) {real, imag} */,
  {32'h3bd4b780, 32'h3c958e1f} /* (2, 9, 12) {real, imag} */,
  {32'h3d33ad69, 32'hbd1c7ea7} /* (2, 9, 11) {real, imag} */,
  {32'h3d0dde69, 32'hbd4a39e8} /* (2, 9, 10) {real, imag} */,
  {32'hbd29bc8a, 32'hbdc61285} /* (2, 9, 9) {real, imag} */,
  {32'h3e0eaa2f, 32'h3d9f5462} /* (2, 9, 8) {real, imag} */,
  {32'h3d0c0d7c, 32'hbe1e9eb6} /* (2, 9, 7) {real, imag} */,
  {32'h3c7b74ec, 32'hbd57740e} /* (2, 9, 6) {real, imag} */,
  {32'h3ddf47ea, 32'h3ce0d7c0} /* (2, 9, 5) {real, imag} */,
  {32'hbdb5d0f1, 32'h3d61e420} /* (2, 9, 4) {real, imag} */,
  {32'h3cd64db4, 32'h3e45f5dd} /* (2, 9, 3) {real, imag} */,
  {32'h3eb98166, 32'h3e84c700} /* (2, 9, 2) {real, imag} */,
  {32'hbf82dc4e, 32'hbe58bc01} /* (2, 9, 1) {real, imag} */,
  {32'hbf475199, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'hbfad4633, 32'h3e39539d} /* (2, 8, 31) {real, imag} */,
  {32'h3f3322b0, 32'hbd8393f8} /* (2, 8, 30) {real, imag} */,
  {32'hbd446779, 32'hbd951b40} /* (2, 8, 29) {real, imag} */,
  {32'hbdc800dc, 32'h3d7eba14} /* (2, 8, 28) {real, imag} */,
  {32'h3e592968, 32'hbd839472} /* (2, 8, 27) {real, imag} */,
  {32'h3d9b1451, 32'h3de7552c} /* (2, 8, 26) {real, imag} */,
  {32'hbbc25794, 32'h3e3620a5} /* (2, 8, 25) {real, imag} */,
  {32'h3dbf205e, 32'hbca48a1e} /* (2, 8, 24) {real, imag} */,
  {32'h3d5bf477, 32'h3d9b6259} /* (2, 8, 23) {real, imag} */,
  {32'h3d164847, 32'h3cfbae84} /* (2, 8, 22) {real, imag} */,
  {32'hbd5beb67, 32'hbd402cbc} /* (2, 8, 21) {real, imag} */,
  {32'h3dc2e672, 32'hbc7bbccb} /* (2, 8, 20) {real, imag} */,
  {32'hbcfd875f, 32'hbdb608ac} /* (2, 8, 19) {real, imag} */,
  {32'h3b33da60, 32'h3bc6d334} /* (2, 8, 18) {real, imag} */,
  {32'hbd16ca7e, 32'hbd4d9621} /* (2, 8, 17) {real, imag} */,
  {32'h3c8b86df, 32'h00000000} /* (2, 8, 16) {real, imag} */,
  {32'hbd16ca7e, 32'h3d4d9621} /* (2, 8, 15) {real, imag} */,
  {32'h3b33da60, 32'hbbc6d334} /* (2, 8, 14) {real, imag} */,
  {32'hbcfd875f, 32'h3db608ac} /* (2, 8, 13) {real, imag} */,
  {32'h3dc2e672, 32'h3c7bbccb} /* (2, 8, 12) {real, imag} */,
  {32'hbd5beb67, 32'h3d402cbc} /* (2, 8, 11) {real, imag} */,
  {32'h3d164847, 32'hbcfbae84} /* (2, 8, 10) {real, imag} */,
  {32'h3d5bf477, 32'hbd9b6259} /* (2, 8, 9) {real, imag} */,
  {32'h3dbf205e, 32'h3ca48a1e} /* (2, 8, 8) {real, imag} */,
  {32'hbbc25794, 32'hbe3620a5} /* (2, 8, 7) {real, imag} */,
  {32'h3d9b1451, 32'hbde7552c} /* (2, 8, 6) {real, imag} */,
  {32'h3e592968, 32'h3d839472} /* (2, 8, 5) {real, imag} */,
  {32'hbdc800dc, 32'hbd7eba14} /* (2, 8, 4) {real, imag} */,
  {32'hbd446779, 32'h3d951b40} /* (2, 8, 3) {real, imag} */,
  {32'h3f3322b0, 32'h3d8393f8} /* (2, 8, 2) {real, imag} */,
  {32'hbfad4633, 32'hbe39539d} /* (2, 8, 1) {real, imag} */,
  {32'hbf8991fc, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'hbfc9b112, 32'h3ec83912} /* (2, 7, 31) {real, imag} */,
  {32'h3f4ee35c, 32'hbd406f5a} /* (2, 7, 30) {real, imag} */,
  {32'h3d957f00, 32'hbde54d1f} /* (2, 7, 29) {real, imag} */,
  {32'hbdaef829, 32'hbe201cd4} /* (2, 7, 28) {real, imag} */,
  {32'h3e132b18, 32'h3d2608c8} /* (2, 7, 27) {real, imag} */,
  {32'h3dcb5b98, 32'hbdb65e67} /* (2, 7, 26) {real, imag} */,
  {32'hbd42a644, 32'hbd4ca314} /* (2, 7, 25) {real, imag} */,
  {32'h3d4e2c10, 32'hbdd78940} /* (2, 7, 24) {real, imag} */,
  {32'hbd78e180, 32'hbca93724} /* (2, 7, 23) {real, imag} */,
  {32'hbdc20f31, 32'h3c2ed9e0} /* (2, 7, 22) {real, imag} */,
  {32'h3c06eb24, 32'hbe26eeec} /* (2, 7, 21) {real, imag} */,
  {32'hbe05613b, 32'hbc8a9be3} /* (2, 7, 20) {real, imag} */,
  {32'h3e078fc0, 32'h3ddf9077} /* (2, 7, 19) {real, imag} */,
  {32'h3d00b031, 32'hbd8a5118} /* (2, 7, 18) {real, imag} */,
  {32'h3cb44004, 32'hbc95d424} /* (2, 7, 17) {real, imag} */,
  {32'h3dca90c0, 32'h00000000} /* (2, 7, 16) {real, imag} */,
  {32'h3cb44004, 32'h3c95d424} /* (2, 7, 15) {real, imag} */,
  {32'h3d00b031, 32'h3d8a5118} /* (2, 7, 14) {real, imag} */,
  {32'h3e078fc0, 32'hbddf9077} /* (2, 7, 13) {real, imag} */,
  {32'hbe05613b, 32'h3c8a9be3} /* (2, 7, 12) {real, imag} */,
  {32'h3c06eb24, 32'h3e26eeec} /* (2, 7, 11) {real, imag} */,
  {32'hbdc20f31, 32'hbc2ed9e0} /* (2, 7, 10) {real, imag} */,
  {32'hbd78e180, 32'h3ca93724} /* (2, 7, 9) {real, imag} */,
  {32'h3d4e2c10, 32'h3dd78940} /* (2, 7, 8) {real, imag} */,
  {32'hbd42a644, 32'h3d4ca314} /* (2, 7, 7) {real, imag} */,
  {32'h3dcb5b98, 32'h3db65e67} /* (2, 7, 6) {real, imag} */,
  {32'h3e132b18, 32'hbd2608c8} /* (2, 7, 5) {real, imag} */,
  {32'hbdaef829, 32'h3e201cd4} /* (2, 7, 4) {real, imag} */,
  {32'h3d957f00, 32'h3de54d1f} /* (2, 7, 3) {real, imag} */,
  {32'h3f4ee35c, 32'h3d406f5a} /* (2, 7, 2) {real, imag} */,
  {32'hbfc9b112, 32'hbec83912} /* (2, 7, 1) {real, imag} */,
  {32'hbfa53e92, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'hbfbde0e9, 32'h3f48b732} /* (2, 6, 31) {real, imag} */,
  {32'h3f1ed100, 32'hbdd9a35a} /* (2, 6, 30) {real, imag} */,
  {32'h3e8da6dd, 32'h3d0bc094} /* (2, 6, 29) {real, imag} */,
  {32'hbdeaf458, 32'hbe1895da} /* (2, 6, 28) {real, imag} */,
  {32'h3e03109c, 32'hbde7bb76} /* (2, 6, 27) {real, imag} */,
  {32'h3dd3cdde, 32'h3c44fd18} /* (2, 6, 26) {real, imag} */,
  {32'hbd4697cd, 32'hbaa57800} /* (2, 6, 25) {real, imag} */,
  {32'h3dc50392, 32'hbd1337a0} /* (2, 6, 24) {real, imag} */,
  {32'hbaf75964, 32'h3d408871} /* (2, 6, 23) {real, imag} */,
  {32'h3db59b90, 32'h3bdde648} /* (2, 6, 22) {real, imag} */,
  {32'h3c986186, 32'hbd110d7d} /* (2, 6, 21) {real, imag} */,
  {32'hbd70362a, 32'h3d958b68} /* (2, 6, 20) {real, imag} */,
  {32'hbcd8a489, 32'hbd0e5495} /* (2, 6, 19) {real, imag} */,
  {32'h3cc7127f, 32'h3d021b54} /* (2, 6, 18) {real, imag} */,
  {32'hbd9c895a, 32'hbc714992} /* (2, 6, 17) {real, imag} */,
  {32'h3d3f49b4, 32'h00000000} /* (2, 6, 16) {real, imag} */,
  {32'hbd9c895a, 32'h3c714992} /* (2, 6, 15) {real, imag} */,
  {32'h3cc7127f, 32'hbd021b54} /* (2, 6, 14) {real, imag} */,
  {32'hbcd8a489, 32'h3d0e5495} /* (2, 6, 13) {real, imag} */,
  {32'hbd70362a, 32'hbd958b68} /* (2, 6, 12) {real, imag} */,
  {32'h3c986186, 32'h3d110d7d} /* (2, 6, 11) {real, imag} */,
  {32'h3db59b90, 32'hbbdde648} /* (2, 6, 10) {real, imag} */,
  {32'hbaf75964, 32'hbd408871} /* (2, 6, 9) {real, imag} */,
  {32'h3dc50392, 32'h3d1337a0} /* (2, 6, 8) {real, imag} */,
  {32'hbd4697cd, 32'h3aa57800} /* (2, 6, 7) {real, imag} */,
  {32'h3dd3cdde, 32'hbc44fd18} /* (2, 6, 6) {real, imag} */,
  {32'h3e03109c, 32'h3de7bb76} /* (2, 6, 5) {real, imag} */,
  {32'hbdeaf458, 32'h3e1895da} /* (2, 6, 4) {real, imag} */,
  {32'h3e8da6dd, 32'hbd0bc094} /* (2, 6, 3) {real, imag} */,
  {32'h3f1ed100, 32'h3dd9a35a} /* (2, 6, 2) {real, imag} */,
  {32'hbfbde0e9, 32'hbf48b732} /* (2, 6, 1) {real, imag} */,
  {32'hbf8b89d4, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hbf967b12, 32'h3f95996f} /* (2, 5, 31) {real, imag} */,
  {32'h3e0d7946, 32'hbe889242} /* (2, 5, 30) {real, imag} */,
  {32'h3eae0444, 32'hbc66e338} /* (2, 5, 29) {real, imag} */,
  {32'hbe336e5c, 32'hbde7ccb8} /* (2, 5, 28) {real, imag} */,
  {32'h3e04c706, 32'hbac75100} /* (2, 5, 27) {real, imag} */,
  {32'hbc65add6, 32'h3dfa1aa2} /* (2, 5, 26) {real, imag} */,
  {32'hbda236b2, 32'h3c9fa9e5} /* (2, 5, 25) {real, imag} */,
  {32'h3cbbea28, 32'h3d455210} /* (2, 5, 24) {real, imag} */,
  {32'hbd16a4ea, 32'h3d90a478} /* (2, 5, 23) {real, imag} */,
  {32'hbd3f53c2, 32'hbd2c6360} /* (2, 5, 22) {real, imag} */,
  {32'h3dbc3cf3, 32'hb95baa00} /* (2, 5, 21) {real, imag} */,
  {32'hba077fc0, 32'hbcf89724} /* (2, 5, 20) {real, imag} */,
  {32'h3d0cb5da, 32'h3c69d941} /* (2, 5, 19) {real, imag} */,
  {32'hbd8e31fb, 32'h3d70f648} /* (2, 5, 18) {real, imag} */,
  {32'h3daf75aa, 32'h3d14f5a2} /* (2, 5, 17) {real, imag} */,
  {32'hbd317fcf, 32'h00000000} /* (2, 5, 16) {real, imag} */,
  {32'h3daf75aa, 32'hbd14f5a2} /* (2, 5, 15) {real, imag} */,
  {32'hbd8e31fb, 32'hbd70f648} /* (2, 5, 14) {real, imag} */,
  {32'h3d0cb5da, 32'hbc69d941} /* (2, 5, 13) {real, imag} */,
  {32'hba077fc0, 32'h3cf89724} /* (2, 5, 12) {real, imag} */,
  {32'h3dbc3cf3, 32'h395baa00} /* (2, 5, 11) {real, imag} */,
  {32'hbd3f53c2, 32'h3d2c6360} /* (2, 5, 10) {real, imag} */,
  {32'hbd16a4ea, 32'hbd90a478} /* (2, 5, 9) {real, imag} */,
  {32'h3cbbea28, 32'hbd455210} /* (2, 5, 8) {real, imag} */,
  {32'hbda236b2, 32'hbc9fa9e5} /* (2, 5, 7) {real, imag} */,
  {32'hbc65add6, 32'hbdfa1aa2} /* (2, 5, 6) {real, imag} */,
  {32'h3e04c706, 32'h3ac75100} /* (2, 5, 5) {real, imag} */,
  {32'hbe336e5c, 32'h3de7ccb8} /* (2, 5, 4) {real, imag} */,
  {32'h3eae0444, 32'h3c66e338} /* (2, 5, 3) {real, imag} */,
  {32'h3e0d7946, 32'h3e889242} /* (2, 5, 2) {real, imag} */,
  {32'hbf967b12, 32'hbf95996f} /* (2, 5, 1) {real, imag} */,
  {32'hbf8444f0, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hbf7d6f5e, 32'h3fde33f6} /* (2, 4, 31) {real, imag} */,
  {32'hbe8d8048, 32'hbe92136b} /* (2, 4, 30) {real, imag} */,
  {32'h3e66ec8c, 32'hbbae3ba0} /* (2, 4, 29) {real, imag} */,
  {32'hbcf193e8, 32'hbe0f416a} /* (2, 4, 28) {real, imag} */,
  {32'h3d88ff70, 32'h3d998269} /* (2, 4, 27) {real, imag} */,
  {32'h3becaa7c, 32'h3dc2e23d} /* (2, 4, 26) {real, imag} */,
  {32'h3e28ab32, 32'h3ddb92be} /* (2, 4, 25) {real, imag} */,
  {32'hbc270918, 32'hbdb46aea} /* (2, 4, 24) {real, imag} */,
  {32'h3dc7cecc, 32'hbbacfdc0} /* (2, 4, 23) {real, imag} */,
  {32'h3bef9b36, 32'hbe0a073e} /* (2, 4, 22) {real, imag} */,
  {32'hbba1d4d8, 32'hbca66b48} /* (2, 4, 21) {real, imag} */,
  {32'hbda5846f, 32'hbd0d6961} /* (2, 4, 20) {real, imag} */,
  {32'h3d951d84, 32'hbc063f3c} /* (2, 4, 19) {real, imag} */,
  {32'hbd6b9f2c, 32'h3d104d89} /* (2, 4, 18) {real, imag} */,
  {32'h3da1af84, 32'hbd2e9e62} /* (2, 4, 17) {real, imag} */,
  {32'hbd84d047, 32'h00000000} /* (2, 4, 16) {real, imag} */,
  {32'h3da1af84, 32'h3d2e9e62} /* (2, 4, 15) {real, imag} */,
  {32'hbd6b9f2c, 32'hbd104d89} /* (2, 4, 14) {real, imag} */,
  {32'h3d951d84, 32'h3c063f3c} /* (2, 4, 13) {real, imag} */,
  {32'hbda5846f, 32'h3d0d6961} /* (2, 4, 12) {real, imag} */,
  {32'hbba1d4d8, 32'h3ca66b48} /* (2, 4, 11) {real, imag} */,
  {32'h3bef9b36, 32'h3e0a073e} /* (2, 4, 10) {real, imag} */,
  {32'h3dc7cecc, 32'h3bacfdc0} /* (2, 4, 9) {real, imag} */,
  {32'hbc270918, 32'h3db46aea} /* (2, 4, 8) {real, imag} */,
  {32'h3e28ab32, 32'hbddb92be} /* (2, 4, 7) {real, imag} */,
  {32'h3becaa7c, 32'hbdc2e23d} /* (2, 4, 6) {real, imag} */,
  {32'h3d88ff70, 32'hbd998269} /* (2, 4, 5) {real, imag} */,
  {32'hbcf193e8, 32'h3e0f416a} /* (2, 4, 4) {real, imag} */,
  {32'h3e66ec8c, 32'h3bae3ba0} /* (2, 4, 3) {real, imag} */,
  {32'hbe8d8048, 32'h3e92136b} /* (2, 4, 2) {real, imag} */,
  {32'hbf7d6f5e, 32'hbfde33f6} /* (2, 4, 1) {real, imag} */,
  {32'hbf8cc5ce, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hbf636f08, 32'h3fd837eb} /* (2, 3, 31) {real, imag} */,
  {32'hbed108c1, 32'hbef695c7} /* (2, 3, 30) {real, imag} */,
  {32'h3e82edaa, 32'h3cd4eac8} /* (2, 3, 29) {real, imag} */,
  {32'h3c8b6622, 32'hbe3b67b8} /* (2, 3, 28) {real, imag} */,
  {32'h3e30cd5e, 32'h3d8b2652} /* (2, 3, 27) {real, imag} */,
  {32'h3d2ecfda, 32'h3dcf0082} /* (2, 3, 26) {real, imag} */,
  {32'h3d826ba0, 32'h3d9035cc} /* (2, 3, 25) {real, imag} */,
  {32'hbd0d996a, 32'hbd45736c} /* (2, 3, 24) {real, imag} */,
  {32'h3e456ca4, 32'hbd329082} /* (2, 3, 23) {real, imag} */,
  {32'hbc797aa0, 32'hbcfc59f1} /* (2, 3, 22) {real, imag} */,
  {32'h3d6960da, 32'hbbf32fd0} /* (2, 3, 21) {real, imag} */,
  {32'hbd02bda0, 32'hbd2f9a90} /* (2, 3, 20) {real, imag} */,
  {32'hbd6dec4c, 32'h3c44c840} /* (2, 3, 19) {real, imag} */,
  {32'hbbc7e1d0, 32'hbd9f0d7a} /* (2, 3, 18) {real, imag} */,
  {32'hbb503150, 32'hbc934032} /* (2, 3, 17) {real, imag} */,
  {32'h3d6abc02, 32'h00000000} /* (2, 3, 16) {real, imag} */,
  {32'hbb503150, 32'h3c934032} /* (2, 3, 15) {real, imag} */,
  {32'hbbc7e1d0, 32'h3d9f0d7a} /* (2, 3, 14) {real, imag} */,
  {32'hbd6dec4c, 32'hbc44c840} /* (2, 3, 13) {real, imag} */,
  {32'hbd02bda0, 32'h3d2f9a90} /* (2, 3, 12) {real, imag} */,
  {32'h3d6960da, 32'h3bf32fd0} /* (2, 3, 11) {real, imag} */,
  {32'hbc797aa0, 32'h3cfc59f1} /* (2, 3, 10) {real, imag} */,
  {32'h3e456ca4, 32'h3d329082} /* (2, 3, 9) {real, imag} */,
  {32'hbd0d996a, 32'h3d45736c} /* (2, 3, 8) {real, imag} */,
  {32'h3d826ba0, 32'hbd9035cc} /* (2, 3, 7) {real, imag} */,
  {32'h3d2ecfda, 32'hbdcf0082} /* (2, 3, 6) {real, imag} */,
  {32'h3e30cd5e, 32'hbd8b2652} /* (2, 3, 5) {real, imag} */,
  {32'h3c8b6622, 32'h3e3b67b8} /* (2, 3, 4) {real, imag} */,
  {32'h3e82edaa, 32'hbcd4eac8} /* (2, 3, 3) {real, imag} */,
  {32'hbed108c1, 32'h3ef695c7} /* (2, 3, 2) {real, imag} */,
  {32'hbf636f08, 32'hbfd837eb} /* (2, 3, 1) {real, imag} */,
  {32'hbf701ed4, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hbf5ea864, 32'h3fcedacb} /* (2, 2, 31) {real, imag} */,
  {32'hbee1d8c7, 32'hbf4dd26a} /* (2, 2, 30) {real, imag} */,
  {32'h3e5e7844, 32'h3d920072} /* (2, 2, 29) {real, imag} */,
  {32'h3e3f1150, 32'hbea26c70} /* (2, 2, 28) {real, imag} */,
  {32'h3da7fe43, 32'h3d79c092} /* (2, 2, 27) {real, imag} */,
  {32'h3d46656c, 32'h3d533ba4} /* (2, 2, 26) {real, imag} */,
  {32'h3d66b8c6, 32'hbb8eb698} /* (2, 2, 25) {real, imag} */,
  {32'hbd814da1, 32'hbdf3a16e} /* (2, 2, 24) {real, imag} */,
  {32'hbca2fff3, 32'h3c4bf4fd} /* (2, 2, 23) {real, imag} */,
  {32'hbc9289bf, 32'hbd849128} /* (2, 2, 22) {real, imag} */,
  {32'h3c7d6360, 32'hbc8d3c0e} /* (2, 2, 21) {real, imag} */,
  {32'h3c96ddf2, 32'hbcf3ecbb} /* (2, 2, 20) {real, imag} */,
  {32'hbd8fa238, 32'hbd19fc5a} /* (2, 2, 19) {real, imag} */,
  {32'h3d583145, 32'hbdf017a1} /* (2, 2, 18) {real, imag} */,
  {32'h3ddef736, 32'h3d459416} /* (2, 2, 17) {real, imag} */,
  {32'h3ce77754, 32'h00000000} /* (2, 2, 16) {real, imag} */,
  {32'h3ddef736, 32'hbd459416} /* (2, 2, 15) {real, imag} */,
  {32'h3d583145, 32'h3df017a1} /* (2, 2, 14) {real, imag} */,
  {32'hbd8fa238, 32'h3d19fc5a} /* (2, 2, 13) {real, imag} */,
  {32'h3c96ddf2, 32'h3cf3ecbb} /* (2, 2, 12) {real, imag} */,
  {32'h3c7d6360, 32'h3c8d3c0e} /* (2, 2, 11) {real, imag} */,
  {32'hbc9289bf, 32'h3d849128} /* (2, 2, 10) {real, imag} */,
  {32'hbca2fff3, 32'hbc4bf4fd} /* (2, 2, 9) {real, imag} */,
  {32'hbd814da1, 32'h3df3a16e} /* (2, 2, 8) {real, imag} */,
  {32'h3d66b8c6, 32'h3b8eb698} /* (2, 2, 7) {real, imag} */,
  {32'h3d46656c, 32'hbd533ba4} /* (2, 2, 6) {real, imag} */,
  {32'h3da7fe43, 32'hbd79c092} /* (2, 2, 5) {real, imag} */,
  {32'h3e3f1150, 32'h3ea26c70} /* (2, 2, 4) {real, imag} */,
  {32'h3e5e7844, 32'hbd920072} /* (2, 2, 3) {real, imag} */,
  {32'hbee1d8c7, 32'h3f4dd26a} /* (2, 2, 2) {real, imag} */,
  {32'hbf5ea864, 32'hbfcedacb} /* (2, 2, 1) {real, imag} */,
  {32'hbf65f67e, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hbf6c95e2, 32'h3fb469fc} /* (2, 1, 31) {real, imag} */,
  {32'hbeb017a3, 32'hbf2c29d0} /* (2, 1, 30) {real, imag} */,
  {32'h3dffe39e, 32'hbae6d810} /* (2, 1, 29) {real, imag} */,
  {32'h3d74f81c, 32'hbe985e8c} /* (2, 1, 28) {real, imag} */,
  {32'h3d89e2be, 32'h3dba21c8} /* (2, 1, 27) {real, imag} */,
  {32'h3ccceed7, 32'h3d96314e} /* (2, 1, 26) {real, imag} */,
  {32'hbd79db1b, 32'h3dbe54a8} /* (2, 1, 25) {real, imag} */,
  {32'hbd7a6246, 32'h3b4bd660} /* (2, 1, 24) {real, imag} */,
  {32'hbda7bb42, 32'hbe0450ae} /* (2, 1, 23) {real, imag} */,
  {32'h3cb718c5, 32'hbe032ea4} /* (2, 1, 22) {real, imag} */,
  {32'h3e0558db, 32'hbc569338} /* (2, 1, 21) {real, imag} */,
  {32'h3d2be5c8, 32'h3d13b4d6} /* (2, 1, 20) {real, imag} */,
  {32'h3bdd7180, 32'hbc84a6bd} /* (2, 1, 19) {real, imag} */,
  {32'hbc0a90a6, 32'hba9b12d0} /* (2, 1, 18) {real, imag} */,
  {32'h3cfa81a0, 32'hbd22dd12} /* (2, 1, 17) {real, imag} */,
  {32'hbd892994, 32'h00000000} /* (2, 1, 16) {real, imag} */,
  {32'h3cfa81a0, 32'h3d22dd12} /* (2, 1, 15) {real, imag} */,
  {32'hbc0a90a6, 32'h3a9b12d0} /* (2, 1, 14) {real, imag} */,
  {32'h3bdd7180, 32'h3c84a6bd} /* (2, 1, 13) {real, imag} */,
  {32'h3d2be5c8, 32'hbd13b4d6} /* (2, 1, 12) {real, imag} */,
  {32'h3e0558db, 32'h3c569338} /* (2, 1, 11) {real, imag} */,
  {32'h3cb718c5, 32'h3e032ea4} /* (2, 1, 10) {real, imag} */,
  {32'hbda7bb42, 32'h3e0450ae} /* (2, 1, 9) {real, imag} */,
  {32'hbd7a6246, 32'hbb4bd660} /* (2, 1, 8) {real, imag} */,
  {32'hbd79db1b, 32'hbdbe54a8} /* (2, 1, 7) {real, imag} */,
  {32'h3ccceed7, 32'hbd96314e} /* (2, 1, 6) {real, imag} */,
  {32'h3d89e2be, 32'hbdba21c8} /* (2, 1, 5) {real, imag} */,
  {32'h3d74f81c, 32'h3e985e8c} /* (2, 1, 4) {real, imag} */,
  {32'h3dffe39e, 32'h3ae6d810} /* (2, 1, 3) {real, imag} */,
  {32'hbeb017a3, 32'h3f2c29d0} /* (2, 1, 2) {real, imag} */,
  {32'hbf6c95e2, 32'hbfb469fc} /* (2, 1, 1) {real, imag} */,
  {32'hbedd49b2, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hbf5a1c5c, 32'h3f72038b} /* (2, 0, 31) {real, imag} */,
  {32'hbdb71410, 32'hbee25ce0} /* (2, 0, 30) {real, imag} */,
  {32'h3cb118e2, 32'hbd93e7c7} /* (2, 0, 29) {real, imag} */,
  {32'hbcfdd1c8, 32'hbe3a9b03} /* (2, 0, 28) {real, imag} */,
  {32'h3e26e388, 32'h3cc92c64} /* (2, 0, 27) {real, imag} */,
  {32'h3d8939a1, 32'h3cae8e92} /* (2, 0, 26) {real, imag} */,
  {32'hbdf9432a, 32'h3d751f2d} /* (2, 0, 25) {real, imag} */,
  {32'hbd950453, 32'h3d1fd9ae} /* (2, 0, 24) {real, imag} */,
  {32'hbcecb9c5, 32'hbde869fd} /* (2, 0, 23) {real, imag} */,
  {32'h3dc0a5a0, 32'hbdd814ad} /* (2, 0, 22) {real, imag} */,
  {32'h3d464faa, 32'h3dade000} /* (2, 0, 21) {real, imag} */,
  {32'h3cef2a66, 32'h3d2e2ebd} /* (2, 0, 20) {real, imag} */,
  {32'hbd090fb6, 32'hbaa55dd0} /* (2, 0, 19) {real, imag} */,
  {32'hbd84a8c1, 32'h3bab6200} /* (2, 0, 18) {real, imag} */,
  {32'hbc340cbb, 32'hbd317a3c} /* (2, 0, 17) {real, imag} */,
  {32'hbbef11cc, 32'h00000000} /* (2, 0, 16) {real, imag} */,
  {32'hbc340cbb, 32'h3d317a3c} /* (2, 0, 15) {real, imag} */,
  {32'hbd84a8c1, 32'hbbab6200} /* (2, 0, 14) {real, imag} */,
  {32'hbd090fb6, 32'h3aa55dd0} /* (2, 0, 13) {real, imag} */,
  {32'h3cef2a66, 32'hbd2e2ebd} /* (2, 0, 12) {real, imag} */,
  {32'h3d464faa, 32'hbdade000} /* (2, 0, 11) {real, imag} */,
  {32'h3dc0a5a0, 32'h3dd814ad} /* (2, 0, 10) {real, imag} */,
  {32'hbcecb9c5, 32'h3de869fd} /* (2, 0, 9) {real, imag} */,
  {32'hbd950453, 32'hbd1fd9ae} /* (2, 0, 8) {real, imag} */,
  {32'hbdf9432a, 32'hbd751f2d} /* (2, 0, 7) {real, imag} */,
  {32'h3d8939a1, 32'hbcae8e92} /* (2, 0, 6) {real, imag} */,
  {32'h3e26e388, 32'hbcc92c64} /* (2, 0, 5) {real, imag} */,
  {32'hbcfdd1c8, 32'h3e3a9b03} /* (2, 0, 4) {real, imag} */,
  {32'h3cb118e2, 32'h3d93e7c7} /* (2, 0, 3) {real, imag} */,
  {32'hbdb71410, 32'h3ee25ce0} /* (2, 0, 2) {real, imag} */,
  {32'hbf5a1c5c, 32'hbf72038b} /* (2, 0, 1) {real, imag} */,
  {32'hbea3cf8f, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hbf68585e, 32'h3ee20071} /* (1, 31, 31) {real, imag} */,
  {32'h3ea47fec, 32'hbe62088f} /* (1, 31, 30) {real, imag} */,
  {32'h3d809d40, 32'h3d0475b4} /* (1, 31, 29) {real, imag} */,
  {32'h3aef6d30, 32'h3cdaa6f0} /* (1, 31, 28) {real, imag} */,
  {32'h3e36690d, 32'hbce211fc} /* (1, 31, 27) {real, imag} */,
  {32'hbd2b61bc, 32'hbd94faf0} /* (1, 31, 26) {real, imag} */,
  {32'hbcaf03a8, 32'h3cc2b31e} /* (1, 31, 25) {real, imag} */,
  {32'hbd17d5b5, 32'hbdc3610a} /* (1, 31, 24) {real, imag} */,
  {32'h3c8ac1bc, 32'h3d3a61c4} /* (1, 31, 23) {real, imag} */,
  {32'h3d46d4fa, 32'hbcb6db9a} /* (1, 31, 22) {real, imag} */,
  {32'h3da540f6, 32'hbcf2893c} /* (1, 31, 21) {real, imag} */,
  {32'h3d1e530a, 32'h3c9a655f} /* (1, 31, 20) {real, imag} */,
  {32'hbd0cbab5, 32'h3ccbd0f0} /* (1, 31, 19) {real, imag} */,
  {32'h3ca3a20e, 32'hbd509d42} /* (1, 31, 18) {real, imag} */,
  {32'hbd083fa9, 32'hbcc6743c} /* (1, 31, 17) {real, imag} */,
  {32'hbaf24f00, 32'h00000000} /* (1, 31, 16) {real, imag} */,
  {32'hbd083fa9, 32'h3cc6743c} /* (1, 31, 15) {real, imag} */,
  {32'h3ca3a20e, 32'h3d509d42} /* (1, 31, 14) {real, imag} */,
  {32'hbd0cbab5, 32'hbccbd0f0} /* (1, 31, 13) {real, imag} */,
  {32'h3d1e530a, 32'hbc9a655f} /* (1, 31, 12) {real, imag} */,
  {32'h3da540f6, 32'h3cf2893c} /* (1, 31, 11) {real, imag} */,
  {32'h3d46d4fa, 32'h3cb6db9a} /* (1, 31, 10) {real, imag} */,
  {32'h3c8ac1bc, 32'hbd3a61c4} /* (1, 31, 9) {real, imag} */,
  {32'hbd17d5b5, 32'h3dc3610a} /* (1, 31, 8) {real, imag} */,
  {32'hbcaf03a8, 32'hbcc2b31e} /* (1, 31, 7) {real, imag} */,
  {32'hbd2b61bc, 32'h3d94faf0} /* (1, 31, 6) {real, imag} */,
  {32'h3e36690d, 32'h3ce211fc} /* (1, 31, 5) {real, imag} */,
  {32'h3aef6d30, 32'hbcdaa6f0} /* (1, 31, 4) {real, imag} */,
  {32'h3d809d40, 32'hbd0475b4} /* (1, 31, 3) {real, imag} */,
  {32'h3ea47fec, 32'h3e62088f} /* (1, 31, 2) {real, imag} */,
  {32'hbf68585e, 32'hbee20071} /* (1, 31, 1) {real, imag} */,
  {32'hbf028506, 32'h00000000} /* (1, 31, 0) {real, imag} */,
  {32'hbf93059a, 32'h3e4b15b0} /* (1, 30, 31) {real, imag} */,
  {32'h3f16f75b, 32'hbe551c14} /* (1, 30, 30) {real, imag} */,
  {32'h3ddd1033, 32'hbb395d20} /* (1, 30, 29) {real, imag} */,
  {32'h3d576eca, 32'h3d780570} /* (1, 30, 28) {real, imag} */,
  {32'h3e020744, 32'hbe02f2ad} /* (1, 30, 27) {real, imag} */,
  {32'h3cfaee26, 32'hbdfc2341} /* (1, 30, 26) {real, imag} */,
  {32'hbe053feb, 32'h3da555b8} /* (1, 30, 25) {real, imag} */,
  {32'h3ce2668c, 32'hbd4bd587} /* (1, 30, 24) {real, imag} */,
  {32'hbda260db, 32'h3d9de8b1} /* (1, 30, 23) {real, imag} */,
  {32'hbd8550d2, 32'h3e15b2b8} /* (1, 30, 22) {real, imag} */,
  {32'h3bd0a060, 32'hbcacb2ae} /* (1, 30, 21) {real, imag} */,
  {32'h3c55d47c, 32'hbce6d732} /* (1, 30, 20) {real, imag} */,
  {32'h3b6378e8, 32'h3d06797a} /* (1, 30, 19) {real, imag} */,
  {32'hbbe24ce8, 32'hbd96b4cb} /* (1, 30, 18) {real, imag} */,
  {32'hbd97c4a2, 32'h3c3449ac} /* (1, 30, 17) {real, imag} */,
  {32'h3cc59562, 32'h00000000} /* (1, 30, 16) {real, imag} */,
  {32'hbd97c4a2, 32'hbc3449ac} /* (1, 30, 15) {real, imag} */,
  {32'hbbe24ce8, 32'h3d96b4cb} /* (1, 30, 14) {real, imag} */,
  {32'h3b6378e8, 32'hbd06797a} /* (1, 30, 13) {real, imag} */,
  {32'h3c55d47c, 32'h3ce6d732} /* (1, 30, 12) {real, imag} */,
  {32'h3bd0a060, 32'h3cacb2ae} /* (1, 30, 11) {real, imag} */,
  {32'hbd8550d2, 32'hbe15b2b8} /* (1, 30, 10) {real, imag} */,
  {32'hbda260db, 32'hbd9de8b1} /* (1, 30, 9) {real, imag} */,
  {32'h3ce2668c, 32'h3d4bd587} /* (1, 30, 8) {real, imag} */,
  {32'hbe053feb, 32'hbda555b8} /* (1, 30, 7) {real, imag} */,
  {32'h3cfaee26, 32'h3dfc2341} /* (1, 30, 6) {real, imag} */,
  {32'h3e020744, 32'h3e02f2ad} /* (1, 30, 5) {real, imag} */,
  {32'h3d576eca, 32'hbd780570} /* (1, 30, 4) {real, imag} */,
  {32'h3ddd1033, 32'h3b395d20} /* (1, 30, 3) {real, imag} */,
  {32'h3f16f75b, 32'h3e551c14} /* (1, 30, 2) {real, imag} */,
  {32'hbf93059a, 32'hbe4b15b0} /* (1, 30, 1) {real, imag} */,
  {32'hbf23405f, 32'h00000000} /* (1, 30, 0) {real, imag} */,
  {32'hbfb50e2b, 32'h3cd0f5c0} /* (1, 29, 31) {real, imag} */,
  {32'h3f3f7aa2, 32'hbe62fb75} /* (1, 29, 30) {real, imag} */,
  {32'h3d13721e, 32'hbd4538d7} /* (1, 29, 29) {real, imag} */,
  {32'h3baa29d0, 32'h3d83b664} /* (1, 29, 28) {real, imag} */,
  {32'h3e98464e, 32'hbc9b2a80} /* (1, 29, 27) {real, imag} */,
  {32'h3c83d7ee, 32'h3c366bfa} /* (1, 29, 26) {real, imag} */,
  {32'hbdf582ae, 32'h3dac1a8a} /* (1, 29, 25) {real, imag} */,
  {32'h3cd2dc94, 32'hbd7eb8bb} /* (1, 29, 24) {real, imag} */,
  {32'hbc5d2f18, 32'hbdc029de} /* (1, 29, 23) {real, imag} */,
  {32'hbd8d7e25, 32'h3d4d537e} /* (1, 29, 22) {real, imag} */,
  {32'h3d3dd078, 32'hbc8391d0} /* (1, 29, 21) {real, imag} */,
  {32'h3cafd642, 32'h3d243957} /* (1, 29, 20) {real, imag} */,
  {32'h3ba9be20, 32'h3b8ccc36} /* (1, 29, 19) {real, imag} */,
  {32'h3c99b69e, 32'h3c72eea8} /* (1, 29, 18) {real, imag} */,
  {32'hbb94a55a, 32'h3c91cad6} /* (1, 29, 17) {real, imag} */,
  {32'hbc042fcc, 32'h00000000} /* (1, 29, 16) {real, imag} */,
  {32'hbb94a55a, 32'hbc91cad6} /* (1, 29, 15) {real, imag} */,
  {32'h3c99b69e, 32'hbc72eea8} /* (1, 29, 14) {real, imag} */,
  {32'h3ba9be20, 32'hbb8ccc36} /* (1, 29, 13) {real, imag} */,
  {32'h3cafd642, 32'hbd243957} /* (1, 29, 12) {real, imag} */,
  {32'h3d3dd078, 32'h3c8391d0} /* (1, 29, 11) {real, imag} */,
  {32'hbd8d7e25, 32'hbd4d537e} /* (1, 29, 10) {real, imag} */,
  {32'hbc5d2f18, 32'h3dc029de} /* (1, 29, 9) {real, imag} */,
  {32'h3cd2dc94, 32'h3d7eb8bb} /* (1, 29, 8) {real, imag} */,
  {32'hbdf582ae, 32'hbdac1a8a} /* (1, 29, 7) {real, imag} */,
  {32'h3c83d7ee, 32'hbc366bfa} /* (1, 29, 6) {real, imag} */,
  {32'h3e98464e, 32'h3c9b2a80} /* (1, 29, 5) {real, imag} */,
  {32'h3baa29d0, 32'hbd83b664} /* (1, 29, 4) {real, imag} */,
  {32'h3d13721e, 32'h3d4538d7} /* (1, 29, 3) {real, imag} */,
  {32'h3f3f7aa2, 32'h3e62fb75} /* (1, 29, 2) {real, imag} */,
  {32'hbfb50e2b, 32'hbcd0f5c0} /* (1, 29, 1) {real, imag} */,
  {32'hbf49ea6b, 32'h00000000} /* (1, 29, 0) {real, imag} */,
  {32'hbfc40ace, 32'h3e102880} /* (1, 28, 31) {real, imag} */,
  {32'h3f3be20a, 32'hbd11c0b8} /* (1, 28, 30) {real, imag} */,
  {32'h3cfb73d0, 32'hbd44409c} /* (1, 28, 29) {real, imag} */,
  {32'hbe362b3b, 32'h3e16165d} /* (1, 28, 28) {real, imag} */,
  {32'h3e6754ad, 32'hbd782426} /* (1, 28, 27) {real, imag} */,
  {32'hbce9af26, 32'h3d2443bb} /* (1, 28, 26) {real, imag} */,
  {32'h3b9a8b30, 32'h3d7ead96} /* (1, 28, 25) {real, imag} */,
  {32'h3df2bc74, 32'hbdbe18ac} /* (1, 28, 24) {real, imag} */,
  {32'hbdbc4a2e, 32'hbccc6208} /* (1, 28, 23) {real, imag} */,
  {32'hbd3c033a, 32'hbdb99ea0} /* (1, 28, 22) {real, imag} */,
  {32'hbcb23e6e, 32'hbd82b69d} /* (1, 28, 21) {real, imag} */,
  {32'hbc37cefa, 32'h3d9a552a} /* (1, 28, 20) {real, imag} */,
  {32'hbcdee6a0, 32'h3cad4061} /* (1, 28, 19) {real, imag} */,
  {32'hbc52bee8, 32'hbbff6864} /* (1, 28, 18) {real, imag} */,
  {32'h3c7621d4, 32'hbc923df5} /* (1, 28, 17) {real, imag} */,
  {32'h3b66f6e8, 32'h00000000} /* (1, 28, 16) {real, imag} */,
  {32'h3c7621d4, 32'h3c923df5} /* (1, 28, 15) {real, imag} */,
  {32'hbc52bee8, 32'h3bff6864} /* (1, 28, 14) {real, imag} */,
  {32'hbcdee6a0, 32'hbcad4061} /* (1, 28, 13) {real, imag} */,
  {32'hbc37cefa, 32'hbd9a552a} /* (1, 28, 12) {real, imag} */,
  {32'hbcb23e6e, 32'h3d82b69d} /* (1, 28, 11) {real, imag} */,
  {32'hbd3c033a, 32'h3db99ea0} /* (1, 28, 10) {real, imag} */,
  {32'hbdbc4a2e, 32'h3ccc6208} /* (1, 28, 9) {real, imag} */,
  {32'h3df2bc74, 32'h3dbe18ac} /* (1, 28, 8) {real, imag} */,
  {32'h3b9a8b30, 32'hbd7ead96} /* (1, 28, 7) {real, imag} */,
  {32'hbce9af26, 32'hbd2443bb} /* (1, 28, 6) {real, imag} */,
  {32'h3e6754ad, 32'h3d782426} /* (1, 28, 5) {real, imag} */,
  {32'hbe362b3b, 32'hbe16165d} /* (1, 28, 4) {real, imag} */,
  {32'h3cfb73d0, 32'h3d44409c} /* (1, 28, 3) {real, imag} */,
  {32'h3f3be20a, 32'h3d11c0b8} /* (1, 28, 2) {real, imag} */,
  {32'hbfc40ace, 32'hbe102880} /* (1, 28, 1) {real, imag} */,
  {32'hbf460cd1, 32'h00000000} /* (1, 28, 0) {real, imag} */,
  {32'hbfd559aa, 32'h3e01d9cc} /* (1, 27, 31) {real, imag} */,
  {32'h3f27b2bb, 32'h3d50dbf8} /* (1, 27, 30) {real, imag} */,
  {32'h3d8c4f58, 32'hbd9749c3} /* (1, 27, 29) {real, imag} */,
  {32'hbe10a81d, 32'h3e473848} /* (1, 27, 28) {real, imag} */,
  {32'h3ea83587, 32'hbd7966f7} /* (1, 27, 27) {real, imag} */,
  {32'h3dbe8d07, 32'hbddd6439} /* (1, 27, 26) {real, imag} */,
  {32'h3cf68b3a, 32'hbc3414b0} /* (1, 27, 25) {real, imag} */,
  {32'h3d5b6df1, 32'hbdf0e8e6} /* (1, 27, 24) {real, imag} */,
  {32'hbd11f298, 32'hbd3d341b} /* (1, 27, 23) {real, imag} */,
  {32'hbc18470e, 32'h3c593c02} /* (1, 27, 22) {real, imag} */,
  {32'h3cc1e870, 32'h3d0aa1f2} /* (1, 27, 21) {real, imag} */,
  {32'hbca3e1ba, 32'h3d8f18ae} /* (1, 27, 20) {real, imag} */,
  {32'hbce18b80, 32'hbd073ef7} /* (1, 27, 19) {real, imag} */,
  {32'hbd88c491, 32'hbd2dfd2e} /* (1, 27, 18) {real, imag} */,
  {32'hbc39fa6a, 32'h3d8f25f8} /* (1, 27, 17) {real, imag} */,
  {32'h3d8b913e, 32'h00000000} /* (1, 27, 16) {real, imag} */,
  {32'hbc39fa6a, 32'hbd8f25f8} /* (1, 27, 15) {real, imag} */,
  {32'hbd88c491, 32'h3d2dfd2e} /* (1, 27, 14) {real, imag} */,
  {32'hbce18b80, 32'h3d073ef7} /* (1, 27, 13) {real, imag} */,
  {32'hbca3e1ba, 32'hbd8f18ae} /* (1, 27, 12) {real, imag} */,
  {32'h3cc1e870, 32'hbd0aa1f2} /* (1, 27, 11) {real, imag} */,
  {32'hbc18470e, 32'hbc593c02} /* (1, 27, 10) {real, imag} */,
  {32'hbd11f298, 32'h3d3d341b} /* (1, 27, 9) {real, imag} */,
  {32'h3d5b6df1, 32'h3df0e8e6} /* (1, 27, 8) {real, imag} */,
  {32'h3cf68b3a, 32'h3c3414b0} /* (1, 27, 7) {real, imag} */,
  {32'h3dbe8d07, 32'h3ddd6439} /* (1, 27, 6) {real, imag} */,
  {32'h3ea83587, 32'h3d7966f7} /* (1, 27, 5) {real, imag} */,
  {32'hbe10a81d, 32'hbe473848} /* (1, 27, 4) {real, imag} */,
  {32'h3d8c4f58, 32'h3d9749c3} /* (1, 27, 3) {real, imag} */,
  {32'h3f27b2bb, 32'hbd50dbf8} /* (1, 27, 2) {real, imag} */,
  {32'hbfd559aa, 32'hbe01d9cc} /* (1, 27, 1) {real, imag} */,
  {32'hbf11db1a, 32'h00000000} /* (1, 27, 0) {real, imag} */,
  {32'hbfce6c52, 32'h3dce283a} /* (1, 26, 31) {real, imag} */,
  {32'h3f09fd6b, 32'hbc70d040} /* (1, 26, 30) {real, imag} */,
  {32'hbd4d3202, 32'hbdd30f30} /* (1, 26, 29) {real, imag} */,
  {32'hbe05353a, 32'h3da3a4f2} /* (1, 26, 28) {real, imag} */,
  {32'h3e624dba, 32'hbe0822f9} /* (1, 26, 27) {real, imag} */,
  {32'h3e0e3c5a, 32'h3cf8b26c} /* (1, 26, 26) {real, imag} */,
  {32'hbd1066e9, 32'h3c1e29b0} /* (1, 26, 25) {real, imag} */,
  {32'h3d924d57, 32'hbdfb220a} /* (1, 26, 24) {real, imag} */,
  {32'h3d7b89c4, 32'hbd905d69} /* (1, 26, 23) {real, imag} */,
  {32'hbbeee088, 32'h3d66f5b9} /* (1, 26, 22) {real, imag} */,
  {32'hbd93261c, 32'hbd4ceb08} /* (1, 26, 21) {real, imag} */,
  {32'h3ca92f24, 32'hbb914bf8} /* (1, 26, 20) {real, imag} */,
  {32'hbb9778c0, 32'hbc2d8b14} /* (1, 26, 19) {real, imag} */,
  {32'h3ba403b0, 32'h3d5b3d28} /* (1, 26, 18) {real, imag} */,
  {32'hbc7597ae, 32'hbc04660c} /* (1, 26, 17) {real, imag} */,
  {32'hbd3b56fa, 32'h00000000} /* (1, 26, 16) {real, imag} */,
  {32'hbc7597ae, 32'h3c04660c} /* (1, 26, 15) {real, imag} */,
  {32'h3ba403b0, 32'hbd5b3d28} /* (1, 26, 14) {real, imag} */,
  {32'hbb9778c0, 32'h3c2d8b14} /* (1, 26, 13) {real, imag} */,
  {32'h3ca92f24, 32'h3b914bf8} /* (1, 26, 12) {real, imag} */,
  {32'hbd93261c, 32'h3d4ceb08} /* (1, 26, 11) {real, imag} */,
  {32'hbbeee088, 32'hbd66f5b9} /* (1, 26, 10) {real, imag} */,
  {32'h3d7b89c4, 32'h3d905d69} /* (1, 26, 9) {real, imag} */,
  {32'h3d924d57, 32'h3dfb220a} /* (1, 26, 8) {real, imag} */,
  {32'hbd1066e9, 32'hbc1e29b0} /* (1, 26, 7) {real, imag} */,
  {32'h3e0e3c5a, 32'hbcf8b26c} /* (1, 26, 6) {real, imag} */,
  {32'h3e624dba, 32'h3e0822f9} /* (1, 26, 5) {real, imag} */,
  {32'hbe05353a, 32'hbda3a4f2} /* (1, 26, 4) {real, imag} */,
  {32'hbd4d3202, 32'h3dd30f30} /* (1, 26, 3) {real, imag} */,
  {32'h3f09fd6b, 32'h3c70d040} /* (1, 26, 2) {real, imag} */,
  {32'hbfce6c52, 32'hbdce283a} /* (1, 26, 1) {real, imag} */,
  {32'hbf38ac70, 32'h00000000} /* (1, 26, 0) {real, imag} */,
  {32'hbfd6fd9d, 32'h3c0ff680} /* (1, 25, 31) {real, imag} */,
  {32'h3f19a775, 32'h3df9e4c5} /* (1, 25, 30) {real, imag} */,
  {32'h3c01a8c7, 32'hbd831e7b} /* (1, 25, 29) {real, imag} */,
  {32'hbe9ad8d3, 32'h3d6305e8} /* (1, 25, 28) {real, imag} */,
  {32'h3e1ba5ed, 32'hbda21bc8} /* (1, 25, 27) {real, imag} */,
  {32'h3d8257a9, 32'hbcedd0d7} /* (1, 25, 26) {real, imag} */,
  {32'hbd9f2eaf, 32'h3e2fa948} /* (1, 25, 25) {real, imag} */,
  {32'h3bd522a0, 32'hbe35205b} /* (1, 25, 24) {real, imag} */,
  {32'hbca0c8a0, 32'hbd49f2ce} /* (1, 25, 23) {real, imag} */,
  {32'hbd27a526, 32'hbd33e940} /* (1, 25, 22) {real, imag} */,
  {32'hbc971b00, 32'hbde1d6d6} /* (1, 25, 21) {real, imag} */,
  {32'h3d0d9c9d, 32'hbddcdc50} /* (1, 25, 20) {real, imag} */,
  {32'h3da56a03, 32'h3c60f647} /* (1, 25, 19) {real, imag} */,
  {32'h3bb57b44, 32'h3c5fddf4} /* (1, 25, 18) {real, imag} */,
  {32'h3c1a8c34, 32'hbad155d8} /* (1, 25, 17) {real, imag} */,
  {32'h3da77bfb, 32'h00000000} /* (1, 25, 16) {real, imag} */,
  {32'h3c1a8c34, 32'h3ad155d8} /* (1, 25, 15) {real, imag} */,
  {32'h3bb57b44, 32'hbc5fddf4} /* (1, 25, 14) {real, imag} */,
  {32'h3da56a03, 32'hbc60f647} /* (1, 25, 13) {real, imag} */,
  {32'h3d0d9c9d, 32'h3ddcdc50} /* (1, 25, 12) {real, imag} */,
  {32'hbc971b00, 32'h3de1d6d6} /* (1, 25, 11) {real, imag} */,
  {32'hbd27a526, 32'h3d33e940} /* (1, 25, 10) {real, imag} */,
  {32'hbca0c8a0, 32'h3d49f2ce} /* (1, 25, 9) {real, imag} */,
  {32'h3bd522a0, 32'h3e35205b} /* (1, 25, 8) {real, imag} */,
  {32'hbd9f2eaf, 32'hbe2fa948} /* (1, 25, 7) {real, imag} */,
  {32'h3d8257a9, 32'h3cedd0d7} /* (1, 25, 6) {real, imag} */,
  {32'h3e1ba5ed, 32'h3da21bc8} /* (1, 25, 5) {real, imag} */,
  {32'hbe9ad8d3, 32'hbd6305e8} /* (1, 25, 4) {real, imag} */,
  {32'h3c01a8c7, 32'h3d831e7b} /* (1, 25, 3) {real, imag} */,
  {32'h3f19a775, 32'hbdf9e4c5} /* (1, 25, 2) {real, imag} */,
  {32'hbfd6fd9d, 32'hbc0ff680} /* (1, 25, 1) {real, imag} */,
  {32'hbf31851b, 32'h00000000} /* (1, 25, 0) {real, imag} */,
  {32'hbfc7d44c, 32'hbd87782e} /* (1, 24, 31) {real, imag} */,
  {32'h3f34db74, 32'h3e1c89ed} /* (1, 24, 30) {real, imag} */,
  {32'hbbf81630, 32'hbd979591} /* (1, 24, 29) {real, imag} */,
  {32'hbea653a1, 32'hbc91c83c} /* (1, 24, 28) {real, imag} */,
  {32'h3e5f35e2, 32'h3be0c080} /* (1, 24, 27) {real, imag} */,
  {32'hbd18968c, 32'h3c7a5990} /* (1, 24, 26) {real, imag} */,
  {32'hbd377582, 32'h3dd27f67} /* (1, 24, 25) {real, imag} */,
  {32'h3d4eb65a, 32'hbd5abff7} /* (1, 24, 24) {real, imag} */,
  {32'h3d8619e0, 32'hbcb3fd08} /* (1, 24, 23) {real, imag} */,
  {32'hbd3936d5, 32'h3d98c915} /* (1, 24, 22) {real, imag} */,
  {32'h3d897136, 32'hbd9789d9} /* (1, 24, 21) {real, imag} */,
  {32'hbdb6b54a, 32'h3daaa458} /* (1, 24, 20) {real, imag} */,
  {32'h3a49b2e0, 32'h3d2db16a} /* (1, 24, 19) {real, imag} */,
  {32'h3c9e788a, 32'hbdb1fff0} /* (1, 24, 18) {real, imag} */,
  {32'hbd00edb6, 32'h3c4f87a3} /* (1, 24, 17) {real, imag} */,
  {32'hbc960126, 32'h00000000} /* (1, 24, 16) {real, imag} */,
  {32'hbd00edb6, 32'hbc4f87a3} /* (1, 24, 15) {real, imag} */,
  {32'h3c9e788a, 32'h3db1fff0} /* (1, 24, 14) {real, imag} */,
  {32'h3a49b2e0, 32'hbd2db16a} /* (1, 24, 13) {real, imag} */,
  {32'hbdb6b54a, 32'hbdaaa458} /* (1, 24, 12) {real, imag} */,
  {32'h3d897136, 32'h3d9789d9} /* (1, 24, 11) {real, imag} */,
  {32'hbd3936d5, 32'hbd98c915} /* (1, 24, 10) {real, imag} */,
  {32'h3d8619e0, 32'h3cb3fd08} /* (1, 24, 9) {real, imag} */,
  {32'h3d4eb65a, 32'h3d5abff7} /* (1, 24, 8) {real, imag} */,
  {32'hbd377582, 32'hbdd27f67} /* (1, 24, 7) {real, imag} */,
  {32'hbd18968c, 32'hbc7a5990} /* (1, 24, 6) {real, imag} */,
  {32'h3e5f35e2, 32'hbbe0c080} /* (1, 24, 5) {real, imag} */,
  {32'hbea653a1, 32'h3c91c83c} /* (1, 24, 4) {real, imag} */,
  {32'hbbf81630, 32'h3d979591} /* (1, 24, 3) {real, imag} */,
  {32'h3f34db74, 32'hbe1c89ed} /* (1, 24, 2) {real, imag} */,
  {32'hbfc7d44c, 32'h3d87782e} /* (1, 24, 1) {real, imag} */,
  {32'hbf030b24, 32'h00000000} /* (1, 24, 0) {real, imag} */,
  {32'hbfae59d3, 32'h3d473e7e} /* (1, 23, 31) {real, imag} */,
  {32'h3eecad30, 32'h3db3e9f1} /* (1, 23, 30) {real, imag} */,
  {32'h3dcac1c8, 32'h3ccf6dc6} /* (1, 23, 29) {real, imag} */,
  {32'hbe77f5ae, 32'h3bafe114} /* (1, 23, 28) {real, imag} */,
  {32'h3d8370d5, 32'hbde7fb71} /* (1, 23, 27) {real, imag} */,
  {32'h3d237838, 32'h3d695115} /* (1, 23, 26) {real, imag} */,
  {32'hbcda04cc, 32'h3d8bf520} /* (1, 23, 25) {real, imag} */,
  {32'h3c423270, 32'hbd936ce2} /* (1, 23, 24) {real, imag} */,
  {32'h3c890571, 32'hbd5f2e9c} /* (1, 23, 23) {real, imag} */,
  {32'h3cec3781, 32'hbd32fac7} /* (1, 23, 22) {real, imag} */,
  {32'h3d39c8f5, 32'hbd85fa54} /* (1, 23, 21) {real, imag} */,
  {32'h3cdf917c, 32'h3d6ccb33} /* (1, 23, 20) {real, imag} */,
  {32'hbc38578e, 32'h3cdff9c6} /* (1, 23, 19) {real, imag} */,
  {32'h3d0ad3b6, 32'hbdcb671e} /* (1, 23, 18) {real, imag} */,
  {32'h3d5411d3, 32'h3db54013} /* (1, 23, 17) {real, imag} */,
  {32'h3bed7046, 32'h00000000} /* (1, 23, 16) {real, imag} */,
  {32'h3d5411d3, 32'hbdb54013} /* (1, 23, 15) {real, imag} */,
  {32'h3d0ad3b6, 32'h3dcb671e} /* (1, 23, 14) {real, imag} */,
  {32'hbc38578e, 32'hbcdff9c6} /* (1, 23, 13) {real, imag} */,
  {32'h3cdf917c, 32'hbd6ccb33} /* (1, 23, 12) {real, imag} */,
  {32'h3d39c8f5, 32'h3d85fa54} /* (1, 23, 11) {real, imag} */,
  {32'h3cec3781, 32'h3d32fac7} /* (1, 23, 10) {real, imag} */,
  {32'h3c890571, 32'h3d5f2e9c} /* (1, 23, 9) {real, imag} */,
  {32'h3c423270, 32'h3d936ce2} /* (1, 23, 8) {real, imag} */,
  {32'hbcda04cc, 32'hbd8bf520} /* (1, 23, 7) {real, imag} */,
  {32'h3d237838, 32'hbd695115} /* (1, 23, 6) {real, imag} */,
  {32'h3d8370d5, 32'h3de7fb71} /* (1, 23, 5) {real, imag} */,
  {32'hbe77f5ae, 32'hbbafe114} /* (1, 23, 4) {real, imag} */,
  {32'h3dcac1c8, 32'hbccf6dc6} /* (1, 23, 3) {real, imag} */,
  {32'h3eecad30, 32'hbdb3e9f1} /* (1, 23, 2) {real, imag} */,
  {32'hbfae59d3, 32'hbd473e7e} /* (1, 23, 1) {real, imag} */,
  {32'hbe9f8856, 32'h00000000} /* (1, 23, 0) {real, imag} */,
  {32'hbf8a61c2, 32'h3dae4d6e} /* (1, 22, 31) {real, imag} */,
  {32'h3edadfde, 32'h3d8bee02} /* (1, 22, 30) {real, imag} */,
  {32'h3dd639c5, 32'h3d9ecac8} /* (1, 22, 29) {real, imag} */,
  {32'hbdff5d78, 32'hbdc2daf8} /* (1, 22, 28) {real, imag} */,
  {32'h3da3b576, 32'hbe30f0b0} /* (1, 22, 27) {real, imag} */,
  {32'hbd22ddea, 32'h3ba330f6} /* (1, 22, 26) {real, imag} */,
  {32'hbe1348b4, 32'h3d7ffc2b} /* (1, 22, 25) {real, imag} */,
  {32'h3d65d528, 32'hbd1a6e71} /* (1, 22, 24) {real, imag} */,
  {32'hbd8e4f60, 32'h3cbccd2d} /* (1, 22, 23) {real, imag} */,
  {32'h3dbd85ad, 32'h3e0d8bb4} /* (1, 22, 22) {real, imag} */,
  {32'h3cdc4ebe, 32'hbd5afe8a} /* (1, 22, 21) {real, imag} */,
  {32'h3cd087d1, 32'h3d065f5c} /* (1, 22, 20) {real, imag} */,
  {32'h3c86f24b, 32'hbc34d51c} /* (1, 22, 19) {real, imag} */,
  {32'h3c6df7e0, 32'hbcc9ba6c} /* (1, 22, 18) {real, imag} */,
  {32'hbcd087f1, 32'h3c90c1be} /* (1, 22, 17) {real, imag} */,
  {32'h3da0bf8e, 32'h00000000} /* (1, 22, 16) {real, imag} */,
  {32'hbcd087f1, 32'hbc90c1be} /* (1, 22, 15) {real, imag} */,
  {32'h3c6df7e0, 32'h3cc9ba6c} /* (1, 22, 14) {real, imag} */,
  {32'h3c86f24b, 32'h3c34d51c} /* (1, 22, 13) {real, imag} */,
  {32'h3cd087d1, 32'hbd065f5c} /* (1, 22, 12) {real, imag} */,
  {32'h3cdc4ebe, 32'h3d5afe8a} /* (1, 22, 11) {real, imag} */,
  {32'h3dbd85ad, 32'hbe0d8bb4} /* (1, 22, 10) {real, imag} */,
  {32'hbd8e4f60, 32'hbcbccd2d} /* (1, 22, 9) {real, imag} */,
  {32'h3d65d528, 32'h3d1a6e71} /* (1, 22, 8) {real, imag} */,
  {32'hbe1348b4, 32'hbd7ffc2b} /* (1, 22, 7) {real, imag} */,
  {32'hbd22ddea, 32'hbba330f6} /* (1, 22, 6) {real, imag} */,
  {32'h3da3b576, 32'h3e30f0b0} /* (1, 22, 5) {real, imag} */,
  {32'hbdff5d78, 32'h3dc2daf8} /* (1, 22, 4) {real, imag} */,
  {32'h3dd639c5, 32'hbd9ecac8} /* (1, 22, 3) {real, imag} */,
  {32'h3edadfde, 32'hbd8bee02} /* (1, 22, 2) {real, imag} */,
  {32'hbf8a61c2, 32'hbdae4d6e} /* (1, 22, 1) {real, imag} */,
  {32'hbe600bf6, 32'h00000000} /* (1, 22, 0) {real, imag} */,
  {32'hbee6dfd4, 32'h3c933588} /* (1, 21, 31) {real, imag} */,
  {32'h3e00e04c, 32'h3b833600} /* (1, 21, 30) {real, imag} */,
  {32'hbcb1a0b7, 32'h3df0397b} /* (1, 21, 29) {real, imag} */,
  {32'hbdd19bd6, 32'h3ca06bc0} /* (1, 21, 28) {real, imag} */,
  {32'h3d62ec50, 32'hbd61b87f} /* (1, 21, 27) {real, imag} */,
  {32'hbd4200a8, 32'h3a8cf040} /* (1, 21, 26) {real, imag} */,
  {32'hbd23742d, 32'h3d50f97e} /* (1, 21, 25) {real, imag} */,
  {32'hbd9e1288, 32'hbd0f3287} /* (1, 21, 24) {real, imag} */,
  {32'h3d4b1d70, 32'h3dcc97ac} /* (1, 21, 23) {real, imag} */,
  {32'h3d5602e4, 32'h3ccd8904} /* (1, 21, 22) {real, imag} */,
  {32'h3da2813e, 32'h3dadfcc7} /* (1, 21, 21) {real, imag} */,
  {32'h3d67b6ad, 32'hbd676b67} /* (1, 21, 20) {real, imag} */,
  {32'h3d3bea8a, 32'h3cb969e8} /* (1, 21, 19) {real, imag} */,
  {32'h3c215b2f, 32'hbd217a5f} /* (1, 21, 18) {real, imag} */,
  {32'hbcdfd983, 32'hbbe0297c} /* (1, 21, 17) {real, imag} */,
  {32'hbd5c51b7, 32'h00000000} /* (1, 21, 16) {real, imag} */,
  {32'hbcdfd983, 32'h3be0297c} /* (1, 21, 15) {real, imag} */,
  {32'h3c215b2f, 32'h3d217a5f} /* (1, 21, 14) {real, imag} */,
  {32'h3d3bea8a, 32'hbcb969e8} /* (1, 21, 13) {real, imag} */,
  {32'h3d67b6ad, 32'h3d676b67} /* (1, 21, 12) {real, imag} */,
  {32'h3da2813e, 32'hbdadfcc7} /* (1, 21, 11) {real, imag} */,
  {32'h3d5602e4, 32'hbccd8904} /* (1, 21, 10) {real, imag} */,
  {32'h3d4b1d70, 32'hbdcc97ac} /* (1, 21, 9) {real, imag} */,
  {32'hbd9e1288, 32'h3d0f3287} /* (1, 21, 8) {real, imag} */,
  {32'hbd23742d, 32'hbd50f97e} /* (1, 21, 7) {real, imag} */,
  {32'hbd4200a8, 32'hba8cf040} /* (1, 21, 6) {real, imag} */,
  {32'h3d62ec50, 32'h3d61b87f} /* (1, 21, 5) {real, imag} */,
  {32'hbdd19bd6, 32'hbca06bc0} /* (1, 21, 4) {real, imag} */,
  {32'hbcb1a0b7, 32'hbdf0397b} /* (1, 21, 3) {real, imag} */,
  {32'h3e00e04c, 32'hbb833600} /* (1, 21, 2) {real, imag} */,
  {32'hbee6dfd4, 32'hbc933588} /* (1, 21, 1) {real, imag} */,
  {32'hbcce0f30, 32'h00000000} /* (1, 21, 0) {real, imag} */,
  {32'h3f0e253e, 32'hbe7f4662} /* (1, 20, 31) {real, imag} */,
  {32'hbed3f884, 32'h3d54f71f} /* (1, 20, 30) {real, imag} */,
  {32'h3d0a913c, 32'h3e097154} /* (1, 20, 29) {real, imag} */,
  {32'hbc0f99a0, 32'hbd873e53} /* (1, 20, 28) {real, imag} */,
  {32'hbe00d642, 32'h3cfd5a2c} /* (1, 20, 27) {real, imag} */,
  {32'hbde54076, 32'h3d6ba22b} /* (1, 20, 26) {real, imag} */,
  {32'hbdb228d0, 32'h3a673f10} /* (1, 20, 25) {real, imag} */,
  {32'hbd5524c8, 32'h3dec63b1} /* (1, 20, 24) {real, imag} */,
  {32'h3c7f6824, 32'hbda5349c} /* (1, 20, 23) {real, imag} */,
  {32'hbc9961c2, 32'hbd637b65} /* (1, 20, 22) {real, imag} */,
  {32'hbd78cad8, 32'hbd8b2442} /* (1, 20, 21) {real, imag} */,
  {32'hbc988273, 32'h3d5f0aa6} /* (1, 20, 20) {real, imag} */,
  {32'h3cd0f7e2, 32'hbd85d476} /* (1, 20, 19) {real, imag} */,
  {32'h3c913bb8, 32'hbd4b843c} /* (1, 20, 18) {real, imag} */,
  {32'hbd0a25f1, 32'hbcaf65bc} /* (1, 20, 17) {real, imag} */,
  {32'h3cc59bce, 32'h00000000} /* (1, 20, 16) {real, imag} */,
  {32'hbd0a25f1, 32'h3caf65bc} /* (1, 20, 15) {real, imag} */,
  {32'h3c913bb8, 32'h3d4b843c} /* (1, 20, 14) {real, imag} */,
  {32'h3cd0f7e2, 32'h3d85d476} /* (1, 20, 13) {real, imag} */,
  {32'hbc988273, 32'hbd5f0aa6} /* (1, 20, 12) {real, imag} */,
  {32'hbd78cad8, 32'h3d8b2442} /* (1, 20, 11) {real, imag} */,
  {32'hbc9961c2, 32'h3d637b65} /* (1, 20, 10) {real, imag} */,
  {32'h3c7f6824, 32'h3da5349c} /* (1, 20, 9) {real, imag} */,
  {32'hbd5524c8, 32'hbdec63b1} /* (1, 20, 8) {real, imag} */,
  {32'hbdb228d0, 32'hba673f10} /* (1, 20, 7) {real, imag} */,
  {32'hbde54076, 32'hbd6ba22b} /* (1, 20, 6) {real, imag} */,
  {32'hbe00d642, 32'hbcfd5a2c} /* (1, 20, 5) {real, imag} */,
  {32'hbc0f99a0, 32'h3d873e53} /* (1, 20, 4) {real, imag} */,
  {32'h3d0a913c, 32'hbe097154} /* (1, 20, 3) {real, imag} */,
  {32'hbed3f884, 32'hbd54f71f} /* (1, 20, 2) {real, imag} */,
  {32'h3f0e253e, 32'h3e7f4662} /* (1, 20, 1) {real, imag} */,
  {32'h3f111036, 32'h00000000} /* (1, 20, 0) {real, imag} */,
  {32'h3f836bc5, 32'hbe9a26bc} /* (1, 19, 31) {real, imag} */,
  {32'hbf0ff06a, 32'h3e7f9082} /* (1, 19, 30) {real, imag} */,
  {32'hbbc81d08, 32'h3e035c07} /* (1, 19, 29) {real, imag} */,
  {32'h3de818a7, 32'hbe1a54e0} /* (1, 19, 28) {real, imag} */,
  {32'hbe1453e6, 32'h3d6cbe24} /* (1, 19, 27) {real, imag} */,
  {32'hbd68768f, 32'hbcca4963} /* (1, 19, 26) {real, imag} */,
  {32'h3cb167b3, 32'hbd8d828a} /* (1, 19, 25) {real, imag} */,
  {32'hbd0ebebd, 32'hbc72b4dc} /* (1, 19, 24) {real, imag} */,
  {32'h3d3de9b4, 32'h3caa027e} /* (1, 19, 23) {real, imag} */,
  {32'h3d36de56, 32'h3c8cc30f} /* (1, 19, 22) {real, imag} */,
  {32'hbca8677e, 32'h3d034898} /* (1, 19, 21) {real, imag} */,
  {32'h3c628404, 32'h3d78e4fa} /* (1, 19, 20) {real, imag} */,
  {32'hbc7989e8, 32'h3d30e8d2} /* (1, 19, 19) {real, imag} */,
  {32'hbc857b5d, 32'h3cdbe43e} /* (1, 19, 18) {real, imag} */,
  {32'hbd363627, 32'hbd06380e} /* (1, 19, 17) {real, imag} */,
  {32'hbe1902e2, 32'h00000000} /* (1, 19, 16) {real, imag} */,
  {32'hbd363627, 32'h3d06380e} /* (1, 19, 15) {real, imag} */,
  {32'hbc857b5d, 32'hbcdbe43e} /* (1, 19, 14) {real, imag} */,
  {32'hbc7989e8, 32'hbd30e8d2} /* (1, 19, 13) {real, imag} */,
  {32'h3c628404, 32'hbd78e4fa} /* (1, 19, 12) {real, imag} */,
  {32'hbca8677e, 32'hbd034898} /* (1, 19, 11) {real, imag} */,
  {32'h3d36de56, 32'hbc8cc30f} /* (1, 19, 10) {real, imag} */,
  {32'h3d3de9b4, 32'hbcaa027e} /* (1, 19, 9) {real, imag} */,
  {32'hbd0ebebd, 32'h3c72b4dc} /* (1, 19, 8) {real, imag} */,
  {32'h3cb167b3, 32'h3d8d828a} /* (1, 19, 7) {real, imag} */,
  {32'hbd68768f, 32'h3cca4963} /* (1, 19, 6) {real, imag} */,
  {32'hbe1453e6, 32'hbd6cbe24} /* (1, 19, 5) {real, imag} */,
  {32'h3de818a7, 32'h3e1a54e0} /* (1, 19, 4) {real, imag} */,
  {32'hbbc81d08, 32'hbe035c07} /* (1, 19, 3) {real, imag} */,
  {32'hbf0ff06a, 32'hbe7f9082} /* (1, 19, 2) {real, imag} */,
  {32'h3f836bc5, 32'h3e9a26bc} /* (1, 19, 1) {real, imag} */,
  {32'h3f6f3bd3, 32'h00000000} /* (1, 19, 0) {real, imag} */,
  {32'h3f8fe388, 32'hbe53e288} /* (1, 18, 31) {real, imag} */,
  {32'hbf342999, 32'h3e005f76} /* (1, 18, 30) {real, imag} */,
  {32'hbd57d53e, 32'h3c9a54af} /* (1, 18, 29) {real, imag} */,
  {32'h3e429720, 32'h3cbdc0d6} /* (1, 18, 28) {real, imag} */,
  {32'hbdb5ef13, 32'h3d39919f} /* (1, 18, 27) {real, imag} */,
  {32'h3d41d45c, 32'h3b324f90} /* (1, 18, 26) {real, imag} */,
  {32'hbd0b69d5, 32'hbd4ce911} /* (1, 18, 25) {real, imag} */,
  {32'hbd8e58d0, 32'hbe0697f7} /* (1, 18, 24) {real, imag} */,
  {32'hbc0cbeb0, 32'h3cc97012} /* (1, 18, 23) {real, imag} */,
  {32'h3d06ec3a, 32'h3c9c1ccf} /* (1, 18, 22) {real, imag} */,
  {32'hbb7f9bf8, 32'h3d7ae7fe} /* (1, 18, 21) {real, imag} */,
  {32'h3c0d1fae, 32'hbd21ebac} /* (1, 18, 20) {real, imag} */,
  {32'h3e0ef2a9, 32'hbd95fc0c} /* (1, 18, 19) {real, imag} */,
  {32'h3d9ce1d4, 32'h3ce682e4} /* (1, 18, 18) {real, imag} */,
  {32'h3c78335c, 32'h3d8add3c} /* (1, 18, 17) {real, imag} */,
  {32'h3d568417, 32'h00000000} /* (1, 18, 16) {real, imag} */,
  {32'h3c78335c, 32'hbd8add3c} /* (1, 18, 15) {real, imag} */,
  {32'h3d9ce1d4, 32'hbce682e4} /* (1, 18, 14) {real, imag} */,
  {32'h3e0ef2a9, 32'h3d95fc0c} /* (1, 18, 13) {real, imag} */,
  {32'h3c0d1fae, 32'h3d21ebac} /* (1, 18, 12) {real, imag} */,
  {32'hbb7f9bf8, 32'hbd7ae7fe} /* (1, 18, 11) {real, imag} */,
  {32'h3d06ec3a, 32'hbc9c1ccf} /* (1, 18, 10) {real, imag} */,
  {32'hbc0cbeb0, 32'hbcc97012} /* (1, 18, 9) {real, imag} */,
  {32'hbd8e58d0, 32'h3e0697f7} /* (1, 18, 8) {real, imag} */,
  {32'hbd0b69d5, 32'h3d4ce911} /* (1, 18, 7) {real, imag} */,
  {32'h3d41d45c, 32'hbb324f90} /* (1, 18, 6) {real, imag} */,
  {32'hbdb5ef13, 32'hbd39919f} /* (1, 18, 5) {real, imag} */,
  {32'h3e429720, 32'hbcbdc0d6} /* (1, 18, 4) {real, imag} */,
  {32'hbd57d53e, 32'hbc9a54af} /* (1, 18, 3) {real, imag} */,
  {32'hbf342999, 32'hbe005f76} /* (1, 18, 2) {real, imag} */,
  {32'h3f8fe388, 32'h3e53e288} /* (1, 18, 1) {real, imag} */,
  {32'h3f82a12b, 32'h00000000} /* (1, 18, 0) {real, imag} */,
  {32'h3fa434e2, 32'hbe802c4b} /* (1, 17, 31) {real, imag} */,
  {32'hbf54b398, 32'h3d5b086c} /* (1, 17, 30) {real, imag} */,
  {32'hbd23422d, 32'hbd83d1ed} /* (1, 17, 29) {real, imag} */,
  {32'h3e415f48, 32'hbe01e2b4} /* (1, 17, 28) {real, imag} */,
  {32'hbdc15ba3, 32'h3d5f9782} /* (1, 17, 27) {real, imag} */,
  {32'h3d280145, 32'hbcf1daac} /* (1, 17, 26) {real, imag} */,
  {32'h3dd8c955, 32'h3cb90418} /* (1, 17, 25) {real, imag} */,
  {32'hbe291aae, 32'hb9eba000} /* (1, 17, 24) {real, imag} */,
  {32'hbd8d2327, 32'hbc66bfe8} /* (1, 17, 23) {real, imag} */,
  {32'h3d050a41, 32'hbd58189e} /* (1, 17, 22) {real, imag} */,
  {32'hbb5a46c8, 32'hbd9fc8ec} /* (1, 17, 21) {real, imag} */,
  {32'hbda96cf2, 32'h3dd34791} /* (1, 17, 20) {real, imag} */,
  {32'h3bc548e0, 32'h3dba4be9} /* (1, 17, 19) {real, imag} */,
  {32'hbd3475fa, 32'hbc6c0aef} /* (1, 17, 18) {real, imag} */,
  {32'hbca61bae, 32'hbd854aeb} /* (1, 17, 17) {real, imag} */,
  {32'h3da12d8d, 32'h00000000} /* (1, 17, 16) {real, imag} */,
  {32'hbca61bae, 32'h3d854aeb} /* (1, 17, 15) {real, imag} */,
  {32'hbd3475fa, 32'h3c6c0aef} /* (1, 17, 14) {real, imag} */,
  {32'h3bc548e0, 32'hbdba4be9} /* (1, 17, 13) {real, imag} */,
  {32'hbda96cf2, 32'hbdd34791} /* (1, 17, 12) {real, imag} */,
  {32'hbb5a46c8, 32'h3d9fc8ec} /* (1, 17, 11) {real, imag} */,
  {32'h3d050a41, 32'h3d58189e} /* (1, 17, 10) {real, imag} */,
  {32'hbd8d2327, 32'h3c66bfe8} /* (1, 17, 9) {real, imag} */,
  {32'hbe291aae, 32'h39eba000} /* (1, 17, 8) {real, imag} */,
  {32'h3dd8c955, 32'hbcb90418} /* (1, 17, 7) {real, imag} */,
  {32'h3d280145, 32'h3cf1daac} /* (1, 17, 6) {real, imag} */,
  {32'hbdc15ba3, 32'hbd5f9782} /* (1, 17, 5) {real, imag} */,
  {32'h3e415f48, 32'h3e01e2b4} /* (1, 17, 4) {real, imag} */,
  {32'hbd23422d, 32'h3d83d1ed} /* (1, 17, 3) {real, imag} */,
  {32'hbf54b398, 32'hbd5b086c} /* (1, 17, 2) {real, imag} */,
  {32'h3fa434e2, 32'h3e802c4b} /* (1, 17, 1) {real, imag} */,
  {32'h3f934e21, 32'h00000000} /* (1, 17, 0) {real, imag} */,
  {32'h3faa108c, 32'hbe64ace8} /* (1, 16, 31) {real, imag} */,
  {32'hbf546434, 32'h3df37dc4} /* (1, 16, 30) {real, imag} */,
  {32'h3d8bb28e, 32'hbe02ba4b} /* (1, 16, 29) {real, imag} */,
  {32'h3e17fee8, 32'hbe0bfb73} /* (1, 16, 28) {real, imag} */,
  {32'hbdc3b84e, 32'h3e4fec0c} /* (1, 16, 27) {real, imag} */,
  {32'h3d8a3583, 32'h3d863507} /* (1, 16, 26) {real, imag} */,
  {32'h3d92639c, 32'hbccc4d6a} /* (1, 16, 25) {real, imag} */,
  {32'hbd9c1be8, 32'h3e01831e} /* (1, 16, 24) {real, imag} */,
  {32'hba2b26c0, 32'h3d56aa1d} /* (1, 16, 23) {real, imag} */,
  {32'h3dcc64f6, 32'hbd65d2ef} /* (1, 16, 22) {real, imag} */,
  {32'h3c018bba, 32'h3d984e96} /* (1, 16, 21) {real, imag} */,
  {32'hbcb02530, 32'h3d850c8f} /* (1, 16, 20) {real, imag} */,
  {32'hbcbb0266, 32'h3cf934de} /* (1, 16, 19) {real, imag} */,
  {32'h3cf20280, 32'hbd04e9ac} /* (1, 16, 18) {real, imag} */,
  {32'hbbf5a8de, 32'hbc7173db} /* (1, 16, 17) {real, imag} */,
  {32'hbd219806, 32'h00000000} /* (1, 16, 16) {real, imag} */,
  {32'hbbf5a8de, 32'h3c7173db} /* (1, 16, 15) {real, imag} */,
  {32'h3cf20280, 32'h3d04e9ac} /* (1, 16, 14) {real, imag} */,
  {32'hbcbb0266, 32'hbcf934de} /* (1, 16, 13) {real, imag} */,
  {32'hbcb02530, 32'hbd850c8f} /* (1, 16, 12) {real, imag} */,
  {32'h3c018bba, 32'hbd984e96} /* (1, 16, 11) {real, imag} */,
  {32'h3dcc64f6, 32'h3d65d2ef} /* (1, 16, 10) {real, imag} */,
  {32'hba2b26c0, 32'hbd56aa1d} /* (1, 16, 9) {real, imag} */,
  {32'hbd9c1be8, 32'hbe01831e} /* (1, 16, 8) {real, imag} */,
  {32'h3d92639c, 32'h3ccc4d6a} /* (1, 16, 7) {real, imag} */,
  {32'h3d8a3583, 32'hbd863507} /* (1, 16, 6) {real, imag} */,
  {32'hbdc3b84e, 32'hbe4fec0c} /* (1, 16, 5) {real, imag} */,
  {32'h3e17fee8, 32'h3e0bfb73} /* (1, 16, 4) {real, imag} */,
  {32'h3d8bb28e, 32'h3e02ba4b} /* (1, 16, 3) {real, imag} */,
  {32'hbf546434, 32'hbdf37dc4} /* (1, 16, 2) {real, imag} */,
  {32'h3faa108c, 32'h3e64ace8} /* (1, 16, 1) {real, imag} */,
  {32'h3f8c1a27, 32'h00000000} /* (1, 16, 0) {real, imag} */,
  {32'h3fc2f082, 32'hbe5ad89a} /* (1, 15, 31) {real, imag} */,
  {32'hbf26349c, 32'h3e2fcbe5} /* (1, 15, 30) {real, imag} */,
  {32'hbd8e058a, 32'hbdad3069} /* (1, 15, 29) {real, imag} */,
  {32'h3e0a64b0, 32'hbda281a1} /* (1, 15, 28) {real, imag} */,
  {32'hbe2d4514, 32'h3e21aaac} /* (1, 15, 27) {real, imag} */,
  {32'h3cd7d1ea, 32'h3d5c5072} /* (1, 15, 26) {real, imag} */,
  {32'h3cbab43c, 32'h3c39e9a4} /* (1, 15, 25) {real, imag} */,
  {32'hbdd31243, 32'h3e13f86c} /* (1, 15, 24) {real, imag} */,
  {32'h3dba7ae5, 32'h3d5679b6} /* (1, 15, 23) {real, imag} */,
  {32'hbd4d8c7d, 32'h3c90a11f} /* (1, 15, 22) {real, imag} */,
  {32'h3cbce23d, 32'h3dbf9e44} /* (1, 15, 21) {real, imag} */,
  {32'hbcbb82ee, 32'h3c204aa8} /* (1, 15, 20) {real, imag} */,
  {32'hbd5324f2, 32'hbd97d233} /* (1, 15, 19) {real, imag} */,
  {32'hbd221516, 32'hbca3293a} /* (1, 15, 18) {real, imag} */,
  {32'h3c6f8974, 32'hbbf0c634} /* (1, 15, 17) {real, imag} */,
  {32'hbd1db93a, 32'h00000000} /* (1, 15, 16) {real, imag} */,
  {32'h3c6f8974, 32'h3bf0c634} /* (1, 15, 15) {real, imag} */,
  {32'hbd221516, 32'h3ca3293a} /* (1, 15, 14) {real, imag} */,
  {32'hbd5324f2, 32'h3d97d233} /* (1, 15, 13) {real, imag} */,
  {32'hbcbb82ee, 32'hbc204aa8} /* (1, 15, 12) {real, imag} */,
  {32'h3cbce23d, 32'hbdbf9e44} /* (1, 15, 11) {real, imag} */,
  {32'hbd4d8c7d, 32'hbc90a11f} /* (1, 15, 10) {real, imag} */,
  {32'h3dba7ae5, 32'hbd5679b6} /* (1, 15, 9) {real, imag} */,
  {32'hbdd31243, 32'hbe13f86c} /* (1, 15, 8) {real, imag} */,
  {32'h3cbab43c, 32'hbc39e9a4} /* (1, 15, 7) {real, imag} */,
  {32'h3cd7d1ea, 32'hbd5c5072} /* (1, 15, 6) {real, imag} */,
  {32'hbe2d4514, 32'hbe21aaac} /* (1, 15, 5) {real, imag} */,
  {32'h3e0a64b0, 32'h3da281a1} /* (1, 15, 4) {real, imag} */,
  {32'hbd8e058a, 32'h3dad3069} /* (1, 15, 3) {real, imag} */,
  {32'hbf26349c, 32'hbe2fcbe5} /* (1, 15, 2) {real, imag} */,
  {32'h3fc2f082, 32'h3e5ad89a} /* (1, 15, 1) {real, imag} */,
  {32'h3f8e3dc1, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'h3fd10e34, 32'hbe8a0872} /* (1, 14, 31) {real, imag} */,
  {32'hbf33b965, 32'h3d97c60c} /* (1, 14, 30) {real, imag} */,
  {32'hbd226d0a, 32'hbd7f401c} /* (1, 14, 29) {real, imag} */,
  {32'h3de3b0f7, 32'hbd878ea4} /* (1, 14, 28) {real, imag} */,
  {32'hbe771f06, 32'h3de2d778} /* (1, 14, 27) {real, imag} */,
  {32'h3d418064, 32'hbd9f894c} /* (1, 14, 26) {real, imag} */,
  {32'hbdb427cc, 32'h397f2500} /* (1, 14, 25) {real, imag} */,
  {32'hbd98d844, 32'hbc6e7494} /* (1, 14, 24) {real, imag} */,
  {32'hbdb56556, 32'h3d684687} /* (1, 14, 23) {real, imag} */,
  {32'h3bb9cfc0, 32'hbbc02c94} /* (1, 14, 22) {real, imag} */,
  {32'hbd68b4dc, 32'h3cd5c018} /* (1, 14, 21) {real, imag} */,
  {32'h3d4f7d5e, 32'h3d1ff73e} /* (1, 14, 20) {real, imag} */,
  {32'hbc750990, 32'h3bcbc600} /* (1, 14, 19) {real, imag} */,
  {32'h3ca983f6, 32'h3c1065e0} /* (1, 14, 18) {real, imag} */,
  {32'hbd9659b8, 32'hbbbb2ec0} /* (1, 14, 17) {real, imag} */,
  {32'h3dbd908c, 32'h00000000} /* (1, 14, 16) {real, imag} */,
  {32'hbd9659b8, 32'h3bbb2ec0} /* (1, 14, 15) {real, imag} */,
  {32'h3ca983f6, 32'hbc1065e0} /* (1, 14, 14) {real, imag} */,
  {32'hbc750990, 32'hbbcbc600} /* (1, 14, 13) {real, imag} */,
  {32'h3d4f7d5e, 32'hbd1ff73e} /* (1, 14, 12) {real, imag} */,
  {32'hbd68b4dc, 32'hbcd5c018} /* (1, 14, 11) {real, imag} */,
  {32'h3bb9cfc0, 32'h3bc02c94} /* (1, 14, 10) {real, imag} */,
  {32'hbdb56556, 32'hbd684687} /* (1, 14, 9) {real, imag} */,
  {32'hbd98d844, 32'h3c6e7494} /* (1, 14, 8) {real, imag} */,
  {32'hbdb427cc, 32'hb97f2500} /* (1, 14, 7) {real, imag} */,
  {32'h3d418064, 32'h3d9f894c} /* (1, 14, 6) {real, imag} */,
  {32'hbe771f06, 32'hbde2d778} /* (1, 14, 5) {real, imag} */,
  {32'h3de3b0f7, 32'h3d878ea4} /* (1, 14, 4) {real, imag} */,
  {32'hbd226d0a, 32'h3d7f401c} /* (1, 14, 3) {real, imag} */,
  {32'hbf33b965, 32'hbd97c60c} /* (1, 14, 2) {real, imag} */,
  {32'h3fd10e34, 32'h3e8a0872} /* (1, 14, 1) {real, imag} */,
  {32'h3f76427b, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'h3fcf8c97, 32'hbe8e6f30} /* (1, 13, 31) {real, imag} */,
  {32'hbf390aa6, 32'hbd1b1cc0} /* (1, 13, 30) {real, imag} */,
  {32'hbd34ee3d, 32'h3cfe7df8} /* (1, 13, 29) {real, imag} */,
  {32'h3db77749, 32'hbda41721} /* (1, 13, 28) {real, imag} */,
  {32'hbde9130f, 32'h3e94af30} /* (1, 13, 27) {real, imag} */,
  {32'hbdcadbfe, 32'hbcf36c99} /* (1, 13, 26) {real, imag} */,
  {32'h3ccdf32d, 32'hbd8c258c} /* (1, 13, 25) {real, imag} */,
  {32'hbdbd3be2, 32'h3dcab50e} /* (1, 13, 24) {real, imag} */,
  {32'h3d6bc4ba, 32'h3d9d3a40} /* (1, 13, 23) {real, imag} */,
  {32'hbcf4f6c4, 32'hbcbe4c41} /* (1, 13, 22) {real, imag} */,
  {32'h3d38fd05, 32'hbcfecea8} /* (1, 13, 21) {real, imag} */,
  {32'h3cb79ad2, 32'hbdf3b1dd} /* (1, 13, 20) {real, imag} */,
  {32'h3e1cd578, 32'hbc1f0466} /* (1, 13, 19) {real, imag} */,
  {32'hbc1657fe, 32'hbd1598a9} /* (1, 13, 18) {real, imag} */,
  {32'h3aed0260, 32'h3c1e3d8e} /* (1, 13, 17) {real, imag} */,
  {32'hbce57d50, 32'h00000000} /* (1, 13, 16) {real, imag} */,
  {32'h3aed0260, 32'hbc1e3d8e} /* (1, 13, 15) {real, imag} */,
  {32'hbc1657fe, 32'h3d1598a9} /* (1, 13, 14) {real, imag} */,
  {32'h3e1cd578, 32'h3c1f0466} /* (1, 13, 13) {real, imag} */,
  {32'h3cb79ad2, 32'h3df3b1dd} /* (1, 13, 12) {real, imag} */,
  {32'h3d38fd05, 32'h3cfecea8} /* (1, 13, 11) {real, imag} */,
  {32'hbcf4f6c4, 32'h3cbe4c41} /* (1, 13, 10) {real, imag} */,
  {32'h3d6bc4ba, 32'hbd9d3a40} /* (1, 13, 9) {real, imag} */,
  {32'hbdbd3be2, 32'hbdcab50e} /* (1, 13, 8) {real, imag} */,
  {32'h3ccdf32d, 32'h3d8c258c} /* (1, 13, 7) {real, imag} */,
  {32'hbdcadbfe, 32'h3cf36c99} /* (1, 13, 6) {real, imag} */,
  {32'hbde9130f, 32'hbe94af30} /* (1, 13, 5) {real, imag} */,
  {32'h3db77749, 32'h3da41721} /* (1, 13, 4) {real, imag} */,
  {32'hbd34ee3d, 32'hbcfe7df8} /* (1, 13, 3) {real, imag} */,
  {32'hbf390aa6, 32'h3d1b1cc0} /* (1, 13, 2) {real, imag} */,
  {32'h3fcf8c97, 32'h3e8e6f30} /* (1, 13, 1) {real, imag} */,
  {32'h3f5b1b69, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'h3fa5c934, 32'hbe81e1f3} /* (1, 12, 31) {real, imag} */,
  {32'hbf2fd606, 32'h3dbeda28} /* (1, 12, 30) {real, imag} */,
  {32'h3cc93e6c, 32'h3e210d70} /* (1, 12, 29) {real, imag} */,
  {32'h3deb9b40, 32'hbe5fcfe4} /* (1, 12, 28) {real, imag} */,
  {32'hbe2b5470, 32'h3e1258f2} /* (1, 12, 27) {real, imag} */,
  {32'hbd0e38a4, 32'h3d92fadf} /* (1, 12, 26) {real, imag} */,
  {32'h3e21aa2a, 32'h3c934ef8} /* (1, 12, 25) {real, imag} */,
  {32'hbd8ef25b, 32'h3d16fb46} /* (1, 12, 24) {real, imag} */,
  {32'h3cf69656, 32'h3b658e10} /* (1, 12, 23) {real, imag} */,
  {32'h3c9ed070, 32'hbcc9b2de} /* (1, 12, 22) {real, imag} */,
  {32'h3d9a11b0, 32'h3e01b501} /* (1, 12, 21) {real, imag} */,
  {32'hbd010f75, 32'hbdc1583d} /* (1, 12, 20) {real, imag} */,
  {32'h3cb0dda2, 32'h3d5e18a9} /* (1, 12, 19) {real, imag} */,
  {32'h3be18860, 32'h3d4156cc} /* (1, 12, 18) {real, imag} */,
  {32'hbc869086, 32'h3cbf94f0} /* (1, 12, 17) {real, imag} */,
  {32'h3cad50f8, 32'h00000000} /* (1, 12, 16) {real, imag} */,
  {32'hbc869086, 32'hbcbf94f0} /* (1, 12, 15) {real, imag} */,
  {32'h3be18860, 32'hbd4156cc} /* (1, 12, 14) {real, imag} */,
  {32'h3cb0dda2, 32'hbd5e18a9} /* (1, 12, 13) {real, imag} */,
  {32'hbd010f75, 32'h3dc1583d} /* (1, 12, 12) {real, imag} */,
  {32'h3d9a11b0, 32'hbe01b501} /* (1, 12, 11) {real, imag} */,
  {32'h3c9ed070, 32'h3cc9b2de} /* (1, 12, 10) {real, imag} */,
  {32'h3cf69656, 32'hbb658e10} /* (1, 12, 9) {real, imag} */,
  {32'hbd8ef25b, 32'hbd16fb46} /* (1, 12, 8) {real, imag} */,
  {32'h3e21aa2a, 32'hbc934ef8} /* (1, 12, 7) {real, imag} */,
  {32'hbd0e38a4, 32'hbd92fadf} /* (1, 12, 6) {real, imag} */,
  {32'hbe2b5470, 32'hbe1258f2} /* (1, 12, 5) {real, imag} */,
  {32'h3deb9b40, 32'h3e5fcfe4} /* (1, 12, 4) {real, imag} */,
  {32'h3cc93e6c, 32'hbe210d70} /* (1, 12, 3) {real, imag} */,
  {32'hbf2fd606, 32'hbdbeda28} /* (1, 12, 2) {real, imag} */,
  {32'h3fa5c934, 32'h3e81e1f3} /* (1, 12, 1) {real, imag} */,
  {32'h3f563a52, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'h3f526876, 32'hbe4cab0f} /* (1, 11, 31) {real, imag} */,
  {32'hbef58278, 32'h3e17e0cc} /* (1, 11, 30) {real, imag} */,
  {32'hbd64f7a2, 32'hbd13a4ca} /* (1, 11, 29) {real, imag} */,
  {32'h3dbf4186, 32'hbe3bda64} /* (1, 11, 28) {real, imag} */,
  {32'hbd3f5f78, 32'h3c620f04} /* (1, 11, 27) {real, imag} */,
  {32'h3b9d2190, 32'h3d6ae0a8} /* (1, 11, 26) {real, imag} */,
  {32'h3d9cdc5c, 32'h3d216b2a} /* (1, 11, 25) {real, imag} */,
  {32'hbd014e7f, 32'hbd02db71} /* (1, 11, 24) {real, imag} */,
  {32'hbd9120f6, 32'hbd46dc38} /* (1, 11, 23) {real, imag} */,
  {32'h3c31b2f2, 32'h3d1a1eaa} /* (1, 11, 22) {real, imag} */,
  {32'hbd813586, 32'h3d479326} /* (1, 11, 21) {real, imag} */,
  {32'h3ddb3f2e, 32'hbd58e401} /* (1, 11, 20) {real, imag} */,
  {32'hbdb01b75, 32'h3c88c344} /* (1, 11, 19) {real, imag} */,
  {32'h3c68258b, 32'hbb01b690} /* (1, 11, 18) {real, imag} */,
  {32'h3c42f1fe, 32'hbd0903fc} /* (1, 11, 17) {real, imag} */,
  {32'hbc6d10b4, 32'h00000000} /* (1, 11, 16) {real, imag} */,
  {32'h3c42f1fe, 32'h3d0903fc} /* (1, 11, 15) {real, imag} */,
  {32'h3c68258b, 32'h3b01b690} /* (1, 11, 14) {real, imag} */,
  {32'hbdb01b75, 32'hbc88c344} /* (1, 11, 13) {real, imag} */,
  {32'h3ddb3f2e, 32'h3d58e401} /* (1, 11, 12) {real, imag} */,
  {32'hbd813586, 32'hbd479326} /* (1, 11, 11) {real, imag} */,
  {32'h3c31b2f2, 32'hbd1a1eaa} /* (1, 11, 10) {real, imag} */,
  {32'hbd9120f6, 32'h3d46dc38} /* (1, 11, 9) {real, imag} */,
  {32'hbd014e7f, 32'h3d02db71} /* (1, 11, 8) {real, imag} */,
  {32'h3d9cdc5c, 32'hbd216b2a} /* (1, 11, 7) {real, imag} */,
  {32'h3b9d2190, 32'hbd6ae0a8} /* (1, 11, 6) {real, imag} */,
  {32'hbd3f5f78, 32'hbc620f04} /* (1, 11, 5) {real, imag} */,
  {32'h3dbf4186, 32'h3e3bda64} /* (1, 11, 4) {real, imag} */,
  {32'hbd64f7a2, 32'h3d13a4ca} /* (1, 11, 3) {real, imag} */,
  {32'hbef58278, 32'hbe17e0cc} /* (1, 11, 2) {real, imag} */,
  {32'h3f526876, 32'h3e4cab0f} /* (1, 11, 1) {real, imag} */,
  {32'h3ec2300f, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'hbcf3d020, 32'h3a2a6100} /* (1, 10, 31) {real, imag} */,
  {32'h3d0a342c, 32'h3d975d78} /* (1, 10, 30) {real, imag} */,
  {32'hbb89a090, 32'hbda2b410} /* (1, 10, 29) {real, imag} */,
  {32'hbd82f9f0, 32'hbde49640} /* (1, 10, 28) {real, imag} */,
  {32'h3d64e923, 32'hbe10281a} /* (1, 10, 27) {real, imag} */,
  {32'hbdba7035, 32'hbb367e1c} /* (1, 10, 26) {real, imag} */,
  {32'h3cc7a4a4, 32'h3d6e9953} /* (1, 10, 25) {real, imag} */,
  {32'h3d1aa68e, 32'hbc1388e3} /* (1, 10, 24) {real, imag} */,
  {32'h3c426492, 32'hbc97db71} /* (1, 10, 23) {real, imag} */,
  {32'h3dcea7e7, 32'h3cfbba4e} /* (1, 10, 22) {real, imag} */,
  {32'hbd5ea1a9, 32'hbd4cc57a} /* (1, 10, 21) {real, imag} */,
  {32'h3d3120c4, 32'hbcc9a298} /* (1, 10, 20) {real, imag} */,
  {32'hbd1cd692, 32'h3da873f2} /* (1, 10, 19) {real, imag} */,
  {32'hbca2d78c, 32'hbc2fcea8} /* (1, 10, 18) {real, imag} */,
  {32'hbd09db58, 32'hbc2fd1ad} /* (1, 10, 17) {real, imag} */,
  {32'h3d8424bc, 32'h00000000} /* (1, 10, 16) {real, imag} */,
  {32'hbd09db58, 32'h3c2fd1ad} /* (1, 10, 15) {real, imag} */,
  {32'hbca2d78c, 32'h3c2fcea8} /* (1, 10, 14) {real, imag} */,
  {32'hbd1cd692, 32'hbda873f2} /* (1, 10, 13) {real, imag} */,
  {32'h3d3120c4, 32'h3cc9a298} /* (1, 10, 12) {real, imag} */,
  {32'hbd5ea1a9, 32'h3d4cc57a} /* (1, 10, 11) {real, imag} */,
  {32'h3dcea7e7, 32'hbcfbba4e} /* (1, 10, 10) {real, imag} */,
  {32'h3c426492, 32'h3c97db71} /* (1, 10, 9) {real, imag} */,
  {32'h3d1aa68e, 32'h3c1388e3} /* (1, 10, 8) {real, imag} */,
  {32'h3cc7a4a4, 32'hbd6e9953} /* (1, 10, 7) {real, imag} */,
  {32'hbdba7035, 32'h3b367e1c} /* (1, 10, 6) {real, imag} */,
  {32'h3d64e923, 32'h3e10281a} /* (1, 10, 5) {real, imag} */,
  {32'hbd82f9f0, 32'h3de49640} /* (1, 10, 4) {real, imag} */,
  {32'hbb89a090, 32'h3da2b410} /* (1, 10, 3) {real, imag} */,
  {32'h3d0a342c, 32'hbd975d78} /* (1, 10, 2) {real, imag} */,
  {32'hbcf3d020, 32'hba2a6100} /* (1, 10, 1) {real, imag} */,
  {32'hbe5e3766, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'hbf3d90c2, 32'h3e421f38} /* (1, 9, 31) {real, imag} */,
  {32'h3ec23948, 32'hbe07a6bc} /* (1, 9, 30) {real, imag} */,
  {32'hbd178059, 32'hbdc63b24} /* (1, 9, 29) {real, imag} */,
  {32'hbe222b1e, 32'hbd0c3c6e} /* (1, 9, 28) {real, imag} */,
  {32'h3e193dd6, 32'hbdd7bbe9} /* (1, 9, 27) {real, imag} */,
  {32'h3c6be4c2, 32'hbd38cc5f} /* (1, 9, 26) {real, imag} */,
  {32'hbbddf3ae, 32'h3e213d54} /* (1, 9, 25) {real, imag} */,
  {32'h3dce8a86, 32'hbe1310ec} /* (1, 9, 24) {real, imag} */,
  {32'h3d37e68a, 32'h3dc84a50} /* (1, 9, 23) {real, imag} */,
  {32'h3d1ce4d6, 32'hbcd89f9a} /* (1, 9, 22) {real, imag} */,
  {32'h3d73f2df, 32'h3c0f44e0} /* (1, 9, 21) {real, imag} */,
  {32'hbbd53020, 32'h3dd16d9c} /* (1, 9, 20) {real, imag} */,
  {32'h3ab74154, 32'h3b44093c} /* (1, 9, 19) {real, imag} */,
  {32'hbdec723d, 32'hbd6ca635} /* (1, 9, 18) {real, imag} */,
  {32'h3aec6640, 32'hbd509f06} /* (1, 9, 17) {real, imag} */,
  {32'hbced7306, 32'h00000000} /* (1, 9, 16) {real, imag} */,
  {32'h3aec6640, 32'h3d509f06} /* (1, 9, 15) {real, imag} */,
  {32'hbdec723d, 32'h3d6ca635} /* (1, 9, 14) {real, imag} */,
  {32'h3ab74154, 32'hbb44093c} /* (1, 9, 13) {real, imag} */,
  {32'hbbd53020, 32'hbdd16d9c} /* (1, 9, 12) {real, imag} */,
  {32'h3d73f2df, 32'hbc0f44e0} /* (1, 9, 11) {real, imag} */,
  {32'h3d1ce4d6, 32'h3cd89f9a} /* (1, 9, 10) {real, imag} */,
  {32'h3d37e68a, 32'hbdc84a50} /* (1, 9, 9) {real, imag} */,
  {32'h3dce8a86, 32'h3e1310ec} /* (1, 9, 8) {real, imag} */,
  {32'hbbddf3ae, 32'hbe213d54} /* (1, 9, 7) {real, imag} */,
  {32'h3c6be4c2, 32'h3d38cc5f} /* (1, 9, 6) {real, imag} */,
  {32'h3e193dd6, 32'h3dd7bbe9} /* (1, 9, 5) {real, imag} */,
  {32'hbe222b1e, 32'h3d0c3c6e} /* (1, 9, 4) {real, imag} */,
  {32'hbd178059, 32'h3dc63b24} /* (1, 9, 3) {real, imag} */,
  {32'h3ec23948, 32'h3e07a6bc} /* (1, 9, 2) {real, imag} */,
  {32'hbf3d90c2, 32'hbe421f38} /* (1, 9, 1) {real, imag} */,
  {32'hbf3f94c9, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'hbf732e91, 32'h3e8c30ac} /* (1, 8, 31) {real, imag} */,
  {32'h3f0dc88c, 32'hbe328475} /* (1, 8, 30) {real, imag} */,
  {32'hbdae6bcb, 32'hbe1aed1e} /* (1, 8, 29) {real, imag} */,
  {32'hbde1ec15, 32'hbd062be6} /* (1, 8, 28) {real, imag} */,
  {32'h3e432e04, 32'h3c4d1f48} /* (1, 8, 27) {real, imag} */,
  {32'h3d83c030, 32'hbd57185e} /* (1, 8, 26) {real, imag} */,
  {32'hbd3b83ae, 32'hbc852fb0} /* (1, 8, 25) {real, imag} */,
  {32'h3dc6359f, 32'hbd9b7096} /* (1, 8, 24) {real, imag} */,
  {32'hbc3bad50, 32'hbab5bcc0} /* (1, 8, 23) {real, imag} */,
  {32'h3d0e51b5, 32'h3d0ae782} /* (1, 8, 22) {real, imag} */,
  {32'h3de36eee, 32'hbd830649} /* (1, 8, 21) {real, imag} */,
  {32'h3d670225, 32'h3e191361} /* (1, 8, 20) {real, imag} */,
  {32'hbd6b4fb4, 32'h3d74a8cc} /* (1, 8, 19) {real, imag} */,
  {32'h3c88330a, 32'h3d665630} /* (1, 8, 18) {real, imag} */,
  {32'h3cb1fa86, 32'h3cb8b896} /* (1, 8, 17) {real, imag} */,
  {32'hbcb14df4, 32'h00000000} /* (1, 8, 16) {real, imag} */,
  {32'h3cb1fa86, 32'hbcb8b896} /* (1, 8, 15) {real, imag} */,
  {32'h3c88330a, 32'hbd665630} /* (1, 8, 14) {real, imag} */,
  {32'hbd6b4fb4, 32'hbd74a8cc} /* (1, 8, 13) {real, imag} */,
  {32'h3d670225, 32'hbe191361} /* (1, 8, 12) {real, imag} */,
  {32'h3de36eee, 32'h3d830649} /* (1, 8, 11) {real, imag} */,
  {32'h3d0e51b5, 32'hbd0ae782} /* (1, 8, 10) {real, imag} */,
  {32'hbc3bad50, 32'h3ab5bcc0} /* (1, 8, 9) {real, imag} */,
  {32'h3dc6359f, 32'h3d9b7096} /* (1, 8, 8) {real, imag} */,
  {32'hbd3b83ae, 32'h3c852fb0} /* (1, 8, 7) {real, imag} */,
  {32'h3d83c030, 32'h3d57185e} /* (1, 8, 6) {real, imag} */,
  {32'h3e432e04, 32'hbc4d1f48} /* (1, 8, 5) {real, imag} */,
  {32'hbde1ec15, 32'h3d062be6} /* (1, 8, 4) {real, imag} */,
  {32'hbdae6bcb, 32'h3e1aed1e} /* (1, 8, 3) {real, imag} */,
  {32'h3f0dc88c, 32'h3e328475} /* (1, 8, 2) {real, imag} */,
  {32'hbf732e91, 32'hbe8c30ac} /* (1, 8, 1) {real, imag} */,
  {32'hbf5e71ac, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'hbfa3aa57, 32'h3eb5fff0} /* (1, 7, 31) {real, imag} */,
  {32'h3f344bf3, 32'hbdfb8e7b} /* (1, 7, 30) {real, imag} */,
  {32'h3b99c4be, 32'hbe17e2b4} /* (1, 7, 29) {real, imag} */,
  {32'hbd6ec4fa, 32'hbe2c32e6} /* (1, 7, 28) {real, imag} */,
  {32'h3e306f01, 32'h3d880928} /* (1, 7, 27) {real, imag} */,
  {32'hbc6deb08, 32'hbd147e80} /* (1, 7, 26) {real, imag} */,
  {32'hbc2b8728, 32'hbcd10fa0} /* (1, 7, 25) {real, imag} */,
  {32'h3dfd77b6, 32'hbcc24de0} /* (1, 7, 24) {real, imag} */,
  {32'h3d5fc218, 32'hbd8ca8a7} /* (1, 7, 23) {real, imag} */,
  {32'h3d0fb492, 32'h3cae4bb1} /* (1, 7, 22) {real, imag} */,
  {32'h3e1ca136, 32'h3cc9faf8} /* (1, 7, 21) {real, imag} */,
  {32'h3d78155f, 32'hbc9e9dca} /* (1, 7, 20) {real, imag} */,
  {32'h3d4c0e5a, 32'h3d2dc515} /* (1, 7, 19) {real, imag} */,
  {32'hbc861f63, 32'h3d4ad1d9} /* (1, 7, 18) {real, imag} */,
  {32'hbd383f4e, 32'hbabe9958} /* (1, 7, 17) {real, imag} */,
  {32'hbd2b767e, 32'h00000000} /* (1, 7, 16) {real, imag} */,
  {32'hbd383f4e, 32'h3abe9958} /* (1, 7, 15) {real, imag} */,
  {32'hbc861f63, 32'hbd4ad1d9} /* (1, 7, 14) {real, imag} */,
  {32'h3d4c0e5a, 32'hbd2dc515} /* (1, 7, 13) {real, imag} */,
  {32'h3d78155f, 32'h3c9e9dca} /* (1, 7, 12) {real, imag} */,
  {32'h3e1ca136, 32'hbcc9faf8} /* (1, 7, 11) {real, imag} */,
  {32'h3d0fb492, 32'hbcae4bb1} /* (1, 7, 10) {real, imag} */,
  {32'h3d5fc218, 32'h3d8ca8a7} /* (1, 7, 9) {real, imag} */,
  {32'h3dfd77b6, 32'h3cc24de0} /* (1, 7, 8) {real, imag} */,
  {32'hbc2b8728, 32'h3cd10fa0} /* (1, 7, 7) {real, imag} */,
  {32'hbc6deb08, 32'h3d147e80} /* (1, 7, 6) {real, imag} */,
  {32'h3e306f01, 32'hbd880928} /* (1, 7, 5) {real, imag} */,
  {32'hbd6ec4fa, 32'h3e2c32e6} /* (1, 7, 4) {real, imag} */,
  {32'h3b99c4be, 32'h3e17e2b4} /* (1, 7, 3) {real, imag} */,
  {32'h3f344bf3, 32'h3dfb8e7b} /* (1, 7, 2) {real, imag} */,
  {32'hbfa3aa57, 32'hbeb5fff0} /* (1, 7, 1) {real, imag} */,
  {32'hbf86b938, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'hbf906a42, 32'h3f0bb469} /* (1, 6, 31) {real, imag} */,
  {32'h3f2b783b, 32'hbde67bf6} /* (1, 6, 30) {real, imag} */,
  {32'h3db9ff45, 32'h3a4a67c0} /* (1, 6, 29) {real, imag} */,
  {32'hbde70981, 32'hbe1917eb} /* (1, 6, 28) {real, imag} */,
  {32'h3e0bbce8, 32'hbc2b56d4} /* (1, 6, 27) {real, imag} */,
  {32'h3c1ff058, 32'h3d9455e5} /* (1, 6, 26) {real, imag} */,
  {32'hbd63756b, 32'h3df7bcb2} /* (1, 6, 25) {real, imag} */,
  {32'h3ddd333d, 32'hbe1f7e5f} /* (1, 6, 24) {real, imag} */,
  {32'hbe0b600e, 32'hbd200c0c} /* (1, 6, 23) {real, imag} */,
  {32'h3bd7d9e8, 32'h3e0c2074} /* (1, 6, 22) {real, imag} */,
  {32'hbd074a1e, 32'hbd48dfb4} /* (1, 6, 21) {real, imag} */,
  {32'hbdb45165, 32'hbb52fbb8} /* (1, 6, 20) {real, imag} */,
  {32'h3e051c58, 32'h3d86c13e} /* (1, 6, 19) {real, imag} */,
  {32'hbd5fc3ee, 32'hbdbcc82a} /* (1, 6, 18) {real, imag} */,
  {32'hbd41d39e, 32'hbc52a80a} /* (1, 6, 17) {real, imag} */,
  {32'h3dc13ec3, 32'h00000000} /* (1, 6, 16) {real, imag} */,
  {32'hbd41d39e, 32'h3c52a80a} /* (1, 6, 15) {real, imag} */,
  {32'hbd5fc3ee, 32'h3dbcc82a} /* (1, 6, 14) {real, imag} */,
  {32'h3e051c58, 32'hbd86c13e} /* (1, 6, 13) {real, imag} */,
  {32'hbdb45165, 32'h3b52fbb8} /* (1, 6, 12) {real, imag} */,
  {32'hbd074a1e, 32'h3d48dfb4} /* (1, 6, 11) {real, imag} */,
  {32'h3bd7d9e8, 32'hbe0c2074} /* (1, 6, 10) {real, imag} */,
  {32'hbe0b600e, 32'h3d200c0c} /* (1, 6, 9) {real, imag} */,
  {32'h3ddd333d, 32'h3e1f7e5f} /* (1, 6, 8) {real, imag} */,
  {32'hbd63756b, 32'hbdf7bcb2} /* (1, 6, 7) {real, imag} */,
  {32'h3c1ff058, 32'hbd9455e5} /* (1, 6, 6) {real, imag} */,
  {32'h3e0bbce8, 32'h3c2b56d4} /* (1, 6, 5) {real, imag} */,
  {32'hbde70981, 32'h3e1917eb} /* (1, 6, 4) {real, imag} */,
  {32'h3db9ff45, 32'hba4a67c0} /* (1, 6, 3) {real, imag} */,
  {32'h3f2b783b, 32'h3de67bf6} /* (1, 6, 2) {real, imag} */,
  {32'hbf906a42, 32'hbf0bb469} /* (1, 6, 1) {real, imag} */,
  {32'hbf7ce040, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'hbf60b8f4, 32'h3f7e147b} /* (1, 5, 31) {real, imag} */,
  {32'h3dd5c1c0, 32'hbe5c8d72} /* (1, 5, 30) {real, imag} */,
  {32'h3e3c1752, 32'hbcad8f5b} /* (1, 5, 29) {real, imag} */,
  {32'hbe0aa347, 32'hbcf4eb60} /* (1, 5, 28) {real, imag} */,
  {32'h3e3f2a7a, 32'hbd2c07e7} /* (1, 5, 27) {real, imag} */,
  {32'hbbf57820, 32'hbbad5f00} /* (1, 5, 26) {real, imag} */,
  {32'hbbb7a578, 32'h3df47826} /* (1, 5, 25) {real, imag} */,
  {32'h3e2c48d4, 32'hbd652ff5} /* (1, 5, 24) {real, imag} */,
  {32'hbd40aaac, 32'hbd7d6e89} /* (1, 5, 23) {real, imag} */,
  {32'hbd0ba544, 32'hbcf908d7} /* (1, 5, 22) {real, imag} */,
  {32'h3cef9650, 32'h3cc7fa57} /* (1, 5, 21) {real, imag} */,
  {32'h3d116a47, 32'h3ce8781a} /* (1, 5, 20) {real, imag} */,
  {32'h3d7026d0, 32'h3ca87a42} /* (1, 5, 19) {real, imag} */,
  {32'h3d5d5842, 32'hbdbbd289} /* (1, 5, 18) {real, imag} */,
  {32'hbd3cc4a6, 32'h3cf26377} /* (1, 5, 17) {real, imag} */,
  {32'hbd80deb2, 32'h00000000} /* (1, 5, 16) {real, imag} */,
  {32'hbd3cc4a6, 32'hbcf26377} /* (1, 5, 15) {real, imag} */,
  {32'h3d5d5842, 32'h3dbbd289} /* (1, 5, 14) {real, imag} */,
  {32'h3d7026d0, 32'hbca87a42} /* (1, 5, 13) {real, imag} */,
  {32'h3d116a47, 32'hbce8781a} /* (1, 5, 12) {real, imag} */,
  {32'h3cef9650, 32'hbcc7fa57} /* (1, 5, 11) {real, imag} */,
  {32'hbd0ba544, 32'h3cf908d7} /* (1, 5, 10) {real, imag} */,
  {32'hbd40aaac, 32'h3d7d6e89} /* (1, 5, 9) {real, imag} */,
  {32'h3e2c48d4, 32'h3d652ff5} /* (1, 5, 8) {real, imag} */,
  {32'hbbb7a578, 32'hbdf47826} /* (1, 5, 7) {real, imag} */,
  {32'hbbf57820, 32'h3bad5f00} /* (1, 5, 6) {real, imag} */,
  {32'h3e3f2a7a, 32'h3d2c07e7} /* (1, 5, 5) {real, imag} */,
  {32'hbe0aa347, 32'h3cf4eb60} /* (1, 5, 4) {real, imag} */,
  {32'h3e3c1752, 32'h3cad8f5b} /* (1, 5, 3) {real, imag} */,
  {32'h3dd5c1c0, 32'h3e5c8d72} /* (1, 5, 2) {real, imag} */,
  {32'hbf60b8f4, 32'hbf7e147b} /* (1, 5, 1) {real, imag} */,
  {32'hbf95a8fc, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'hbf462304, 32'h3fa25e3c} /* (1, 4, 31) {real, imag} */,
  {32'hbe896f0c, 32'hbe8c3bc5} /* (1, 4, 30) {real, imag} */,
  {32'h3e5f5c22, 32'hbe0f3ec1} /* (1, 4, 29) {real, imag} */,
  {32'h3ac96780, 32'hbe6e66c3} /* (1, 4, 28) {real, imag} */,
  {32'h3da9a29a, 32'h3cc5fc44} /* (1, 4, 27) {real, imag} */,
  {32'h3d2e4f31, 32'hbb0a9d50} /* (1, 4, 26) {real, imag} */,
  {32'h3da8ee32, 32'hbc125978} /* (1, 4, 25) {real, imag} */,
  {32'hbd4b99c9, 32'hbc84b836} /* (1, 4, 24) {real, imag} */,
  {32'h3db534b2, 32'h3b988c5c} /* (1, 4, 23) {real, imag} */,
  {32'hbc4a8dee, 32'hbd7dc711} /* (1, 4, 22) {real, imag} */,
  {32'h3d731bc1, 32'h3d877d07} /* (1, 4, 21) {real, imag} */,
  {32'h3b582142, 32'hbd0290ab} /* (1, 4, 20) {real, imag} */,
  {32'hbd12b90a, 32'hbd0f7ba6} /* (1, 4, 19) {real, imag} */,
  {32'h3d890c95, 32'h3c83277f} /* (1, 4, 18) {real, imag} */,
  {32'h3d06458d, 32'h3cdc0fff} /* (1, 4, 17) {real, imag} */,
  {32'h3ce35905, 32'h00000000} /* (1, 4, 16) {real, imag} */,
  {32'h3d06458d, 32'hbcdc0fff} /* (1, 4, 15) {real, imag} */,
  {32'h3d890c95, 32'hbc83277f} /* (1, 4, 14) {real, imag} */,
  {32'hbd12b90a, 32'h3d0f7ba6} /* (1, 4, 13) {real, imag} */,
  {32'h3b582142, 32'h3d0290ab} /* (1, 4, 12) {real, imag} */,
  {32'h3d731bc1, 32'hbd877d07} /* (1, 4, 11) {real, imag} */,
  {32'hbc4a8dee, 32'h3d7dc711} /* (1, 4, 10) {real, imag} */,
  {32'h3db534b2, 32'hbb988c5c} /* (1, 4, 9) {real, imag} */,
  {32'hbd4b99c9, 32'h3c84b836} /* (1, 4, 8) {real, imag} */,
  {32'h3da8ee32, 32'h3c125978} /* (1, 4, 7) {real, imag} */,
  {32'h3d2e4f31, 32'h3b0a9d50} /* (1, 4, 6) {real, imag} */,
  {32'h3da9a29a, 32'hbcc5fc44} /* (1, 4, 5) {real, imag} */,
  {32'h3ac96780, 32'h3e6e66c3} /* (1, 4, 4) {real, imag} */,
  {32'h3e5f5c22, 32'h3e0f3ec1} /* (1, 4, 3) {real, imag} */,
  {32'hbe896f0c, 32'h3e8c3bc5} /* (1, 4, 2) {real, imag} */,
  {32'hbf462304, 32'hbfa25e3c} /* (1, 4, 1) {real, imag} */,
  {32'hbf9f4694, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hbf2af1c2, 32'h3fb1a81e} /* (1, 3, 31) {real, imag} */,
  {32'hbe81fe95, 32'hbeff2a62} /* (1, 3, 30) {real, imag} */,
  {32'h3e8563eb, 32'h3b559710} /* (1, 3, 29) {real, imag} */,
  {32'h3d5f15e6, 32'hbe254ecf} /* (1, 3, 28) {real, imag} */,
  {32'h3d56d51a, 32'h3e295118} /* (1, 3, 27) {real, imag} */,
  {32'h3dd57b12, 32'hbd3cc858} /* (1, 3, 26) {real, imag} */,
  {32'hbd3c365c, 32'h3c4537fc} /* (1, 3, 25) {real, imag} */,
  {32'hbcc7c8a8, 32'h3cea140e} /* (1, 3, 24) {real, imag} */,
  {32'h3db1407c, 32'hbd865de2} /* (1, 3, 23) {real, imag} */,
  {32'h3d66cc1e, 32'h3d81ab5f} /* (1, 3, 22) {real, imag} */,
  {32'hbd90de06, 32'h3ca3dfb4} /* (1, 3, 21) {real, imag} */,
  {32'hbde664a0, 32'h3c05500c} /* (1, 3, 20) {real, imag} */,
  {32'hbb961ce0, 32'h3c8b91f2} /* (1, 3, 19) {real, imag} */,
  {32'hbcff5bf8, 32'hbd435aee} /* (1, 3, 18) {real, imag} */,
  {32'h3c5b1c83, 32'hbc94abd8} /* (1, 3, 17) {real, imag} */,
  {32'h3d7e5f7d, 32'h00000000} /* (1, 3, 16) {real, imag} */,
  {32'h3c5b1c83, 32'h3c94abd8} /* (1, 3, 15) {real, imag} */,
  {32'hbcff5bf8, 32'h3d435aee} /* (1, 3, 14) {real, imag} */,
  {32'hbb961ce0, 32'hbc8b91f2} /* (1, 3, 13) {real, imag} */,
  {32'hbde664a0, 32'hbc05500c} /* (1, 3, 12) {real, imag} */,
  {32'hbd90de06, 32'hbca3dfb4} /* (1, 3, 11) {real, imag} */,
  {32'h3d66cc1e, 32'hbd81ab5f} /* (1, 3, 10) {real, imag} */,
  {32'h3db1407c, 32'h3d865de2} /* (1, 3, 9) {real, imag} */,
  {32'hbcc7c8a8, 32'hbcea140e} /* (1, 3, 8) {real, imag} */,
  {32'hbd3c365c, 32'hbc4537fc} /* (1, 3, 7) {real, imag} */,
  {32'h3dd57b12, 32'h3d3cc858} /* (1, 3, 6) {real, imag} */,
  {32'h3d56d51a, 32'hbe295118} /* (1, 3, 5) {real, imag} */,
  {32'h3d5f15e6, 32'h3e254ecf} /* (1, 3, 4) {real, imag} */,
  {32'h3e8563eb, 32'hbb559710} /* (1, 3, 3) {real, imag} */,
  {32'hbe81fe95, 32'h3eff2a62} /* (1, 3, 2) {real, imag} */,
  {32'hbf2af1c2, 32'hbfb1a81e} /* (1, 3, 1) {real, imag} */,
  {32'hbf90a92e, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hbf65c8b5, 32'h3fa92c60} /* (1, 2, 31) {real, imag} */,
  {32'hbeebb10a, 32'hbf0fb3a0} /* (1, 2, 30) {real, imag} */,
  {32'h3e81f710, 32'h3d12f3ef} /* (1, 2, 29) {real, imag} */,
  {32'h3b0e2ba0, 32'hbe80db88} /* (1, 2, 28) {real, imag} */,
  {32'h3e34d18c, 32'h3db631f6} /* (1, 2, 27) {real, imag} */,
  {32'h3b257a10, 32'hbd4680fe} /* (1, 2, 26) {real, imag} */,
  {32'hbd04fc1f, 32'h3c9a7bae} /* (1, 2, 25) {real, imag} */,
  {32'hbdcf7467, 32'h39e47f80} /* (1, 2, 24) {real, imag} */,
  {32'hbe219510, 32'hbe07a5d8} /* (1, 2, 23) {real, imag} */,
  {32'h3dabd29e, 32'hbd4d394e} /* (1, 2, 22) {real, imag} */,
  {32'h3dc93eac, 32'hbc224534} /* (1, 2, 21) {real, imag} */,
  {32'h3de1eb50, 32'hbd91069a} /* (1, 2, 20) {real, imag} */,
  {32'hbc6215e6, 32'h3b4f385c} /* (1, 2, 19) {real, imag} */,
  {32'hbd95a670, 32'hbdee53c9} /* (1, 2, 18) {real, imag} */,
  {32'h3cf1354c, 32'hbcb61fea} /* (1, 2, 17) {real, imag} */,
  {32'hbc1d5804, 32'h00000000} /* (1, 2, 16) {real, imag} */,
  {32'h3cf1354c, 32'h3cb61fea} /* (1, 2, 15) {real, imag} */,
  {32'hbd95a670, 32'h3dee53c9} /* (1, 2, 14) {real, imag} */,
  {32'hbc6215e6, 32'hbb4f385c} /* (1, 2, 13) {real, imag} */,
  {32'h3de1eb50, 32'h3d91069a} /* (1, 2, 12) {real, imag} */,
  {32'h3dc93eac, 32'h3c224534} /* (1, 2, 11) {real, imag} */,
  {32'h3dabd29e, 32'h3d4d394e} /* (1, 2, 10) {real, imag} */,
  {32'hbe219510, 32'h3e07a5d8} /* (1, 2, 9) {real, imag} */,
  {32'hbdcf7467, 32'hb9e47f80} /* (1, 2, 8) {real, imag} */,
  {32'hbd04fc1f, 32'hbc9a7bae} /* (1, 2, 7) {real, imag} */,
  {32'h3b257a10, 32'h3d4680fe} /* (1, 2, 6) {real, imag} */,
  {32'h3e34d18c, 32'hbdb631f6} /* (1, 2, 5) {real, imag} */,
  {32'h3b0e2ba0, 32'h3e80db88} /* (1, 2, 4) {real, imag} */,
  {32'h3e81f710, 32'hbd12f3ef} /* (1, 2, 3) {real, imag} */,
  {32'hbeebb10a, 32'h3f0fb3a0} /* (1, 2, 2) {real, imag} */,
  {32'hbf65c8b5, 32'hbfa92c60} /* (1, 2, 1) {real, imag} */,
  {32'hbf6e94e9, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hbf5a7438, 32'h3f8d5d3a} /* (1, 1, 31) {real, imag} */,
  {32'hbeaaea9c, 32'hbf236a54} /* (1, 1, 30) {real, imag} */,
  {32'h3e6eb8da, 32'hbcf57be9} /* (1, 1, 29) {real, imag} */,
  {32'h3d01b0ca, 32'hbe72e8ce} /* (1, 1, 28) {real, imag} */,
  {32'h3e8628cc, 32'h3e42b51a} /* (1, 1, 27) {real, imag} */,
  {32'h3d06682e, 32'h3dc483f8} /* (1, 1, 26) {real, imag} */,
  {32'hbd866f60, 32'h3cfbf318} /* (1, 1, 25) {real, imag} */,
  {32'hbd806a02, 32'h3ce2573a} /* (1, 1, 24) {real, imag} */,
  {32'hbd6815f2, 32'hbdcc8220} /* (1, 1, 23) {real, imag} */,
  {32'h3b0ae480, 32'hbd725a9b} /* (1, 1, 22) {real, imag} */,
  {32'h3c3a61d4, 32'hbd88e3fb} /* (1, 1, 21) {real, imag} */,
  {32'h3daadc4d, 32'h3cb69f19} /* (1, 1, 20) {real, imag} */,
  {32'h3c638184, 32'h3b84d8b0} /* (1, 1, 19) {real, imag} */,
  {32'hbbf68a82, 32'h3af251d0} /* (1, 1, 18) {real, imag} */,
  {32'h3a8168e0, 32'h3d1e676e} /* (1, 1, 17) {real, imag} */,
  {32'hbdcafe9e, 32'h00000000} /* (1, 1, 16) {real, imag} */,
  {32'h3a8168e0, 32'hbd1e676e} /* (1, 1, 15) {real, imag} */,
  {32'hbbf68a82, 32'hbaf251d0} /* (1, 1, 14) {real, imag} */,
  {32'h3c638184, 32'hbb84d8b0} /* (1, 1, 13) {real, imag} */,
  {32'h3daadc4d, 32'hbcb69f19} /* (1, 1, 12) {real, imag} */,
  {32'h3c3a61d4, 32'h3d88e3fb} /* (1, 1, 11) {real, imag} */,
  {32'h3b0ae480, 32'h3d725a9b} /* (1, 1, 10) {real, imag} */,
  {32'hbd6815f2, 32'h3dcc8220} /* (1, 1, 9) {real, imag} */,
  {32'hbd806a02, 32'hbce2573a} /* (1, 1, 8) {real, imag} */,
  {32'hbd866f60, 32'hbcfbf318} /* (1, 1, 7) {real, imag} */,
  {32'h3d06682e, 32'hbdc483f8} /* (1, 1, 6) {real, imag} */,
  {32'h3e8628cc, 32'hbe42b51a} /* (1, 1, 5) {real, imag} */,
  {32'h3d01b0ca, 32'h3e72e8ce} /* (1, 1, 4) {real, imag} */,
  {32'h3e6eb8da, 32'h3cf57be9} /* (1, 1, 3) {real, imag} */,
  {32'hbeaaea9c, 32'h3f236a54} /* (1, 1, 2) {real, imag} */,
  {32'hbf5a7438, 32'hbf8d5d3a} /* (1, 1, 1) {real, imag} */,
  {32'hbf1b44da, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hbf39d1e3, 32'h3f3c5560} /* (1, 0, 31) {real, imag} */,
  {32'hbdea4aa0, 32'hbed59685} /* (1, 0, 30) {real, imag} */,
  {32'h3d5e0f24, 32'hbd5b6ffc} /* (1, 0, 29) {real, imag} */,
  {32'h3a07f300, 32'hbdcb3860} /* (1, 0, 28) {real, imag} */,
  {32'h3de6bf5a, 32'h3d2a7042} /* (1, 0, 27) {real, imag} */,
  {32'h3c207f60, 32'hbd5eaa06} /* (1, 0, 26) {real, imag} */,
  {32'hbd8d7372, 32'h3d758db3} /* (1, 0, 25) {real, imag} */,
  {32'h3ca1a23e, 32'h3d57197c} /* (1, 0, 24) {real, imag} */,
  {32'h3de50854, 32'hbdee28ce} /* (1, 0, 23) {real, imag} */,
  {32'hbd2fad34, 32'h3d7f15ff} /* (1, 0, 22) {real, imag} */,
  {32'hbd3755c6, 32'h3d564520} /* (1, 0, 21) {real, imag} */,
  {32'h3b20b670, 32'h3cde09fd} /* (1, 0, 20) {real, imag} */,
  {32'h3c124aa8, 32'hbd729dd9} /* (1, 0, 19) {real, imag} */,
  {32'hbcaaabd4, 32'h3accd848} /* (1, 0, 18) {real, imag} */,
  {32'h3c977076, 32'h3c3518e1} /* (1, 0, 17) {real, imag} */,
  {32'h3c8ca216, 32'h00000000} /* (1, 0, 16) {real, imag} */,
  {32'h3c977076, 32'hbc3518e1} /* (1, 0, 15) {real, imag} */,
  {32'hbcaaabd4, 32'hbaccd848} /* (1, 0, 14) {real, imag} */,
  {32'h3c124aa8, 32'h3d729dd9} /* (1, 0, 13) {real, imag} */,
  {32'h3b20b670, 32'hbcde09fd} /* (1, 0, 12) {real, imag} */,
  {32'hbd3755c6, 32'hbd564520} /* (1, 0, 11) {real, imag} */,
  {32'hbd2fad34, 32'hbd7f15ff} /* (1, 0, 10) {real, imag} */,
  {32'h3de50854, 32'h3dee28ce} /* (1, 0, 9) {real, imag} */,
  {32'h3ca1a23e, 32'hbd57197c} /* (1, 0, 8) {real, imag} */,
  {32'hbd8d7372, 32'hbd758db3} /* (1, 0, 7) {real, imag} */,
  {32'h3c207f60, 32'h3d5eaa06} /* (1, 0, 6) {real, imag} */,
  {32'h3de6bf5a, 32'hbd2a7042} /* (1, 0, 5) {real, imag} */,
  {32'h3a07f300, 32'h3dcb3860} /* (1, 0, 4) {real, imag} */,
  {32'h3d5e0f24, 32'h3d5b6ffc} /* (1, 0, 3) {real, imag} */,
  {32'hbdea4aa0, 32'h3ed59685} /* (1, 0, 2) {real, imag} */,
  {32'hbf39d1e3, 32'hbf3c5560} /* (1, 0, 1) {real, imag} */,
  {32'hbeec9a39, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hbec7693c, 32'h3e1c1ee2} /* (0, 31, 31) {real, imag} */,
  {32'hbb07d080, 32'hbcf251bc} /* (0, 31, 30) {real, imag} */,
  {32'h3ded8fce, 32'h3d74e5df} /* (0, 31, 29) {real, imag} */,
  {32'h3d8a77aa, 32'h3cb4377c} /* (0, 31, 28) {real, imag} */,
  {32'h3ded7b1e, 32'hbc26e4fa} /* (0, 31, 27) {real, imag} */,
  {32'h3c97f6ee, 32'hbd9f0477} /* (0, 31, 26) {real, imag} */,
  {32'hbd290855, 32'hbc0af7d8} /* (0, 31, 25) {real, imag} */,
  {32'hbd911129, 32'hbd502d4f} /* (0, 31, 24) {real, imag} */,
  {32'hbce4010a, 32'hbcb7c129} /* (0, 31, 23) {real, imag} */,
  {32'hbd41b0d7, 32'h3d4f5c56} /* (0, 31, 22) {real, imag} */,
  {32'hbbb5c2ac, 32'h3c749336} /* (0, 31, 21) {real, imag} */,
  {32'h3cd40672, 32'h3d458a7c} /* (0, 31, 20) {real, imag} */,
  {32'hbb1812e0, 32'hbcec5e0f} /* (0, 31, 19) {real, imag} */,
  {32'h3c8e0bf6, 32'hbc82e8a4} /* (0, 31, 18) {real, imag} */,
  {32'h3b793ce0, 32'hb9a3be80} /* (0, 31, 17) {real, imag} */,
  {32'hbc082c30, 32'h00000000} /* (0, 31, 16) {real, imag} */,
  {32'h3b793ce0, 32'h39a3be80} /* (0, 31, 15) {real, imag} */,
  {32'h3c8e0bf6, 32'h3c82e8a4} /* (0, 31, 14) {real, imag} */,
  {32'hbb1812e0, 32'h3cec5e0f} /* (0, 31, 13) {real, imag} */,
  {32'h3cd40672, 32'hbd458a7c} /* (0, 31, 12) {real, imag} */,
  {32'hbbb5c2ac, 32'hbc749336} /* (0, 31, 11) {real, imag} */,
  {32'hbd41b0d7, 32'hbd4f5c56} /* (0, 31, 10) {real, imag} */,
  {32'hbce4010a, 32'h3cb7c129} /* (0, 31, 9) {real, imag} */,
  {32'hbd911129, 32'h3d502d4f} /* (0, 31, 8) {real, imag} */,
  {32'hbd290855, 32'h3c0af7d8} /* (0, 31, 7) {real, imag} */,
  {32'h3c97f6ee, 32'h3d9f0477} /* (0, 31, 6) {real, imag} */,
  {32'h3ded7b1e, 32'h3c26e4fa} /* (0, 31, 5) {real, imag} */,
  {32'h3d8a77aa, 32'hbcb4377c} /* (0, 31, 4) {real, imag} */,
  {32'h3ded8fce, 32'hbd74e5df} /* (0, 31, 3) {real, imag} */,
  {32'hbb07d080, 32'h3cf251bc} /* (0, 31, 2) {real, imag} */,
  {32'hbec7693c, 32'hbe1c1ee2} /* (0, 31, 1) {real, imag} */,
  {32'hbe9199ed, 32'h00000000} /* (0, 31, 0) {real, imag} */,
  {32'hbf01f914, 32'h3d2fa970} /* (0, 30, 31) {real, imag} */,
  {32'h3e2d56bd, 32'hbc9a74c4} /* (0, 30, 30) {real, imag} */,
  {32'h3dcf9ffc, 32'hbca9842e} /* (0, 30, 29) {real, imag} */,
  {32'h3dabca0c, 32'h3cf4cf7e} /* (0, 30, 28) {real, imag} */,
  {32'h3dced7b0, 32'h3d2bce3e} /* (0, 30, 27) {real, imag} */,
  {32'h3d6c35b3, 32'hbd12b3e2} /* (0, 30, 26) {real, imag} */,
  {32'hbd85a5ae, 32'h3c2277d0} /* (0, 30, 25) {real, imag} */,
  {32'hbd1433b8, 32'h3c8238dc} /* (0, 30, 24) {real, imag} */,
  {32'hbd24fcf6, 32'h3d30fb17} /* (0, 30, 23) {real, imag} */,
  {32'h3d762d8c, 32'h3d85f620} /* (0, 30, 22) {real, imag} */,
  {32'h3cdfd5a3, 32'h3cd101f0} /* (0, 30, 21) {real, imag} */,
  {32'h3a966f48, 32'h3ddadf9c} /* (0, 30, 20) {real, imag} */,
  {32'hbcbd8169, 32'h3c4ea566} /* (0, 30, 19) {real, imag} */,
  {32'h3d0479e1, 32'h3bda2e28} /* (0, 30, 18) {real, imag} */,
  {32'h3bce6c30, 32'h3c6c23f2} /* (0, 30, 17) {real, imag} */,
  {32'h3cad90a7, 32'h00000000} /* (0, 30, 16) {real, imag} */,
  {32'h3bce6c30, 32'hbc6c23f2} /* (0, 30, 15) {real, imag} */,
  {32'h3d0479e1, 32'hbbda2e28} /* (0, 30, 14) {real, imag} */,
  {32'hbcbd8169, 32'hbc4ea566} /* (0, 30, 13) {real, imag} */,
  {32'h3a966f48, 32'hbddadf9c} /* (0, 30, 12) {real, imag} */,
  {32'h3cdfd5a3, 32'hbcd101f0} /* (0, 30, 11) {real, imag} */,
  {32'h3d762d8c, 32'hbd85f620} /* (0, 30, 10) {real, imag} */,
  {32'hbd24fcf6, 32'hbd30fb17} /* (0, 30, 9) {real, imag} */,
  {32'hbd1433b8, 32'hbc8238dc} /* (0, 30, 8) {real, imag} */,
  {32'hbd85a5ae, 32'hbc2277d0} /* (0, 30, 7) {real, imag} */,
  {32'h3d6c35b3, 32'h3d12b3e2} /* (0, 30, 6) {real, imag} */,
  {32'h3dced7b0, 32'hbd2bce3e} /* (0, 30, 5) {real, imag} */,
  {32'h3dabca0c, 32'hbcf4cf7e} /* (0, 30, 4) {real, imag} */,
  {32'h3dcf9ffc, 32'h3ca9842e} /* (0, 30, 3) {real, imag} */,
  {32'h3e2d56bd, 32'h3c9a74c4} /* (0, 30, 2) {real, imag} */,
  {32'hbf01f914, 32'hbd2fa970} /* (0, 30, 1) {real, imag} */,
  {32'hbec59b17, 32'h00000000} /* (0, 30, 0) {real, imag} */,
  {32'hbf1fb971, 32'h3d0cbcc0} /* (0, 29, 31) {real, imag} */,
  {32'h3e8eccbc, 32'hbd25f8b6} /* (0, 29, 30) {real, imag} */,
  {32'h3ccc8f7c, 32'h3d1ecc6e} /* (0, 29, 29) {real, imag} */,
  {32'hbd08d5b2, 32'h3d21ed47} /* (0, 29, 28) {real, imag} */,
  {32'h3d6b195e, 32'h39030c00} /* (0, 29, 27) {real, imag} */,
  {32'h3d674c56, 32'h3cf79e71} /* (0, 29, 26) {real, imag} */,
  {32'hbd297c0f, 32'hbd21bbec} /* (0, 29, 25) {real, imag} */,
  {32'h38f12800, 32'hbc179292} /* (0, 29, 24) {real, imag} */,
  {32'hbb10c63c, 32'h3c659160} /* (0, 29, 23) {real, imag} */,
  {32'hbca32771, 32'h3db024e7} /* (0, 29, 22) {real, imag} */,
  {32'hbbecb038, 32'hbc88d813} /* (0, 29, 21) {real, imag} */,
  {32'h3cf655fa, 32'h3da8dd5a} /* (0, 29, 20) {real, imag} */,
  {32'hbc5769e4, 32'h3d2b09f4} /* (0, 29, 19) {real, imag} */,
  {32'h3c9f2260, 32'hbc7e1d0a} /* (0, 29, 18) {real, imag} */,
  {32'hbc807490, 32'hbaedd800} /* (0, 29, 17) {real, imag} */,
  {32'h3d2363c4, 32'h00000000} /* (0, 29, 16) {real, imag} */,
  {32'hbc807490, 32'h3aedd800} /* (0, 29, 15) {real, imag} */,
  {32'h3c9f2260, 32'h3c7e1d0a} /* (0, 29, 14) {real, imag} */,
  {32'hbc5769e4, 32'hbd2b09f4} /* (0, 29, 13) {real, imag} */,
  {32'h3cf655fa, 32'hbda8dd5a} /* (0, 29, 12) {real, imag} */,
  {32'hbbecb038, 32'h3c88d813} /* (0, 29, 11) {real, imag} */,
  {32'hbca32771, 32'hbdb024e7} /* (0, 29, 10) {real, imag} */,
  {32'hbb10c63c, 32'hbc659160} /* (0, 29, 9) {real, imag} */,
  {32'h38f12800, 32'h3c179292} /* (0, 29, 8) {real, imag} */,
  {32'hbd297c0f, 32'h3d21bbec} /* (0, 29, 7) {real, imag} */,
  {32'h3d674c56, 32'hbcf79e71} /* (0, 29, 6) {real, imag} */,
  {32'h3d6b195e, 32'hb9030c00} /* (0, 29, 5) {real, imag} */,
  {32'hbd08d5b2, 32'hbd21ed47} /* (0, 29, 4) {real, imag} */,
  {32'h3ccc8f7c, 32'hbd1ecc6e} /* (0, 29, 3) {real, imag} */,
  {32'h3e8eccbc, 32'h3d25f8b6} /* (0, 29, 2) {real, imag} */,
  {32'hbf1fb971, 32'hbd0cbcc0} /* (0, 29, 1) {real, imag} */,
  {32'hbec1ca78, 32'h00000000} /* (0, 29, 0) {real, imag} */,
  {32'hbf325e9e, 32'hbc2a2c80} /* (0, 28, 31) {real, imag} */,
  {32'h3e519199, 32'h3c21866c} /* (0, 28, 30) {real, imag} */,
  {32'h3b53b670, 32'h3b729570} /* (0, 28, 29) {real, imag} */,
  {32'hbd4e88e3, 32'h3dfaf8d9} /* (0, 28, 28) {real, imag} */,
  {32'h3e2dd147, 32'hbd39116e} /* (0, 28, 27) {real, imag} */,
  {32'h3a896008, 32'h3d2c43b0} /* (0, 28, 26) {real, imag} */,
  {32'hbcc4acaa, 32'hbc16ddcf} /* (0, 28, 25) {real, imag} */,
  {32'h3d22fe04, 32'hbdcdda7b} /* (0, 28, 24) {real, imag} */,
  {32'hbaf97960, 32'hbae1cd54} /* (0, 28, 23) {real, imag} */,
  {32'hbcb55427, 32'h3c29972d} /* (0, 28, 22) {real, imag} */,
  {32'hbcc86dd0, 32'h3d76e3ea} /* (0, 28, 21) {real, imag} */,
  {32'hba1ef610, 32'h3d29b12c} /* (0, 28, 20) {real, imag} */,
  {32'hbc9ff3ae, 32'hbd48e538} /* (0, 28, 19) {real, imag} */,
  {32'h3c248dd8, 32'hbd6f3a6d} /* (0, 28, 18) {real, imag} */,
  {32'hbc253012, 32'hbc51f96a} /* (0, 28, 17) {real, imag} */,
  {32'h3bab76ae, 32'h00000000} /* (0, 28, 16) {real, imag} */,
  {32'hbc253012, 32'h3c51f96a} /* (0, 28, 15) {real, imag} */,
  {32'h3c248dd8, 32'h3d6f3a6d} /* (0, 28, 14) {real, imag} */,
  {32'hbc9ff3ae, 32'h3d48e538} /* (0, 28, 13) {real, imag} */,
  {32'hba1ef610, 32'hbd29b12c} /* (0, 28, 12) {real, imag} */,
  {32'hbcc86dd0, 32'hbd76e3ea} /* (0, 28, 11) {real, imag} */,
  {32'hbcb55427, 32'hbc29972d} /* (0, 28, 10) {real, imag} */,
  {32'hbaf97960, 32'h3ae1cd54} /* (0, 28, 9) {real, imag} */,
  {32'h3d22fe04, 32'h3dcdda7b} /* (0, 28, 8) {real, imag} */,
  {32'hbcc4acaa, 32'h3c16ddcf} /* (0, 28, 7) {real, imag} */,
  {32'h3a896008, 32'hbd2c43b0} /* (0, 28, 6) {real, imag} */,
  {32'h3e2dd147, 32'h3d39116e} /* (0, 28, 5) {real, imag} */,
  {32'hbd4e88e3, 32'hbdfaf8d9} /* (0, 28, 4) {real, imag} */,
  {32'h3b53b670, 32'hbb729570} /* (0, 28, 3) {real, imag} */,
  {32'h3e519199, 32'hbc21866c} /* (0, 28, 2) {real, imag} */,
  {32'hbf325e9e, 32'h3c2a2c80} /* (0, 28, 1) {real, imag} */,
  {32'hbe915680, 32'h00000000} /* (0, 28, 0) {real, imag} */,
  {32'hbf2b8939, 32'h3d8acae0} /* (0, 27, 31) {real, imag} */,
  {32'h3e3a8d1e, 32'h3d6d0a00} /* (0, 27, 30) {real, imag} */,
  {32'h3bddf218, 32'hbd6adaf9} /* (0, 27, 29) {real, imag} */,
  {32'hbcb6bdd2, 32'h3e0155ba} /* (0, 27, 28) {real, imag} */,
  {32'h3db51949, 32'hbceb3028} /* (0, 27, 27) {real, imag} */,
  {32'h3c10ff94, 32'h3c90e5d2} /* (0, 27, 26) {real, imag} */,
  {32'hbd468046, 32'hbc8b9926} /* (0, 27, 25) {real, imag} */,
  {32'hbbe8fc76, 32'h3bb3a2bc} /* (0, 27, 24) {real, imag} */,
  {32'h3c7ce8c4, 32'hbdae8e96} /* (0, 27, 23) {real, imag} */,
  {32'hbd4eab14, 32'hbb7a0c00} /* (0, 27, 22) {real, imag} */,
  {32'h3d50ba80, 32'hbb18ef00} /* (0, 27, 21) {real, imag} */,
  {32'hbc98ad5a, 32'h3b0efaa0} /* (0, 27, 20) {real, imag} */,
  {32'h3cc31608, 32'hbcc6d1b6} /* (0, 27, 19) {real, imag} */,
  {32'hbaeebd20, 32'hbd1c57bd} /* (0, 27, 18) {real, imag} */,
  {32'hbbbf58fe, 32'h3d0bf8e4} /* (0, 27, 17) {real, imag} */,
  {32'hbda084a2, 32'h00000000} /* (0, 27, 16) {real, imag} */,
  {32'hbbbf58fe, 32'hbd0bf8e4} /* (0, 27, 15) {real, imag} */,
  {32'hbaeebd20, 32'h3d1c57bd} /* (0, 27, 14) {real, imag} */,
  {32'h3cc31608, 32'h3cc6d1b6} /* (0, 27, 13) {real, imag} */,
  {32'hbc98ad5a, 32'hbb0efaa0} /* (0, 27, 12) {real, imag} */,
  {32'h3d50ba80, 32'h3b18ef00} /* (0, 27, 11) {real, imag} */,
  {32'hbd4eab14, 32'h3b7a0c00} /* (0, 27, 10) {real, imag} */,
  {32'h3c7ce8c4, 32'h3dae8e96} /* (0, 27, 9) {real, imag} */,
  {32'hbbe8fc76, 32'hbbb3a2bc} /* (0, 27, 8) {real, imag} */,
  {32'hbd468046, 32'h3c8b9926} /* (0, 27, 7) {real, imag} */,
  {32'h3c10ff94, 32'hbc90e5d2} /* (0, 27, 6) {real, imag} */,
  {32'h3db51949, 32'h3ceb3028} /* (0, 27, 5) {real, imag} */,
  {32'hbcb6bdd2, 32'hbe0155ba} /* (0, 27, 4) {real, imag} */,
  {32'h3bddf218, 32'h3d6adaf9} /* (0, 27, 3) {real, imag} */,
  {32'h3e3a8d1e, 32'hbd6d0a00} /* (0, 27, 2) {real, imag} */,
  {32'hbf2b8939, 32'hbd8acae0} /* (0, 27, 1) {real, imag} */,
  {32'hbe88f38b, 32'h00000000} /* (0, 27, 0) {real, imag} */,
  {32'hbf496816, 32'h3d7bd300} /* (0, 26, 31) {real, imag} */,
  {32'h3e3c427b, 32'h3daec14d} /* (0, 26, 30) {real, imag} */,
  {32'hbd12b92c, 32'hbd29c27f} /* (0, 26, 29) {real, imag} */,
  {32'hbdfa53e6, 32'h3de19571} /* (0, 26, 28) {real, imag} */,
  {32'h3e11c5c2, 32'hbd0018cf} /* (0, 26, 27) {real, imag} */,
  {32'h3cca84b3, 32'hbba2f3c0} /* (0, 26, 26) {real, imag} */,
  {32'h3ce0f145, 32'h3d8be12f} /* (0, 26, 25) {real, imag} */,
  {32'h3d55470a, 32'hbdc1d792} /* (0, 26, 24) {real, imag} */,
  {32'h3db4f015, 32'hbc07cb40} /* (0, 26, 23) {real, imag} */,
  {32'hbd8e4698, 32'hbc522d78} /* (0, 26, 22) {real, imag} */,
  {32'hbd215500, 32'hbd3f011b} /* (0, 26, 21) {real, imag} */,
  {32'h3cb6bdde, 32'hbc1358c8} /* (0, 26, 20) {real, imag} */,
  {32'hba863dc0, 32'hbcde6f78} /* (0, 26, 19) {real, imag} */,
  {32'hbb073030, 32'hbc7d313e} /* (0, 26, 18) {real, imag} */,
  {32'h3ba6365c, 32'h3bf75e34} /* (0, 26, 17) {real, imag} */,
  {32'hbb868e48, 32'h00000000} /* (0, 26, 16) {real, imag} */,
  {32'h3ba6365c, 32'hbbf75e34} /* (0, 26, 15) {real, imag} */,
  {32'hbb073030, 32'h3c7d313e} /* (0, 26, 14) {real, imag} */,
  {32'hba863dc0, 32'h3cde6f78} /* (0, 26, 13) {real, imag} */,
  {32'h3cb6bdde, 32'h3c1358c8} /* (0, 26, 12) {real, imag} */,
  {32'hbd215500, 32'h3d3f011b} /* (0, 26, 11) {real, imag} */,
  {32'hbd8e4698, 32'h3c522d78} /* (0, 26, 10) {real, imag} */,
  {32'h3db4f015, 32'h3c07cb40} /* (0, 26, 9) {real, imag} */,
  {32'h3d55470a, 32'h3dc1d792} /* (0, 26, 8) {real, imag} */,
  {32'h3ce0f145, 32'hbd8be12f} /* (0, 26, 7) {real, imag} */,
  {32'h3cca84b3, 32'h3ba2f3c0} /* (0, 26, 6) {real, imag} */,
  {32'h3e11c5c2, 32'h3d0018cf} /* (0, 26, 5) {real, imag} */,
  {32'hbdfa53e6, 32'hbde19571} /* (0, 26, 4) {real, imag} */,
  {32'hbd12b92c, 32'h3d29c27f} /* (0, 26, 3) {real, imag} */,
  {32'h3e3c427b, 32'hbdaec14d} /* (0, 26, 2) {real, imag} */,
  {32'hbf496816, 32'hbd7bd300} /* (0, 26, 1) {real, imag} */,
  {32'hbe92af36, 32'h00000000} /* (0, 26, 0) {real, imag} */,
  {32'hbf65e3ba, 32'hbe494f78} /* (0, 25, 31) {real, imag} */,
  {32'h3e8060fb, 32'h3e42b451} /* (0, 25, 30) {real, imag} */,
  {32'hbdc0a8f9, 32'h3c8ad2c8} /* (0, 25, 29) {real, imag} */,
  {32'hbe0cdbf4, 32'h3cf93a00} /* (0, 25, 28) {real, imag} */,
  {32'h3e4f5b8a, 32'hbe044082} /* (0, 25, 27) {real, imag} */,
  {32'h3de882e8, 32'hbc881342} /* (0, 25, 26) {real, imag} */,
  {32'hbc07bb3e, 32'h3de3efc8} /* (0, 25, 25) {real, imag} */,
  {32'h3cc2320d, 32'hbe27d723} /* (0, 25, 24) {real, imag} */,
  {32'hbd978c53, 32'hbd64e13f} /* (0, 25, 23) {real, imag} */,
  {32'h3d19b63f, 32'hbd4714e6} /* (0, 25, 22) {real, imag} */,
  {32'hbd9254a6, 32'h3c95b51c} /* (0, 25, 21) {real, imag} */,
  {32'h3c885bec, 32'hbd0c42a6} /* (0, 25, 20) {real, imag} */,
  {32'hbc43f4c6, 32'hbbfc45b8} /* (0, 25, 19) {real, imag} */,
  {32'hbc87c30d, 32'h3c203879} /* (0, 25, 18) {real, imag} */,
  {32'hbd02d125, 32'hbd4d6543} /* (0, 25, 17) {real, imag} */,
  {32'h3d4ab017, 32'h00000000} /* (0, 25, 16) {real, imag} */,
  {32'hbd02d125, 32'h3d4d6543} /* (0, 25, 15) {real, imag} */,
  {32'hbc87c30d, 32'hbc203879} /* (0, 25, 14) {real, imag} */,
  {32'hbc43f4c6, 32'h3bfc45b8} /* (0, 25, 13) {real, imag} */,
  {32'h3c885bec, 32'h3d0c42a6} /* (0, 25, 12) {real, imag} */,
  {32'hbd9254a6, 32'hbc95b51c} /* (0, 25, 11) {real, imag} */,
  {32'h3d19b63f, 32'h3d4714e6} /* (0, 25, 10) {real, imag} */,
  {32'hbd978c53, 32'h3d64e13f} /* (0, 25, 9) {real, imag} */,
  {32'h3cc2320d, 32'h3e27d723} /* (0, 25, 8) {real, imag} */,
  {32'hbc07bb3e, 32'hbde3efc8} /* (0, 25, 7) {real, imag} */,
  {32'h3de882e8, 32'h3c881342} /* (0, 25, 6) {real, imag} */,
  {32'h3e4f5b8a, 32'h3e044082} /* (0, 25, 5) {real, imag} */,
  {32'hbe0cdbf4, 32'hbcf93a00} /* (0, 25, 4) {real, imag} */,
  {32'hbdc0a8f9, 32'hbc8ad2c8} /* (0, 25, 3) {real, imag} */,
  {32'h3e8060fb, 32'hbe42b451} /* (0, 25, 2) {real, imag} */,
  {32'hbf65e3ba, 32'h3e494f78} /* (0, 25, 1) {real, imag} */,
  {32'hbe9102c1, 32'h00000000} /* (0, 25, 0) {real, imag} */,
  {32'hbf28e684, 32'hbd55784c} /* (0, 24, 31) {real, imag} */,
  {32'h3e3ad7e5, 32'h3db51054} /* (0, 24, 30) {real, imag} */,
  {32'hbcd93086, 32'h3ce27866} /* (0, 24, 29) {real, imag} */,
  {32'hbe230d0c, 32'hbd06a040} /* (0, 24, 28) {real, imag} */,
  {32'h3dcfdd8c, 32'hbdae7034} /* (0, 24, 27) {real, imag} */,
  {32'hbcd94dbe, 32'h39191a00} /* (0, 24, 26) {real, imag} */,
  {32'h3bb7a2a0, 32'h3d0fcff4} /* (0, 24, 25) {real, imag} */,
  {32'hbc7fe01c, 32'hbc9c468e} /* (0, 24, 24) {real, imag} */,
  {32'h3c15a7e8, 32'hbd8b6822} /* (0, 24, 23) {real, imag} */,
  {32'h3d82e808, 32'h3d959f62} /* (0, 24, 22) {real, imag} */,
  {32'hbd507fda, 32'hbc676f1e} /* (0, 24, 21) {real, imag} */,
  {32'hbd03f76e, 32'h3b7ef254} /* (0, 24, 20) {real, imag} */,
  {32'hbd3d6c31, 32'h3c7c96da} /* (0, 24, 19) {real, imag} */,
  {32'h3d268cf8, 32'hbd2e4a31} /* (0, 24, 18) {real, imag} */,
  {32'hbd01b96a, 32'h3d26f5b3} /* (0, 24, 17) {real, imag} */,
  {32'hbc630497, 32'h00000000} /* (0, 24, 16) {real, imag} */,
  {32'hbd01b96a, 32'hbd26f5b3} /* (0, 24, 15) {real, imag} */,
  {32'h3d268cf8, 32'h3d2e4a31} /* (0, 24, 14) {real, imag} */,
  {32'hbd3d6c31, 32'hbc7c96da} /* (0, 24, 13) {real, imag} */,
  {32'hbd03f76e, 32'hbb7ef254} /* (0, 24, 12) {real, imag} */,
  {32'hbd507fda, 32'h3c676f1e} /* (0, 24, 11) {real, imag} */,
  {32'h3d82e808, 32'hbd959f62} /* (0, 24, 10) {real, imag} */,
  {32'h3c15a7e8, 32'h3d8b6822} /* (0, 24, 9) {real, imag} */,
  {32'hbc7fe01c, 32'h3c9c468e} /* (0, 24, 8) {real, imag} */,
  {32'h3bb7a2a0, 32'hbd0fcff4} /* (0, 24, 7) {real, imag} */,
  {32'hbcd94dbe, 32'hb9191a00} /* (0, 24, 6) {real, imag} */,
  {32'h3dcfdd8c, 32'h3dae7034} /* (0, 24, 5) {real, imag} */,
  {32'hbe230d0c, 32'h3d06a040} /* (0, 24, 4) {real, imag} */,
  {32'hbcd93086, 32'hbce27866} /* (0, 24, 3) {real, imag} */,
  {32'h3e3ad7e5, 32'hbdb51054} /* (0, 24, 2) {real, imag} */,
  {32'hbf28e684, 32'h3d55784c} /* (0, 24, 1) {real, imag} */,
  {32'hbd442210, 32'h00000000} /* (0, 24, 0) {real, imag} */,
  {32'hbf149373, 32'h3d4a0f22} /* (0, 23, 31) {real, imag} */,
  {32'h3db3c324, 32'h3de6bf66} /* (0, 23, 30) {real, imag} */,
  {32'h3ddc5787, 32'h3d05e1d4} /* (0, 23, 29) {real, imag} */,
  {32'hbd82d814, 32'hbc7d6156} /* (0, 23, 28) {real, imag} */,
  {32'h3dd8faec, 32'hbd7423aa} /* (0, 23, 27) {real, imag} */,
  {32'hbd14eae2, 32'hbc2a94a1} /* (0, 23, 26) {real, imag} */,
  {32'hbd79b577, 32'h3d66087d} /* (0, 23, 25) {real, imag} */,
  {32'h3d8e1f99, 32'h3c1417a0} /* (0, 23, 24) {real, imag} */,
  {32'hbc3b846e, 32'hbce57dbf} /* (0, 23, 23) {real, imag} */,
  {32'hbc913fd4, 32'hbd03a6f1} /* (0, 23, 22) {real, imag} */,
  {32'h3d65c1c5, 32'hbca34e38} /* (0, 23, 21) {real, imag} */,
  {32'h3caa2ea1, 32'h3c1787fc} /* (0, 23, 20) {real, imag} */,
  {32'h3c174272, 32'h3ba3bca2} /* (0, 23, 19) {real, imag} */,
  {32'h3d0872b5, 32'hbd095eb8} /* (0, 23, 18) {real, imag} */,
  {32'hbd67c1ea, 32'hbcf6d19b} /* (0, 23, 17) {real, imag} */,
  {32'hbd2155db, 32'h00000000} /* (0, 23, 16) {real, imag} */,
  {32'hbd67c1ea, 32'h3cf6d19b} /* (0, 23, 15) {real, imag} */,
  {32'h3d0872b5, 32'h3d095eb8} /* (0, 23, 14) {real, imag} */,
  {32'h3c174272, 32'hbba3bca2} /* (0, 23, 13) {real, imag} */,
  {32'h3caa2ea1, 32'hbc1787fc} /* (0, 23, 12) {real, imag} */,
  {32'h3d65c1c5, 32'h3ca34e38} /* (0, 23, 11) {real, imag} */,
  {32'hbc913fd4, 32'h3d03a6f1} /* (0, 23, 10) {real, imag} */,
  {32'hbc3b846e, 32'h3ce57dbf} /* (0, 23, 9) {real, imag} */,
  {32'h3d8e1f99, 32'hbc1417a0} /* (0, 23, 8) {real, imag} */,
  {32'hbd79b577, 32'hbd66087d} /* (0, 23, 7) {real, imag} */,
  {32'hbd14eae2, 32'h3c2a94a1} /* (0, 23, 6) {real, imag} */,
  {32'h3dd8faec, 32'h3d7423aa} /* (0, 23, 5) {real, imag} */,
  {32'hbd82d814, 32'h3c7d6156} /* (0, 23, 4) {real, imag} */,
  {32'h3ddc5787, 32'hbd05e1d4} /* (0, 23, 3) {real, imag} */,
  {32'h3db3c324, 32'hbde6bf66} /* (0, 23, 2) {real, imag} */,
  {32'hbf149373, 32'hbd4a0f22} /* (0, 23, 1) {real, imag} */,
  {32'hbb41d100, 32'h00000000} /* (0, 23, 0) {real, imag} */,
  {32'hbef7a3d4, 32'h3e139836} /* (0, 22, 31) {real, imag} */,
  {32'h3de44362, 32'h3d20c64e} /* (0, 22, 30) {real, imag} */,
  {32'h3e170bca, 32'h3d9c06ca} /* (0, 22, 29) {real, imag} */,
  {32'hbdd55b81, 32'hbd3660b9} /* (0, 22, 28) {real, imag} */,
  {32'h3dc9833b, 32'hbda29d9a} /* (0, 22, 27) {real, imag} */,
  {32'hbceec9ac, 32'hbb8c1b1c} /* (0, 22, 26) {real, imag} */,
  {32'hbdd00e68, 32'hbbecb3a0} /* (0, 22, 25) {real, imag} */,
  {32'h3d6d69b8, 32'hbb27cc86} /* (0, 22, 24) {real, imag} */,
  {32'hbc9ead3d, 32'h3c6b227a} /* (0, 22, 23) {real, imag} */,
  {32'h3d274051, 32'hbc0aa346} /* (0, 22, 22) {real, imag} */,
  {32'hbc93aba9, 32'h3c7f7860} /* (0, 22, 21) {real, imag} */,
  {32'h3d48c54b, 32'hbc8e64d1} /* (0, 22, 20) {real, imag} */,
  {32'hbb071f54, 32'h3d9b18de} /* (0, 22, 19) {real, imag} */,
  {32'hbd526b2a, 32'h3cfc5ad2} /* (0, 22, 18) {real, imag} */,
  {32'h39593bc0, 32'h3cb3f14c} /* (0, 22, 17) {real, imag} */,
  {32'hbd4cbe82, 32'h00000000} /* (0, 22, 16) {real, imag} */,
  {32'h39593bc0, 32'hbcb3f14c} /* (0, 22, 15) {real, imag} */,
  {32'hbd526b2a, 32'hbcfc5ad2} /* (0, 22, 14) {real, imag} */,
  {32'hbb071f54, 32'hbd9b18de} /* (0, 22, 13) {real, imag} */,
  {32'h3d48c54b, 32'h3c8e64d1} /* (0, 22, 12) {real, imag} */,
  {32'hbc93aba9, 32'hbc7f7860} /* (0, 22, 11) {real, imag} */,
  {32'h3d274051, 32'h3c0aa346} /* (0, 22, 10) {real, imag} */,
  {32'hbc9ead3d, 32'hbc6b227a} /* (0, 22, 9) {real, imag} */,
  {32'h3d6d69b8, 32'h3b27cc86} /* (0, 22, 8) {real, imag} */,
  {32'hbdd00e68, 32'h3becb3a0} /* (0, 22, 7) {real, imag} */,
  {32'hbceec9ac, 32'h3b8c1b1c} /* (0, 22, 6) {real, imag} */,
  {32'h3dc9833b, 32'h3da29d9a} /* (0, 22, 5) {real, imag} */,
  {32'hbdd55b81, 32'h3d3660b9} /* (0, 22, 4) {real, imag} */,
  {32'h3e170bca, 32'hbd9c06ca} /* (0, 22, 3) {real, imag} */,
  {32'h3de44362, 32'hbd20c64e} /* (0, 22, 2) {real, imag} */,
  {32'hbef7a3d4, 32'hbe139836} /* (0, 22, 1) {real, imag} */,
  {32'hbb968080, 32'h00000000} /* (0, 22, 0) {real, imag} */,
  {32'hbe8a8924, 32'h3dcc8096} /* (0, 21, 31) {real, imag} */,
  {32'h3b303e40, 32'h3cad55b6} /* (0, 21, 30) {real, imag} */,
  {32'h3d85aa18, 32'h3dcbd848} /* (0, 21, 29) {real, imag} */,
  {32'hbd701e51, 32'hbc78b690} /* (0, 21, 28) {real, imag} */,
  {32'h3d06af79, 32'hbd854b02} /* (0, 21, 27) {real, imag} */,
  {32'hbd4a0881, 32'h3c8a9ebf} /* (0, 21, 26) {real, imag} */,
  {32'hbcbe8666, 32'hbe02c042} /* (0, 21, 25) {real, imag} */,
  {32'hbd1e7927, 32'h3c42dc50} /* (0, 21, 24) {real, imag} */,
  {32'hbc8e4e97, 32'h3db636f6} /* (0, 21, 23) {real, imag} */,
  {32'hbb092208, 32'h3d37d58f} /* (0, 21, 22) {real, imag} */,
  {32'h3d12ced0, 32'hbd69cc9a} /* (0, 21, 21) {real, imag} */,
  {32'h3d88acbf, 32'hbd304856} /* (0, 21, 20) {real, imag} */,
  {32'hbb8af83a, 32'h3ceefe02} /* (0, 21, 19) {real, imag} */,
  {32'hbcde1ba8, 32'hbda01f1c} /* (0, 21, 18) {real, imag} */,
  {32'h3c008ca6, 32'hbc9abcb8} /* (0, 21, 17) {real, imag} */,
  {32'hbca0d4df, 32'h00000000} /* (0, 21, 16) {real, imag} */,
  {32'h3c008ca6, 32'h3c9abcb8} /* (0, 21, 15) {real, imag} */,
  {32'hbcde1ba8, 32'h3da01f1c} /* (0, 21, 14) {real, imag} */,
  {32'hbb8af83a, 32'hbceefe02} /* (0, 21, 13) {real, imag} */,
  {32'h3d88acbf, 32'h3d304856} /* (0, 21, 12) {real, imag} */,
  {32'h3d12ced0, 32'h3d69cc9a} /* (0, 21, 11) {real, imag} */,
  {32'hbb092208, 32'hbd37d58f} /* (0, 21, 10) {real, imag} */,
  {32'hbc8e4e97, 32'hbdb636f6} /* (0, 21, 9) {real, imag} */,
  {32'hbd1e7927, 32'hbc42dc50} /* (0, 21, 8) {real, imag} */,
  {32'hbcbe8666, 32'h3e02c042} /* (0, 21, 7) {real, imag} */,
  {32'hbd4a0881, 32'hbc8a9ebf} /* (0, 21, 6) {real, imag} */,
  {32'h3d06af79, 32'h3d854b02} /* (0, 21, 5) {real, imag} */,
  {32'hbd701e51, 32'h3c78b690} /* (0, 21, 4) {real, imag} */,
  {32'h3d85aa18, 32'hbdcbd848} /* (0, 21, 3) {real, imag} */,
  {32'h3b303e40, 32'hbcad55b6} /* (0, 21, 2) {real, imag} */,
  {32'hbe8a8924, 32'hbdcc8096} /* (0, 21, 1) {real, imag} */,
  {32'h3cc72f00, 32'h00000000} /* (0, 21, 0) {real, imag} */,
  {32'h3dd86d78, 32'hbdaea494} /* (0, 20, 31) {real, imag} */,
  {32'hbe76523f, 32'h3cb3d514} /* (0, 20, 30) {real, imag} */,
  {32'hbd336daf, 32'h3de9b033} /* (0, 20, 29) {real, imag} */,
  {32'h3d273987, 32'hbd01f5cb} /* (0, 20, 28) {real, imag} */,
  {32'hbd0a2e2e, 32'hbdb98f28} /* (0, 20, 27) {real, imag} */,
  {32'hbcc6ff2e, 32'h3d5d654a} /* (0, 20, 26) {real, imag} */,
  {32'hbda34d31, 32'hbd37cd54} /* (0, 20, 25) {real, imag} */,
  {32'h3d1b988b, 32'h3d213af0} /* (0, 20, 24) {real, imag} */,
  {32'h3cecdee5, 32'h3b547320} /* (0, 20, 23) {real, imag} */,
  {32'hbd091f60, 32'hbd4f401f} /* (0, 20, 22) {real, imag} */,
  {32'h3c9a618b, 32'h3cda8d1a} /* (0, 20, 21) {real, imag} */,
  {32'h3d637d6d, 32'h3c9b04c4} /* (0, 20, 20) {real, imag} */,
  {32'hbd85ffa4, 32'hbc235a88} /* (0, 20, 19) {real, imag} */,
  {32'h3d57fdb0, 32'hbd2a86a0} /* (0, 20, 18) {real, imag} */,
  {32'hbd0e46d1, 32'hbcd5241c} /* (0, 20, 17) {real, imag} */,
  {32'h3ca19b74, 32'h00000000} /* (0, 20, 16) {real, imag} */,
  {32'hbd0e46d1, 32'h3cd5241c} /* (0, 20, 15) {real, imag} */,
  {32'h3d57fdb0, 32'h3d2a86a0} /* (0, 20, 14) {real, imag} */,
  {32'hbd85ffa4, 32'h3c235a88} /* (0, 20, 13) {real, imag} */,
  {32'h3d637d6d, 32'hbc9b04c4} /* (0, 20, 12) {real, imag} */,
  {32'h3c9a618b, 32'hbcda8d1a} /* (0, 20, 11) {real, imag} */,
  {32'hbd091f60, 32'h3d4f401f} /* (0, 20, 10) {real, imag} */,
  {32'h3cecdee5, 32'hbb547320} /* (0, 20, 9) {real, imag} */,
  {32'h3d1b988b, 32'hbd213af0} /* (0, 20, 8) {real, imag} */,
  {32'hbda34d31, 32'h3d37cd54} /* (0, 20, 7) {real, imag} */,
  {32'hbcc6ff2e, 32'hbd5d654a} /* (0, 20, 6) {real, imag} */,
  {32'hbd0a2e2e, 32'h3db98f28} /* (0, 20, 5) {real, imag} */,
  {32'h3d273987, 32'h3d01f5cb} /* (0, 20, 4) {real, imag} */,
  {32'hbd336daf, 32'hbde9b033} /* (0, 20, 3) {real, imag} */,
  {32'hbe76523f, 32'hbcb3d514} /* (0, 20, 2) {real, imag} */,
  {32'h3dd86d78, 32'h3daea494} /* (0, 20, 1) {real, imag} */,
  {32'h3e99354e, 32'h00000000} /* (0, 20, 0) {real, imag} */,
  {32'h3e930610, 32'hbde121fc} /* (0, 19, 31) {real, imag} */,
  {32'hbe5c738b, 32'h3c3891c8} /* (0, 19, 30) {real, imag} */,
  {32'hbd73aed3, 32'h3d033c96} /* (0, 19, 29) {real, imag} */,
  {32'hbbf3e798, 32'hbd8d94d6} /* (0, 19, 28) {real, imag} */,
  {32'h3a80e400, 32'hbbbed990} /* (0, 19, 27) {real, imag} */,
  {32'hbd90d589, 32'hbd8bddf2} /* (0, 19, 26) {real, imag} */,
  {32'hbd16eb00, 32'hbd3ada10} /* (0, 19, 25) {real, imag} */,
  {32'h3c425f56, 32'h3da1f3d4} /* (0, 19, 24) {real, imag} */,
  {32'hbd0346cc, 32'h3c91d3ca} /* (0, 19, 23) {real, imag} */,
  {32'h3c9d9e80, 32'h3d275e2b} /* (0, 19, 22) {real, imag} */,
  {32'hbd0491c6, 32'h3de27822} /* (0, 19, 21) {real, imag} */,
  {32'hbd2116e8, 32'h3c35e7d8} /* (0, 19, 20) {real, imag} */,
  {32'h3caf05f7, 32'hbc201752} /* (0, 19, 19) {real, imag} */,
  {32'h3cdf83b4, 32'hbb1b0902} /* (0, 19, 18) {real, imag} */,
  {32'h3c202915, 32'h3b02dbec} /* (0, 19, 17) {real, imag} */,
  {32'hbc3943fc, 32'h00000000} /* (0, 19, 16) {real, imag} */,
  {32'h3c202915, 32'hbb02dbec} /* (0, 19, 15) {real, imag} */,
  {32'h3cdf83b4, 32'h3b1b0902} /* (0, 19, 14) {real, imag} */,
  {32'h3caf05f7, 32'h3c201752} /* (0, 19, 13) {real, imag} */,
  {32'hbd2116e8, 32'hbc35e7d8} /* (0, 19, 12) {real, imag} */,
  {32'hbd0491c6, 32'hbde27822} /* (0, 19, 11) {real, imag} */,
  {32'h3c9d9e80, 32'hbd275e2b} /* (0, 19, 10) {real, imag} */,
  {32'hbd0346cc, 32'hbc91d3ca} /* (0, 19, 9) {real, imag} */,
  {32'h3c425f56, 32'hbda1f3d4} /* (0, 19, 8) {real, imag} */,
  {32'hbd16eb00, 32'h3d3ada10} /* (0, 19, 7) {real, imag} */,
  {32'hbd90d589, 32'h3d8bddf2} /* (0, 19, 6) {real, imag} */,
  {32'h3a80e400, 32'h3bbed990} /* (0, 19, 5) {real, imag} */,
  {32'hbbf3e798, 32'h3d8d94d6} /* (0, 19, 4) {real, imag} */,
  {32'hbd73aed3, 32'hbd033c96} /* (0, 19, 3) {real, imag} */,
  {32'hbe5c738b, 32'hbc3891c8} /* (0, 19, 2) {real, imag} */,
  {32'h3e930610, 32'h3de121fc} /* (0, 19, 1) {real, imag} */,
  {32'h3efa9a1e, 32'h00000000} /* (0, 19, 0) {real, imag} */,
  {32'h3ed59edf, 32'hbe27a5de} /* (0, 18, 31) {real, imag} */,
  {32'hbe916d98, 32'h3dfc2471} /* (0, 18, 30) {real, imag} */,
  {32'hbdcd0ad0, 32'h3d724364} /* (0, 18, 29) {real, imag} */,
  {32'h3dc0e467, 32'hbdb3d5cb} /* (0, 18, 28) {real, imag} */,
  {32'hbd7b866e, 32'h3c865d4d} /* (0, 18, 27) {real, imag} */,
  {32'hbbe7f62e, 32'hbd8add85} /* (0, 18, 26) {real, imag} */,
  {32'hbd7a7e24, 32'h3dbfd66a} /* (0, 18, 25) {real, imag} */,
  {32'hbd0e2ba7, 32'hbca66d03} /* (0, 18, 24) {real, imag} */,
  {32'hbd04f41d, 32'h3c16e61c} /* (0, 18, 23) {real, imag} */,
  {32'hbcf1107c, 32'h3d4e7f31} /* (0, 18, 22) {real, imag} */,
  {32'hbc0d4245, 32'h3cf76682} /* (0, 18, 21) {real, imag} */,
  {32'h3cfac042, 32'hbd0bc3e8} /* (0, 18, 20) {real, imag} */,
  {32'hbd2137a8, 32'hbc833210} /* (0, 18, 19) {real, imag} */,
  {32'hbd1dc45f, 32'h3d3784a4} /* (0, 18, 18) {real, imag} */,
  {32'hbd15800c, 32'h3c2834b0} /* (0, 18, 17) {real, imag} */,
  {32'h3a9f5f95, 32'h00000000} /* (0, 18, 16) {real, imag} */,
  {32'hbd15800c, 32'hbc2834b0} /* (0, 18, 15) {real, imag} */,
  {32'hbd1dc45f, 32'hbd3784a4} /* (0, 18, 14) {real, imag} */,
  {32'hbd2137a8, 32'h3c833210} /* (0, 18, 13) {real, imag} */,
  {32'h3cfac042, 32'h3d0bc3e8} /* (0, 18, 12) {real, imag} */,
  {32'hbc0d4245, 32'hbcf76682} /* (0, 18, 11) {real, imag} */,
  {32'hbcf1107c, 32'hbd4e7f31} /* (0, 18, 10) {real, imag} */,
  {32'hbd04f41d, 32'hbc16e61c} /* (0, 18, 9) {real, imag} */,
  {32'hbd0e2ba7, 32'h3ca66d03} /* (0, 18, 8) {real, imag} */,
  {32'hbd7a7e24, 32'hbdbfd66a} /* (0, 18, 7) {real, imag} */,
  {32'hbbe7f62e, 32'h3d8add85} /* (0, 18, 6) {real, imag} */,
  {32'hbd7b866e, 32'hbc865d4d} /* (0, 18, 5) {real, imag} */,
  {32'h3dc0e467, 32'h3db3d5cb} /* (0, 18, 4) {real, imag} */,
  {32'hbdcd0ad0, 32'hbd724364} /* (0, 18, 3) {real, imag} */,
  {32'hbe916d98, 32'hbdfc2471} /* (0, 18, 2) {real, imag} */,
  {32'h3ed59edf, 32'h3e27a5de} /* (0, 18, 1) {real, imag} */,
  {32'h3ed00180, 32'h00000000} /* (0, 18, 0) {real, imag} */,
  {32'h3ecfe619, 32'hbe44ede8} /* (0, 17, 31) {real, imag} */,
  {32'hbeb45ad0, 32'hbc82ee14} /* (0, 17, 30) {real, imag} */,
  {32'hbc725cdc, 32'hbc997124} /* (0, 17, 29) {real, imag} */,
  {32'h3d358aaf, 32'hbcb1c08e} /* (0, 17, 28) {real, imag} */,
  {32'hba10cc00, 32'h3d78c733} /* (0, 17, 27) {real, imag} */,
  {32'h3caa6e61, 32'hbd292b4c} /* (0, 17, 26) {real, imag} */,
  {32'h3c90e5be, 32'h3d7fe156} /* (0, 17, 25) {real, imag} */,
  {32'hbc095478, 32'h3b0c1370} /* (0, 17, 24) {real, imag} */,
  {32'h3bf45068, 32'hbd0d999e} /* (0, 17, 23) {real, imag} */,
  {32'h3d8d8486, 32'hbc417cee} /* (0, 17, 22) {real, imag} */,
  {32'hbdb1e4d3, 32'h3cfbf8a8} /* (0, 17, 21) {real, imag} */,
  {32'h3cabf3bb, 32'h3be49f70} /* (0, 17, 20) {real, imag} */,
  {32'hbd12e14a, 32'hbc23a052} /* (0, 17, 19) {real, imag} */,
  {32'hbb9c5890, 32'h3d318469} /* (0, 17, 18) {real, imag} */,
  {32'hbb592322, 32'h3c56db13} /* (0, 17, 17) {real, imag} */,
  {32'h3d215d93, 32'h00000000} /* (0, 17, 16) {real, imag} */,
  {32'hbb592322, 32'hbc56db13} /* (0, 17, 15) {real, imag} */,
  {32'hbb9c5890, 32'hbd318469} /* (0, 17, 14) {real, imag} */,
  {32'hbd12e14a, 32'h3c23a052} /* (0, 17, 13) {real, imag} */,
  {32'h3cabf3bb, 32'hbbe49f70} /* (0, 17, 12) {real, imag} */,
  {32'hbdb1e4d3, 32'hbcfbf8a8} /* (0, 17, 11) {real, imag} */,
  {32'h3d8d8486, 32'h3c417cee} /* (0, 17, 10) {real, imag} */,
  {32'h3bf45068, 32'h3d0d999e} /* (0, 17, 9) {real, imag} */,
  {32'hbc095478, 32'hbb0c1370} /* (0, 17, 8) {real, imag} */,
  {32'h3c90e5be, 32'hbd7fe156} /* (0, 17, 7) {real, imag} */,
  {32'h3caa6e61, 32'h3d292b4c} /* (0, 17, 6) {real, imag} */,
  {32'hba10cc00, 32'hbd78c733} /* (0, 17, 5) {real, imag} */,
  {32'h3d358aaf, 32'h3cb1c08e} /* (0, 17, 4) {real, imag} */,
  {32'hbc725cdc, 32'h3c997124} /* (0, 17, 3) {real, imag} */,
  {32'hbeb45ad0, 32'h3c82ee14} /* (0, 17, 2) {real, imag} */,
  {32'h3ecfe619, 32'h3e44ede8} /* (0, 17, 1) {real, imag} */,
  {32'h3ed0829d, 32'h00000000} /* (0, 17, 0) {real, imag} */,
  {32'h3eff9562, 32'hbe353312} /* (0, 16, 31) {real, imag} */,
  {32'hbee303b1, 32'h3c4d824e} /* (0, 16, 30) {real, imag} */,
  {32'hbd07b097, 32'hbe5a41a8} /* (0, 16, 29) {real, imag} */,
  {32'h3db6ae6a, 32'h3c446fb8} /* (0, 16, 28) {real, imag} */,
  {32'hbd8da400, 32'h3e046e1b} /* (0, 16, 27) {real, imag} */,
  {32'hbd11b5a4, 32'hbc8a8da8} /* (0, 16, 26) {real, imag} */,
  {32'h3d9de84d, 32'h3ccbab40} /* (0, 16, 25) {real, imag} */,
  {32'hbd526bac, 32'h3d2be942} /* (0, 16, 24) {real, imag} */,
  {32'h3ca2604d, 32'h3d171b0b} /* (0, 16, 23) {real, imag} */,
  {32'hbb0ed288, 32'hbd711194} /* (0, 16, 22) {real, imag} */,
  {32'h3cedf9d5, 32'h3d2af2ec} /* (0, 16, 21) {real, imag} */,
  {32'h3c5dd7e9, 32'h3da031b5} /* (0, 16, 20) {real, imag} */,
  {32'h3c0447f4, 32'h3c270580} /* (0, 16, 19) {real, imag} */,
  {32'h3d73030a, 32'hbd740036} /* (0, 16, 18) {real, imag} */,
  {32'hbcb004dc, 32'h3d0d669b} /* (0, 16, 17) {real, imag} */,
  {32'h3c8564a1, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hbcb004dc, 32'hbd0d669b} /* (0, 16, 15) {real, imag} */,
  {32'h3d73030a, 32'h3d740036} /* (0, 16, 14) {real, imag} */,
  {32'h3c0447f4, 32'hbc270580} /* (0, 16, 13) {real, imag} */,
  {32'h3c5dd7e9, 32'hbda031b5} /* (0, 16, 12) {real, imag} */,
  {32'h3cedf9d5, 32'hbd2af2ec} /* (0, 16, 11) {real, imag} */,
  {32'hbb0ed288, 32'h3d711194} /* (0, 16, 10) {real, imag} */,
  {32'h3ca2604d, 32'hbd171b0b} /* (0, 16, 9) {real, imag} */,
  {32'hbd526bac, 32'hbd2be942} /* (0, 16, 8) {real, imag} */,
  {32'h3d9de84d, 32'hbccbab40} /* (0, 16, 7) {real, imag} */,
  {32'hbd11b5a4, 32'h3c8a8da8} /* (0, 16, 6) {real, imag} */,
  {32'hbd8da400, 32'hbe046e1b} /* (0, 16, 5) {real, imag} */,
  {32'h3db6ae6a, 32'hbc446fb8} /* (0, 16, 4) {real, imag} */,
  {32'hbd07b097, 32'h3e5a41a8} /* (0, 16, 3) {real, imag} */,
  {32'hbee303b1, 32'hbc4d824e} /* (0, 16, 2) {real, imag} */,
  {32'h3eff9562, 32'h3e353312} /* (0, 16, 1) {real, imag} */,
  {32'h3f0487c7, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h3f346e38, 32'hbe6629d8} /* (0, 15, 31) {real, imag} */,
  {32'hbe6241c8, 32'h3e690fde} /* (0, 15, 30) {real, imag} */,
  {32'hbdfd9cbc, 32'hbe00145c} /* (0, 15, 29) {real, imag} */,
  {32'h3d2bcd99, 32'h3c285800} /* (0, 15, 28) {real, imag} */,
  {32'hbdfadce1, 32'h3d89b428} /* (0, 15, 27) {real, imag} */,
  {32'h3cb04047, 32'hbcd46bb8} /* (0, 15, 26) {real, imag} */,
  {32'h3d11d716, 32'h3d83a84f} /* (0, 15, 25) {real, imag} */,
  {32'hbda32795, 32'h3d7e69c5} /* (0, 15, 24) {real, imag} */,
  {32'hbd7a939d, 32'hbd552158} /* (0, 15, 23) {real, imag} */,
  {32'h3c35b25c, 32'h3d096540} /* (0, 15, 22) {real, imag} */,
  {32'hbc96f2b4, 32'hbcad0bd4} /* (0, 15, 21) {real, imag} */,
  {32'hbcdc7e5d, 32'hbc42983c} /* (0, 15, 20) {real, imag} */,
  {32'hbda6e389, 32'hbcffcccf} /* (0, 15, 19) {real, imag} */,
  {32'h3c85c13d, 32'hbd90b172} /* (0, 15, 18) {real, imag} */,
  {32'h3b96a1a1, 32'hbca61e3a} /* (0, 15, 17) {real, imag} */,
  {32'hbce3b9f2, 32'h00000000} /* (0, 15, 16) {real, imag} */,
  {32'h3b96a1a1, 32'h3ca61e3a} /* (0, 15, 15) {real, imag} */,
  {32'h3c85c13d, 32'h3d90b172} /* (0, 15, 14) {real, imag} */,
  {32'hbda6e389, 32'h3cffcccf} /* (0, 15, 13) {real, imag} */,
  {32'hbcdc7e5d, 32'h3c42983c} /* (0, 15, 12) {real, imag} */,
  {32'hbc96f2b4, 32'h3cad0bd4} /* (0, 15, 11) {real, imag} */,
  {32'h3c35b25c, 32'hbd096540} /* (0, 15, 10) {real, imag} */,
  {32'hbd7a939d, 32'h3d552158} /* (0, 15, 9) {real, imag} */,
  {32'hbda32795, 32'hbd7e69c5} /* (0, 15, 8) {real, imag} */,
  {32'h3d11d716, 32'hbd83a84f} /* (0, 15, 7) {real, imag} */,
  {32'h3cb04047, 32'h3cd46bb8} /* (0, 15, 6) {real, imag} */,
  {32'hbdfadce1, 32'hbd89b428} /* (0, 15, 5) {real, imag} */,
  {32'h3d2bcd99, 32'hbc285800} /* (0, 15, 4) {real, imag} */,
  {32'hbdfd9cbc, 32'h3e00145c} /* (0, 15, 3) {real, imag} */,
  {32'hbe6241c8, 32'hbe690fde} /* (0, 15, 2) {real, imag} */,
  {32'h3f346e38, 32'h3e6629d8} /* (0, 15, 1) {real, imag} */,
  {32'h3e941f2b, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h3f2bd902, 32'hbe18296e} /* (0, 14, 31) {real, imag} */,
  {32'hbe54b40e, 32'h3da4c60f} /* (0, 14, 30) {real, imag} */,
  {32'hbda9169e, 32'h3db876c4} /* (0, 14, 29) {real, imag} */,
  {32'hbcfc8244, 32'hbd11aa18} /* (0, 14, 28) {real, imag} */,
  {32'hbda0a341, 32'h3d8e2c1b} /* (0, 14, 27) {real, imag} */,
  {32'h3bfe4642, 32'hbd007fe6} /* (0, 14, 26) {real, imag} */,
  {32'h3d10b898, 32'h3c11dfe8} /* (0, 14, 25) {real, imag} */,
  {32'hbc3c2cbc, 32'hbbd49944} /* (0, 14, 24) {real, imag} */,
  {32'hb9a36680, 32'h3d51504a} /* (0, 14, 23) {real, imag} */,
  {32'h3c90e45a, 32'hba802da0} /* (0, 14, 22) {real, imag} */,
  {32'hbd0a4927, 32'hbc2a59cc} /* (0, 14, 21) {real, imag} */,
  {32'h3d139931, 32'hbd24ff16} /* (0, 14, 20) {real, imag} */,
  {32'hbceb5ba0, 32'h3cbf2b02} /* (0, 14, 19) {real, imag} */,
  {32'h3d09f7e1, 32'h3cca6b28} /* (0, 14, 18) {real, imag} */,
  {32'hbc4336c6, 32'h3b848e9c} /* (0, 14, 17) {real, imag} */,
  {32'hb92bb358, 32'h00000000} /* (0, 14, 16) {real, imag} */,
  {32'hbc4336c6, 32'hbb848e9c} /* (0, 14, 15) {real, imag} */,
  {32'h3d09f7e1, 32'hbcca6b28} /* (0, 14, 14) {real, imag} */,
  {32'hbceb5ba0, 32'hbcbf2b02} /* (0, 14, 13) {real, imag} */,
  {32'h3d139931, 32'h3d24ff16} /* (0, 14, 12) {real, imag} */,
  {32'hbd0a4927, 32'h3c2a59cc} /* (0, 14, 11) {real, imag} */,
  {32'h3c90e45a, 32'h3a802da0} /* (0, 14, 10) {real, imag} */,
  {32'hb9a36680, 32'hbd51504a} /* (0, 14, 9) {real, imag} */,
  {32'hbc3c2cbc, 32'h3bd49944} /* (0, 14, 8) {real, imag} */,
  {32'h3d10b898, 32'hbc11dfe8} /* (0, 14, 7) {real, imag} */,
  {32'h3bfe4642, 32'h3d007fe6} /* (0, 14, 6) {real, imag} */,
  {32'hbda0a341, 32'hbd8e2c1b} /* (0, 14, 5) {real, imag} */,
  {32'hbcfc8244, 32'h3d11aa18} /* (0, 14, 4) {real, imag} */,
  {32'hbda9169e, 32'hbdb876c4} /* (0, 14, 3) {real, imag} */,
  {32'hbe54b40e, 32'hbda4c60f} /* (0, 14, 2) {real, imag} */,
  {32'h3f2bd902, 32'h3e18296e} /* (0, 14, 1) {real, imag} */,
  {32'h3e819e2c, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h3f2afca0, 32'hbe045110} /* (0, 13, 31) {real, imag} */,
  {32'hbe75592d, 32'hbc0e08c8} /* (0, 13, 30) {real, imag} */,
  {32'hbdbac1a0, 32'h3daef856} /* (0, 13, 29) {real, imag} */,
  {32'h3d953186, 32'hbdc61ea6} /* (0, 13, 28) {real, imag} */,
  {32'hbcf884bc, 32'h3de556e3} /* (0, 13, 27) {real, imag} */,
  {32'hbce2c599, 32'h3d6805fc} /* (0, 13, 26) {real, imag} */,
  {32'hbc57b8fc, 32'hbc36f330} /* (0, 13, 25) {real, imag} */,
  {32'hbd6b9362, 32'h3b23c250} /* (0, 13, 24) {real, imag} */,
  {32'h3d238e22, 32'h3d89bc62} /* (0, 13, 23) {real, imag} */,
  {32'h3cfe5340, 32'h3c142254} /* (0, 13, 22) {real, imag} */,
  {32'hbd2fd8ba, 32'h3c00e84c} /* (0, 13, 21) {real, imag} */,
  {32'hbc2cbf45, 32'h3d3f5c16} /* (0, 13, 20) {real, imag} */,
  {32'h3c9836cd, 32'hbd2fead0} /* (0, 13, 19) {real, imag} */,
  {32'h3c02b405, 32'hbbb64d29} /* (0, 13, 18) {real, imag} */,
  {32'hbc2a7797, 32'h3ceebac4} /* (0, 13, 17) {real, imag} */,
  {32'hbd569639, 32'h00000000} /* (0, 13, 16) {real, imag} */,
  {32'hbc2a7797, 32'hbceebac4} /* (0, 13, 15) {real, imag} */,
  {32'h3c02b405, 32'h3bb64d29} /* (0, 13, 14) {real, imag} */,
  {32'h3c9836cd, 32'h3d2fead0} /* (0, 13, 13) {real, imag} */,
  {32'hbc2cbf45, 32'hbd3f5c16} /* (0, 13, 12) {real, imag} */,
  {32'hbd2fd8ba, 32'hbc00e84c} /* (0, 13, 11) {real, imag} */,
  {32'h3cfe5340, 32'hbc142254} /* (0, 13, 10) {real, imag} */,
  {32'h3d238e22, 32'hbd89bc62} /* (0, 13, 9) {real, imag} */,
  {32'hbd6b9362, 32'hbb23c250} /* (0, 13, 8) {real, imag} */,
  {32'hbc57b8fc, 32'h3c36f330} /* (0, 13, 7) {real, imag} */,
  {32'hbce2c599, 32'hbd6805fc} /* (0, 13, 6) {real, imag} */,
  {32'hbcf884bc, 32'hbde556e3} /* (0, 13, 5) {real, imag} */,
  {32'h3d953186, 32'h3dc61ea6} /* (0, 13, 4) {real, imag} */,
  {32'hbdbac1a0, 32'hbdaef856} /* (0, 13, 3) {real, imag} */,
  {32'hbe75592d, 32'h3c0e08c8} /* (0, 13, 2) {real, imag} */,
  {32'h3f2afca0, 32'h3e045110} /* (0, 13, 1) {real, imag} */,
  {32'h3e477f6b, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'h3f05d1ff, 32'hbdfee4dc} /* (0, 12, 31) {real, imag} */,
  {32'hbe5eed75, 32'h3d8da948} /* (0, 12, 30) {real, imag} */,
  {32'hbd28a15b, 32'h3c9d63c4} /* (0, 12, 29) {real, imag} */,
  {32'h3caaf036, 32'hbdcba6e2} /* (0, 12, 28) {real, imag} */,
  {32'h3cee1560, 32'h3d6d6d1c} /* (0, 12, 27) {real, imag} */,
  {32'h3d10435b, 32'h3d084c9a} /* (0, 12, 26) {real, imag} */,
  {32'hbc5ff468, 32'h3b0725b8} /* (0, 12, 25) {real, imag} */,
  {32'hbcacf29e, 32'h3cee23a1} /* (0, 12, 24) {real, imag} */,
  {32'h3d260008, 32'h3cc16a00} /* (0, 12, 23) {real, imag} */,
  {32'hbdb18909, 32'h3c21b77c} /* (0, 12, 22) {real, imag} */,
  {32'hbd12fbca, 32'h3d1389d5} /* (0, 12, 21) {real, imag} */,
  {32'hbdb2a0d0, 32'hbc2c9183} /* (0, 12, 20) {real, imag} */,
  {32'h3ca4c6de, 32'h3cbee5ec} /* (0, 12, 19) {real, imag} */,
  {32'hbd018664, 32'h3d0a18fc} /* (0, 12, 18) {real, imag} */,
  {32'h3d2ccfcf, 32'h3c1bddac} /* (0, 12, 17) {real, imag} */,
  {32'hbcecb6c2, 32'h00000000} /* (0, 12, 16) {real, imag} */,
  {32'h3d2ccfcf, 32'hbc1bddac} /* (0, 12, 15) {real, imag} */,
  {32'hbd018664, 32'hbd0a18fc} /* (0, 12, 14) {real, imag} */,
  {32'h3ca4c6de, 32'hbcbee5ec} /* (0, 12, 13) {real, imag} */,
  {32'hbdb2a0d0, 32'h3c2c9183} /* (0, 12, 12) {real, imag} */,
  {32'hbd12fbca, 32'hbd1389d5} /* (0, 12, 11) {real, imag} */,
  {32'hbdb18909, 32'hbc21b77c} /* (0, 12, 10) {real, imag} */,
  {32'h3d260008, 32'hbcc16a00} /* (0, 12, 9) {real, imag} */,
  {32'hbcacf29e, 32'hbcee23a1} /* (0, 12, 8) {real, imag} */,
  {32'hbc5ff468, 32'hbb0725b8} /* (0, 12, 7) {real, imag} */,
  {32'h3d10435b, 32'hbd084c9a} /* (0, 12, 6) {real, imag} */,
  {32'h3cee1560, 32'hbd6d6d1c} /* (0, 12, 5) {real, imag} */,
  {32'h3caaf036, 32'h3dcba6e2} /* (0, 12, 4) {real, imag} */,
  {32'hbd28a15b, 32'hbc9d63c4} /* (0, 12, 3) {real, imag} */,
  {32'hbe5eed75, 32'hbd8da948} /* (0, 12, 2) {real, imag} */,
  {32'h3f05d1ff, 32'h3dfee4dc} /* (0, 12, 1) {real, imag} */,
  {32'h3e65b1bc, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h3ec56c44, 32'hbd733e44} /* (0, 11, 31) {real, imag} */,
  {32'hbe6695ef, 32'h3db2079e} /* (0, 11, 30) {real, imag} */,
  {32'hbc6fa73c, 32'hbc4459a4} /* (0, 11, 29) {real, imag} */,
  {32'hbced9a5e, 32'hbe15a451} /* (0, 11, 28) {real, imag} */,
  {32'hbb975228, 32'h3c2c3710} /* (0, 11, 27) {real, imag} */,
  {32'h3ba4f898, 32'hbbe2c6fc} /* (0, 11, 26) {real, imag} */,
  {32'h39285b40, 32'h3d236a8e} /* (0, 11, 25) {real, imag} */,
  {32'h3c77313b, 32'h3c408494} /* (0, 11, 24) {real, imag} */,
  {32'h3cad0341, 32'h3d209e2c} /* (0, 11, 23) {real, imag} */,
  {32'hbd493922, 32'hbdb7d0f0} /* (0, 11, 22) {real, imag} */,
  {32'hbd97ba4a, 32'h3db47295} /* (0, 11, 21) {real, imag} */,
  {32'h3d7f959a, 32'hbd3ed354} /* (0, 11, 20) {real, imag} */,
  {32'h3c8ff65e, 32'hbcc928e6} /* (0, 11, 19) {real, imag} */,
  {32'h3cc11e14, 32'h3b78b290} /* (0, 11, 18) {real, imag} */,
  {32'hbc9bba2d, 32'h3ca081a0} /* (0, 11, 17) {real, imag} */,
  {32'hbcb8db17, 32'h00000000} /* (0, 11, 16) {real, imag} */,
  {32'hbc9bba2d, 32'hbca081a0} /* (0, 11, 15) {real, imag} */,
  {32'h3cc11e14, 32'hbb78b290} /* (0, 11, 14) {real, imag} */,
  {32'h3c8ff65e, 32'h3cc928e6} /* (0, 11, 13) {real, imag} */,
  {32'h3d7f959a, 32'h3d3ed354} /* (0, 11, 12) {real, imag} */,
  {32'hbd97ba4a, 32'hbdb47295} /* (0, 11, 11) {real, imag} */,
  {32'hbd493922, 32'h3db7d0f0} /* (0, 11, 10) {real, imag} */,
  {32'h3cad0341, 32'hbd209e2c} /* (0, 11, 9) {real, imag} */,
  {32'h3c77313b, 32'hbc408494} /* (0, 11, 8) {real, imag} */,
  {32'h39285b40, 32'hbd236a8e} /* (0, 11, 7) {real, imag} */,
  {32'h3ba4f898, 32'h3be2c6fc} /* (0, 11, 6) {real, imag} */,
  {32'hbb975228, 32'hbc2c3710} /* (0, 11, 5) {real, imag} */,
  {32'hbced9a5e, 32'h3e15a451} /* (0, 11, 4) {real, imag} */,
  {32'hbc6fa73c, 32'h3c4459a4} /* (0, 11, 3) {real, imag} */,
  {32'hbe6695ef, 32'hbdb2079e} /* (0, 11, 2) {real, imag} */,
  {32'h3ec56c44, 32'h3d733e44} /* (0, 11, 1) {real, imag} */,
  {32'h3d208620, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h3d6f3904, 32'h3d071956} /* (0, 10, 31) {real, imag} */,
  {32'h3dd8c5ea, 32'h3daede09} /* (0, 10, 30) {real, imag} */,
  {32'hbd852448, 32'hbd73bd8f} /* (0, 10, 29) {real, imag} */,
  {32'hbd12f00a, 32'hbc931898} /* (0, 10, 28) {real, imag} */,
  {32'h3d6ca2ae, 32'hbd99dfce} /* (0, 10, 27) {real, imag} */,
  {32'hbd478ece, 32'hbce1b279} /* (0, 10, 26) {real, imag} */,
  {32'hbcc77988, 32'h3da4c536} /* (0, 10, 25) {real, imag} */,
  {32'h3dd178ac, 32'hbc3d756e} /* (0, 10, 24) {real, imag} */,
  {32'h3d2ba17e, 32'hbc899d3c} /* (0, 10, 23) {real, imag} */,
  {32'h3dea34b8, 32'h3c3982aa} /* (0, 10, 22) {real, imag} */,
  {32'h3c160a4e, 32'hbd784646} /* (0, 10, 21) {real, imag} */,
  {32'hbc966992, 32'h3d45ec58} /* (0, 10, 20) {real, imag} */,
  {32'hbaeb0d68, 32'hbca22146} /* (0, 10, 19) {real, imag} */,
  {32'hbdcda4c7, 32'hbd3eff91} /* (0, 10, 18) {real, imag} */,
  {32'hbc978cfa, 32'h3b3cc840} /* (0, 10, 17) {real, imag} */,
  {32'h3dc2355b, 32'h00000000} /* (0, 10, 16) {real, imag} */,
  {32'hbc978cfa, 32'hbb3cc840} /* (0, 10, 15) {real, imag} */,
  {32'hbdcda4c7, 32'h3d3eff91} /* (0, 10, 14) {real, imag} */,
  {32'hbaeb0d68, 32'h3ca22146} /* (0, 10, 13) {real, imag} */,
  {32'hbc966992, 32'hbd45ec58} /* (0, 10, 12) {real, imag} */,
  {32'h3c160a4e, 32'h3d784646} /* (0, 10, 11) {real, imag} */,
  {32'h3dea34b8, 32'hbc3982aa} /* (0, 10, 10) {real, imag} */,
  {32'h3d2ba17e, 32'h3c899d3c} /* (0, 10, 9) {real, imag} */,
  {32'h3dd178ac, 32'h3c3d756e} /* (0, 10, 8) {real, imag} */,
  {32'hbcc77988, 32'hbda4c536} /* (0, 10, 7) {real, imag} */,
  {32'hbd478ece, 32'h3ce1b279} /* (0, 10, 6) {real, imag} */,
  {32'h3d6ca2ae, 32'h3d99dfce} /* (0, 10, 5) {real, imag} */,
  {32'hbd12f00a, 32'h3c931898} /* (0, 10, 4) {real, imag} */,
  {32'hbd852448, 32'h3d73bd8f} /* (0, 10, 3) {real, imag} */,
  {32'h3dd8c5ea, 32'hbdaede09} /* (0, 10, 2) {real, imag} */,
  {32'h3d6f3904, 32'hbd071956} /* (0, 10, 1) {real, imag} */,
  {32'hbe95ee72, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'hbe328cb8, 32'h3e173d1a} /* (0, 9, 31) {real, imag} */,
  {32'h3e10dd07, 32'hbcab9f16} /* (0, 9, 30) {real, imag} */,
  {32'h39c7b500, 32'h3b1c0a18} /* (0, 9, 29) {real, imag} */,
  {32'hbd39e70f, 32'h3d6d0f3e} /* (0, 9, 28) {real, imag} */,
  {32'h3d335af7, 32'hbe002be2} /* (0, 9, 27) {real, imag} */,
  {32'hbcf961b4, 32'h3ca87cc6} /* (0, 9, 26) {real, imag} */,
  {32'hbd3f8e45, 32'h3c3173c4} /* (0, 9, 25) {real, imag} */,
  {32'h3d1e7296, 32'hbd24917c} /* (0, 9, 24) {real, imag} */,
  {32'hb99d6540, 32'hbc8f731d} /* (0, 9, 23) {real, imag} */,
  {32'hbd0c636a, 32'hbcade4be} /* (0, 9, 22) {real, imag} */,
  {32'h3dbb8a76, 32'hbd46a202} /* (0, 9, 21) {real, imag} */,
  {32'h3cc8fa21, 32'h3c694884} /* (0, 9, 20) {real, imag} */,
  {32'hbd7a0bf0, 32'hbc1b369f} /* (0, 9, 19) {real, imag} */,
  {32'h3d3d11ef, 32'hb8d96700} /* (0, 9, 18) {real, imag} */,
  {32'hbc832db0, 32'hbd1f4e38} /* (0, 9, 17) {real, imag} */,
  {32'h3b545210, 32'h00000000} /* (0, 9, 16) {real, imag} */,
  {32'hbc832db0, 32'h3d1f4e38} /* (0, 9, 15) {real, imag} */,
  {32'h3d3d11ef, 32'h38d96700} /* (0, 9, 14) {real, imag} */,
  {32'hbd7a0bf0, 32'h3c1b369f} /* (0, 9, 13) {real, imag} */,
  {32'h3cc8fa21, 32'hbc694884} /* (0, 9, 12) {real, imag} */,
  {32'h3dbb8a76, 32'h3d46a202} /* (0, 9, 11) {real, imag} */,
  {32'hbd0c636a, 32'h3cade4be} /* (0, 9, 10) {real, imag} */,
  {32'hb99d6540, 32'h3c8f731d} /* (0, 9, 9) {real, imag} */,
  {32'h3d1e7296, 32'h3d24917c} /* (0, 9, 8) {real, imag} */,
  {32'hbd3f8e45, 32'hbc3173c4} /* (0, 9, 7) {real, imag} */,
  {32'hbcf961b4, 32'hbca87cc6} /* (0, 9, 6) {real, imag} */,
  {32'h3d335af7, 32'h3e002be2} /* (0, 9, 5) {real, imag} */,
  {32'hbd39e70f, 32'hbd6d0f3e} /* (0, 9, 4) {real, imag} */,
  {32'h39c7b500, 32'hbb1c0a18} /* (0, 9, 3) {real, imag} */,
  {32'h3e10dd07, 32'h3cab9f16} /* (0, 9, 2) {real, imag} */,
  {32'hbe328cb8, 32'hbe173d1a} /* (0, 9, 1) {real, imag} */,
  {32'hbeb681ee, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'hbe99c9a0, 32'h3e6368c3} /* (0, 8, 31) {real, imag} */,
  {32'h3e58b519, 32'hbbb75240} /* (0, 8, 30) {real, imag} */,
  {32'hbd32ffc5, 32'hbd85e444} /* (0, 8, 29) {real, imag} */,
  {32'hbd3d2488, 32'hbd4e1e18} /* (0, 8, 28) {real, imag} */,
  {32'h3d44d291, 32'hbcecff0a} /* (0, 8, 27) {real, imag} */,
  {32'hbc8324b4, 32'hbd8c3a13} /* (0, 8, 26) {real, imag} */,
  {32'hbcf94048, 32'h3ba75aec} /* (0, 8, 25) {real, imag} */,
  {32'h3d05b75b, 32'hbd5120d3} /* (0, 8, 24) {real, imag} */,
  {32'hbbe78a50, 32'h3be4a640} /* (0, 8, 23) {real, imag} */,
  {32'hbd35222a, 32'hbba06848} /* (0, 8, 22) {real, imag} */,
  {32'h3b5f2d40, 32'h3cc1e599} /* (0, 8, 21) {real, imag} */,
  {32'hbc1b6a62, 32'hbc4d33e1} /* (0, 8, 20) {real, imag} */,
  {32'h3cfd7255, 32'h3ca6cd89} /* (0, 8, 19) {real, imag} */,
  {32'h3bea1f2c, 32'h3b5ad660} /* (0, 8, 18) {real, imag} */,
  {32'hbc01751e, 32'hbd0ac3f7} /* (0, 8, 17) {real, imag} */,
  {32'hbc0dd17b, 32'h00000000} /* (0, 8, 16) {real, imag} */,
  {32'hbc01751e, 32'h3d0ac3f7} /* (0, 8, 15) {real, imag} */,
  {32'h3bea1f2c, 32'hbb5ad660} /* (0, 8, 14) {real, imag} */,
  {32'h3cfd7255, 32'hbca6cd89} /* (0, 8, 13) {real, imag} */,
  {32'hbc1b6a62, 32'h3c4d33e1} /* (0, 8, 12) {real, imag} */,
  {32'h3b5f2d40, 32'hbcc1e599} /* (0, 8, 11) {real, imag} */,
  {32'hbd35222a, 32'h3ba06848} /* (0, 8, 10) {real, imag} */,
  {32'hbbe78a50, 32'hbbe4a640} /* (0, 8, 9) {real, imag} */,
  {32'h3d05b75b, 32'h3d5120d3} /* (0, 8, 8) {real, imag} */,
  {32'hbcf94048, 32'hbba75aec} /* (0, 8, 7) {real, imag} */,
  {32'hbc8324b4, 32'h3d8c3a13} /* (0, 8, 6) {real, imag} */,
  {32'h3d44d291, 32'h3cecff0a} /* (0, 8, 5) {real, imag} */,
  {32'hbd3d2488, 32'h3d4e1e18} /* (0, 8, 4) {real, imag} */,
  {32'hbd32ffc5, 32'h3d85e444} /* (0, 8, 3) {real, imag} */,
  {32'h3e58b519, 32'h3bb75240} /* (0, 8, 2) {real, imag} */,
  {32'hbe99c9a0, 32'hbe6368c3} /* (0, 8, 1) {real, imag} */,
  {32'hbeb2bb57, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'hbed95da4, 32'h3e4252e2} /* (0, 7, 31) {real, imag} */,
  {32'h3e7a708e, 32'h3c9bd0e8} /* (0, 7, 30) {real, imag} */,
  {32'h3be01550, 32'hbcc2524c} /* (0, 7, 29) {real, imag} */,
  {32'hbd7a416f, 32'hbde3c718} /* (0, 7, 28) {real, imag} */,
  {32'h3dafc4c4, 32'h3d735e6b} /* (0, 7, 27) {real, imag} */,
  {32'hbd8c6170, 32'hbd80ec00} /* (0, 7, 26) {real, imag} */,
  {32'h3ccf35dd, 32'hbd6da2ec} /* (0, 7, 25) {real, imag} */,
  {32'h3d88e301, 32'hbd0c8238} /* (0, 7, 24) {real, imag} */,
  {32'h3d6e8e9a, 32'h3d103279} /* (0, 7, 23) {real, imag} */,
  {32'h3c35fb43, 32'hbb81be00} /* (0, 7, 22) {real, imag} */,
  {32'h3d270d86, 32'hbc7b2c58} /* (0, 7, 21) {real, imag} */,
  {32'h3d0cfcf5, 32'h3d8ed8dc} /* (0, 7, 20) {real, imag} */,
  {32'h3d1016ca, 32'hbd668ce7} /* (0, 7, 19) {real, imag} */,
  {32'h3ca673a3, 32'hbb975c26} /* (0, 7, 18) {real, imag} */,
  {32'h3a84c4e0, 32'h3c96621a} /* (0, 7, 17) {real, imag} */,
  {32'h3c96b696, 32'h00000000} /* (0, 7, 16) {real, imag} */,
  {32'h3a84c4e0, 32'hbc96621a} /* (0, 7, 15) {real, imag} */,
  {32'h3ca673a3, 32'h3b975c26} /* (0, 7, 14) {real, imag} */,
  {32'h3d1016ca, 32'h3d668ce7} /* (0, 7, 13) {real, imag} */,
  {32'h3d0cfcf5, 32'hbd8ed8dc} /* (0, 7, 12) {real, imag} */,
  {32'h3d270d86, 32'h3c7b2c58} /* (0, 7, 11) {real, imag} */,
  {32'h3c35fb43, 32'h3b81be00} /* (0, 7, 10) {real, imag} */,
  {32'h3d6e8e9a, 32'hbd103279} /* (0, 7, 9) {real, imag} */,
  {32'h3d88e301, 32'h3d0c8238} /* (0, 7, 8) {real, imag} */,
  {32'h3ccf35dd, 32'h3d6da2ec} /* (0, 7, 7) {real, imag} */,
  {32'hbd8c6170, 32'h3d80ec00} /* (0, 7, 6) {real, imag} */,
  {32'h3dafc4c4, 32'hbd735e6b} /* (0, 7, 5) {real, imag} */,
  {32'hbd7a416f, 32'h3de3c718} /* (0, 7, 4) {real, imag} */,
  {32'h3be01550, 32'h3cc2524c} /* (0, 7, 3) {real, imag} */,
  {32'h3e7a708e, 32'hbc9bd0e8} /* (0, 7, 2) {real, imag} */,
  {32'hbed95da4, 32'hbe4252e2} /* (0, 7, 1) {real, imag} */,
  {32'hbee4a1ff, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'hbec39e14, 32'h3e84d214} /* (0, 6, 31) {real, imag} */,
  {32'h3eb0ed1e, 32'h3dc8de3b} /* (0, 6, 30) {real, imag} */,
  {32'h3db20232, 32'hbcf46dee} /* (0, 6, 29) {real, imag} */,
  {32'hbdb12354, 32'hbca9b674} /* (0, 6, 28) {real, imag} */,
  {32'h3dad97ea, 32'h3c1f27f4} /* (0, 6, 27) {real, imag} */,
  {32'hbcd417f9, 32'hbd115142} /* (0, 6, 26) {real, imag} */,
  {32'hbd08a6f6, 32'h3d193832} /* (0, 6, 25) {real, imag} */,
  {32'hbb3356a0, 32'hbd756198} /* (0, 6, 24) {real, imag} */,
  {32'h3c8ecd7c, 32'hbc1e9a26} /* (0, 6, 23) {real, imag} */,
  {32'hbcbce11e, 32'h3df9a577} /* (0, 6, 22) {real, imag} */,
  {32'h3d8d86d0, 32'hbcdbaca2} /* (0, 6, 21) {real, imag} */,
  {32'hbd84123a, 32'h3ccec01c} /* (0, 6, 20) {real, imag} */,
  {32'h3d301b92, 32'h3d1dc658} /* (0, 6, 19) {real, imag} */,
  {32'h3d66d4a0, 32'h3b6f965e} /* (0, 6, 18) {real, imag} */,
  {32'hbd207ada, 32'hbd15445a} /* (0, 6, 17) {real, imag} */,
  {32'hbd233935, 32'h00000000} /* (0, 6, 16) {real, imag} */,
  {32'hbd207ada, 32'h3d15445a} /* (0, 6, 15) {real, imag} */,
  {32'h3d66d4a0, 32'hbb6f965e} /* (0, 6, 14) {real, imag} */,
  {32'h3d301b92, 32'hbd1dc658} /* (0, 6, 13) {real, imag} */,
  {32'hbd84123a, 32'hbccec01c} /* (0, 6, 12) {real, imag} */,
  {32'h3d8d86d0, 32'h3cdbaca2} /* (0, 6, 11) {real, imag} */,
  {32'hbcbce11e, 32'hbdf9a577} /* (0, 6, 10) {real, imag} */,
  {32'h3c8ecd7c, 32'h3c1e9a26} /* (0, 6, 9) {real, imag} */,
  {32'hbb3356a0, 32'h3d756198} /* (0, 6, 8) {real, imag} */,
  {32'hbd08a6f6, 32'hbd193832} /* (0, 6, 7) {real, imag} */,
  {32'hbcd417f9, 32'h3d115142} /* (0, 6, 6) {real, imag} */,
  {32'h3dad97ea, 32'hbc1f27f4} /* (0, 6, 5) {real, imag} */,
  {32'hbdb12354, 32'h3ca9b674} /* (0, 6, 4) {real, imag} */,
  {32'h3db20232, 32'h3cf46dee} /* (0, 6, 3) {real, imag} */,
  {32'h3eb0ed1e, 32'hbdc8de3b} /* (0, 6, 2) {real, imag} */,
  {32'hbec39e14, 32'hbe84d214} /* (0, 6, 1) {real, imag} */,
  {32'hbf07327b, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hbe8feea2, 32'h3ef730f0} /* (0, 5, 31) {real, imag} */,
  {32'h3d361de8, 32'h3db4c4c0} /* (0, 5, 30) {real, imag} */,
  {32'h3deec432, 32'h3bbe72f8} /* (0, 5, 29) {real, imag} */,
  {32'hbc9417f6, 32'hbc9c4000} /* (0, 5, 28) {real, imag} */,
  {32'h3dcdaccd, 32'h3c920572} /* (0, 5, 27) {real, imag} */,
  {32'hbd2a187f, 32'hbdceb9bc} /* (0, 5, 26) {real, imag} */,
  {32'h3c2df3b8, 32'hbcf9d8ca} /* (0, 5, 25) {real, imag} */,
  {32'hbce686e6, 32'h3cd55cab} /* (0, 5, 24) {real, imag} */,
  {32'h3d5b052b, 32'h3dad5d4a} /* (0, 5, 23) {real, imag} */,
  {32'h3cb8c385, 32'hbc4d5ff8} /* (0, 5, 22) {real, imag} */,
  {32'h3b32eb78, 32'hbd1d60d3} /* (0, 5, 21) {real, imag} */,
  {32'h3d8e9720, 32'hbd705738} /* (0, 5, 20) {real, imag} */,
  {32'h3be1ae56, 32'hbcb8a10e} /* (0, 5, 19) {real, imag} */,
  {32'h3d076219, 32'h3ce10fd6} /* (0, 5, 18) {real, imag} */,
  {32'hbc10cc82, 32'h3b2cb040} /* (0, 5, 17) {real, imag} */,
  {32'h3d801440, 32'h00000000} /* (0, 5, 16) {real, imag} */,
  {32'hbc10cc82, 32'hbb2cb040} /* (0, 5, 15) {real, imag} */,
  {32'h3d076219, 32'hbce10fd6} /* (0, 5, 14) {real, imag} */,
  {32'h3be1ae56, 32'h3cb8a10e} /* (0, 5, 13) {real, imag} */,
  {32'h3d8e9720, 32'h3d705738} /* (0, 5, 12) {real, imag} */,
  {32'h3b32eb78, 32'h3d1d60d3} /* (0, 5, 11) {real, imag} */,
  {32'h3cb8c385, 32'h3c4d5ff8} /* (0, 5, 10) {real, imag} */,
  {32'h3d5b052b, 32'hbdad5d4a} /* (0, 5, 9) {real, imag} */,
  {32'hbce686e6, 32'hbcd55cab} /* (0, 5, 8) {real, imag} */,
  {32'h3c2df3b8, 32'h3cf9d8ca} /* (0, 5, 7) {real, imag} */,
  {32'hbd2a187f, 32'h3dceb9bc} /* (0, 5, 6) {real, imag} */,
  {32'h3dcdaccd, 32'hbc920572} /* (0, 5, 5) {real, imag} */,
  {32'hbc9417f6, 32'h3c9c4000} /* (0, 5, 4) {real, imag} */,
  {32'h3deec432, 32'hbbbe72f8} /* (0, 5, 3) {real, imag} */,
  {32'h3d361de8, 32'hbdb4c4c0} /* (0, 5, 2) {real, imag} */,
  {32'hbe8feea2, 32'hbef730f0} /* (0, 5, 1) {real, imag} */,
  {32'hbf5143bc, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hbe973c29, 32'h3f1b355f} /* (0, 4, 31) {real, imag} */,
  {32'hbde6090a, 32'hbcffde1e} /* (0, 4, 30) {real, imag} */,
  {32'h3dba47e8, 32'h3d461bcf} /* (0, 4, 29) {real, imag} */,
  {32'h3d582505, 32'hbde57123} /* (0, 4, 28) {real, imag} */,
  {32'h3daa81e6, 32'h3da55a43} /* (0, 4, 27) {real, imag} */,
  {32'hbc8cb7a0, 32'hbdac4c22} /* (0, 4, 26) {real, imag} */,
  {32'hb74c2c00, 32'hbc356755} /* (0, 4, 25) {real, imag} */,
  {32'hbdccbed6, 32'h3ac7a340} /* (0, 4, 24) {real, imag} */,
  {32'h3dc175aa, 32'hbc0722d6} /* (0, 4, 23) {real, imag} */,
  {32'hbcfcc1f5, 32'h3c859eda} /* (0, 4, 22) {real, imag} */,
  {32'h3de34640, 32'h3d31d8b4} /* (0, 4, 21) {real, imag} */,
  {32'hbca05e9e, 32'h3c667dd8} /* (0, 4, 20) {real, imag} */,
  {32'h3bff31f8, 32'hb9e93e00} /* (0, 4, 19) {real, imag} */,
  {32'h3d7ea882, 32'hbd9dd3db} /* (0, 4, 18) {real, imag} */,
  {32'hbb9d164d, 32'hbcf4ac3b} /* (0, 4, 17) {real, imag} */,
  {32'hbce0631a, 32'h00000000} /* (0, 4, 16) {real, imag} */,
  {32'hbb9d164d, 32'h3cf4ac3b} /* (0, 4, 15) {real, imag} */,
  {32'h3d7ea882, 32'h3d9dd3db} /* (0, 4, 14) {real, imag} */,
  {32'h3bff31f8, 32'h39e93e00} /* (0, 4, 13) {real, imag} */,
  {32'hbca05e9e, 32'hbc667dd8} /* (0, 4, 12) {real, imag} */,
  {32'h3de34640, 32'hbd31d8b4} /* (0, 4, 11) {real, imag} */,
  {32'hbcfcc1f5, 32'hbc859eda} /* (0, 4, 10) {real, imag} */,
  {32'h3dc175aa, 32'h3c0722d6} /* (0, 4, 9) {real, imag} */,
  {32'hbdccbed6, 32'hbac7a340} /* (0, 4, 8) {real, imag} */,
  {32'hb74c2c00, 32'h3c356755} /* (0, 4, 7) {real, imag} */,
  {32'hbc8cb7a0, 32'h3dac4c22} /* (0, 4, 6) {real, imag} */,
  {32'h3daa81e6, 32'hbda55a43} /* (0, 4, 5) {real, imag} */,
  {32'h3d582505, 32'h3de57123} /* (0, 4, 4) {real, imag} */,
  {32'h3dba47e8, 32'hbd461bcf} /* (0, 4, 3) {real, imag} */,
  {32'hbde6090a, 32'h3cffde1e} /* (0, 4, 2) {real, imag} */,
  {32'hbe973c29, 32'hbf1b355f} /* (0, 4, 1) {real, imag} */,
  {32'hbf38b5b0, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hbe74df4b, 32'h3f1edb82} /* (0, 3, 31) {real, imag} */,
  {32'hbda0216d, 32'hbe414ad2} /* (0, 3, 30) {real, imag} */,
  {32'h3de36777, 32'h3cc20278} /* (0, 3, 29) {real, imag} */,
  {32'hbdbd3ea3, 32'hbe1d38a0} /* (0, 3, 28) {real, imag} */,
  {32'h3d9a4f81, 32'h3dc5eb6e} /* (0, 3, 27) {real, imag} */,
  {32'h3d55ef14, 32'hbc94666f} /* (0, 3, 26) {real, imag} */,
  {32'hbcb526aa, 32'hbbdb72a0} /* (0, 3, 25) {real, imag} */,
  {32'h3ad15620, 32'hbca08f65} /* (0, 3, 24) {real, imag} */,
  {32'hbbc535ae, 32'h3c9c0590} /* (0, 3, 23) {real, imag} */,
  {32'h3c789ea6, 32'h3ced1f54} /* (0, 3, 22) {real, imag} */,
  {32'h3d3b9708, 32'hbd1d4bf4} /* (0, 3, 21) {real, imag} */,
  {32'h3c9a6544, 32'hbc74f320} /* (0, 3, 20) {real, imag} */,
  {32'h3cf523f2, 32'hbd041ce0} /* (0, 3, 19) {real, imag} */,
  {32'h3c8579e2, 32'h3d02e222} /* (0, 3, 18) {real, imag} */,
  {32'h3b315c6c, 32'hbcff2680} /* (0, 3, 17) {real, imag} */,
  {32'hbca162f3, 32'h00000000} /* (0, 3, 16) {real, imag} */,
  {32'h3b315c6c, 32'h3cff2680} /* (0, 3, 15) {real, imag} */,
  {32'h3c8579e2, 32'hbd02e222} /* (0, 3, 14) {real, imag} */,
  {32'h3cf523f2, 32'h3d041ce0} /* (0, 3, 13) {real, imag} */,
  {32'h3c9a6544, 32'h3c74f320} /* (0, 3, 12) {real, imag} */,
  {32'h3d3b9708, 32'h3d1d4bf4} /* (0, 3, 11) {real, imag} */,
  {32'h3c789ea6, 32'hbced1f54} /* (0, 3, 10) {real, imag} */,
  {32'hbbc535ae, 32'hbc9c0590} /* (0, 3, 9) {real, imag} */,
  {32'h3ad15620, 32'h3ca08f65} /* (0, 3, 8) {real, imag} */,
  {32'hbcb526aa, 32'h3bdb72a0} /* (0, 3, 7) {real, imag} */,
  {32'h3d55ef14, 32'h3c94666f} /* (0, 3, 6) {real, imag} */,
  {32'h3d9a4f81, 32'hbdc5eb6e} /* (0, 3, 5) {real, imag} */,
  {32'hbdbd3ea3, 32'h3e1d38a0} /* (0, 3, 4) {real, imag} */,
  {32'h3de36777, 32'hbcc20278} /* (0, 3, 3) {real, imag} */,
  {32'hbda0216d, 32'h3e414ad2} /* (0, 3, 2) {real, imag} */,
  {32'hbe74df4b, 32'hbf1edb82} /* (0, 3, 1) {real, imag} */,
  {32'hbf35cbf0, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hbe93601c, 32'h3f0893be} /* (0, 2, 31) {real, imag} */,
  {32'hbe38e96b, 32'hbe3a2778} /* (0, 2, 30) {real, imag} */,
  {32'h3e3799cc, 32'h3d0f5f63} /* (0, 2, 29) {real, imag} */,
  {32'hbdaaceac, 32'hbdb51238} /* (0, 2, 28) {real, imag} */,
  {32'h3d4bd838, 32'h3d956507} /* (0, 2, 27) {real, imag} */,
  {32'hb9d34f80, 32'h3c194974} /* (0, 2, 26) {real, imag} */,
  {32'hbd69b9f0, 32'h3dc7db0f} /* (0, 2, 25) {real, imag} */,
  {32'hbb417a98, 32'h3c82bc84} /* (0, 2, 24) {real, imag} */,
  {32'h3cf007b4, 32'hbd28ecf1} /* (0, 2, 23) {real, imag} */,
  {32'hbc9e0558, 32'h3c6e0990} /* (0, 2, 22) {real, imag} */,
  {32'hbb745ff0, 32'hbc67cd70} /* (0, 2, 21) {real, imag} */,
  {32'h3cbdcc2e, 32'h3c858286} /* (0, 2, 20) {real, imag} */,
  {32'hbd318da0, 32'h3d2332b6} /* (0, 2, 19) {real, imag} */,
  {32'hbccc2006, 32'h3cd41492} /* (0, 2, 18) {real, imag} */,
  {32'h3d00aa96, 32'h3c10172c} /* (0, 2, 17) {real, imag} */,
  {32'hbcdb4f51, 32'h00000000} /* (0, 2, 16) {real, imag} */,
  {32'h3d00aa96, 32'hbc10172c} /* (0, 2, 15) {real, imag} */,
  {32'hbccc2006, 32'hbcd41492} /* (0, 2, 14) {real, imag} */,
  {32'hbd318da0, 32'hbd2332b6} /* (0, 2, 13) {real, imag} */,
  {32'h3cbdcc2e, 32'hbc858286} /* (0, 2, 12) {real, imag} */,
  {32'hbb745ff0, 32'h3c67cd70} /* (0, 2, 11) {real, imag} */,
  {32'hbc9e0558, 32'hbc6e0990} /* (0, 2, 10) {real, imag} */,
  {32'h3cf007b4, 32'h3d28ecf1} /* (0, 2, 9) {real, imag} */,
  {32'hbb417a98, 32'hbc82bc84} /* (0, 2, 8) {real, imag} */,
  {32'hbd69b9f0, 32'hbdc7db0f} /* (0, 2, 7) {real, imag} */,
  {32'hb9d34f80, 32'hbc194974} /* (0, 2, 6) {real, imag} */,
  {32'h3d4bd838, 32'hbd956507} /* (0, 2, 5) {real, imag} */,
  {32'hbdaaceac, 32'h3db51238} /* (0, 2, 4) {real, imag} */,
  {32'h3e3799cc, 32'hbd0f5f63} /* (0, 2, 3) {real, imag} */,
  {32'hbe38e96b, 32'h3e3a2778} /* (0, 2, 2) {real, imag} */,
  {32'hbe93601c, 32'hbf0893be} /* (0, 2, 1) {real, imag} */,
  {32'hbee75dbd, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hbeaaab64, 32'h3f051d4e} /* (0, 1, 31) {real, imag} */,
  {32'hbe94214d, 32'hbe30e42e} /* (0, 1, 30) {real, imag} */,
  {32'h3e1871ed, 32'hbd6d5f25} /* (0, 1, 29) {real, imag} */,
  {32'h3d401d3b, 32'hbde1d84b} /* (0, 1, 28) {real, imag} */,
  {32'h3e07a697, 32'h3d933747} /* (0, 1, 27) {real, imag} */,
  {32'hbca6dc20, 32'h3cfb7c9f} /* (0, 1, 26) {real, imag} */,
  {32'hbd3f75e7, 32'h3d919701} /* (0, 1, 25) {real, imag} */,
  {32'h3ade3b40, 32'hbd8cbce1} /* (0, 1, 24) {real, imag} */,
  {32'h3d072930, 32'hbbbed78c} /* (0, 1, 23) {real, imag} */,
  {32'hbcf8d176, 32'h3d072126} /* (0, 1, 22) {real, imag} */,
  {32'h3d602b36, 32'hbb7cb512} /* (0, 1, 21) {real, imag} */,
  {32'hbd0a73ed, 32'h3d441240} /* (0, 1, 20) {real, imag} */,
  {32'hbd828243, 32'hbc9e310d} /* (0, 1, 19) {real, imag} */,
  {32'hbd2f7255, 32'hbd4845a4} /* (0, 1, 18) {real, imag} */,
  {32'h3d2e61f0, 32'hbd36fc0d} /* (0, 1, 17) {real, imag} */,
  {32'h3d2dd2ab, 32'h00000000} /* (0, 1, 16) {real, imag} */,
  {32'h3d2e61f0, 32'h3d36fc0d} /* (0, 1, 15) {real, imag} */,
  {32'hbd2f7255, 32'h3d4845a4} /* (0, 1, 14) {real, imag} */,
  {32'hbd828243, 32'h3c9e310d} /* (0, 1, 13) {real, imag} */,
  {32'hbd0a73ed, 32'hbd441240} /* (0, 1, 12) {real, imag} */,
  {32'h3d602b36, 32'h3b7cb512} /* (0, 1, 11) {real, imag} */,
  {32'hbcf8d176, 32'hbd072126} /* (0, 1, 10) {real, imag} */,
  {32'h3d072930, 32'h3bbed78c} /* (0, 1, 9) {real, imag} */,
  {32'h3ade3b40, 32'h3d8cbce1} /* (0, 1, 8) {real, imag} */,
  {32'hbd3f75e7, 32'hbd919701} /* (0, 1, 7) {real, imag} */,
  {32'hbca6dc20, 32'hbcfb7c9f} /* (0, 1, 6) {real, imag} */,
  {32'h3e07a697, 32'hbd933747} /* (0, 1, 5) {real, imag} */,
  {32'h3d401d3b, 32'h3de1d84b} /* (0, 1, 4) {real, imag} */,
  {32'h3e1871ed, 32'h3d6d5f25} /* (0, 1, 3) {real, imag} */,
  {32'hbe94214d, 32'h3e30e42e} /* (0, 1, 2) {real, imag} */,
  {32'hbeaaab64, 32'hbf051d4e} /* (0, 1, 1) {real, imag} */,
  {32'hbe89dbcb, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hbeb70e86, 32'h3eab0c49} /* (0, 0, 31) {real, imag} */,
  {32'hbe0917e2, 32'hbd580336} /* (0, 0, 30) {real, imag} */,
  {32'h3d77f3d7, 32'h3d210366} /* (0, 0, 29) {real, imag} */,
  {32'h3d3ca4e4, 32'hbd9538dd} /* (0, 0, 28) {real, imag} */,
  {32'h3e01daf9, 32'h3cf04d7e} /* (0, 0, 27) {real, imag} */,
  {32'hbc82e4a6, 32'h3c251c9b} /* (0, 0, 26) {real, imag} */,
  {32'h3d0e55d6, 32'h3cb1a050} /* (0, 0, 25) {real, imag} */,
  {32'h3c2a9dba, 32'hbb782400} /* (0, 0, 24) {real, imag} */,
  {32'h3d517b5a, 32'hbb3c65d0} /* (0, 0, 23) {real, imag} */,
  {32'hbd5d6380, 32'hbcb9e944} /* (0, 0, 22) {real, imag} */,
  {32'h3c180d26, 32'hbce228d1} /* (0, 0, 21) {real, imag} */,
  {32'hbcba4f48, 32'h3cba516d} /* (0, 0, 20) {real, imag} */,
  {32'h3d09db67, 32'h3d6b51e4} /* (0, 0, 19) {real, imag} */,
  {32'hbc96b7a5, 32'h3d2bda54} /* (0, 0, 18) {real, imag} */,
  {32'h3c0f4220, 32'h3b26c440} /* (0, 0, 17) {real, imag} */,
  {32'h3c479af4, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'h3c0f4220, 32'hbb26c440} /* (0, 0, 15) {real, imag} */,
  {32'hbc96b7a5, 32'hbd2bda54} /* (0, 0, 14) {real, imag} */,
  {32'h3d09db67, 32'hbd6b51e4} /* (0, 0, 13) {real, imag} */,
  {32'hbcba4f48, 32'hbcba516d} /* (0, 0, 12) {real, imag} */,
  {32'h3c180d26, 32'h3ce228d1} /* (0, 0, 11) {real, imag} */,
  {32'hbd5d6380, 32'h3cb9e944} /* (0, 0, 10) {real, imag} */,
  {32'h3d517b5a, 32'h3b3c65d0} /* (0, 0, 9) {real, imag} */,
  {32'h3c2a9dba, 32'h3b782400} /* (0, 0, 8) {real, imag} */,
  {32'h3d0e55d6, 32'hbcb1a050} /* (0, 0, 7) {real, imag} */,
  {32'hbc82e4a6, 32'hbc251c9b} /* (0, 0, 6) {real, imag} */,
  {32'h3e01daf9, 32'hbcf04d7e} /* (0, 0, 5) {real, imag} */,
  {32'h3d3ca4e4, 32'h3d9538dd} /* (0, 0, 4) {real, imag} */,
  {32'h3d77f3d7, 32'hbd210366} /* (0, 0, 3) {real, imag} */,
  {32'hbe0917e2, 32'h3d580336} /* (0, 0, 2) {real, imag} */,
  {32'hbeb70e86, 32'hbeab0c49} /* (0, 0, 1) {real, imag} */,
  {32'hbe72fd9b, 32'h00000000} /* (0, 0, 0) {real, imag} */};
