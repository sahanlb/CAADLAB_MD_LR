-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1U0Mb4eQ7rhboH0VlJVPRrlw4hdKWFSCtSzhutx3EK3Ch5lSJnMul9W6k1l91iKN
jV2Q+pkTWnxft+jCzmIkbdE5lXbM3Aug+SkTmPUw8eYYWgaceuYwHnZXNKE2sH5r
Iqy13WjyhnWPG+Oje3OAEwpNbUTHaDR5UR7S3ZUtA/c=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6832)
`protect data_block
dUbRD+O74e8HMXuzXX/PLWdaiH6y35ZgDLb9gY7siBpIzZwer6GbbT4sHJ62ELCU
wMM4XRxXIsjm0HOcavoAy9R5OdIC1rIeHozAU7iQfGcQBEK3XPShF5CKAwXz8NFr
jsJTl7ifAU60cmqGTu0N91D4lha1GDKB8CK0gYIStwJljkzoZpwD/mbMqwB7XGfn
CRuMuVKN1hnjp4FGiOfeGlm1pdNb8WNiQZeNY5by9LAhHLVXU0FFbAicYUbUPSPz
K6NenL+Le5uOQ/8nvhxKhoIcd3959Hhj78chDokLO4N14eUY1Vyld3+keFDEZqu4
e2P74BS/bXbJBi6RcJHDTstUwX59o5m1TVJwgmOZxcmAz+Mseyw9pcTNVVfzXt4x
yJ5cEWsc+o6xS9LpOgP+nBRJflg/rKrGcbFx98MFLnq/xZ7UFYCnAKYI5pCIsYJW
+kKfexV3h8VWV7N9F1uNkdf/XVSn0u+Q1daHFO4ix5C2fAwDHv2/TgI7LLcNVrBE
gL/prXTBKMiHCX0SsjCIcJY/86Z4pFRB6j1dfutVlUqddtT7qtRzacRR5upJbN1l
FBJP6sejfINFNKFZ+aiG912bUHvL3PGQEfsrm4I3kxI7L3iN/94qAhd1/ko3/Y17
6roUwd1TUWUHGrqGPi5mwwzqdVARyckxfuuWwQmxLKU0fun717UIahU2Q1d7vFiZ
6BcGcluPdhQBkO6CbGdgFU/Fqq82Kvhp3+lcCNh5eAYe7yFze97KFsCpC++nLiV5
sM3IK2znf0Tn77vRnn70VZOWAu+jnRM0K9Ww031OXHdXL+uvuFOjBWCTDWu6hp7f
JzHzWxMukPNZ6+03zqdHbYipNl/2m6q7PiPOSCFmb/kzdrKvm+dcytTHFr9TBQpP
IrdlKCOHoR5Vrp6J6TlOF0aAlg70hR3ykqhnf2sH7cICxVom98atZNy/cZQ6f/dL
E//vJTD/HObcI8ytloXNuwe4il6DghmQ9PuMCDZxaefh/DmBeX9k0I1Fd3gx8K85
/octsoxvPbIDDosm1dsKi/3Im6dZNYwhhJInP/FR5Vdc0fWL9dsXcZlkN6DXCaq4
dktEwP4XJpqCOAFuqLzWd7oHKkH26h0uo1hiMy8XRvj6JhEET/Q2JjOIr2C7Kat8
HBP2+5cbEBIGxm1f1iBcUCFETmgis3jzn0S1zKroE6FBSoPq4LGlgiYa9M6411y5
/C8r+IW5ebq3VFAAfOEWHQ2E0syAOR4hfGLdbE79DMTlMjBX2TFG+XRYWL7DwgD5
yo9Y+0fsBPDTWwV0n8eB47vwqqKeDxRaJWRIiKdCtL8YSRb/fUKuNWOGQQDRiWDd
Kur2FAuCo8CLDJoehLBdG01PyFpYrXD63F4UQLEKZAFGDypMneMSkx1IYRm/3w7B
Do0358AyuM9Jzik9rlHPQ3n+NbMf4gS2qRMvR4tmoG7IECt+UCKr7zQ2eikZsYop
zzTqCO3DXLmbIyvB0GRm+P7g9f/Zv0KUIXgzr/R3oXjWKZXwG/hH7NAa97ZVp+eb
5DTAu7FgVmeOFYERU4n6BF7yxN5d2LMl+ioS4j0ky4oy1qs5o+ySIg9Mf9/5GPXB
B99yTciL6hWx/011Ly7FL7wyi00Zcf++aAeWT6LVCNP3IQuFXbEDFV+p5u3Itlr4
euctBdmQj6Vr+OhJN1XJZuTtcBYGkOmVUn0yMLnOM1Rw5ZkubamH5pYzBYfeDovb
4rMpZi+iCt8JID7/s7Zx2b4H+czyOqgfmbaG1TDgJuggfvQDX+CypSe1hvTXTGJS
aQwEucbnmg1N33JuEF+MobhkaCym/0H5elKJH6gQ2vWwnHoC8pTduoFYNWt26mEU
++h1d2dkzCUb2HySZ28rv9ThWYRdYmdghZ1nc/fDLMVrIJVLoPyg1ooS8NVENz6c
givKNFYgjgbOsYTixlLPsLDNJFwSVXGDZhRSCku2aeRtoJPpkVX32/Xg0Yrf0nhU
W0f+qpG/m1uT2FaJfFO7GmirPeGEa8uRxw5QRWSWDmUhAtmjJ6QRJ8m2TCfvSODp
++R+pNtXz9TirDIoGgKcuVDim2di2NyKs2odFehyOCT7rw7B5T3vzqIfUDp5kYBJ
S+/tAq5+EzX+Dpmev8InlZlzYWbx6+Z9Z9KG4JZ8qH2wgSJmZMWVDbZW9YkO3zNO
s7MDN3Ok7bHA8RrE2A24RPX4iGlSskxOCZ37f7dcxzufWsEnbKL5vgTkwtTUnA1P
XbJkwH98Hjq+xEekp5PGma2Cq3deLhTmAYeb/kxLeZxhh1h6Se+3jVxUIISw9ksr
8/AJm5AtBkvZuxmVUfRkIgwfREHISA/kPz5cYH6uDKTOL1fBa4rY74KAZHxsc2Lj
U5diywOOLgA3MkruiAyPgYVsBAm/r/JYobkC3r/ufd21xsajTAcYPDc7mInN1tQR
7Lpzyzd0wGDEeuQtMYTT3y/qE2K9oBQD5RxXowtwEEa2iOJcyixD/eaD2ms+LK4e
PrvaIBVdMSKQ5WU5wEeHrXo//sOpXTHl7WgmVoI/ZeO7j3tYk6Pang1HOKLioTS8
9Eak5V/5gPHRSjJUP7gW2mTedu1K9ouf4+c1BGEPcdHrr/VY2QR5UfC2+GMrtp5p
G2uHROx2jNolPSXGSg4rRgNfykKBQBsv7Q7MNorEG5sK1/DwqHiAVvsBxFaMuYl1
yGv6VTPAYpbRmrV0h1aLl/a8GRP/I2pBixr4UZCdx9M1jPwWpI3XJ8C/Fg+M3xAB
cSuZN9hoTjp7WTEhmTMVn6JsaKsEzLpjxXWY/D9C1fFkIdPBgy0Icmf4q0xrczPs
wKHeeufuSUuowQ1Ku9yWKpEV07+QDQ2fNaWggv9xdBbPRsDYncPvz2n13ioLFcCH
IpCAzzWDCJDsBuMVI8RUYaI0CNd1Wy7wZnP44emhIfMI8AlFVgoDQBkG5Fv6Ds7I
W5mokePXPaJ5ej2CsdaNAoeP60cRxPhQvqVjFT3Y/wHrPr6Hh+CEKiWVwyibjJ47
VH91/LGFNQxCPsXOglqZs+9+UFQ6Aj/0BR6yV+1fKEKdfFyWD1rtl4of87yp9jLE
fEbY/7y1q6e7n2nV89UdUnEWc7gzjXG8e/Z+ThfoV4B/j/thP18qhNGBPG7ts8ZJ
+uOKCgLp1YIfefvu6pfoaWd26ByO4rH/5Q9OnDudSr2NEg6OpryjhJFc4vDPHVJI
PAThExzVN9ZyNblkK4wd4bPXtVY0SLsEJuRWy0RIhHfls0TKTq5YxalomP0ip8MQ
T+BEl8EwhlR4rs0gsqavwQh+wX3AnxVZm3FHc7kkE/4DtfQk902JeERCygIpx4gV
NzyNsOBoDp10i5IhDQdH4n5n8VJi5hRAKvYHifTxpuf5/sLlzr+X6v2NDgW3B0il
EjAsU8FmxCNrbiDXrOH6zXvH2V6yj2ziG3vkhqzGKiKyx3Qy9aHOSmmLtSCcv12T
xuup8Gxit8zdAMtvLZn3SuS8cCGQcH3AznBaifHx0K1eh7DoFU4f16XmhHomq5pK
3pDX7gC2O1mOIvcxCkUChMSa2MZyoAswL3+6tX6eHsqlR8hzQs5RkNZKpOvnwYd2
9EpU8NUGgkJb1De7ocKWpTTzYg2g6DYvPSfvRznHEfEHffa4YWeXjoARz1S/hNz0
zI/fKAm/jr2LJQ0o8PEH/feklvXUBTBko0xrWlzdk09MtvNRJq7GrotytBS8rKNy
2PClJW5nU1zUvOOI98GAEsPrS1KYy1G2a4xkG7T4ZtpTYRe7GbS/qgPdvgo72ZXe
QUkuhJcpuOm75Sxm9BCI8/dEOvfBofyj7iTlxnjoNuOCM3Zgc9tAx/bZi3OGrtG+
DjGx+mgzoRqs7owMDDrylSr8dyhYjZjxSM5u7jwW6uNuG2MjWDVeFXsB02AkRdoo
l7Qjf+EhozbCmJTIB6XZRnPoP4BUn2/IOqj2HLd+01PClaQK29qDZgyyBZ+Lrm6G
Z0Ffqr+5OnQTtd8OcHfHPywrDfDdtOjP1mDvpQMHjPACp3s2rquFyw7zgK3hqovQ
pDbKR/3mRikRbB8V/ErH3wYa+1rJjW22GVUmxnoICVzMsDeGkEOdaKT4A75OWsao
xjJB5CfPBzLuhxHKhisgpb/o+Dy2n80vhpfy0ETHryXPiJ9R8h1yqyt/ISzRaP3W
s3ixQIx6KhiSz11lm16o4+/WFdxSPL4YG+LQDkEe1lWzwkAAbjXmFXl1pHAhe9Ys
UuHeNVOe/OZIWsVksc04bodjHIy5gqduYfzrBDwoz0eTzLVxwJQuxzOLiP/DPawJ
p7+kfS9lTbX71v2wlmAlol6C/ZYCUJudWdNaHUnB/zvomvNrr+cc1usxFX+dS8K6
kFBbpcEWy+gosye097H39wBO+N5Bvl494LCVtxMrpQ/Dj+jHndb6nWCQ8RyufoCl
CIqKlAqSqx7Wc7c2RqKy8G6PomF0mIkH3Sl2j6Ptprn/kdIi3KFkKngapEQwe7ES
+Ggt7SHMPmFWjHwnWTEEoan8umqu4HuTuTb3iy9aAajmiPRetwmBalMmiqWpzjqR
rkTuNYu6pyg8MVizaK0DeJXFXs9kPrh1MLtq7KcynbAK8ltbQ1mbsTpjqF0nPF0P
ITepcwTsUgI+F5nXZsn5VMLkzdKld038ZAjXYlKaMiGZkPuP3XubcJFjwyYooF9G
VVhxUxqN3USCrhgruYHYVEqk1AMjHJD/SqZVtIYrl+60QRli+7R83eq4bpjGM3mM
B71o9PbqYGvPGtFh7HD7Ly2H3MqbMXF67AYyiVzJLJUjYrH5JFCIv/Zu0WnHFAAK
2SsEaNKWDS7kQvVw1pEQ83l0Z/IocEDy9PhYqPaNtoON9s37ZjaXSewcweA670t7
UySkTFoxMxQ+CaUir2iK19xrv8EkkoBJRUv4hIJLiN9YvpsL2raEuK23Y38Pck3U
zlm1O1xlpbtDHROhq96qM7VPNjY7M9GTZLzN2cgb5+Wcbrdkyy5psX0nRRgWBuwP
uZL8cnwSN4Az88uUdDvcvTFw1A2tI/yDH+xcoc1etxMeyYcWdIBahokTpUOs1RiQ
MMUTNxCA2vxQ7LCwvE2Y9DFLJygbXD961vbaR73srcz5kafeTLcI6A69PDOTUWvZ
A6UOeE/GSECHKMa8UxiXx7IO/mRks23S3aR/rAAsxeCg7gf0b9VHTk7/LjJoPeWv
zkdjZJB2aFZteuiqcHxjsKZSmI1n6vvSaqX0X++G5UJ2rJ4K+aHfJqC37JUeqKpQ
ep+TnPZq/a0/Nsem9vEm+44HfhKQfB/DesbTfP6gzB24lWyGNaEL5xaMfxSrSQ4Q
DKw7EnA81jPsFs+FTg20WLRg+HslCxicZbf6NEPwP9j0MMxQsFpTfm8SgFT7p7dk
r/RfqnxzpupDZ2HyNS2z8fCB4dqYcesdEj/1oqb3Pw4YqDdVCdjgqa3BK38yHrHx
7nOG1vR/cvr+u/IIHAY+WTdHvxj7AgHZ4cN9k0of0DXashA5bhmTEBp+bJ9NPR7+
IqkBdkUnW9Dc5cujrRtzu//eFv30rV5CtsrSa1mYYxH4J/nfLmeRbhx09p3LkVnz
CtBQARah9T/qrk1F6Lb+DE18SQOo6TVPi/aBd0jXjNjVaGY+VaDtAu/xqFKVtQFk
Ws6vhmWtKNqZjGLkauenl0sMtCDoUjhCJmnfYOthTwj8pj+5tMoq1LU5SVNbT0vN
SpQPqWvrUAMWuLfLrgYMtEVPDqy4ujzM3S9sCFMs7/fyG/QFp4Arsc/hyJdJWM46
rF/AiIrs7dboV4lSM7BNO1TKdp8TJYKLC33YGnZ025FUJUyj1suYMszHlaFeSnH6
RNwuNnFPDmqSgtcJiupkHWisTCwICwFgj5D2mSiu5mpy2t7/JRtp5RU6WOMojS8F
Z1kP8C8pkT0nD0TAijZKm8NRkbjwGLe4WpO4Qmuy9tJysLHJczd002Abg0rVC0mD
iSz8MY9Kbsf/Ev9E4xPAElZuJHMVe8SqGXg9k91feIHdUeF3zrW9R9s2r57AQ5uC
yyijNHngROH720HQkZebm9qAOg/P9O+IVavOOZjcPzhGvo6w4DO8Diz2n5/gpfD1
uxQicHr+HJfwmxPnu58edlJt8lXqCWy0YJcLTYkHbPfc0kYGRhsQ/aeY/pR9jFVN
/eHVBWYkfWFN+MnjeH3XCt2FwGFhYotmPkUKkr/kXEh64i/MJeZU9zhjpVGa7eEo
ID1EArzS7LAK/VWZD3JSZBnMBGtyXuLWU4kLDBaMiNVrwDIT1o+Ko1AFf2v4XRJu
H//aYz/xmLj6jje0sZq2F3kVriYVbA1UL9h/IFBaYt/fKDulXuGr1x/SwU4/bZ64
ZFYSiNsTwpicMNZMhgtBJ9dqcoNeUEto8LNtREck0/eKtHStVvfo0M4UnSEsmRFD
cyJ+IG/OdC4wDG0+f1S5t4lmqskBTyuDPMQqbo2vFnSYRoeQPPVh4H73XePnjZJU
kUBP8pGbyGnsXXTE7tx2VTY9aVNdnWo2yadqQ8c6xyeIgsDwAk34JPn/nlHRltPZ
xdItuHuSBq2GHMj1BnRmVGyZdYjlhWXLb93rrigozjYOidBNneDRChJ4ykgOx0qt
NThGYmtqm/tEZO6hL31x19ZbB/HRREeuAkymqltuYBLQIzeT17zRL/ndnNOnMc9E
P0o44+n9ukawa/YXZ7WX4db9cT9YK3lAwPQES2RVGLfKWhcjN3cgiRyhQW6wvoXb
D5d13ibrqtSiaBNDjNmpgvRsXipX5TaJzmKfim9nEjadGNNciL5uIV3OtzovAXrG
gKOnA7n7KtQmpbGt/sjTGHRzB0t8tCvBc6N0ToumBDu2uFYTgFfh7dy0fNpdRVPx
NFYvsaw3CRIUlQZaicY9ZW8tT+Kk+VwdvqK6yT0tRvCtgJK4Bq6/9ppjf6NpB9Fc
a1uQy2Sg+eMX6u1KYqNToKdvu/Qim1R3t3HVUnCBiMLyw7NUyQNErsolhyq5SpUa
uyYJoFEzKlNpDE4fv5xMihbWwx+YJoVCFkes7dAwsaZ+B7Sk6KPX2Mz2rkMKz+I2
Jvhss2mnEspo71CJWSMtRLy9+dkVpNETad70B0nWDorBjBcEo26sNI32NqcmueBV
aCHxQMPf3SgEZGE2XAxHtU5dB/oUvpPpnl3PeR8lqqlnPqkC3akM1N8p8m0I3EDH
6grqvouTQJ67DtGlsXsE3djtrjzcuYket3vYD3u7+Hr1J4s1DbuVR4hnvp7ePrR+
L1xWPZhpqEAPkm+lAStScg8iIsAB3cQKonErE22dBOHPDAEn7UhRfn5n7pebdeXo
9avcVtk7fLhQO846rZAk9sSf+SY8pQsoldqNGmDGtGvrH80fAqwak+ROzGQU2DEn
xBVskZRCsD/VsqBiezOn8qfg5aLkFVPcojnCYmX7Y3bzW1panqtHr9V/4W9NdDvO
J/9D3jG5JPkQNx1aYUaowfG9c9c0o04VCrJz1MXdZK1iL/0IJFTAIW3uriAeyLqJ
1QiVWFsKgfdS965VDKqk2lOnxcL85FLALKHc2Rpo8en+95Gzoa4I/bvbnPsDTx2d
X+aZ7Sg0g06UzwLR2uXt7veP2K2CEnaeDF9/Zf2OtXbM6nHU4W8SJiSdD7juvDBI
z0qjNSHuNMoPyX71pCZphmxc2STcNRbuUlci3jzDxlLjYZybfE8eH0z0Vru2RzSj
pGI+Nrs1aHuxN75HImLJopA+0dYSlq1ADKaFvPgJSMBcUyY6+nzNfih8pSVxpDdR
qgPHRi0wWwqtpINQYt2Bn2QTK8l1GMJIYZW/YsPKjOhnw52DpT5x081Nu37ZJCrj
ADwPTfAkhpygjdS+nAXMKE3LKB9xY3gnjzPXq0kvDDzCb7X0Z+YO7NVfHRt07ckG
3ETKl+7Th+cq2ixOElwi0ORT5TjFsLbnFQds2I2dy/gHYKibh15oZUxKkTPwmIev
tp6q2QnJuRiv8so1AFb0VLjbJZbHxCk17gqM1/GW7L9oQETQTqaGHW40a1MFysVL
9XhzRG+Ml+RK1o50reIXA8oTitnONv4GgStKk7dMM2n+IlkQLjbtGHq2W762FuF8
IvlkHe+HE47F3CFts8FkCq3AsuZkwA3C4+QKfOrYSxCcNiW+UgDcwXJ6ccAbB++i
okfNBalqDS1ejNzpUu22o8tBRZSr1Ix5de4FMfEwPiuumHgZbo3ghw8T+cCM8CAP
7r02vvl6M1XcPZ0tOdL2Xpwiff4KtpoPaHUJMfzrvQDZx4Mo8dDXaTYFfg6REzyc
+phz/RgSZgAOeDrYE30HCnrYOqOeuJsYiOuRk4Hskl9XQjpKn1dgtlLpeiS2QvWa
9MRgMjtYAnf0VWDKIeww83UA3FUSyNa71ceOQbML1d5FLdI88IBc3MlZJ9xDKiXB
6lb0QtXsevWxGim5NjICotM8sakPj+IXj6aOwW9G50AKBdfZc0xQPh9aqFuMtN/S
wwxZ2YJlmRh8t1kIfUNUyHPv+K4BnaY5ghadLjqXDzrX3DkVVmfEtw8A1qxSRR42
MOte3cpgEqZFt+MioDyZDzBPUIKihRA1aY+YxyZAJGbAM6PPd/Ev/k6H+8tANIyT
qDFJTb9+hnchDglong8ZybCx9ArIDE4dkukGHp2cTWZHRFq0HQhumSsU4MF//MCJ
jKmP2Oeg7yYZZQcGSDuvZ0Zvz3GVCiFa3/QcOl5JP9G9yMyHfZkkLZraqV2GBLD+
QEu0iRz6WJIm0p9qxgjgMIRYA5D8mGsfAKGGTjqtaHX0eLDAH8XIr9Pv1hOqYgx0
p1pIlTjmqX3gcV+ReOhuQ8/KSStnEJQhBlByvyB/PON7a83MGxK40qSiT/5VP10j
h0CXR7NskhyAg/eJi42duaqZC6oGr+SvGg6qTklpyjJAYYtZBWHM7k+Z05co3cGS
ZwNopBcrKIdpPFQyn627ZxvmQwzRaOXrEfTYZyAcHqp8+COefMYQ2Wc6cieM/KCn
bHYAkBUfzmBV/1ej3AaQ19yBWqoJCGoouDR6OqIBIEArMA0zYRXtM3giDloBaNdZ
WVu4hW012Pj6D8iC49LfYTdF+7yWTo1TZIE6cE++hxTb72lUvr1Cj8l3iUmgDDV5
rpYtkqSx40WhCZLpsaS9Ow==
`protect end_protected
