-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
doUJZ3FMKS5pxNoNM3v+iIrL/dKQiJLBHMYW1qqtRS2m6xOsnwNF8RbCbjwoEvGG
8oq6L/iS1xuQw/KU9apZUpuRpOZwL4Pv9kOT8kIuF1hZBUo9ORlOKmhf8fMiTEOG
vL/RsSL43KSrWu8k3XS9ZYYBE82duakrUPP2akiv0hE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9260)

`protect DATA_BLOCK
3oG++llcIUycHKi+WCHybvKGjSWiQxa9CSHcWKMXSEjHSdFsorzEY1NW5I+HEPqx
7XAbqaTO4cL0h4r2Jp07pHTPSeZRqkCzYSPZFxLqilH5ZM+vJhCMp3gWn/k+a3NE
fv+uG751TzYWciGRoTxO6PdBfIW6toLb6PF9PjZk+82vZ0SADzu1sPsRv9GsA6le
e/s2TzCRAU6o0SQyffyYV6z04V0FmSeRw1bIianwdDARFyq4rCO2R/aq7KzLC5cT
Ie2PceH89tPNZMzDmndb94PowG+YMIumtPFn5FCc1wE6QLmgn5fIWN1lumZb1WPA
egvzyZX07WNnaZnZyM+/Bp3ElWonQ3J8oX1caV6qzG4x8RI+IIr0e12U66sa6bZL
RRhBaKUuCGNZ1Asv+soNmGNVPnsV9u1KEI+IZyLA2qnYu57/k3J4by6ZVesSP4f3
Rfy6se19BY+QSbsIO3Sat89K7oc0k52ZHwvuFJYnmCeMnfotKuyvQVxJGC3Dsgk5
ToDwecfF3D7OGkw5hw+ie33c8R/cNNWgpZFzqzC21KTGGApbu1jljTuCgyMc3mH8
h8uJGfN0YckybA6JaAOpS9IODUqzf6ok5fLW24/eIABmuqn2k4eNfDkXRA0vqKZn
/qmpLsw907iithACfE1d+9gVFDKg1Dv7+/xfBtuNy05JZ5UF+OJZH6l6xAEfofqt
RQiu1WKG8fhruUTsfp4o9WuyMEZA//D5Lf9ZnRt/EOG6NHKuc2l3eH+MMCE+OULE
9cbWRvXuBln43tgvJkHSkc7vB11s3HfyFv54EwyKkroX35e20Pc/ItG4NuF0Ld2t
ummstAuVr9mUWpbk1ZE44AwsS4aVHfFWejxH8s4iVx58JpNmRyz92D97/CmAAZwB
GmllAVdCPAmx/cIK6iAwDrkNZQDKhvi0Jtj3FeuZf63g4QTkLhqcP1zbeuOjz/0+
WN8SIbLn5BPkejsiP5VlSk4nzpWxOVC7R6Rrc/DGr5JqkjmGOL7VvIkIA+xEX3SW
iE51PLClYW2oz/TtsiAYbPRx66o8C0csy44AXGuYnBM3KGPpYz2T9iJjDmW5Djxy
TdK+8UNNe/I1hEjHyO8fyCZH0Tap/8bgSq2k31EtYhz3ht2dwZRxmPOl93bAkEyD
ANdFh1V+WfoammFIBdlZH05JZzAmVoVX7Q3fAHyu2hqg/c4ubsw2q1B5u5unncKq
pp7C1hwFE9Fto9z+BYdmHVsteDLDUUDKCq361adCnbBUCKdSMG+MHUpu/QeGoO8d
5KgMwoTTkaW5TJNFIIwGyF5nPfJCvxkz/UAYXL40K3DtJceYAuxqicF2ewn50fBC
duCyp220ZWf2iHB1i4PBYEgLVZM/fbz/Zle7bQ0jnczomdzd7E+5fLi1eZUDRNv+
BJSbOdWN2aDBQwS7cQSxemFKwbL7zJHoLat0BVNoNFOlG2KKP6R4WVASf6Cci82r
YqIBJpLAYQUxCkNRBWmSXaYWu7ZUW8WVOmQpzxPMdZAnGRjUdOrLO/my15L1kFKV
BE/KHWkOmAXsTcSMDrS/IbKsClkMpt6ng0LZLHEu6yvJ2VuKf+NQDcJU1bif27Rh
qt2DG0PX/TFNx6iAFnvx7HZblfSMFLg7dAIGNCReqfA2RwgQbAHoiOc88rEP+4tE
WS36CWo0UCSZ8/KqPruihhUi8e2EvfylMgiBGDK4Uwo7k/j1fm5WlwhA//AqXFTH
Wdw/eOcyOIqKzii9SmmD1yoCUGNiujajp0t3ORiR8jHCBmyKmmVEYGKgEbhGt3Rq
FrL/Mqj5qFJp7gQeBnWe3MENXrxvDWdut92w5mlzaxImoB4+iK6u5peilUK5itk+
9rp0nco11ZKjub5rzpQ7OBR8eQ7SRSftI4UzpTnuksCDpOBy4+RVnIi2IBZeHH+X
QxJCVdk9mC+eayFDXv4KGu+T2KVbfiZ63THOXdCj5Z75XCW9r64CKBygdlLPgYWC
tdOjfgP2aRtFFlWiVqu8COMARx9V4Q8kJHijfHTWvduBtFK5rLNLUvrRQPwuyFCl
bmJh0akhL84bEOSFVl9RgdvyeTcJRiW1xLxv8wBw909czOHB4zA74XM7FMLV/I/J
fMlT4rvmojBWI2hCIkjCbDkw1nMp3wzewJK+67RU2psRyD8/n/cqRUUXt41Hayml
aa0SMuyu0DjGNEtxqo+So9g690p2d67rJVzVUdiA9VTXHrXshNrYGbaxvgPRGZpA
ZWia+NmaLXt6V94v2psrFgTp4KgO2cAkyNp77SwZEiDdosAxvRLRJ2MTrnP5Lrff
go0Gu3f5yH03UM5gdTJ1q9FoGdfC7CBXDE2NOV9+NnaHpddK9Y1P+PJTF2ekK4hO
28itompHGAgtiF5Brok/MgbFlifO+KODo2StwLMwK3yoYz8MHGyAVYRpKS8tSpNx
jGGIFp5c5lr2iLUK7q44Y7vqPdrdguWbdn2ZH0JhkVyafPbpUjYmEXWra31jbOtV
okbFPVeTvkBqTkY8D/01uzY7WfSQ1OxTstmvR8GJvWJITmp7xdWvZuAU9nwQd1uH
Ye8p+GGqBODquytyR17cesKcxDK+TWb5yGvTtmBJgmX+xdg6WrLxRKykj7DMCUfx
i0H6gqN2FqE6O37Jk8jR5+RSKPiIKs2iZG51I1pkZ7fy4gl6Ht0GYa5dEXSCCe/s
/F6nExy+TD0nrxHRNzfJgl5AqGKDKwrexQ7TlNS1Lly5EOrsHRtzCkFrxvFAV30h
V/jU4q1QKWaTIAV7dGT8jjXTgv1PHtSaW+Or2/MY7Z8guuNAusUb9lSFYwS6bJ86
UIZX1gDLeqogWUuMmcPtztpWbJC47Tv+PtKTI/V0+h/8W/djYjhExFmS4Aj+BDkE
FEjOX8xyjql1Vh6AnoWashqFCR9sYZvpy/tDP6TIat0rqziRtJct01mzMXoxTt6/
KHu0i1fQpUoMrvxM0ve2JRUkC5XXuzAycMbaKrXbz5we14fJGBeR7aI8MasFzqKe
A9gFjwlG6WGJjmAYYRhiCD1/fxOO3X/iRW6T+FKcI/kpjhuyVyTDfMtcO980lM7n
SpQUrXKJYPtSLZEpd7V7YRMYimoz84M1rUAvqRfTXcVVfJ5+sE/P1/DY4T1xbOp8
FKG/Bc57TqDOBXe2OBP5DoUN9LJkFmRPJgZk3BorxeO0csB07zKvIu366EgqxGZx
IEXK+E5T1cdUL3hUXyTW9yMcoO7roSBVrSLFeAvfyzikrBdPcw2t6+hpeJdX0ytV
1NzxCX5i4OkQHHBMOC3ZqEV3tM+6NMCGtpwUwMjT3q2GdmOVLdiRkq6D2MPRuWno
tC9EqP/KGYX4AyRoCqpHLy/Inrp7tC1kBhdXLz5Wh6LKnAJ6fjnpT0gw2WFqRg4Q
Uq5PmG9fsaxQa1nTiAR4gYXJr5MVZzgh1OQeAjbORvBWwzHDuB8THwUBKKXdcgKS
zGRJMvSfGs8y4a2/Rod0k9RumGkfq+SXBKrFB7KKV8M00C1Fb56WN/YTMqfK4A9w
P3WYSWey6+MrsSR6Ggd9obUJ4xhZjUamWT4RCI68T57L+nz6eaQGk7hqk9dv6Z7T
pfEeIFO8t6NO7wVZPvVQW1whOQiJofX/Qh3vYB+j+MAvToGpgLbmaIjLm/gq/deW
78Y1UWVolnDQN+5oUnvja/m3wWpzvqRMvtcHRtsOHmeMq/kDo/c7bBxDTkfvx9gn
B9KDvNq77Hoz17uRG8EMWT7heJSSYoZY8CvX8zDpi02fYR9WZQk56Ls7cW5u5zRF
nNDu8Fbz4qyiGtpbMrEtdAf8BmOjh6ZVE+hJChvg6sBcHQRWMMT+V/8JgjzOuNTl
4FJ2AXJUn8UnAzRIoIgF+w/eULVE136xU4NHaW7fALIN4lMH1S4mdYE+CmoBkHpM
kDKLjFnbUPR8Ei1wowlstIdATlZJYyNN+RZgPQIp1naSe9ScWoki6OcZL6268peU
aBT1xZyggAmusQiemUoHpcxTcjjKx+ykNcPVYSF9HcDxqmpFJ52XXhl6r4JYteUi
7V6Ln/j6ZOex8zK+l6WknxWZspwMuzGRpqGvXZtHi1PVmnMgmukR/qYBTOpqgGpP
8NdOzDd2zFvK02O1s3vCPO/re2p2tK1y4IXG4jtZO6lWWk1+R3YZpGaPxFBpBdLp
QJosHBXA0GCrfn9tMoUbfdxk8VfVlwgiik2eJexZ3SVHOb5eliTx4nTVhV4dsrVk
F+92nvNIEumtZiYfXpb9XdR6fmj0npGS0AIPF7E5/mmM2iaoOYTNKp/rg2/5TLAE
kq9TmPZUHGpPjCmqNcfzL88MzvMOvAJOgw1S5nirHB+l9NGIoeOMjuODwJhIIZD7
s4yFdvOw9D50hQvZfCSzjTUp/g8tz0KVSFaHLsAaX/fGhEauIUFKzLgUHeOb6pv6
/UGVaVTf5yoHihevFDJwT741CpKgeiXrbLeaBxK9xHyxpUnhfXz7+00Y7gkz3FAO
LewBCom248i4QjgVvXD/TbEU7g02mW3FWQwgcdWpMnjP8S+AQegiZCS0ymhjQUiE
nAQVipzhytmUmG/1UV2SMA6zy5s6YiPZVtx+/zM6IrToYkgESB7J7+IbszPE1AKO
fVSsY3J6lOXlbUlNMgA8na469ufxALJzDxd22OqdJueHLXy5Dmuvl3iOUHNxeh8b
i9sxKx5qK3nyu2ZPHPvpNqMCwRmIfpzjxeKGqGanp48TSMXCDAe2D6ZUPtrPdJTo
CPRqHVj91+DmduCCv2URxB008hGkJxkLLOiPhXvoFa/sKC9Reaj/aVYkGwOTKCSr
ekXVDJQfs+tivA2ZfBR2W8L0pII2+BFN7PhIw5wYxF9Q69wDnU3qJZoCNWuyB1qw
GY/DFdBa4p2boIhcdB0TUVn23ZywFBtUlZxP+X5OqF74EqEuta/wkKq9mQz0Pwh2
9PDmFxJGyXqk8b6BreQh4AtE78yaJJymXG3IRqdhZGO+TOLNUUJhu6fXv1k11a/J
sKMDOA1KXxjdXL+HzVkME8cf0HbwUcycMUBfX5X06uz4oZp2jNwHU4p7ofIm1Epu
QEvN4Hn4opgL3ZDDkR8siDkvgGwlRBw7rVxKYTj3RIYoxtMSI/1FPZCyrBiAz3Pm
DCZIyebbh/veaTreUunuDBMD4qRfpi2nY1zygPkEaMBy4tb15jwNBwiqVoGUfFaU
NJIAn0wtOkjohiADZH7wUroIfF6HoK0BCMzF1pmsiDNsQnu3nahygn9TgDn8pFgw
81SjLuvclx31Xy/gG9U8kJ8u7jg0cAij9uWNLOVZllrLjYxM783JB/j1IuwjBi9w
tninjJ2RLUWDwoC3kXZACQu+TSlEBRu5gfUymthc/Nn+3xCGAKoxGMBf+v5mG+PV
tSnb9bXf3OyxIebQxGKdxlcDDnvchIVUezc6cSWYT6pAvV3V+5Ai3hDkUjMsIZI4
197ExRNBgXgp4DCTHmyxGQpbdub0N+WWjCXBN0FrglSqUvAxfoTWYJJqXoXV3nTW
eucQN85mwldO5zJ4d5Q83JQdKqWCQOZiCzB2+5NbQmamv7olwXXx6fBcz6sRxHtY
AF6sjR9wqpDhQQI/02FEy8gqAFSpDusdCOeZ71AyZo4zOdDS3ARq3u1DPh65n2Ai
Lisu8zAVL44sAg7twM30aOc6pLs/iwxbPGUBtQwlDAASRMyqvXJb5p4CJ4MqQELf
mG2/nwHLtYoGRBLpeGrVBVenxuSWu8p4wOLyxRNAeh/mAWG85qBtqS/sTN0dsb7R
ury57wnSzlw9Csp5VJgLwII8sKbgr9+J8+RzoXYLzoTi6tgBnjqpg+K/1qvQ61/b
4MGXlqq6aDOoJ25eaKjbAqBE5aoH1A6uzlLe6m6VvwY8zEJQ2K8p/+jIzq/XqrlO
Y0jFcYPHVDetHRDlmLVBJGdZ9ucv6sn6xoxkfiGqw93JKDAcngvRs2LjrA5oPi7+
TPoWTGfpKcNpVFuU5nthNxdo6l2PKwlaHSN/FxERo5PGg2JuDVcEEkQdg8QdbQB3
S3jIXHRP2muG1kopmf+uKYUdnvTniC6RgU/Nd7xwcANCbgZRedDWshE+SbF6bELZ
3GuZnghJwLVl0z4h/vU39/PpUKXKqld0qqAE3QQ2vzIDmnfPNDN7Oqu6OLOdGQ1l
Nt1ppX6gOdXvn1AALSAFmh/BkQmH0lR0zGOJ/wsh4XsKZzV/WoNvGbUOG9EA47Q7
yG+vSl4ngPNbY29Titxwc9F53dG5Y/neDR0ir9fi4MkGwSR8pLFhLXUeXxkhz0q0
D3EC+vsYtwvPb7Q3/AvZyGm6h8rdlGXekNRbMQYV/HAOUbTplOLUCXq/9HGi0JtR
ah8ySNPlNVYvYr8Y+YubPRyiRHBxwvxO9TXbwDtit75RBoTeuvchGgoTIXYy1Fl9
BByUs7gfUVwJDT8PCs1HgZzrTnc3sEbk8I0Oy9iUV1mt5QlNXj8qOTrVnOovAoOr
BOwdc873EmPR0vPS0T3pVK1huq+4PHO15URRbOfx8LC/PJDFWo4b29aiMih90kID
TM31uMe8xdeoDoDZp+lt2M1tbJzJa0T6SquyP47us88gMdc/uWpupz4O+r8ydjgQ
JDAq9McNgcGGZvH9zLyZUbPVSkAOUZUZOjKJ+tLDZZJ6tftled/VJ0l1WWYEq0GZ
8pbHiFiBcqYlMLdbiDdDIwDmWAjF4ifs1DkxkoTpRiWcq/ixcrrNjOUyPzdAmfzi
xy4bf/PASwDJHcb9YSmc4UlMnnxJZuIdiLLK9zvQDtaTFdbI//jYqu6jW+D5b5cj
jSLcBTCwp7vyHX8IaWCs29e38tjgGUSPMDnxYJtkprG69w22xkFtyRWbOe+sCZUi
iKqpSTgbhPtIiqH50MzGbAfpIRrARY6qZL06waN6q3IxFf3XTz8agbyJOLg5tqBK
ZAk0aXxSk43Pn2SD2K9gsxh+1DWNfR1Wy0SWjJXLaGBBnpKZP1PordiXAqyNgWVI
cH+ogAszg0TrGP2m5CxB6oBPD365ijtsVuCpZmO7mbdb2CHJFQiac8n1dUahVz/e
2/ZOB3sLWHjuGDtHe/ze2h1oQl2KGCDcVflySP4j69s49REOL5S6+suuawfFNKlp
raskEZnfq4Rxd/OpnE3TJJjQ7nImtQaIpJtBpvcoWOG+FkqKw8KHNXzgK//OC11C
7qmvQAtEpNKMfGy4rkqASAlnH72g4WpUrSzC0HV81RNfGI0U8X8ez9wz3nJ1z28k
+zMfwo/oIfWbBe4QosFwYX5q3K4ReQEGArprLsBxLE1x45BABRE/gsp0ChITYdin
NJ58HckDTWcXBjJc9gcjHg4vJUJbgHVGPIkOzyIxe65IxFIBSZtQZ9WdV5J1jjP+
bAhNG/IHSpqVXYWZzkOCWPiZet81xVvs3ItRaJG937Ym0f61uv+Y+skk9Nu+HGNK
tfgcSHffU0E8WTEgKle2STBuUpPItwyO5FDZewqs8mKJbQhVr0hbUAa80+MWzAXB
eQl7Cxv8ltIWgA1Bs4/6YW1reu0Js8yQ35uGrVWqvOn1kMDmhf6MRMtFtJyTIWiU
I5wE01tpe66sb0meS52Bt4RXyVcVCPJ0TMg8rlC5cYzYqY1m+67jisDXyx3UKAnW
sSRkKP/NwGRa3DDl+2U3EY6DljzhqrcDhwXDSHwICEOioFwijCE2N+Nsd5w9ouDD
JjPeFhqmq70AoycwL7Iap70MhKRPNnMxxNBXuSEXfFowLAaHopfS5d53kYisE75S
Mo3LKFs0GzzKOGducfYEkcpFjOWQ8dYluNXfY4XD/fRZbUKjU2A9jvexNCSfxsSA
OGMYcQZeppFzu57TXXJ9dlkaVHF6/e0xIeYTWO8TsKJKEbg+dsuiuR2epbE0Pdfh
jsmzpGGIrvwbhw0Xs3qr+8XDfpxqDw3ti3aqpAOG0ZosL0O3E57ECXSqDpboLzwz
+AfG0YU7Bc9Fjn34Z1aiamOYCAYM9YQ/vXQmQy6qxxXhrA0O8Dh3En4+7eCV+iAa
XbAWYiI/R9TWI2zrLJhk4ZlXPJ0dOVwJT3s+h5CBMFFp9ECmhXcd1rIpYqIImvrw
Jp5NAAS6fFMDX6VhzguZsQ8Y8zMMlnP3/4ccqAh/173ekwqSxega+NQieqYIIg40
Vmrf2yXDWrwznXgxJIM071eirtv9NRTHyr//ksIs4GX6G/GDl0Pnkn9g6sAyvOEX
7t3ipfmvme8b2xq3HQ2R4BY1uD1UUA8DqtTiT3btoYZotlgDMSbWPumyOU73ycEr
zSd0rnRSwzpHA9P0shRNN+1HmdMk0BLQpEMcEQzOvMybda50H9f28bdC/rHhk/io
XIyhTjYqHInMfKKh08j8csCo+SdqYmOI2j1u4mp54e/OnOLteWdK3tiJUbh7iZm0
JYhjUqIhScssGwLez3rARROaf+qrprmwy13xPw+BHvKyiNsQxH0OPANLM9fEBR9+
YVzCtAtrGYQbjj6Qwz1J4aNq01dkWIFOyiigsZk9oZuTc0fsoZbX1vt1EkPmGeI1
WAC7AIrCUjvpW4Ct2ViqJ1Hfnaq7y6F65uxWn495++lnKE0ljmlrtNLNUyuTioTo
6IpSyC5VBzcdkip2pB6Sv0zzHjK5Hk0cFAK8gyQzBcpqB/oSjo88ckHID+TDKY69
ajWopI/iArmxAa/FC04paWtJkTN+b6ph2xlwZub7VZS6jo5SZRsF+bsF4vWk+Z7s
OUdZW3zJL47M2g1DSLJjpFGfZ+MoyoQj391+F5va8TBLz0yJOcC/aLZEDURqjgQ5
BV4GPxmIpSmJMvnOeKiGc2Felx9iRr9DRO7TpYS23QSxA8b2c87W+DzBTjiIfZqs
+RKcWG6smSljp0/7gAF/4fFMOrb6NdHOfKeHtO6IsrmkfYH7chjXP69HWXOjpMLY
yta0XHTgXk2RvGcrUZxHjXve1LaqpaZyuC8NC4OAHNbAXFlro8FEsXrzxEnvqGfT
x7YlBoewJwjHcoDA16OKFERbjgcB2jAdpImwa8p8xO1mXN04dSI7xpFBTAGnvF9B
aHCt1rxY1L+sYCs77oj1qHDMwHcZK4GFEfiz+ktz3vY+A2bdZrEc5/npG9OWw4oL
Dg24dRA9B6dM9Y3zmF2EA7ylVNkprQVneLT19+DUkbJOXh7yaraQ2VGnj2Sf4oVi
TCSv4oUlZW8KwNpjT/OTJZX0Y6+jm2U/GCcfyjo5d3d2DfK8ApHPZZkG8xGTgGPY
bpp09yVbYTXpmUhXwXe5f75TjSUbDyr8siGzOx4J0hXziaIlZmhcrzSWM8P5UtgN
U0zl+1GAGP9KCTRHmZW0Or/RuRqe/gVBGfLL2TBexWX8Vm7cQ21Mlw2wMhvJqSKJ
I+UByVGEuYxM0jVEaEWrchcj9ypV04668F749YNoeR41aJnGp7vWfJsmsRYG1+gL
rtvy7DxjFUvZ/41WZYYTw9alciQqHvzkr4q/HgY2nYQWP5ZwR0XlMQ7SDFAJLfwg
KnTiWx2ypTxofyWV8ZiAoYhW4XEsWHI381PHjbif/3jlKv0K4GBhFz2tlSs00OIU
DJKWwt5xachYo2nPnXnkR+3/U91+O7Qr33HmPJ9myuMkxTnmaYfIcIbWJJDBIjFe
m3cCKG5yJ4GAD+qq40YZWJ4venCZZhEyZ9Cy+jX2sWk9Ekt7EgDj/DsLaRYP1//H
GXqpxU10BeIEaBbr2Iq81o6gVgWXA/PGIVCI1okPNygaDj1ZvO8uxCVWwPVViYOi
L795NBfQqD+fhtZQIhK2Hc5L493Puet+RroQCjmYHfB6eLhuL+MhS5ekNSHeapOQ
emZzQBYrtFE3WxOtI9EmqdBxjvRwSKZEpXs5qunBgo/OINK6p5pL0jWKLG2QdMVN
XKVYtRVqu2Cki5Z7Dmaa7HANMIO3rlCxChG+YtR7I0X3K8QDFmzUQ30Z4rv5goW4
80uRsQ5vnMVaOJIHlafiOSr4B/X21yCFQuZC8zpzcostDMNq3vnlss9dvI8RLfZ7
xh1JN59YZvmvH/43l79H69cvLJ8NUuH8aLXYIE7sW2sgLvW6T10MwwxtCHo451mj
aHMjDYJ/pgsOsZLwUdg/qrlKdU/eWD1WItLzp5vkmgWzQLfG36F0UQqovE/+nvdo
jRG7M/9Y2d2Py/08AzyJ6CEYfpNjxOC8hozzof4/Zz89f2LRx+doNAwV68wK9Pyy
yY6oEc4UcQMYiHT1yYBTikOl0RXu3+vMoCT9k55gDG7WbccozbiO7pPbxnfuE++y
atqASB3ucszDjF/J7TwZN2LqttexcfvEcv4Q1EztsrUW9UtvpRKSDDTOIGZ/+iof
lOuwa33T2MAE6S7tiLwBHO4ydOxr4AJ0QdvDhZCe0ozRNCS0qIIlrNNYotG7iuoz
3CZOi7lTE92hfHm2VKewJU7d+DCTRUJ4/LyiAESsBAiX7wHyb+U+Q7j757T52hgL
E4K1drHY7LFPWZUI+xCjpPd2ivLeNsIuOsUwSUcZa7sKX0qnc+XCI3Nu9F+pPaHJ
Sq5tPi00D2vxGfxeo9NV6M9O0n17HBjY1xTyC0nbKbhn28Lm+mAHQ9r92PL8IeVq
wqIU1hlTOgUZl/Tn7SEVu9oym85KWcoX3wYubpN442FiuxFDh3jd4dddkfqhej+P
EOCPA4ei20vMYdJKRo8Sl/LYt0pdi6xIiufcttpNqG96zV9ilV5DIOqD3cLEUfrx
LJ9OZBktI7qp+nRu45ZgZk/D1ACPRJvq/6/mu9KCZ018b48R5v+laUiL8ha2Tfua
rYgZG4fsw+keTvlptfVsk3WArafk6zlaA7Eb08wu1zUDwMihGAC3JExq2U4MdkRK
KbPxtKM+lCYkvcZhBY4vudmB1GQwDjFIMj+psgFme0C5km8gQIco30Lv49s6yFPV
InkWchFUH/c3V0q0MWJD4eIacu8oTyf3sR52Fq9iGML/vtMoBwmuZ50Cgfkd9C7d
tvIDTrzIIjJdSapk1lcwWdNlw/NDfozFhWnNLa8Xl/g96Yv3rvk60Rb2RWNByg/t
gvkkomoKHWxKRLTmymksV2dOpGjWmOE02e22EtQXqFRwtLAVkUCQQqvVjLAkuJEK
xtodmCKa67CMdBbWm4MoIOdl4M7FVQvvF+lWIa6g5d1TOSGPoRH1yHu/vc9ObDnl
KW9oSfveKnQijPMYP6igHJlUqgU54lXNFC9fyqj9XTLn96fePhhqXvJc0san7eFY
P/F9+WBG7uq8YQ6k8zhk8x7q+P0e0IDZewt/Bx0DUtM7pD119bUVPw/k/rD36FGr
ExoGsuRRBmM2Mz+wC/I0N0MJ1be3lHrLxBW8BHJn8ug9+dLgq7frTuxz7NPczB9c
e1C1iXI2YAz9ihlyTxu2iI0mIVkZ7mW0k3aweMP9AbZ2nYo60JH++VZNMiFhRGXz
7nRw7oZDOeVsJaMEX3+G6OASmDlS03IwkzLt8EMN0oCCAGwoYD4obVmPxA3QHYY0
UbSQXF7TUxJnmA7CLfYksX25lacAWqF6YcFOFI/qhFcN1DxZnQeq69kdNIWCq8TA
wI1pmYDujgaJlHOk0xHxP4a715fQaCWF1HuKSqNbfDqMnpX+UzeRnwHM6cKNwvsF
ORYJiX8v/20UJTZ5QgKsnMdRKQmGVRODzK5z/pXydw+NyCd53VJpKx6A9v+Nl4RK
fZ9j/+53/eOkTiKNk5GogUTfX/QOPbBOdY9yY7N6SQ2AJluKlkfxcckA5KgfuQoR
yBonIvzQHuzoW57AzCB6oFspxYnGaoqzXNHk+bbhWBy0G8gNPCm52IEgzGU+RyKi
Rlir4cHCjBjvnW43WWdPMDCwMO8JEC+hv4Q7LdSzSSNj7RlwnT4pHOBf0CJt1/1q
8IOfN96QpF7DlnKIaZ/IrBpqz8sc0NAhTd2tdKzovlngiPMTDSfjjS1JJMpy8oxU
FP6vwlRd/FiFYr8Z3UP8bvxcgtt39WbK3M6lGNvDEVEjlVBrfUjmdWdMa/5CkSCv
2SrJdl7gPQJeFkOUf0yAao0LODo2P6TC+cf+eDxcgEMFI2XalangDbx0pSrbunSt
dxs/HANQIR5EqtMqp1eWSJ2SRqjy0Ew1Zupu5pfOTQxQQMFwn0NaC95aGV4jc5dr
Oq3iC5bvEbfsuNLoHmtqvm5xY0o4GvhWfSC7ZgTV4e3iW+fhvxZO3KmNrWrdMY0x
kEiRbVxi7R/403u+uMUjeJoWGvHv+5MQ0NYTBYG8WkCunPV20/AtVlLlEjyVJ3PV
SowxApQhXhoIIvt3i16Bju1r/12KNki1NP2Yx5KbYYoaO9ZEtrD+MbO7A/Q/RQal
/4MsrqgrPCRgzU9EDE/OcYyY8mHMeydJ1pXaNlr1KFBxCFc81WJ39IluYH1Ao1Zd
oownm5MoyHtp7/SGdcXRhA==
`protect END_PROTECTED