-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1rj1GJF5XDCNxwAuiXDPjIvyMeChX5mTdkjtfr6KBSlumw6K9/eaK4tVKS7H5Gbx
NduV/wmj9q7QokG8/23Be452x0pOQ6zhN+PFP5t/TWw9P2Z4YPQbLLEeWX7Z7vpt
PUlRaFAYj+8aLG35Ss6RPZM+L8uQcTgee3o2DXIsslU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9488)
`protect data_block
mFKeWYqT9iMxrOZEyXhOPc/vQ0EB8aR8cOU27fNXGFSU7fe1EFNgMcw8pjJsjRMs
kRkIt5x3h+vSIiQL3f00RInYtizLjzYSu/lY4lAHNWb8sAdj300GURPT/mSc6g9m
FWQf670EnX8Vo3eFqhX+Z5al4DEhVFJA0kl2/QjYm9jlsshFX5zZVxJx7Sbngf1+
dcTVewEG1sgjNT6AOvrLDhwUudHNadg26t/HEVSPiVzLDFqX9d8s7VEpq3m/2JY9
Rm3Vnz87AzW1tH3OVKzdgFJZErwD1O6tD7GKvxcSDUhI6Zdc3q/2T+5AXgPM4Nvc
yz4zFxCB6LAHcgwNWqWlu4mZLzOVUN88KNzuvK1H8v/ezLuiWlW/4klaQrYW5u20
L9spdgvMgItJaf8o+VPSqAPV8ELAq6tZinacbgLhmX9Se9stFdwxhtuu2XrCq8pq
7GHci2Er7fKQUQsfOLOD+MGAzbeQ48FBBEvN62Yvs15adsPF0pqA2P9hgoAmmi22
Coo2WMmiRPYXKM90xbf//HMeah2aZJe86w35YoHxYZPG3J5Jkfocf4z/cjvRAmz0
mQAxx7qYogpByIyS8E3MUyW9GF9Tc/DktQnpn+BCorT503RABMJJNAUd/LjBl+i/
AoHjfuaOAkrH06zVjuZL9vRicxnPWM0bkYiMWC6Yk2PkWq0I6u/B10+05GMU8hru
XJQHwosO6xoTft1agBgeS0ofiAQT74Trl7Qn/4ZpU37T9yvgKjpUDF3Xp5ldeEs1
3CjnJ7wVYuaVzsdq6I8+fOG7X1svS48rq0/q802FtgliZA5X2mg2Jky5BaF/DJ4l
Co4lbJmO2xgrO/fXIcWmCn39t51o4YDSiALj2PVUZMZHtUddZ3sgJ9H3cMGLu3SS
j/NXaI1bYd2OoiRU04b5x5T+6fpzSMj4CDeWiPp7BQfEyNYijMAECyiFLK3WA2Gh
9KGzOHs9/YyAoBPEb+2ksxboXcYTE2xFsxqcXqtEcV+tekmQvuuuEUvZvUnQFHoA
XV+KwwrGZgsKFAUzuX2uZekZB50RZKhPbxkiglj8IHetDwbOG64Su5cKCPfOPlvM
RdnGxV+faIQN7jB0T3dVLQI/yMUjlRso+5V1v9DZqSe4jNFDbYH2hreT9SRpDFmr
+4YfJkBuAlpfX92uhdjYcPKR/MlYQr8XRQImwu4N6Rie0m4EvjaALeAIPQEXcz6e
PTELwGdkGtWgSfdFLZUNIuHXb9cnVU3LZn9c7sMY6wFQZnrO9U4AifWJ9VqBMDcr
nZV0Dvz9nKEwQVC6nLPd+Jk0OV6sKON8jI1x8RxWYkJFuygCRIlx+1inFs9WTLSw
62FezxJ3vUIq564ID/G2gcF4m2W/KqVEYgImmMxr/W83PWDDYs/y/1CSoehUm/7x
U03bkv40//cTwzX7uAa8XpYvRzpvu/JTgKAw2Y2JWOYglHt0WCMQglB2VveedrHE
VxMyLi0iTAM5jbpWjzvLFY1m4Kcovry+RE6nXwx4XJgMXeW49tl9072P2u0Tcke3
5hpPgIngcsazuH6qQgyrllosm2Hr7/7YvWkwF+YLR6T+UjsvrU3tX9whENCcDRUE
Ug4LDU8QNmKU6BKbxkk3Ga+YzG72aVLDu67buOmyKevFfXSG8WWiVGJEQXnF9dVf
4i9+6v8+K0LtqSNZaZAesXsMx0/crl7fxkK9Wc04xgJBJ7gVV5eP7J3EeABb/zHV
y7snwZ0NPk6yLBhg1/dPrPUwdExTV3nBZ9jo9LBDuv7YyTKFHEEbyYFT4JPSYjk7
9I1MS6TfXfEv082dHtKjBTLmdQAHYv1Rb1FGFGtGuXg8sK0NuwopWcKGTiuiev//
W8xonIvcuCZLmPA6kcvKwg8Hyt4Hyi8r7ZX3zxV6j7P7XQ24aUsF4Qd3i1sYjZHs
sGFNIEsgLYsPpQCtU9PWHtd1WT3edEVFz+erX2X+UR2f7HBVE0fSle+q4cHqfIM0
huKn4Gtnk0yrSpM9VYf53dDfRW0cr1371ymXymWT5g0Y6YpLOOrpd8IU7RsEerm3
c5ISi5VBttLUf5chlXt6Dj0FIyCTKqFLK+iUmyPTIPYRwuzZHnGrp4s1hpEbwuEV
p9I84lisegXzQmaaoo0JFXDPXyIeFWhJGU5IXVu+ja6NoxEyBAJ+32IvwtBrsI6T
ZA51wey/bnYiPAZtoiFTkTqRK1CAQ8d5o8K4iEWJ8f3V+rd9v1DrPAxntdOVnU7A
9ZLQvgHVSEucdwGoozXWyfKqgw4HxWHWso9DQY3q19IrDpsORDzeZUQ2CbZ2js+H
UftNDJBsXXvsXGWzVfm6vcGqzf/UHtw1oLycjyFe6ttqbHZIKKq+E1P2hG/TOqdh
lDEPs5DVHV53el/LWSXJwI/nUt4rvpSyUh61/pK2ORyOyrV5HOON9nxkmUK3TUZ0
xVu0etlIjMYoXae/YUV8CzC2VvQxQiecOPCaZsvctlPcy3sgZJDccJGymc/hycwN
o5xiKjCBWQQy7lnrqeEJotYiQf2GmHaAPfcrSZ0miwG1VKn0DSLtM2261PV8nNQF
E02z1JmeCrLCTBRizhr79KB6cc1nhzPRBuqJzdAPWbJseRKRBTEnVC9UHbdx50OP
oWAdSO77ebIU991VK26ZpUw8Xqj8CcToL4b+IMM9n0F+ha93kDFwDYtLHayvRPSO
lvvdk2MO49l4xQJCdWd73WQ7ie+K6bcN9mJ5D3Uh+Itu091rybrXA2SdyZoR/Ag9
QN1eDkMsACf/0bhmD20sFjwR5uoDDkBrSdqNLPHo/nAVVdtC13Y29Vr4DoxWBIRx
FhYsrIj+xhDCKWlXcmke5giZvF3z8tTVdtcPRMMV553ez1K0EIJmK1tgaupJLD1E
IN8m+nVQDuRmRqViM5qjj3petMjoWk5rMyoJtbQyUS7JGack3AmJHv6QPVOJDKno
rZgGgL/4YcHTdF4AriLwAiXffE0S1iRAzoAsyu4jUbj4uyC5o8PqJWAXumtGJSUb
K/HeS1o2+7Lr0hrxlsP5WiY82vkNSyoSaTlo2GbBfRDEGYMqNfF/uMK6R38jjOhh
XVgKhSgw5D/uZOZwlWLwShd7g/TMv4QyY51/TgC8llRkOhJtmSeFB9NoD9tFr7FJ
xUjH72XjNGFGGC+jdsn3k4uyR7FZbAXcK8ftF+zqGREUQvRVppMfoEodsLhA87xD
32ZbIr8MSOHPB7gNa+bkDVVDvNDJ77xrR/yRYvudHV8ZuYxaenRzfysuH+8LNuyK
GDEwR4GoJ0xdvWutQl2Q2cg/aH0NxYDnuL48c4NoDBM+n7tdp0S66WdKIDBJQKoZ
fRcsNoP5xSVaOsbolLHpZB8jKL2lRYeBwwkttJ/+iOzgJXIk6wURYwgFXuYH7JGA
jmimx4OI9JBM8o5Hm8q9FnpkCtaV1x46/sAXeh8chxuTJ1lv1H2/J8KCVQY9hp7R
3SBA9a9aeWeYS09Pm8gEAFBNzsjNxg0xPYVL/h6XHvQE3y9+kCpMQ8y4w15TYiMn
Uvod0TiIM6bG1RWh/QFOs8n9MRrxksKXWvgDXcAav+G8+Rctnm5ylVSSxD5Vg2Ed
4fh0eGNi0gCIkdd1+tH39DDYrLWMHWVlyIgmgP1ua2KDHFLHSDTLGL0O7sjI3Eb5
ozRQxZpYv99Do05LGVAj/2//JH4yOHse2oyTkmDswnPG/WNnsQFCv8xFMcTc8y2s
eNJ0wOsaRHPbHvL1/oqfQgXNxwYrGo++oxR9PA2cgBbG3P3F2Ow7aWnGn2FtUP2d
/t10sUfG8NCO322FXpalWE57MyKE1Y+tJIkfEH02/Fm/kRkmMHtyLueFnAaCvZ5E
fIIZE6EcasGbfjv2mgNGGKynfElMhjilXhrEFtOYpeFxWkhwCbyTM1f4ce61TdIN
LgUWYRsJYROdDNnhqQd1io8o13n+BsgOaRW6/rUp1SQW6Dj7/vKcHMGfCpc/zH2Z
eEwHtJwzVDsHJIT2XH0y0ZW6cVa5N47Fy9LPUT3edpI19JOnAIhGvKrsl+Uei1yQ
KJFrSV5HEsjmJS60yqOQxFQjovy4PLevoZmRkLCSqAVbPVFAXpbXYDESdCUbfUYr
Yyone/xXbPbOYfoSi2AldJM3riRSy7toWmFKf6jOWZrg1EKFRyFHCz5vaiDW3JSm
Ju39xrqHhFMh6ZwtU5nSOuXgsWXjBOZPxrUCUJKLp7y6JEYUZXr75XVFQSUjJa4o
IZlVSXCioWpHov8Nm+R1Z/zBtt/rfOPfakvr3RiV/fhGpzMX8vU8lUqI7ucFfAwc
t4pUfQxB8CG26FW0EnApHkfWfytGD8iui68wbQ7NTjySH+PwCaN52HguC42/oIBP
FPLhu0P7d1WBoAw9XK3Ihnk+kPRDTsZUscrcp232I2KOdVxPaS11PMfq/+XiAXsG
5bWx1pN0KzOOh4/V+YOkQl8S8xyv/jU2qShkmmCBPbWrXqupMAu6tmaSOijK7dnZ
luVE2RqD9e3rcfhf0w0QyZye/0JS1l71G+0GkgS8K53r2a1Cy6AxAbMJ+VuXbnQT
G801s4YBi4ZI+Y0ABXp6ahm8Apju58yKs7xmNs7NZOJmi65l6S0ywa81wThMCaGP
jHDWAiP6jmryn4L3sbEE5G8xBY1t0pTJMPQshBkpTpNDsCwcruyt1jZrGtIvcgXx
/QCtgkZkphrngFzZUV4SKI7TFIOg5BghPY6WMxAFO0JAchtohdiAJJPBVdnJ9R2e
N0Twdgo9QmRKpHafNvCg/rUzNmqOvVTjsHnCyYBJFDrDJSJFqOAhTsR5El7FpAcr
k2JWkxNij1JPwvUcPjUd4S0h+rda19WmhcpNFaLhytiYoWJCuDS3yYergLHxYWpx
itBNsAHQzg8vseSeNRjEcVKRmigh1AaNHzhl0rLyq2+UQR27cbLfcjX2gfWBEV8j
N/HLtV8RSIFjN5HUouFUeCBovJvg+rIGkmcWK3HS4gRXqAOgyNQ1PdJHLDjacxzO
VUYQbtVaLUlp31AJEyYY1ZOPwk1kZbMF6jWGv/qe88ZcUhBjuyL3NKsZthara6MY
aWeDhUIMT0HbR90IKCt8P36f46b0qwSZPU6A5dp+z4rw3MvPn0SQTIgsd7bjBUBG
62kAfhc2J7VDgIftG892RZyg+HagHzYGryQ8PjuMVz98b0V8CvKvpjd9HsSFyrqE
n4cG8Hex6XohkeRTQ99QPmBNnFQ8e3eUJsu0uANBBRfBxpWaQczln1crlwzrmKgF
3UQ2ot2vOB3z1RWVruPAa0+uX3zc00rBfTDFwwUoVMs8nH//lQXIimsd9cgK8yme
cnV7IkAy8KiD4Fxk9MIG7+FHyL4Xv7wlM847g0OCvVPCFxXbEYJnQHuEJryvw0OP
gQkm/XkimyDe2qbwaKLFjn83vX2HWKzmKlwDz0gloSS9FJBB/M8VTnxe949almaW
rg8BD7YUahsBPye0G4GVjXdPazZ86t+HUQLiXbplwcQTswDMQJLhO7zomS5EglYF
u6/nNhakVsT4tcoqoy0ZADpFdhMkfAtXv9f4VSscseKfuv+0CVdC1QKWhVobSidc
1IbefG6KxiwLlJRszPUl25PhnGdkYSp8N2cBENb09F2/AVlPfxvy2dD/5PUC7fzv
P7ELYL7KBVRlmKdnACSooegT/iVkhunRiej3qeS6YlzSdDdOxeY+8VrXkfHjdTXv
rQZ6VOm+QXl2tZiS16XPdIjp2FRr6hlsyZsZL3Sr3CdtLmSB8J5h9g3QjkHDmfmU
iEa73Cs4h0W/UxyGGVK0q9H1x0L3+zlK2BO0d0aoCsBuAc9kprpSDHp+B4PtFXd0
PEo19QpfnIxRhcee2S6ZZCLLTKy+x0A+ZYMNS+z6BWFdKRKvQ9hYvgcr7KWrkDBi
7SfpR4nf1z1rVOZS1VGeFlG/98n7FOfprJbB3CohFnVov/HcidRb6EZzC9chw7H3
Wz+/Cx0E8f+DU5OkTAYz9weWAbGfSOvt0hTvlO2XJfT+xixfT7eGHeMyPrhv5dPn
CAuQd5qSkwTif86xMtIY7gtroNSgF5sME0H6klLrjAxskqgO8P25iXF1f3bsvvAs
9H/uSAFAA18W1O43Rj78sefAxyWK/VD70L1xv+d+Il807oCIP3eveWs4vMiwdxoD
HhxNy4STI020GdxB/up8EhAS4qRqnkZApHkfMfQEqRYPHLDvRkT7P9TCeqiEG6No
uxx59x0HzxBKpr5/A6FXw1ZZUg8M+Y7/u0pg7NbJJX300IjS134ll1vrzDbAJZT1
3Feu4QrLAU1arh2Fxpy8x9hr2t1AE2d0axwvC/YXEdOMXDkoB+brk85skN1oGwKU
B9IrI+BDG67AZYvwkimGjsjp4UfH8UaRz8wUi8axhQXANNDSxxNp3r13tbM4KjD4
w1+FqGtwuIBWs+IHehAniRNl2eYtOdurxc4auxWTB9rvpDp7pn/O/zdAWMY+dqml
sVKlNlomxIvMA7BkbOA8FtIqO2++FMfSWHFANyhgxeUbTyWPXpGY+iZvHQ6y0pPB
aIiHDsO2TKCcQ5IsOpg4kbAkqL8ZuevXXkf2k7lVYMS3HvOE0JYUDQ4mf4QFogFw
ImPmx+eY/VYXWn3GNjgaGhRfZFGwXpCDtKIfn2xL6LeuXsqKJAaLb2Vpi/DUeKsd
Qm/n5bNbEc7iD8Sr20PTZGSrZpRG5FQ8jea4z3DvlavcrdCytOrAT9RpbssAV2lC
uqcew12b/0k88Z+RBbY1Um60wGnqvHGFrjzxgLV2JPSJ5A/49z7+OBZ2X+nMyDxX
v8oaIYyZVHlYAg6rPXr5ET8XWYhq4Bf6VDbrz6le/vDds47t0UUVk8EUluNhp2fP
miOJkrGZQ4AFb0VYaTAVia5Lp/xEcdZB7io4If/bQYU8hipjGNTiUtHi2RZhyLA6
7x/sAuOGFcvB1a7chKsckRdGpC5BG7I5weUHLEMqt0qgcDHwjtcEkf/D6CtW1sCC
meko0fxWNeRxR7k0OVwZsRDgXzYSvCiUmFi7aCz0Euopu54QAdw37pkwcLAh+cUC
AMwm2k18MFZKWoH9vhO+sw3psjeZOczxXbvFoW8vAQOZIpuwfF28MCTgGYi/9Ob9
IuUNfoRogpUhomw7x1/4DLVuk7WfJicxJ6Qg7w0o60OHwLxqo+OOUIkauIsVtC8G
pcmzYi72PK0DrWmPCcvwQbplDUIpykjsh3lS1DKPsVjwCnc+AtuVjzL6LL9XqJGZ
2IGx1kFJzdAVaobG+2vgqweJWOzjbtVrCIFkZhVV2MHv11b3LgICDikTBFKuX4QE
D7E/LmeqHBWzzUxd0PzTLkWNpK99f37jTfIjBPaczzbREKzcxk80ftAPog0ToaRj
u4gClPME3D9l4tobp3Kf/aifhK+jGrTLq8bv6QOK25fwNszXE4M3G9mKwHyVRymG
ccytfHTeJeSp+XUFT4FDDHo/oLatyXXxPO8UMCEeQ15of/J7wnfZkqKhnUSCe95y
XkYd80/K3UOguNXrk3SKOwFA9NHX0F54ID7lLgmq9Y23a4qJw8pR0Uyg+m9gz3rW
vCk3a3Sc8ToVEDqOc8yUxXwI2qMxlMg9Hzir47KTVVH/mVzKYt8nrBBUiojFXhPU
rRWjAGPkZ2YAXkYxuxJNMKM4FILZRdWvTMItmQgin78Cik511lqFMhXsw4aRmQhZ
56VIIfJ3f+W4Vf0gd8EvftDxxDpXd3oehRg8M5ZpQHZv+s+JR00HqybXFsURnTuE
y9tRUslQ/KdBsIF/TdzvPX0+Kw4Tsy/gwcLsDUe6FcUiS3ApafhcWYwRER08QOdH
v0msJM2e/MhlIHmlnL7/Tek6x1oZhD30t6v72+63RGMHEee2BN9Uv9Fgdbjtrpab
/V4MmYRbbWbnd+zYVzEqghXf6ahUkYOwWUHi80ra5AYBrV8uSHL6+5Wcj6QfFVf+
wyq8VcVuLUGx48VO7RZc+WysP7rFqXp9isU9VHyGWW1DbXPAyGNp3Y3xTI6iyQby
dMoZ9IJe9kD8B7vEbwoHZNmwpOn1Q/zA6oBgPdx5TxFwXuVoDQpcTxMwnqFrLcY8
TC7ioDubu3d0Z0V2/QQ2hZApCa+Nk0ew2J3Na0x4vgV7UdGlU0MvJXzq9gcBIHW1
MCv4c0TGxRztBTOHi/v5UCcaC0tnaeDaQXdQ787poWvFk0N8sqJxGevq/HRC6pn8
IDZfhLQq3dKsEumwN8u1x9HYUN5X7zEEOJg1xavjQe9SDkfyQieh+FmE0TSG5uOj
i2YiB94ouBjPHtdk8DX9PTVilP+onfdzWtLX6eoUFu03GB6dSAqQbPSCze6eRB3o
ZlaHvuQqCRtNchfZHCOXKzqWMNF9DacH7X4B4xFYgl7IjxgBPMga9CtzMvbbwgYf
9XpJbYv4KEh5GPwiBBM/M01uUI2cN0Kzp6Zp1eU8gGF8fHo7EcV7HvpkGSNKUMvR
tFtk+H4DWXhoOIkJJsrYT7EMdffPW1gOa3o7ZauwOtweHB+KbJ/Xr/WXy1T0/Odt
PQsGIohh73f2Bh00ia+ZzVp1x1CEgsoM0DsPGnI4MhRrSnV5Nczc2Cwszv+Gtmjh
2iUzVXgGioJVD4Sw9tw3KXn6M4wrgvnBsTYXKm0Klv+q1aNYTzUTW5l6ALj3ZS/K
tv1E++9pRCuW9MTopyjyTE4CCIFHaBC6lH6xdQmhavNuTL95XIT3Ov+syHiXvHKE
862iHo+54mMT/rzoTlogvwjaME0EIOIky5W6Si/NbvPa8MEKndg/ZRpKcwhfA2d6
SbVmkFemjbkr9tl1pMg5IUVMlnLhaea/yD9aMFqDtBz5NrwSt/+bNEkAYLP5lCxC
VJXYgXYswQLYZfJpvXl58SPkGmeGoXzdpqyB3qbhIMiq8vGtEPOe3lSdeHp+rqsp
mKeiYbNfJZoSJnqRix+LRxAvAZtXFLBLXhHPcHRReRIaWoOOlJ/+i/nSRQCb9AGV
VgcU1BXT5wqd/hsg7tfooKAMZW54DYnum8lL9SRkjlpcsUNapftVt+gPATV+OAVX
rkZFydJLQZ0vbAjUVu7wmo/tSiVrpKBgA3FUd3vnYNzRgu4hEvCPI7G7I+TWlo75
YaekuNspMIBgpE9E3Z1UdR3iu5eO8AYrZQT2m5S6xB4xhpshsXteBFoyDNjJ5ast
oUhAX0MvMF8iUUIP6a8oYYc4CHeyU/RlkOBidlBRLDB586yHWuoV3u0P06+5pOQU
RKzlW0IMbUUogAxgreys+HUGy1l28IUvC3rqMyXx2UMl9cF55vpdqGR1ulm4OkNS
WDpU8qQ33vvhYqFB2V8OxL1EGBVNnb7aij7IsyZ3nlIaJ4BSMhN4Dwd1lHonkK3F
4UCoXiMQlg0zPOgapeq3HLzzKiezJxDvtY+ftHl9GG8W0274eRYtXQa80dQFqHHT
ZSZsZ4zii3ZUEMq8ezGp3OPpzyjpSV7Gd7l/mkstFd6hhirac9Hfq9tfdY/m6iNb
5Pp8XM0Gtdg/Bz1dYFv8wF5L0rAKn98x5ZaYQfsDSegiKE9A0FEbQtqia3k2YCNX
0P5/Fi5j5WPBcRTkG9u1vAM94QaB9p+hsohhJ6HvrhCIq0exMQd+FvDA0WqW23CP
Ft5kg4nd+PIidxjPLIPFkXtEFP90Rhf+vNIBMhbAbLsvTNckYnkbx/VPtenzaVTK
N1RWrjYxeX5nN8shPk/rgnDfA9DnIgmNtpuQDAuFOVfZB1ImTbYteLN3ikdAjqk5
EPiTjQsD4kAybYLKWUaMqsn1vJuNqoilMa4r9NRRNkNjPWgbkx9pfEK0ya2/kw6d
5xx/yFj/IwM9GOB8OJuaDDJlic8t5KBOtNVPgx6bAG3JwbpaNk7waiX7gWXmwxxe
/vAddpPlpfGI/T/Fc/yKHa4d6jwbnrq73gZ/c0WPz52N6/wRc5+u6g0gSAYltBGR
dOrQgWqeTptbCDGdq+xz2XGoCbFzwGWSjuGlsMkyBG0Tp0jPbyhG3j2v2muvSd22
jhyzadm4j8RKHTKz/LgMMnPqrBFok/6PVL8Hz8+ydlJiJRhMWPhmmHerhsBAvOsG
GHqjmtIqzijeb1Rm7y9/dmwm07K+ltLtUZwLvHKenQ4wjAVJ0yL7D3wohgaPbSPL
4+5qvdxD3fpKu3Fo/m7LxXiI7oB2nWLEcIKe5y0dvP1OtsSc9VSOQApTdrjdaYdO
aNZvjn+lHz4xnFjQW5zXjZqUt7RO31eCO5b21Ab7+cUya0c9T4uAm3J9jqDwlC6S
/jE2wyKnJADcNEL6yPWr2YwWOUgfDAcWCoLC8y7Cwe1ZCi9qCTeM64qA1duOTR/q
+sWqAvFDEqy0/mIqxsSo9teEO+lMEZ42FQH+aN5SUVtFEQnBpMNvje0DW7JHzYwH
A5/mXjt1yNBNa6AbQFankPaKvvgrVM2okMGWyMLrhxcxvzmjFt2MKz3oqflm03o1
cnb09GbvbBAEPjlxQN46SsVpI8Lqp9eENbHCyjPV+qkIh8e+7FybBR0/SBFlzn0D
ICu2+WZ/BUTbw2vFooxPmFT1tZQUTa9E0+UpHggWg8JeOblkmv+NaMxulHPHGKO6
D3kmdLxk9uFQPLTybG240Cp2nEQ877SeCWsriXeSdG2Kyn52V+STHdJka3nETPYs
10g1vCTr+yqQMBXvSdD/EErHqrCSyvZ21vg7a8x4RXzag3zTuMmfyK8i69FYvWZe
QQCUebCOm5H0Es7UqcBeFq2JtdU+2we6sCfBAfhWsxgRioIGaMkf2UsORAepG+xf
VuHBjp03BK22YTMXiDSeLR60W9gi5IWbeUpW0Dmz6DKDZdqQF7ZS3fiNZqD4kfGo
0rFjXMeqHX7TXV3SlJztXQlyvAN7vDl7FapRxr3FaYguvmOTfFIVAhN2huiNF/3G
SCr9vNe5pBKqsCY3c2vZy67PF8NMRxLRWeCC9NavNdMRkS32/G4cD2maHOf47Zyl
n4xV/CGyXEvfqJh3L1XOP4U2MiBzumuf3FKAlwkEeVMEA3ow/nv6B3J6WsVVGWVS
wXrGetVH9RnjXrtfhFjGA63qONDdoaoHOlir89m8/aSwqD4elzxC4E+KzNjehJ7W
3NbRCrTbkCYS5yhRanvs/eDmwxmu5rGQS8IAGbX7WHvTEYzGKYOv/70j+cKWJ4C1
KtOFHJkoz4NZ+UZr47MynQ3rK5xZc7muMNiCh0XwYSxNtnQDbahCnKEBycPYe2kz
8Qi4yK9kgKVTa0MMvDLFyOlp7UKlc8wAwzPoIfkXIXCgnPYxlPDfqDsM1+T1R62X
0cL7qhQEfhJIkI2VTSnwRMkKggv0k2Q+ph7dxp4WFu5lzFbaLxgAvaEyDX/MVTB3
EOODU5xXV+NykhCmtqZoUaRTJfFgiuM9AyESMnBiN3R/Xs+1EA4WyacBee/j05xt
Oe/IXh4BXfuWrhznSm/mulrAUJNtLT8EUpgrXZ1hAyppZyQYRSHp03+eos8iY0Q6
ncKORynb46wCYA7N3t/bC1bpU0cd7O4i6eRLv2E83EuZ97pxehuIKDFnWKpSrGoc
zpMFfpO+RbeCtPMnt2y+Fle2ZkO6Bqq8A4+ckEI2K4lrT/qJmU09nYzpNclu3S/X
f293KITQF01gJqXtGn1RAt8E2+E0NaaAXsuQp6VwvmBYwU7473sYxCYYHDNRuzEf
LrezYvr77aNTT99bTaG+wKso81LyKcpuCzJ7NaJMT3vx4JsMMItugEe2HZYNN55d
k0/B7tmxcKwWfJf57FSTyipXWf0ipgxCgqESp6yd65R6B0z3o5P1NZxv2wU16e60
IvPl6Zxj4S01PW32ni6Pt6PsZsD1s6dlVantwbnZABCnK1Mev4VRqWAxPe+FjXm0
eC/T+THXn1jICuEBKz3vA5my+UqqVu6uyuw73CZtLJktVkwNm1RWDDjzN93p3aNq
5+roRoiIhqqKLmJ216J/jEIZ3JXuFerl9/Q1RfEnaZ/4BSOJwfiwX3xtj6rEE2nm
cjbBqX4KdkiHhpkvNztPHzF2j5FFyG4aii3NmOMDnb/NaPSeDH0Xu/f6XBUIVenR
iD2dTKljwoqfvTPHc2i96roPnAA4IrmLKZjtnOmE38UgCDshEdVlJC7ACG0QDQOk
9Gqt7SkZy54ziAFdZSZ9niWs7Er98kSPbseOPbAuffEcwAFW1eQIkq5dN6Gustgk
iPj1zgrZXrtENuEygdxJfrMbCJab4WapKV9C9De8RmY6CUqYAZk1Tgp/dj+ql8d4
DCGC3Nsi2QlLmHmRcX2yJ9JbMFltqSS/i8IRdyaE6RQzfN5Iiq8jDPNavVsltILP
Y2td9vaL8qvnrWEIaU+aNAQhFCHKEU6sYMnhZ8Fk2IwuVqpT4hUE3LifTMOqNuc1
nN95zDD5L3mrj6z1r+mo1BUdAidT3rRU38YYqmjSaX/0IHtaVFPqj9bEp3GMMhRX
uURWo/MNfXqKXGQgEiNdt15M2Kdk0cMVWZn1K2o1hfO0kp0aWQQCBKCg9gsJqsTo
Svj6taoJjnfcFMLXcQYVacTDT8SprSYbae/FC5T2Ir5NbVwdvcHToMXdQy9zEHEV
NuN/hbS4rzULM1yJa85xcSgyM8VaNcBGLjfhzvRC4GpTlo1HWJuOFZVM/efb9wpk
B6wkwHxtRyRqruQ9AyUW6W4pmsaxyIxR3XIY2AQyqzM=
`protect end_protected
