-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
mV8+XlMNjn48/vVI5Ok+aCZIMSPV8bzJsQ3HlKs+F3aLTaC8ZaubUSC3zLp9H30o
9kGTEotLoYmanTRqUoxX8zhHCanZU7X6Wb/CWEERTWBZemHauvnVcQUGVk61snIA
T+ly2jDUlz9QBaVa+KwL7d3f/nAGmTnzUPF0Y3PVJ8Oz7T2OF+OUpA==
--pragma protect end_key_block
--pragma protect digest_block
OIUrwitnA34dmbZsAmiHqZSTLWI=
--pragma protect end_digest_block
--pragma protect data_block
SHrNhUPI6RcZ/1RPw6C53YYH7xC6ZJgC8uYkmmKHYPPXTKCxecwwTOtO9INCu4th
f6RClDbiogtzUwugra62a1z1Qo7nCp9te8r0mkLqqHZbVyhYAuxfNCJp2wrnjzFc
Hpv3NKyJ6UKbhBDt0NNO6nF+B8LWg4Sr/osOHezBOsZgcspYc0FRycXv5eRE1hNC
uuCgv55veWohnTL3uvkPAJ78HUoicsArqcyM67jwLGFkJawALFjOtZDFKPxspFp1
GnCJLEeYbyFwAi4fBceQbEwUkFlYRLjhNz0LoXKtqPlUrJ6jeMspGRFpE+Vw0cCB
WrIefaoWo978Ons7jEVUVfxwSHW9L2luaPz9I3NcF40P5UyZRMEZIXGnDV3kWHOp
+JoBAjCI2xjTalTqNyOZDnkmJRhH13GPT+w4QBKQ+YwqJ6bYQe1wOlAgHJ1ScPG5
vtE0T3YTLRyWZ8OXzPXFGnAsnr7ebm08MRriw5ux3hb5b/Tb4dNHAajhu2CICzib
XaTDheOvpb0PEyOlvYVDgNR1SR5yANyBrzQ2dsAMhQ695LWKO69JoMZfAz5pmJvj
/s+9Yg1m/8m1IocDLv9QlLU8L0efu1zRzSdDacd3xU/UiOXUwCnueVatpl6EvXdb
xVKytUSNo8fXVnjwQUeQB8H6Thw7poPlyxaj7+hu+De1PFT7kD6Uaa1LhrEZdYv2
x2mjJfOwx1LsVQc1rgX7u1dp5rN3u4CkhRSeDlVCgNc+Io4o96Nr6WggqK7MA6mt
kpgyj09YkKBcxMspnTw3dg4l5OYNT6sGYj23nQAewupl139HEVM8CYjAsoy3J/FT
XtZJHcJ8NdhlmXgSP9+d0is+3WbJpuRgU9deKAEz/D9uUVK0um3Nh3VhXIAXFgAn
zPo7j2xDnFrybN0EBPD9FpG3wDTy0VbVCp0RZIw1i0K5XhMxT3crs9RJqlcG/nQH
c18Rh97yWi4fhtwVNjxx22hARohXH+ZRRDB6/0RJLZDhLpGMx/1T0X/0AtpHRcmp
+EREFl8Wnh2RSqvg4teFcD2L5ksTaN5XizrvVtR5MvaEubJSidtU5vkqTcxhL8g8
zYGwMHESypw7wyvSq7+UDi8DeUfzLaDSKdOSv42EV5AsRDh34bRCsJUrmx19o1kJ
Q3K92iHL0/zpFInXFVSKWai1ajImwNDp9dL8QsRQVBvSf7du624vcjiSw1Y8yAgh
71RFqywqdrGCD6/P7Ko4HLZbkOJve1ka8Kjtw7eyNHtrSiBhATiuZP7C9q+vNgjO
cSrkmqq/vbPQm1UJQODTIU66zGTi3eQfmkobwywr2xYRDA/h6tQ0O8n6V1R40Cmv
bIV6m1LbuslH33g379EX692vH04sjRs0YaCU7K31sIVrlQSaOiiynldwl06q+2eL
XAcdqG4mslZWnkky2Bwj13B/9YOBhvC3eBnOfY9yibkgldaRVF6fJv0hJzBfUtPB
nzNeyodPoobmSSS7JK2lxJYTKRDbmf//G/nnRFgYlbsc1VBJ2mvV23LnLVQoISJa
PszHQ9fjfPIjnzBeTp10Ofj0EOHURA/I2XInK2i1je0xS3OwUYy6jruOy9BWZGCa
wNbsLWQGn/MVboUMpd6r/XpLYP3G5pQZatBznMBUdFQjXjLhfVXIr3mNFIDRtbIF
3hyww3ph1sHJFhzApjxeUnLUzUQ3gDwnpnbqLHikTU3YmVUcv6neNIi8/hO+EqhH
lIGDHNwWEn94DshxoNkos8Q9wVcE9oThr9RooOWU48Cr7/rg4HCKXJIaB47Yi3XT
t4W+ur4S/0eIT0UuUXt/VDDS3rXet/ETR5svc3ilDZiS/tfvQzjMDcaMeZM1+HUo
lERGTn56ep/+TDUbJDhML2Wd5EzMWU/Be30dkFE/Qoo/JwR89yXV/cc4qtDjfQFD
VapfTqU1yAGz//94/C8Y07menOmrcv3Ho4MF9x3y5ZBkBVEpWlAAg0g0+VJvp5xn
TKadhvT+ay72k287mV8hHbW6OkvHJAjzx1mlhWOc/sWzh3d0tiVz6pUv0lN+waVi
9I194+ydOeRwP5oiAz+UID2/crbvnU5hxBpABjQanbtJWwfkgmkuSW5Ze8qZTWN8
wwnqkmI8bPeE0vljJ2EqfAN/x8W62Kf4DST0mmb3Sg1BFrSxEdGt2R6sWALwHbYH
KiMCXcdp44qI9hxdTp6kN30vnv5jCbwqnQMi1qw9E+EOM2At8ggQXfGslWZF8oF+
WZK8FS4qoUpOojygOLr2Kfti3BW7hwup1ZsVjzAYGAv/ZoGDf9W3itm/cVivjwhA
6+IunGZH6tKimtzlZLDQNpcWO5HsBLKdG18O9FIQmtesa15vrS/ykedkGZVDK+6r
Q1oSmUpeaKGm5lnwfi3UEbUQIWaadYkwjYpv5odtCN+WbUBjm5cmtxaCBMfVr3hR
0dAjKXXZVliqR74q5j9kVPE80E+qqSbYapswIli1SCV6W/2NMS0jWCguz2TahLIp
QqeiIa2xTWgkhZ7sNiHD5BBZo12X+i/Vubp2dgP20CNMcUm7EgRMzF5zoO2FWE+P
xb2PbW3y3aNZ1S5a2eRiJB8MNGJbfEBLOcfbAbLO4AU7xrqi0MW4xmTPNRnNgHdn
D3D0RUWiDNrA8xnTs6d/0Q2FqGygY64xPOgzlkCji9N/vKq6XpJNUI6obTLwUoyN
24P6d/zHUI51IaknzmiS9QjYhO7KiwSzGWv9h7HOF6HT281IRihpzdv3y/QRwCSi
OoddI7LIS7m3nz5paTCYTZJ7R9JiuvoEcTc//Br228uN+j39ksW/MMFOQyUe41i5
kO/ddMXIvx8Fo2nbUT40tJolCtUPZDJgnHlOxIk2uTSE3q9kiwsMcOjd3dC3Iiud
BOzmUkpcnQOK2OCuF8kmd3Jgq7H/x4/ZNW1ov6yd/uAf+f/i//h0CY4RUlJUdYIj
ygJ+FU6/ICC9IelG334K/Y578Hp90bQi68JuJCnVXzE2/dxG7mQQpc4jkY1MOOAG
Svq8ycddiWCX66ShjA1HhQqUVo8gAyeEBPRfnNWdSJFLJAwR0HrxWbQoob7sE1cs
iAfig26lia/e8tVQNPC4MUbIRUdkUjD/riDzaonmrpYhHRfLawKGuQMRx/g+wEsZ
S2qZbgdPr5OcMBokPXGHUZIzm27dkdhz4Q/PNqcg8/sYuCiajUWWUQ6IVUrcp+e6
zQLHS27uG4BpOo9arJWZwWbuVHhIYCu2eN+ELeCglfb1h6ukKgwkvqT4OfTobSJK
bRN09SuSde9OQFuyvg4Ks61J3N1Kne2rg686R//fiUPHYaLfHSWgrH1XEV9VDzk1
Zv8FizP1587tCfWAo+4cGxBvEeh4FF7mLHDDbFqpfLpGPd0omy/ICX+DDoA+ZhHA
IEV/swcxWv+3vYPeiFju7NRb+eakigmiotH0aLIx/sn8dM9m5comKOtqqJB2E0So
cuhYTmcAoPiusL0qDIVIIGz7akdhQSqvBlUvZVosowAE5jDo4Ld2W7ijf13uoB5j
dlggbre80MwVTh+Cj1o7OPKzWv9TGTN7XXOGbRqwwKo/ZyoTy3hz/xylD2Jq3nlX
kNg4Zf5M7hnqWyP7Fpz3PdROEDpY+XdiOjYxXD6++dPn5MRc0aLxyCp9t0VjxlNR
lego13dWo6m2O+KsO3z49QL5hVr1E1oCwVRDqsAAHsF4ypIEA4FX0AJRqDVvZAi3
38DXBDIt/KBijCnWHI+MCmfQk2Z6YVPVZlwxQaZcQi4sM+HF4S+E0tvfjAzK8YQZ
PfkXMflhqYBlApT12RGtyp18cq4Gf4mbDHWqMcqCUCC5v/TJRxk9imR1HZesy1Fl
b1wqtTDQrn7Mja59TNR/GxKg1UM1GUvCPm40/DjwcUm9vvuaJ6H6td0uY1peMqww
T1oE+/BWtjkBbaJvdYDVGOQ7AFShFZ4p1s+yyK+E92X9J7fIyUzXu8+E6cD7uvvR
XdGgfgjHk8qAdiKzImVR3PCKI1uW1TtGTAwWPMlTSUMy1rr0WmKndPaW8ksCfxJw
7EPv5xOQ+92txHo83Nm0zO/0015+qm/uxJr8zXNm6j9wzr1Pqsll1du9EUIkkIlU
w5Md+kHIun5VrWNNAxWJyrwkt4CPzp/P6bF13NEaqLKOgSIi0YSUsO42aiT0rvir
1ZhW0vlx8cnTmN286/tBBoZSYGiIuMx2ifyHpWb5v/hD6LH/U2GgVo+6P8xDfBN6
FDTKeVfJTqWlATxiDKNJHVpMNkAYxP0V69Bz5ssk8qpCa1ed8QKWbrYaPUobvgyN
gROU0FWTfJjKE6hsTkFB+b8bEQQtowxZr14pU3BwXFEQ5qNwXxA9SnaxDusfEUyR
ERPUCF+UraKweTHcaGYDqsaPoMuhNtfM2h9R8PyZspueZYN94looaHdJGZrncDcN
6fF9yJ8LCLq2hcPx3NbRldYQbVnXmDgQdGQorHheE5hSYMnvRVeOTV6WSyU4AZK5
9ZDVF82dMTV7wv7zOmpCov20laUIF06W849oy68zF75Ke3qlIPyjTHYkwBvmEAXe
QjM3484hXWqr1RYAY/QNX/Yo1gejrVaKrfqTUB4xX29Xi/0pqxaXStWFIiv5SowW
InUz0HoWLwU0eAqVYew3uTrakYN6qikGLRKP4XojG4y3LcuUWqAQLbKFSnNlAqKO
p+NhkgkuvSfidnXiMA5oc9/b+xnwzwasFwTHKcuQct3gWbLqPsUKCt7VpWoUAtDy
O2Hywjn7RyzoIBUH6LVdEtem/v/kyEogQgiiFbB1RJi2xPXrJIb8dzkVakX/6ac3
BFlHRAI82gWt3huIPKrfAhCpy+V/H4YhbkEj4PhBXFw0faBxERMvDZqCkHPMfuvG
zKktiLrc7c8GSrqE1BPh+9mz4ORI76IqJG5915A5TtGDin2rXgZ4trghnhUeNQSx
31Z3q1m9j4hd0C8Si6DsLZfb36m2x/7OSc7XAzSvL5i4k5TMxmHM3fBt8Bu6pL/z
WD9W2xFCjEYw2UAIDPxg2xng1cueF+LwkdRF89qql/nYlY7ArFLC5bHrC18cwA4j
h31tzvCXOVOHi5tOzizdoQp32htwZAY7YZJ0tTxA06VW3hY3taD5OuIVHiLTDbl3
r48huzgRwCm1gpfCxlGT1swkkS4Z+DnD87geujEt/0Cv+XRTPYYeUh/WMZzXFwlM
nQnbMr+pn14w7fhfLIpIbqrilvw11BKt5y7cqBMEZH0Iu2g9KceKaKp5aISPNhXm
h8Sy3/Q3ykCkFAnX4VggoVQevY3nRXafxnloJGuyM6m/sAg3Nypnan78pmxhlYOd
i3gSsotP+Ynr0h1S9G1PZ3o58I3do6b1jt4wTqet3xBTC4ZKzqt1RgO5bopyOAF9
iZEoxdD88xkKGow1fRg6ErjU7hBfjehL4yJ8LUXyMDjlaan3go9oThprJwqdJj46
iyiWmzvmPwJ8Fojv+PjMHchM3E2YaTuABg1YkPc3nphVH35iPa3zT6tQnUQoixR7
VLe5rSagmiHq4lhlkSGHcvRFUOsT4N2AlQtLtSbSkwkpR7CEzU7nXjqNX0CDdRdS
HybzCafqQCdM4NkW6b8jRo7ZMYQJuP93zyOvhpHFiYrUQpUIEwAcaJx095NpiKDB
8To4el3UcDyHqvzxJ84wPfwbOAMYELAfBrjDe1VrnyYgTtHOpz05+G+2xd4UX1CY
DzqEsy73nXfLm091sdHUItD9BhrCV3kMvAF5GgHBCipxBoW1bp5/R3L3R2MF3Bgf
JUOdQBJbjidGhoJnV+vLg9ToW6mxr7fo/8N7Ic7USxYppXB+5NEjOxAm3peTerfZ
Q4Ye6dYcvJ16lB/0N6DZc5M4Vz2ptxvhsa2g5b1oLF6crXVBf84kkhk1iudAH0H8
Cwa2OqlcX4WzHU8tvwvUXQMdfxaHLjDoRafzZCWiBifm70Fjy6XTKCr0OdsV0QTD
2zmyMJ7VyUrgjzuRrtVIe0Txr1QRWX/q/tLdEtnE/H2y5oPWYWzb0jlRPKBtQPCX
12q+BTRKmyRmOgJXGG1e3X5CSvNFIgVd26bXDBsl1vyjIAluNHtMiTadL+Lh3g6v
Rlqqnm060kH9pzGG+FnJuX42QaHPmeQs9DHDccLEG+FkWu3ZPXr8OVIjTz2YsI0S
hMgvcJpSWQebheNaKnRtxssd+93AxoMMG2XhWXPKWyvtEoG+Ogyo3vp4ZHSlDeAn
cAjgCR9ln8gcBm63xInE1hbwtjNuGwd8jwC3FZdm7FDA1r9gLNMXQrc7WBBKVLbN
MrxUZs8bFNbi0vJVGCGulC4SrwipBA7KiD34jYbVLtxUer73uirQSESZeA6TbqtU
ewRWq6QHKyV61cmnXlXGgbOB/B9TGoG+bOQuVSb5b8qDlZaLlu7MxSjZIportw8n
fa5cA+YgMWtZl2BTvxi9Y/eBctxbYXZxM2cnjSp+9VhtVZLRTHQxxor+tCeVV0IY
6FfUxVePIJgeCs2xe80tnrObRFy1JmRKRvtJBblmwAZSSBENfXZHBcj9SS3PZWAO
ZhPHvh5iNGqtGCGjOcKtvYwAhl0gfmCexdDH5bXBQZnBmko9TSLmpSQNNQX1v/si
aPETPpVCkZbwSOBqo+GaZ+12+S1Obj/3tvh9x6jIS9IcaOMjuVkK5Iaqwe84gOjv
uxvXbAkqTdlpgXyGUoTPXKyTG8CLz4o9xL8w0OJkucCle30npS1Z+1QF00yhzf4G
vhdQV5El8tsiAwQMmzf58fPNhrDZqef25UXWvSssB0+y91jjYxn5i7NodKV4Z4FX
HyvTYSvDfP1XqHHyNZ8Y4KSA3UBAgnx8l6pZcQ+vznJLA0+zmz5u2vly7p0yOKpn
z8OK3knpnQQBq9kxEZNEMbp7zQRq9xZla0YKEvXM4+hQyVmJwbawxgjCX4I449MN
G3H1L+uri0URLgO0eM+PJptOCZnZtFv8iuKCGQ7JOlEnnQkita0gTeIwhdVOwFNp
2JI2kgy4lt0XgnqH6Wvo+dxE2bV9Cu55rS0NPqhXJIsMa7hdWX2p0GDyYRJi/4wZ
eS/7lWfBySJtf6BZnNrmAsWwJLoK6rUMYK/0Uco+7L+TFFO/SaHA1NUn1WEwVQZ+
o4s6ZhEYWnPsfV+yhT16jr1HN/eje1C+Hf2Zg5b1CH7WtQF4P7vNTUmdlN1Kd8Cm
aam8CA+lJ23wr2OkNw/oWDgAFJa1q8zeOFzF66k4+yHg+fUdEf/P5yuWzo9VDiGz
DaRDrE1zqfqy2GWHhqScC5cQlh3lcdnm7VnDOP/bkKl8Gp4e/5bt4ez+mlZJIhpA
sbKfgpW2N8RJRRbMrVBJ1ckbk6lecybJWVgz70eo7GiAY35k1Cxp4I6vwgLzNesa
noPtXlnrjMr5NND/DtiSRF3Ablq4XMZYxnfSTX9Aagm++hYrN46NHKZSY5jbGdOt
gKyU75ysbhxYABCB1oZP/3+UHwGaiMVIyzjZWFJP6aliaiZDEXklVytdNdFBtzlx
9lzDBCJdludDGLFAX+hHR15xXtn+QiMKJCHBN3HwgcbfdjzB14OkVxCH5N9uiUhI
0lDnTR9r0Qhig9eMMoc2lcp4TwQ9hy9dy63Xjc1ywf6dvccUM2gNtqg+oAM8usj7
eSrkICfUvz0EZZalqbgZqeVIGMm5z0dddUJgXVOw+U/YfXa5AN99xnFm/0aagt/+
N+T6W4lV2nt0MDTUMaA1CPdSeJyF4/IHUSE7xLSxJabmIwm6Brihrahd1dnGw9GS
1AtHua35ERiPj6BJyf0NSEM+rQnxSZKH5B9AegaQ/+7OmhCP+50wY428I1JfJJsK
uUSaJLcvqoWOygP/kyhGuCtUzJeCHINA6lxPz3gv+0s6lgngJa9TD3xyQP4cKUwd
+Nl850t8BF12E3LC70SBVNiEcw9xAMOD0xPxzkY9vekYtEc+EaQNQci2wIok3qI0
DCa54syM8nbGht5EMef0bT/yldUtaZZutBlJeNheXsiythEFGAbOlibXLtf0YR/U
TxaOMlbxtE6Ey27XIgUzXxn1RziH0zWQjg14bk8EJgowpj2iDDajhBHXkUELFKZE
QzsPai7fOcJZpnicXo2mBHZRtF3gTl29h8Qj2Qz4qnxirgRdC7tlIJo9aQoU6ny3
ekXxeaOXjSnRhc6fZbd7nES7cZy8tm/jwKp4BLAKWQ9Z77VDr7RuVCUYI5i4OC0H
fN26iGlbPVX3CxyDsveUb+T/7UoFoV2M2TKXUY+h1hJPbNqGFekFpXYdgkKPIfKh
vPAjupCF79j7C4x1lm7KunrJGd98tRqFNB5wrP6AKBwLPxIqqYU+yl0zkOuA5aus
Lglh7YQakCr1kh982mLlxhK20vUdKZZSx7QNZ6vQkfSQsPJN7I/NTy3kjAbzA4A/
Ga/j/2LAAeKdLclyGI6I2zm1dxM7BVuwmWTnrM2+5ohe7Da9Jron9j9wG8LAHSlS
7zLMkPRtPibJScn5Sr2EHpgqinu4uiPNXTa1yfA3vApYc+evF5xcO6RfPm8Ww+/H
+f2bEEEZPfGp3jZ+fjqutr891jJ9EGvNNLwZL8THhpv9rnr/9to6ditS39tgZ4r5
2qnGBeVdmUSEG+nn5o7rFYvxEaJsJJbt0NArwBgiBa8UGLTxAJibPNhNBqz5uNXv
7sLJfQUUFE9gHaPAlf/9VWW6gyWotEmDMgFjQ555dlOnC8xc6i05Vr/D3U9lfIxa
vc6y93zvLVtdwL+IArl3b5l1wljFJXvZJPpBlu+N3STpqDfYcQWIymY4iRGEcZn5
ehzNRUVnEsdR4ytNvujnYDabMPK0U90ZQedHHp2E8JNpSdkwWImgrbfh9kn5krKl
fxjYBvfNbfNnVkZFSTTJHf9xgrPfpNNkADvoQRA3cJCRAsIp0R+w7t43q39CgJpf
JLq8Yl7tjaK8HGhmMH1IOfVC3pg7CalCWgCpD0NYZyqx0n8m2iMZdrk5DqWxkz6T
V+4Nur5MGUoGKMZYh3jOH1/XLr2jkuLAU1FW/OXYWkWA1UY4cIzZ30jPQFqTh7nx
I4v53h9lJy0MH3tJDezKSWVdp91h8y/hpvaNr+D5o2YjDGCmZ+VNGu6AoEb+1Dwr
yEftwElVemfY7Kr0N13g1c5B5WsXqLzS8gXJNU96KCzJz3+ujrsEpY5+kzoQVtc+
MtxsWEpsrlhz9jgIrN9MxLy5mmyh0cXTj/D9XMDkrsK+GFdbeHWN2LMQAwS0Cna/
NW/QoNQjTl4CMEmekXNNo24VV0s41D+IYYecQJ1mFAmHOVz7KfUhHGw3XaFaFwVB
Ns6InhrMeqs42ky4IK2dy/uTXN/a8qZTNwV5gUF95dNECGQGu16P83kTGNA055+d
RYZyJKN6vL4YIxmm88wNY0NJxN+uV6gui+ZydVRACVUut621tzwc2lmFA/cJG5UH
tO5RKkjV2mdsivJlPIjI+WDta3XqAf3H57dCfg8hyurWu1ggFOB7gUsVUiKYfU2b
kYgHWSEXT3ORz5kDU+6ccJr1j+YfcNH+PT42aQODaW1X+Vu0oI0lc6DC4vElJAxC
CfP0NEMNxC7Cdmg7CX6zQ1GzC90/rSbCMtehyZfoSIGhf+Zqg56m9YJqwnmFEhhn
VL58EJ8Uc6hunhNN31A2X8k4J4vc8nj3speuuQXSHMiX3twvcgzQ4MQMSxf1OfNN
6ftOwEPz52PpGC6PBH6KfId1Uz1UQKIL0gmmZGDjFJWsciucx1JHpN7v8xcroP4J
Apb/RyeClFI1xZXrxR3NvSJQMIF724n1RGd8+YpYXwSjBClqvzantzMxnUBYvvqm
3xKN89M5zLzRcu8x8enDKm/RKOYP0jKyaIke08kn2SqGqs1rsqIeOeWaQE8MpwAP
Eb2gMCVxn4ayBy0cnQP2ke4X8XlGWECj5Uxm/OFT1nFXhFPYtV5evVRAcinM2Wkz
NKFN16r1YmeKUYLl7xJbejprL8AO92K+9iJyn5Edpij6tXXYTeyyYsAAxLN6VcA/
c+fyJp3Jyp7C4Bs/YgxEp+3FtJuxPb1uNIuuQHqHd1/g/6UmLpxOe0FS2MaJt81a
7QKShbJMDbhnaNT721VGQKctR49tdrVwgFZRx54PpAvp3Fh78JsTO7jDWWhQgAWw
f5anB4tJzuE/77Wg9aO8Qj3fBfe9OYBSbtME5xGMEcXWmQVyzPS3BknPbvsnfZp/
KCpMVaWkMDocpJD6gdWl8HXB8QPFlpywMC0SdZQwDujGhsjRPK+gieajnG0Naal1
Fk+jlpBzXTgcNZmpaFMJ3GxPE9YzsqHxfFMzUYZQy9/G8xK0OB6y8PrMJJLvOG+P
uemSKt0pA/WPAVB35rXGdiVCWO2bM7N3ZpVyDijIM+zHXJBKDe79AkanIqfbEKXd
j6PkrFX+PRhjF/PMi3eUOUkjvXFuMocYVvOONBxGKTHwm1ZWhQwwdPE+xHWJ7wqm
sFU+UffqOnGkem1EV4ilD+OszSsxMWii8KIZdBygRIi6RKhHrvyeHL+/lQyy330v
LlZf/FpUsVXxs2qNjqR+NqVuVWdGBR/O27DYsTlx3+BpXxDNiT6NiBPza4x/bubS
+wd4YIopqLG8PW23Dt+Sp2ImOjs2ncBtlxeqUXUbMLsSc7GA4jKY11H8bKzMhMpH
nS54WaEfidIaw2ndqT6Rsg3yTMvpsIVOo9qt8ffaF1i5Ah197S6Ju2trWtqgI6qr
wJbspsEsOCSL2vilvvAKVnOUFf1GC3rV8fAFwdJIyGGK5szfY+1nsKxSzmH/6ej3
DkdXuc05zl/fl6oRi1dKLfObkSW78taC+3NMwJq6P9ahzhknP8zfR0Zk5ysQytK6
pjvoSEdsnN92WMsLAUppmtvpfStRavvnfor+uz1lIOey0Wo90sg5jzxnBmErQ1HA
HZjuzeUZyVRYw0QfmONWZKqDR3sMTjSKaltAkHlkZL11lXb2ZZH2s2rrcGN1jPRu
Y2ZQWPL+uQsibwtwWVwMLS0zhzy/OnQJTi7tg8c27nGIP6drnE7QclxJqxClOrbO
JnAZM5LR/qvnai3iU/BcN3mwVV094C262iD3m3MwojvWbqk38LappcmF/BMceGf+
pbYMS1sftPNjty/ZJp72m7mgiJbVc3ydJt6344B5L22fvbCoFnuXCv0GhqTjZDIK
wAheFfSUboRkQmrwku7jj7HW+q+ohv15hNxNYnVuyDRbDfjTsIQ6jU/KzxA/GxSz
Y+kvtNCGS7/Zum8lzWkr7kXyp1dlTFxC+QR9aaJkLAiiQttfifXMvTC2BcIJCa3E
49/nzPCkeYg6SvONXRrFIGM7at49gJJQlhII9H49uUF0cbJUwm7N56UGcKYh82NJ
CaKMd5RJqoJaVXdAYscYs+3675retnihmrrz2n2mjH4gq7CyGkLRueGACelDtRTl
Vr3fjF1wu+MWc/Edk7Bwh0+ykWGLkUurQCRqMK7I+oTdercaDQl0tHz4Hy1bCXW1
MGFCPudYPSciFy8js3Dz+aHsOUPoN3/wqXEnoBlEiCosvg9aGO+9D97bdA/udeL4
GRFn7Mw1wN/jMgCfFa11dtyd+YqL6sJDGvEllSSFUgxdhJAPbG+0ENeh1QHYO1N3
QzZClfSnq08GJyNPCf77doGH7NeV/MyjiiaaEowlkX9FnLuC4dqtJ1HllObU/jgl
QltB68t5caAkhN62A10naia1UA47AQzV1j8uaxC11BG3kFY2GKdF/XHwYuG8bI/R
FaUEQLaACfQPQHtJ0O5DlYvS6GacB4aI44zkA+2Sh/P2Vx6e3PKPDKB0ygfjgRd0
qJT2w2jErgUh/2lWxs4ILKP9AW/l+AeEIjCcUFlX9p1Zjyk9HbwhIBbpQPLqeYKZ
RVx2aIjkeyIDf7j46t7i64BV49/48OgQkIDWx0+sozKl4jVodrNGQs+j8Vm8T2gd
Z06T2unD6ULgIlVQvh2hxJgINCvSqZx22JArLMkOdD/8n/1WJJckzSxqKR3mwknB
WWqzMYh1PG2p7SR6+RLe+hUseBjvFBUXcOxcyhMNjHoVDIu0RpbBeUZa4NDZagf5
Gkm/QLHaQmin7lCUvyJe2alBFY6OUN5BzGlEOZwZ8Nc31jPuI34z7CHX/HmswcSo
dH7oXcWa9tQFLybDjdmeEdkRZNlP+RgEH/QtUp/e+W6ihm6AGfta6yA9S8VvMtTj
rwrELDkoOavUxTennDHPsb9E57VxtmyoAi7/jzSEWYkhgtfsOmzqPbQK3KHTCWEM
9PlGJed1A9EMijxvz93EpX7/6RoVg9OH+ZldwB6rvpiQR+uVqGsD0B6Zy9qUQPzc
B6T6Le6CT+m+8gB/0c1CKXgwE+ecMoMwTbzEZQwVdFUbDL599amLdZQEesGUBpLd
WJLuqpuhQekp2jRtTy3sGMMnCIEJhQ9sJh1cTCV4YJ+/TkCvUZZGcP/hqs+UHL7R
G6YgjBH8Gr7JE4H5Js+fJwL5KhEjWNDnc5s9354uVP6QEyDDbGLxF5Dr4ThVo9GG
JYNk7bA0HLPn0my49+ZL1Yl/A8+yI6ckOwS1x1PPK0YeJzrrWzBRjIk6eO9yFK3V
rJijdKKopxxMrKP0MR9rafBG2kxvUMIUaqvELfpOOO0/2BjX63ukM15yDB0S7L1B
E7OrvQFAQf7qMBV51l7CPj7AgkK0oardZ2dssecSGt3I1/UP0I77cYRmC9HxDq3O
yTr6qTxDEcaTSai8i1vDFW1Tshi6TTopSYK+Iuqeh99ebHBzNm7vcZKgqEQOjnDB
Iwa/wRtngzFOehuwbF/97hLoNMG4kcCrJd1fvwDGYzSjyF83sOw9NJB5LXe79IGz
W1mbvr0vlPFTnKbLMi1CzoS4hFUtzyU2w17IRnUSvRcUuMJ6eWwuWIjrwmKLPfwC
BEG22SvFntqphtXnXw5uLoOjSlTUEgc+6831A6jLwk3assyBZvaI/zctYiO4oXPB
cueEzIBG9k+Q3909uqTKmlcI7nYDhTc1OASeDTHdA/iAPWyq5Ssu4T2MsCp09PYh
sFPCRkLk0rBkRw0o1u85R49UXnVKLyuCTboKqF2GzKc5lHpC34YdEqtV0jagVxPZ
iEiW3iAn7BaM0+8wtnYoNG2SbGyDkBdmVvoc5yy+1wXFLYUYOz13FLkTdk6YLT4M
p4zMZRnTnN9qJs1Rde/TJ+q+zMhnXbcPha24yF1xTzX7jMYrzAe2PxD4P0/XeWSv
FJnQ0BW5XYydRzrRd/Tkdnu71YHfaSslvu5zBE7cTEDtX3J7kMifYR8d7nIcdd5X
UnuZvEBMxiiLm1dXFRR/WNRmWVMNoDYq6pY3lTilnyMZwEcTz50ug9bShwM5vi8g
eyGwfHTVKXPWU7SC2fhEMsXqZMDS9y/vBXOsigU1kkBDVe/8HP0/ZR1JvraqIclm
COIysHO/JLgkRXX7I8l9wNqjk7Bl8vmb5MJvIsODarljo/qqzOiVpPGv56WDMsU8
NcQYXS9ZTXtv6yGuVHQNPJJ1j2jSUhpWzyoTZr7rsoFDUvHu67sVtOdCxgfsNd20
gHekYfFIqxYAfM2mRPVI2JkBsMDejHX5Iq6yARYOGlzSEg9GyJe1EyLSQrov5Ewv
gW92UDGXQ3rzxSQWHXxIlZjriGB62+lss+3nF7Rupq1qtrY9i/A1+cmPMjrRvpwy
g9otAW/5TBco5gk7iKRhp/8CSdScDTMwM2eMqJKP8Gjh85kZlrRzgyEuN0v5p3He
A6k4XraHwh9BT2Io2xWoXf375REsfnC0GgR37j7gHl+UQ+/r9oRU2X3HWut+Isrv
o4MZqhAnLAN2xOEs7/mozgs/h4rEs08UTFKNiPoqr0OgwBTuhIaLIDVhd2RViU9x
Uw2NdydrhNI5Ohf3cUTaioZ/Et3je4TyX2FGf8ylQcZiFL5Xo0MoHtAzW6aHfmLo
Gs+yyRAnzOKO0HJSkzOzAbhRbHf45vBQgEHJUVM3aXG7jqx5JgykrvVfz4ElxuyB
SMrRhynD741F4YrAga4UU31kJOYQYLwltKxxR/0PtMuXhMqvyqwCqJoh/lVleyGu
qAvPUcHfeJ4jD8bXsSlJBVTlL+cmD6zy8POJgZcJPcqGuiSdWH+7sIcLk4POMaj0
do8tsjqxz9kw2dzjGA+9MiB6EgsmXXOnTl7gZvx3Yw11HbsbaPFyfq6DgcERWjId
x/tXBoFMjHFN7b+HtvS6MntiW6+FBsQXzdHcE7Ev8Prf/zA/RxhaHHMBAM7Ej03K
EZgE7l4CRpn5Vx5DzvCAj12jYLSukqaRGUjmR/TK0BBYWOYNuDH6B2a8+EYWMjo7
Oi5WyjW6bKmpqeN22Ify3k0zCkXWV4ymCnSUsHkf99e/WXEzWhMk5cR6rwBmItqi
Y0AcJC11X5zp+PBJF4p317l8q2I9yLae4WRFxoLcRIjzHGYYcLVSbNVg/ylGLeXZ
JayxJqKdo5tKpJepHmU1E1Pz/+hVjPQjpAMoH1DNPUVZjG8oB0esalA+B88f1fHp
fapLpl+TZ6B22lbNkNCZ/QhZFAyYgxZNkCviBaP06ptsFawLkJCpNQ6LQGOeslI4
vCYipIrZ7gYaDvzlGrhn5+01dz1WhcQg1XMTZ3VOtRJhjV6xU2u+qYa985aWQFf/
fzjGv7zOkL+OMHMxx6LG4AaFMJamGJpig56LdIhn1t6sFl90BOTRKr/jMm1h0y2P
gl/D3RnJ/UOoR3QMQZ8wv1PgAoFXVUyBkC1YTAUI3CMfXJrWVJz7lOIbLmyDjvFm
cxriAN2VQozCD9J0+n0lZCSTA9tO4idO1zmURFZStpT5vhjiiIrGvCtp7QPqhfKK
mvLOT6Rx7hhMpp8nPaJUypkozNgKAIFZvT1ohOYYdOQr617QgwY452gPMHJR5Kqo
pGsty94PbmxuYPLFRXsCech/udFiq0bfuTtG5sa+/K+sAJKV9gX8sVe9icCwlFrb
HyUvfsRhjOAJOP9scSznUPCbknImfeQlfe1PU7jrQuNgplyx2YmWi+I8QknuUIoz
/lYacXQI08d6sax69x96jH7X9K/wS5xPlpk5SfBG6ErRqF0ofwTYQ1U73f+Li1TT
QDS0ra43O2STQ2QAmolS4gC3FB1UTM4bbKKg0/LWhqtheL7T0J7xjV5JppRHTEQ0
TqO2VwMtMPPj1TuABKLMedvmuMsAsNIsEVD8P0r4T9RjMUnq4HpUjP1QUggjL3OZ
ed+DRvvLn1M9N9R8LPQq/Y1fajnWbN738nloHueijPOgHQFgBMitinXNFJLfnCRt
ex/qrBTIUGqD8h0pYJh7ymuekJhvs6QcB1+aklFVetUYmJ2VTeMsEvADIHoLvoO1
+HnwO3L+DCbymzA+z9H5Z6BLCGgRU5a6enN/PrELd99ST5G9F9jLgk3OzhSWX/CU
ISxK/Jt/U5suuwhVqZC+gfmQrrvZ0Jjs1tWVQrjOvjkMsHCeAJnYTJ42b09SzSg6
rYBc3ufIuVVTw62GJtQsFQi6DMORkU382xrd5TPVSkJ6SeasLAQi8Ae8YU/0+rp3
2OxZbe+i9S0SmuNNaGqx/PEQR+qWv1e9q5ZaWLbb+5oxoiYfY9/GvVPnpMTC3m75
AkXQHHSDdGW0mnR9yTZ2laqcLVuTs3VNEkurIQ09cgPM106ybtND+u95RMy8Rp8Y
hG7pN53JewqerRANjkNncb0qa0/hVN2TdmLvDA0vl9GXRts9iJo3PZPAC/t289dq
o4gaBHaI/W5nz2C3y6u9JR5Ng9wL8rLXLXpIid/ul+pFoCFjAXZ+o7gnk2Os4e/F
YAcHT10T5oM/NJoeH2bHJMUtOzZ1SE8yqWzN+X6F58j0lFBxcvwmv3vvEygO2wPB
Fll8qh5oYFv6PM19vNUhXWMT6Hd6JDv4BdDPE9JFsA/0Eynx+7zQiMJoq5T2i+Cc
Er73x+nLui871FYBEIUBt7l/U9qvNYULKoeaLgHIWNXV0ckvmlN/FHTpRv9pon7i
jDtmb46tOZMyaJhRvNZltqwYrcc8x4zN8elyD9hrS1aXRhnweCFgTMhwemUymb5d
x+1bDezHHWO64ji5GJKZPVfwTDDyTCmSblRSPGf+i+2EgMkUzRGeIK64mZQfSsfQ
j+aRdaIK5Z+D/dC9Kgh8XbptqOGWes7q/QqNYYGyfeVTp7Aqx8ztNBB44NeLpbxC
cx5ML7T5xf8ztLii1way6iwWLxfCMXv203w4E8I2Xsl0agI+/tThuWEL+6GvSiqs
JriuwU/h+C5X1z9VOMws36CLYXYhn2DOd2Nk0eu1tYfI9OVrPLxwe5jF1bijoDyd
gg+522UqFDTJkPw4lcdCjRjBBXemRkSMxmlbNfzHBu9zu8Dq3hGdsFokBLdQQuLG
S0lq+m/bQNOZZ/FJ4ScDaagNKhCBXeW+xqGgEb42YZBUrI8TFCnVbyNzBSL+j8F2
UVEl0E7UE7UcLa+4fkJqZD7EyNS/21lVpgGBaRi2q6ObYSLGKrmBcW+YSznMujUB
VSj/zDbvZTJJCUqFPf4vhChHv0GZ22FfuaCcuA+ZySg9wES6YDUydYOHT1ECqzXn
DZV8wKb2DsL5kIlNiU0AT+P2hN05t5YeV4g+D6elOI7XLA7ZuHuTl1NVmfq8lwQp
beRt1UYCevvtgxixmXB4MtNRD5cz2f8m+LBLzbzeFigh7PJHjcVhHMHKIvPMa/hf
jjXdjsHWdeUXj7FFwnsFobNdufPALkWA8OHlXfWjla+8kEcNgSPTmVNZWfpTI36O
d9LuRrcsB3hKhnvbVDpfD+ggz9krKSD+18Wl8tcxluwD+47bxB/hTuIbwb3r2kfS
NnA4xx/Bb3r7x9oZxVqo28eEpTJvFMpG9UvCGyznoXB8GaflHFDZbJGE/YZlV9nv
CQBjlA9S+XXQlNgJPjPfsYdYjOQIT9Q1YyC+bRJaDJbjUnODFWTIG5u+Mn7DQMll
Oa4O0+F9UOvN85idOoXNHd5j4sNESdGBaZA5eOZCBULknifb69eXtO5dLuiGnjjq
diajR2zwpRdJEMwqt8h2ggNsVCi98Yxcl1EiqronNfVPIBPiRLNw2mjUUDiyIj8+
FMW5anmKNDKbisKWVPIbconQEKZ3JTrcQk0bG2yB9Rv/daYCNztQTNwqAIcU5RCu
d02RnxYt9G9URLUrb07LbN4IavTFAUZfnccMk3LNApIcB6kPj/mCTG4IIjxcngRz
OafWj0+PCr58mLrsWtvHtTtqfGdgiTnsWu1rEjHWwDtOIo7H6w+621X3XyhAOzNA
DS00rQxK20AkiKdggSKhUqrUv5cwP6JiMRHOkqIPzePLD8VyaYdRnBTIbnGACs1f
mUxtvrVw47eAdIDgzjmM3PcJyB+FqURBerdlr1dtdvh9cL+jdsFKhNNEmBBuSo01
BK+u4mCzum/Nemqd3GpWRF2IiuecC5dMFO+21D4guZBlL1E8DHVxWXWEklYC4l3f
c/OeMsKHnuFYrslCsDmYkN8gSlj1ZgnZgsSdVHZpxIizInWpjwnVyCrIpp1QIvUZ
4aiz+bVSdjbw9jZkdDISEKCtgoAFE0Sn3lv1dCEdE+3K8Z8u0s++/DtUxFzab+am
T0K0WC8QVSF1ZmXvicbXR5r4a9Ch30xszv2F43QIQV+DmA793ZU09gSfqW86VJfI
HMfxjr7O7OtJI6xDrzMAwMeUqE9gnVv+EfvbEmltRx50dzUMlsiOz8+y3U4QaHUh
HAviEEvGGOd2jQXTbQeMRhlEH8NH1q8YtxmSyHvnF+qpjbVznLCIADH8iwNaCS+J
TfOLSYS0whrNAw6jxGnB8lrUkKsd/wPFPG9j5UwgBgFsi6GP88tvf2QAOy+oAX4w
QQUL5lLSDMDIasMD/8jI0o1X27M7crjDNFfLndciYeAShECNwnNjOkigEVdAEiai
UBkp5YPkbP4ALXBwG3erPaNYga4rLiyDR4REIzyYWpaaeAD5KHEIQDOofPHZtJ2f
NvN2Jb8/SBd0NQqiVztFQzCPsCxDe8ymRMNw49uwmkiS1Qfm4riT2NZj1kv0OnvL
FhR/DwOya9zyjWZMPeUXPi6HRPsFlytFOcpz4BKtNyVjHw8FyBV/k2Wj7VIrCSyq
UXLyoLsHzv2Vqy+ds+430Rl73Vh8aEpxtQq9bzE+NmrXRHD2dEbeEFRThCn9dXg2
YxzhRIf0Fe8nYxRSVN8xsBTAaw/NNMmwn+qHqD6Vhp8LgO90+FNifybOZOIgH8DX
Pk7GrG3YzrOmc9t77emwI7IJ5pOGm74+SLrm4pjNQuo5cTi2SESC0hEamRXHxueg
ExQN1lHRrokH0jNbBcECFPzhG0EcvVqkRQNYPYLse6cY6zIDtDd2WwmudO01aSoM
/EExgZ0+MzeA4OsqonQULUI+PilNdPc0g6A0+cbpjA4u2B8z4lUpgwjFD3QqUswP
Xg+laKG6R0rzQ3c76Hm8vty8Txr+/Qc7O5hrmMNYY2Z4JUxw74f5uYZ+TBKBhA9W
stGcQsnRp+LFWzy3UN6cgoRFRTC5ctBLrxlaKZcSJ37+103uysnxAfeb+28BV8rg
cm3lSmhMY67Q7JLkuYtq2dNXZPxtLr+VMt0h23IRIPK8YjTxIkT7FgNKl9cgDxhE
+VScrcMYNUkWBczl2uwS1Sxw92yVZRbd0RhJDHMk0DjGXLqkTc8ppOorJJxWacOH
mvesxr+h5Hv2mFQi58fS0usSrnw+x8cgjvqLdIIdOJ8+VNhqaUSS0FuUn+JyQZ3D
unsGL8piMyCTOt11+W+lq8+dS1mi5BvWeQEW+etGnSVB+lntH232KKOJfa9ZcTOE
knUhgltpd0kJmOLXsVS5Oya82D9zOIkWNwqhGBrKqbHfExNYsMXQZvp/fDmXYO08
SV7thTtq9baKzWDbxwdNK+FNtDgXwtyThdKyE25r+G6Tj0LrJETFzeR4lqPx2Jvk
3LWATzhoV/PjjyKMKUxMWapvQLiBUDGlcGTGnlB01hEQIY3kP9CLme2NGwjKEtPf
qXVXpb1geZ3/nbhis3UVyyNsE1TzjIcXbBXCAeVoS+LrfvjJWQLPTRMcKUnh8QyT
6s/X4bPwKk69x0Yaw/fhfBdzbDxUplwqDZ1vfnXvrA8RY+L64Ib/G40CaUaI2z/2
k1IDzrl5fdkvteUiyQxWrlEYx8IdOEKRaUxomiRTgfdRKM29l9Gh49AWjylk7yE0
rfVJqDpOP/uP9DrhL5IHnMhgdi5CB1SdN+bmrmPnea7kT35cqqcG6sxOBoxsTVtk
W/XboG0nacJtnvZi0gqAP9nGg5jdAd8hEqOD7Qr7cuedZQkiTA2fBUtcoY2rtr+m
+RNeWLnx9UBwxyFylQgpLapGIABaBXCc0KFfsXslE5DSO2piW95Xfif3nI2e3nJ/
IX0eE6hh7mjlIsAZaHu20/wzCV+xCumkJpdumJztdU56fIQovVxSXxrFxMTHyvDD
gnBt6KK/hocej5ulUHfTyZqijpJ5EN4bT7ItSKOmv4lCMsprVoiJrUEfCCeOeawu
+PzH9SHYWQF0DR8+2m6JLsNIOj5aJiGSNWeOp9YleDK/TRdN5Wk6tWwrFfLJ1u+U
n0picLTgZ0S1QZShDXJG82uIsINseQhqGhO3+IiPeDmYZBsCXR+Ux7sVXvJCeGHD
9DpxdU4xmRorUqd5aW/UJpbGIDNWGCHpNwt13W1HUynJ+sFYxbVQMMzshg1hGiXT
zhnA12dJqMrKsT8x2kukJDw54LXUDzI8b9KYjnTlvfvDtv9TkjQu8BQ79Rd7Kt92
goosvtbOpm4zJJetHslaXNoZIXhynq5AOUNLU+b+4XVoWDO1y7SPkOIgA4ywElTA
tMrdTTIU1BlblUO9xEHDhW4VkICM0LTkEj1oFbGKDRNsPhM22oTWh511hpIGbzLK
qbTeTmUG31Z+kdD0WBI23JFwwmG0AKPlxD/HNoDzKrC9TJXRlbPyGmF7XaDBqRsJ
vmLtNM280pAP6Re7II8Nj4sZICSlvcKulUUWh2oqRbL9QT3aEmHPBv1qxNtyxvzG
tsz0UqX8EcI1ty4SwCE/TqQBGHqsFnD/67hj/zi2E7U6vlx1Pyw8832472MtAw8r
Yp890Wnb7J4X2if1K/GriDw8/tPckUXTZIH0FoQxnwwLsCP/0K6XvUXekKCaiz5/
FgvasDIoi+jxcK8cVB2QgONztbFdx52c5eF6k+5sso/jSORWzF83QB/gKUd6lfO8
+WaNVdSbJF67W7b+IFcmPh/C8p/3OKboUY1mQT6U31amIKKW3tm1rwu6K03AdkzM
d05WyoUZKn+v9ygWV3aHqUyCZ9HZR792BNveeaQe5Lk8DH1sW0MIreBPoLk5oSwT
DRB73oSEp1tz/EtSZsik9XepPaJYoa1Ue7bE5bq2W8oaRfY+NIzc3+8ubkdzmFDV
vXUycbb4A7GgVlQbmK4ngX7aR3b3vYfdEpjlr+XKVUjfrFM8H+i+Z8VGn0JH8Rto
IL1wKxCoaRpKBddzhVK1EC+G9K7AK1RkhkY92m3+YsXdBxoj0ix/6sVVAXYv4oaI
4wBobGUZXu3Aq6BPoiv2c+keAMsndtPwT74En0kXv43agdvJbUdUe3zYnfQGoV1A
OfGpN3LI8B6Y2LDurfIO13QYUuQlTSX+8jaU9l8KEla0Qg8lMjVGptRLfXDw++J6
zPRcOFb4TLDGbjGRqTpmv/bw7yvF4mXB8PKJ0iwhhc+UjrDBn4DE2YWL2nbgerXv
3vW4nMNbAio/i9e05TeOQ3c4KyM3JSTrU1QPCYzmCxuoVHpK1I8NSmBeDyO7BetM
t6ny2DIzcq3FdtoGYN/0ibEVIQc37yNjCdrPiYZhPQe6LV/Uq6WweUH3FXUIyW0X
dSgbPCrMomKROSCQ4409pwzXVDJj4eGzO7C2hvZXfzAjs/EO06ns/A+LwHqDNhGh
Q4K+BiQBE64lXLa9vtodQc5rZnsLz6t2KqkW5Uj+dUiPf7skO+JvOxPaQNgb9/3H
ljjdUYV9XL+2puSRkGK+SXEzfPczTlBEdUegqBPVlbcEvZoHeS+VD6Zg4K+eAtOO
OJEtxediixaPW6GsOCExr3j4jTfP2zKaO7c6p4hCX+LRrY+mwBMK+sOpMPn+eAUH
0XNNZF3fty9CPiVRVW9Zdc6NKprFBwGW1HwqqorrWyNoiK2yOuvg7rzQ+T5ovLyR
0pmsYtwjFhMinhh84/zQlFUQy0nb9XUUlcg/9q/jwvYV7QpV0oE26kEa4LoXbOTU
YO9lAYtb3eZsQuhxpccepe4xhukCvyD465QhKDsZ+X8HkmAhXkFd5I1pvm6Pbw6/
Eh+IwrVzJNLZsrQu0XtLe7CzOKZN/8MN/DwR/mvoFWAs+gwDEnSSuBlKxyknYwKg
8D11fuj+eImfzTRc0vT2JEFDpOEF7bBCdQuN9y+W1K/uddP4t16NgT7mErQYBea9
FH7bcN6zrQAsICVSIqexNXvO5qnumlM70JkuWLDTL8NMiT7VfV1HxskqnpllzpCq
1h3zqyUHZ8JLXG4wHw3v5ooQvl+5lk6mQY+BFqQ4FRAf1rYXLuwpom7C/Wi6CJAp
e+bB+A2qq5CaZVEmbIUrllW9pDjys4ZIVnBaVavZVwQ5JCLY2NSggmrQFsVWUavy
63i4tRfhZ5K6aAjHMPUub4vgrkIh0I0GBhlqZ9elatAIKKLjAp2iuesxcmQsEt6y
amABRyD7/AW68pXjiT/IDi1Tnn7Cm86lr8iafwSI2KggwauNVLL+CN7NDTGN5VDa
vPlkRMEckobOY/jWIi2mLF7iwCth9luboB+lGA86I5j76+selJYX6ebqJWrLxYN9
8ij/zKNG/ts/bfXcL+f53t2E4cMQLpFcHagtAzUaW7YYumsX1pF8SMW5Kow3aQX1
GIxo5jZ9oqoF+N1UoCyuLrl5lc63jexk6AZHEcxy67s/v6QFenLdcoDZpwTlyfQu
w3fxNMW8od0p4vSX7NObhcdkBv8zbKSNLbaANWLUuaHyYI/jI7MbFBp5yYnTA3jl
2Kkg4KcjEFAL3yvTa2OCItY9zh9SKNgHPuRGyvVWVP9fxmEMuxvgLUtkn7FAqeMr
UtDnJbb08CA6Oa+TzqBqYzdGdfky17x5xd+kAM+OlNuZLZmNBSacveWv/Q9LFpuy
kCOXwURePlRq80Rsn5i+exZFT1lmEzuN4ZGLlhf8YccdsXFfIRpjnzcLzT4R8nQ2
F/89cK7+ElR0ZagL4AMYDMRhSQWbHaviRRkqgHUEksG7+bqtwXZYI/gFaGOnr+df
GKfko4i/IW8yn+hdeWliwnMDPGJeMW6IVmsyZF0N4YJwSaZwkr9TASDKHtUMCqL3
KThd3PQYPWIKB52B/Z1neBv2ixhy4Z7GMMO/SQvgOCeVrWViwGi6QHJd3umyIKdS
8zOT8axVmg3JFAF9MSvhFk3lQLcRclHk/dSce7NqV/kDDaPkdyc7wPS0NKLOiNiR
V5M3sf+3ji4/WU46FvHaqYjgmPKQ2u8IV77iz5D++OrDNN1WZD5VZTm9CTH/8uBd
tAojtkyGF0E3bA78oOAq8QD2Gmwgj+SY8zDGfu9bjoO5H2C6HI6bJAt7V0ARDn6h
ZGE8jqHSYIlf48oI1fmrp5pBbIW2PKOptmiZN6CHcl7zPXPV7P4wFHT7SeUhZCZe
IewYQkGFK9P0RHODcohYcnHM1mmfpQrytFq7T+iVHGhvggvPwAqE7XPRfun8yrgh
sduqbBBiqvrDUDJWE8EqIQxLXbepAonaHbelEupVK9QV0hgJvvfZhUIRetTCkbBf
mPpMKQZCXfZsMK8BC1JRTZTWZgsvYTJ+MKBKnPnkjqdvd5SIGpYvtzKd+zduWyK8
de0KO5vUAE3HsIkZKTDHbs9pUyw317vV8SExXJLGR/7m2O2zgZr+24m0GK75aOpz
BtcTs/NTLt0nb0UcGcDUilOX0zB1J63o78vu1qEHs/9orOlLPDIa4QdYRmLMq6kh
LwwJ8uLB/fauJoIlBs8rv43DlEFUhb+1uGa+HYpfS8m2w75HlSS3HMsHGgxbDugt
otREplJBybSgpXK0eikEa99c74bOOsK79pMmsMd6Li9hEvlAPxs460wfhMG1a2Xm
hjmQJIUSVo5hSgZAYkeFpjzwkLT/lCwB6qa9oqrhWbsF70XDRuS7m0i0+cPAJmHc
aErMgZhNXY0Xtjk/aVY7Zxyatw7jbd0/aty8pxBo2h0ThweiR72/YGsLY4rhSk0y
pxBJE5mos9elucCJ4x92p/tPj8G4wDkgiwUkyrrCk86aPcFsrCqzy+rPrTyeWdcK
CEad8REHXZ7wjD34Ea8dFUI8sCvb5L8Gxs/23dVB05S7/6SEbpFeNPNTQRlmuEFv
TAFECqU2YXej/wgzqnreKKtqMoyLYsCxlOof/GmAUnvdL+9mUDyrn8QBgQHrxdVL
PuIAlAYmfh1HJfd2yE9m/uc9c1IMCAVIy23BZOje7NXpgLsfaEwMDatcjIhKzpFV
YV/y8BB1tqvwfVzdQ5mjzZvkuJ8f/IWUoiImrLixGpptjnxZ/ct0+vbJXmxaZbww
Yaa+ND6hCtjcoi5m/etWrp/WceOqqte0cXdVZ0JfeBV/qr3HOmvoZgRnmrv0cewT
FhOsev/AMKjXhlKSBeXzrC5S9SGi3pgdLfbdu0ZtEJ3BpRxObeieBA4/3zzNlIhw
Jv1ugJ+299jNVOj0DXYSy3zwJIfYrpwrb3igf37eAyXYSVtGXTSyYRSgSKQYH2SB
JcUYiNC5Y4i+i8UPp4hio/9BsKMmDcheE+HFsA5Bd54a0F9NdgP/CucSnD2jeW7a
shM0cX54gjm0DlQoZWIL0GDlAMh9sSZyvxNQIbOoC4A5nGxjQoVn5nv+bE3mbn3I
PToubfA0qAbh+EbhfXflfJ5IWLq98YJLB9ApHzAhM9U40+yT3SiplfWj9QXTKmE/
XRxEGLh2id9AvkC8U9dhzNM0lD8ngqEGO24/z33D9lxgc8y+Usm1NjHBoXGnUL15
0DYc2+apYAF/29oIzkNUu4s9suSL/Snyi3H5fIlzPSEbvdxtbpGG7iUklIsUih4v
loseyL2jknhAKVRl1ggweW7r/yUkmvLwodF4bqIuMdB5bv03/G4CG2LNrvBPBQKX
er1DML5K/CimVlgVs4AMHFPQNF38u9EBi8ZeGnUwxeeaxiAE8v2zvgs58glmH3cs
u/lhRr6PJqF1cjgtECWb2orSg07klo9yyR2H1zu1WCxDcjJtAACAd9EC1ZNPY3aC
pTND8L85H9725JKcxGvWyVnhGP2le1V1YqRyzXUqHisNShdJrNILyDaiYi8WSj0f
Lc5QzF+vdNM2n4q2HJGLLkzng4NKrIDahOLFW+k1uErZDpGpwSw2p8LQj/66ySVS
BmXyK+DPjtUhDeLMJiaK5EjVG1HVsz5Mdzlk7/xdfzTIN+s/4p7FVaBUwt65irLp
3JjsIhgkZE+eseiucY8IdyXezw/EAjP9Tsf2bAl4UNfG8vN5CXvF06a+kPmDQM6+
sk+MDb+Kgm1g/Ri/MhxGcnBylgfbILvUio6yAih6f6QfAnvBTkUTnW2XzkqXmfai
1JaLmHfEce6HzJcMs0pT27Bq0NNvTl+g8aUWtaRF5D7sfEUs0ZMFbl1Hur3hSYCo
BLECy8P0ncmKBOZFaPWeyvp+EZy1N+F6gZz62scB3BZuDnHH7qB5g5PKKEBi+Mzd
smPicegdl/0DPfqesr5r1SL8QV8+ah7emp1yD8zK8QerkBzNI6feYW2yoQ40GZB3
L5YPeIkg+U7nW+Z0CyW52JxoxBtuK9SL6fYRQ7CCw0r/jByswfqO1g7ME70hBGxN
fXaqh3AK/Iswjp1tyVxvXEWubH1CaOvJnH5ioaYoDHf0eZiwLEbrxE18G1bPErE/
/lYclD9Juws/0MfEiIdTF/Z+RMewjOKQeAfIjkpM8lIAAoUSD87+K1AcQ/1pyCzN
3BxKc2x/3oz2BNs+SwvVDkCz47t7t9Qqexp/daq25gpkW86qhEJEgtkmwpfcSmrr
Rb97YSToBuW7v9UAXwMkWx2ATnR4YMt4CnQFBCD1In200rBVaBVZhKUcgZWfZUyc
XgbF4T4IyDNDajfxU3jjEepWN9mOZsaiKzN6UK3fnWgcMnMv2/tlRpBomFgiK3SR
dmb8hS6l+GJh11Pqg4D4cy+gLUjVTXbHK4X1+3VZTdNnNw4AQKZAbEsEbNGzFu6x
ElSX6CZzDyI9+ub+QOkJmUcC35T+2UOGg2gnIhuhFdBJeNaGDjJjLi+jyS+WmyiS
4eZLnMDR3ZspEm9xHBFEqWzzUC5OB0rE1kIDMBV/0Bmo88IkkfOsqdN9WVUOCZLd
NpJY8m0sPogykz/xuzalreIddF9M2byBRasTIUYuJ3+a17aKSjIp0v1dXBPjy7G2
UbuK/mD5PKa5qlix3JO51t/lPIID55/l6hD/U0scLFVkhuz17Rhna6X3v3yhJXYB
cs+C7me7Ihak12YHrDPyHYWVldwRKWg0tT03XrxcS+E+GCSVK3Tov1+uXEG6Hay4
ckWx+lh0VvrjMFl2187UgHdu5IHH6nGQj/SG8BuJhWF6+0HCN4v97TIk4AuASVfS
8tVNdBn3R7JHPTS5k8JjzBg+TgDto+SPbDJ53zACnGnli8B0qoBOOMTwpZANJtmY
TxzJm4KM841GRyKXFv+iHx7jj2Mijs3vS14aCdvu7E/MwOpetSBJiXQjcHB32t8V
3yubQ1TPXtV2bQoukR3MIwbWJ6JOIkX5rWMkKlUAQA99G2l6tJ4Fsw+abkDl1Vs9
qRtUTQFKfFIGbtQpZVLxFd7k9oyjTrWqLwPxSLyRRLR4d4zP3ZCmhEBBlYfs+sK5
3hKScWS6D+Z5p1QZlmpJ6kRDkAIUoL8iE5FsIqfklRQe1o9bvoZ5GLCb+GpyCWBL
zb8bCHhVqhlAXrkss9AnDUw+vkO/JpTM36KzQ2Ea8cRq9u0TuSmwcsAMGOzHo2G9
sNqCAGi7K3aBNDol2wDMR5dZ8+vogsnDijULK4hdgl7QkLu0EKstk7KTeer/IPVK
Jb6Gyllmkw7/F6e7sIcmdT5RVNk4ybc8TVVPUkxIoCiPvhWrvmCiwJW8YoawHW4p
OPBjo4OVFUsoIeuuAz7qjV0MHh7XcIiVcwGIvgZZQFa4bUEVNZ1ZK5oNEglfF309
NlBGdaoUsDZlV2ymWnn01bMq1eXt2qLPBV+tlqGw7DaRZ3NM9c9wMKWXQM+KLbxw
CN2fI4YsvijQvEmR6aDFMrKm3uQXIc3MiIUFNO6rTplgnKACenNPXQoZD2KYQPDi
mIcDJgGRlC7dsswpuk+T0lP8nrhko3xIf5kxIShNW3DEPvLuf2V1hzDf73LAPteq
iZUxx8l0fbAvTee31lMOvtYwcHKvo9K6v1KQUH+Plpz4fFGtd8ehhKJz4Ty7LvBW
EVlDREJnifrKOXgPR5oUEDua8Id8wldIthZDGEugCX3o3uCt1j1Cf7FdyH1UvKPV
ZrN3PyhkuvZz+Tv8AeW8s1ET3n2mddmAcvb7M8rX13Uf23/6t7nN8kNvFQmMFARX
onYs7i5j9mCkwL5UG7fykjaoF0cDN32NM3IA8FzCYRxHzNwQKmI9UDKv70e2UFDS
PZEMryPcUBcRUKryynUuLkizclxexrSwkCAV+gE2K3mPS/wJbFm8M6RQ+NbBfwLo
hYfEEuJyK7LLZESLaQnQAsfIT+CrACViI+9gKjQ3Umyn/0aRjlhNzqun6jhEvaPF
Z96fJ+izslToHbGHP6kO+JtnHoICWp+oTs/35/VHrHoKZtcjLrzEN41Hltfw+xBR
MwzlogbuKidiX1PFTobhAPfKieFf2PTHxIzVAPnNYjeihCwgszxKy5hHRBFL088E
aX7MIPJwwzQge0LztDz2G03glkGvBErtihnVEccyKfutjFT1AYzENBE0gngKiGbK
jkpY3HMsbUldxFbSvh/ICWkhYe+s6edc6CH/iB6zRG9SLnSEaAtmDS3V/L44QqCB
ZxAAM0QCZ1ZP314wtDn6er/EQ1N6K9V3jyQ+hT0YuNjRbzHYMuYBYzy/GgGDvARg
zNMG6mt2PBP84xKUJfac9DBHAYIuVQMf3oh6UL8som3q6gj96j774QgflFwm9LHb
8HHIXDIVNSkouvVkx9/2hLujeexjFAdJBvlBXm15qZWRvGj3LtVKmskxx18wxtdp
UuQf2wjnqdn4RxMcP+NQMwhgrSwa5cYbevFhcwLVC8IswvJf+bbuUcUZ2/+e9ptE
9RRYn/RdEMWYdOlcAOPfOANeYeDkrjrbbfk3FLZM0qAY0EGrz46qOn1EgRZ/GgUW
7U2WzYjwIMi766HzYhaAaIZJsWYdA5j7JjDPhuz3+naIsjdOjKAJgIehaVV7VMnC
9X5Ab7Ilp9xJqXl7N07Fw+aV3IvT/+Kf8cFeSShTBXIiqiBldqAADLIK47OCIHKq
hVqtYEBMF3/nuAijMKuan+/etdEOr8WRCLhda+Y0qIpiYfwzmw6XUZn8rNerC338
4Jl3AxfR3Kbvq8+HuYUlvRY1/usOuOK+loLBc7RTI9kEUE0eUXnmVMa9C3OK+uRL
/iZPQTa7yvKTeF5vv+upN9zRSVkKdbsFLGtignGj0rE4+8TbNezFUPbD26pKXsO7
GvFeP4HqPEZ3H3A2pigf0uwgftWii1R3FOTN9bhUmyBRGsln3C1qBM9RSU+bhFCU
jFk2M4pK4V8ZOJrICEflIjc2wuHd3r2uhAh5A+EtcH9OdlTGRs1WgZz9FepkDKDG
DlNLx0WQKq+VDG3aauN9x14lObCu92LR1JdjM2ndbEFl5zJtkR3HNhReJb61XHEB
oum2GEglBzoB+yIRKnSheCb7VxQERZB0lPYvRob9QwvdarvPOCplr7yf5ykEZNth
XUBVu7yf2uzLweXTxj9Zn3MW+wlMNpp1yBiplnx9B1lTasnl1MfrLwhrxM0ciKqN
KHTpOHFiGw/iNCf9/p12LTqT83zfsS/xKnSLrQvQVxDjmzHFlR0JwbULMu+HLOq/
QABdR8NK1HTfn7ur0Mgb6hI2pY2xGqqI4Oh1MeUb4bHOVNNFIDkFnf/RPxNmvtGv
vJgpLyA6rQojdNyOknLxVsHs00e0qwuaee2CIs6bqAMHs5uBcr8cQZrZQwc+9ewi
Jzh9mBW7N0SRx7pOSTq4DIr33+etUrY7b4N+fpPkmllm9v+67TKGZpwpmjxZrcXN
BOm1vzDD4OPooqSsXvX0ho2eYrqiVYhP0T7wEVgL4sXttj0IBF5C2UYdpYUW8hE3
Y3h/5oXa7fSsJDV+JiqhKzfND6ADd4zMXjE+Y+h5N84uEKP0wU+l6CztWsWrx/sa
BZlwGV9LH0coCMMRnByRx/05u3fUZR0p+HHxOGQC/kelf0oCR7a5f3oncyG7+zAi
HFVuLjHiHZY+wP739QepIwq0gRiQBJph+HhaktT+K89M2DcKkdvTRDMQAmeTxROh
8QLk/BG997utTZlxCe2kI+1N0fEhywSrG5MDpR0GqJWNfIjob8M6puAuRiVzXPM1
ABqHsZqBwne9GJmpxfqxwMWOC/Fr7aWQyoK/+0+PuJBBggQKmGPL5APmBZGzyL7k
GDOPgcn9W7HPQo9yxKSSFYXX1AfL2Sj7U2v/MQ5i6D/2mY0zoRsKA5omyc4hlTMr
j8jslDDUg/krUVpiAFWTYwqVBqFtENW3znWtWjk9kiyT8f8QKTvTmpmgroSu3nI2
BABFKhsMSG9sB7CqAA8AhC/jxr3eE12tDkd5Qb/ZANP7fb90YLnn7hBfQ6IUNeXP
efz2ArUdIh8YWAqhpWV2IAkp10OA7cAnGszkfBTUYYzOpaoZRlT0EMt5irFV8SCM
5sNYXbBDmD0FOQM2UOOm4+r9rQW8Opq+/ViXYFdoA15oex2Ykcr+IZYdtZ1qi0yq
/uypTffTAYlyL4JQ5PYHk6xI+ngCKMZxxZt5RgwatO88f5l04RLG8/UABeGAvs2D
GXDGazZmcjTMjI8Ct1zDn1PImANUxYagtjeXEyf6rAuwl9O1v45IqRe1sDrDpwkl
0zIW+ostcWmtDR0LPLn89ehLpemq1lrnbhqM/Vn28o89eiBN6gvCd/zZTFfpnjY+
V/p9LfZ0AHlV1Jqz18ChlDUFTQLZl2abC+3jPuapmjnmEv3q5Ttw/4YFDSoNy5yz
qzIUKBj/Vx/PzctWSPupfahqKdG8groZ5+pJB4p2Mzar310Rjtq5TIRwYpVPrOQV
qOdPN5DeamWA/8FVypQQi9kbhlEMbnAk6pET6zNbznbF+tUuGMYpxsqpaG/sGrRm
hKmP6yrjagOqXkwXZtNed8DFSWpWqs99v3MP0WInDO6A2ejNxxtOfp/j1tPVp5ov
ApzxUtQQg7ExEq+iNCkGX/QCJHrSvwLy4hCyRBiDX4V9CSW0nwl8a3vUADRjC0b2
drcucpklLUds8qwsr+XEGApzXYrKk443yKW4EeSwZXmazAnHpiNR/kwAZ9lZCENb
jY0hX8m43BZjVS7YiN22GvxiPw1cdujWC2bdzv1gNOTM/RcCSuVKHYD3j9T6w7mP
eq/JlctwZf0Nao2znM0NGNgvIO7fm1AE50b18DM7ZBTC5Uszr3LFpvJ2ztku508w
LaV7LG5/XBJNasFGJOr+l5HNeW7jFAgpA6Ya5P8efMDKkk7RdW0amIt3b+sk/YUd
JmQEcq/2w95AMcY9kB+lwVMjKh5dQtoVvVU3Vwgh0QDglNSoplyC8fKgHum5rFp5
/6gqC9lEuHyJw1vZ0ZKT1/ogOuId/jZkWoe45HEuwl86RR1LDujBDep/fW57S3ch
jsPqv1piV2I9uSliLytZquwF974qe63j00OxRfzx19y1HktYbEOen1j0A7ogYrMq
U+5FVY1qpSOtjesRcb7vRdur7XVtJhIHoLW8UW/ze20XTarXFDGJLUlqhyGQ0f6h
bT4LsNB3Td1uoWyGY9AB6YdLPXGNB3BflHq2vp7r5cSYZ7T+TSKnPJAj/5JFTCHB
TfYaGbfDsv0Cm2xuSMISao702Kk7fXKGOrHaBEyZvqMjdTNmls3iCRdYN6RMcQjh
HxmF+BbdqBi7nEQNs5nEiQGB6HoUkE61//AjfS6cseTP9Hdfyhbn24Ot7hjey2cb
Y1zXdTF5uSh5fg0JvXI3qyLTqBkG5xagiarhFOiIheh9qW7CRUOSCJEJa19xAadn
2ReC/heeoQlqiCLHwy2RmZS3wFWyNUZuFoUQuWH0iph6qMEDL5DnX351etoiylmz
2+4URIaVI6gXocnBlZHb4BMQSM7SEmK6TUbOWCX3HfhGOkEPbEF2Kv4bZTwBWsRo
sIQ+MOh1bovAlYfKL3BqCbGy8TWtZtTnw/bpPYj/NVL5ZNI9aK0jKQnPJ5Gp62rO
aA35j+04KLIuyDDJ8GYLDYvF6cCM0G7r7Jv+8j+uEQrJ9vABoYzCqIaLbHdMB/Tx
sIuPKCp57davCCH+2Yqo7fvW9EC5hh2gGZnAchVI24qUMF+xtjGYJSvfc9Vx6PEt
6o4jzka8Vit8crSO80OIstYsih0yo2Vlce96He3L3U8ta4xMZQPGOOjga8ZNLv9b
c+RLUpZoOY7bMwhPFetj6WeeolI4ViccrY3WoIiZwXgOii723/UwB+zvYXvnoCD3
My42khmUK3J5dT8uUuKkYOKQuGUm56l8Hv5DuhHgi4kSKgC0TfHtiLUucwi6L18x
QWoSXJ96Xeifv+2DxrXRttFaD0nqxXzBt0PQvUE1ZLgexmzkPvXC14r98uqPvNrO
WvYQfFN6Fg46GbbnD3AoXoFX+uCw9ZSBsMd9gXUq8PPrlLcsFfIdriPVCq//sbf1
5b+/7RzrNs0zmLuf196L5/+hBnJxcc4DgCk1O4WjvZ8cISR04ApzMlySXw5g4bML
pK+h8xXGHuBMrH5zdzJBKQMg2r9JyYFdALDWK8TXc0cM7wgKF/onmCSgh6ImW2qU
fhudMzXHrN+Nl7Z2BN5oEHsVG5LnjCVeFLgjliSnzlG0/T480HvLqiiDHW1f8EBg
Dq0+lsXl+y5ytcWxUFahgE6tiagaBrd+t7GDxgLrZ/ekeHyMwAgV4eYz3JdNmfQj
hrQvjgioQQF1U+hKDbbh5whQmeYttVuUj63XQsmZJOBNFGkSzJ6Ep6qN51IUjZGM
l/Z/WbkHFhNpbmvRXyToGYJ09ZwLZ3Nl1yqF3jcabcRfZTtTSheWdKzkzQFaonKU
4jc6pZwLmjOJZvZ/30p6uHzbiB0yuZBwDBJ8XL0i/X23CgtrJ0A7dPQbj8s2zRlH
sHHLCRfs7NQB/sLSS3XiXgGeL1CeIpmI+NbdpDcEsIls/aAxo0k9U+CFAeiJuH4l
DBto8EO6cBbefj4b4szeE6al694JiN8kqMgbWW9OsCI7F1CfHCEjmKTaUczaCBEm
dXJwKqcusvC+HDpt6494U4Xfoy/evJpWOwUfU6tKOVPjos3L/mja2/f5FsxXSSkI
h0pU2qHDfMme6bH9zLFmb+qiPrisp39/OuwdvXQLZdUbJz5iuvCPUozyrrKnL25F
nMBhRZfobBnFGw+QbCfLTxN3gu2sd+uTT0cl77mu1V/GLREm9KW6FJ15K2tmVpdi
8N5BQpnYVZB3m8ZpHHa6YD1r3qGyNROJDXniMpN+taLLYdPaQwjd6tFJeB4xkKeO
saoINNzUeNz7e/2ez1PTPkBYejMoPnBb1E66dQS7QbaxAv8yNM3A5CuGOQpbe7ff
ygwWsOXA+oU+pDbhYSf++eCXyTKnOhCzEsy2a+gJdqJPNatdDW/wxjjl/Ruy/Wum
LyjV47m3dVxaGPmL41IpLEv5PYafVzTyyafGGbtBj738mdXIUvxsCLNwtDPCuV08
DuvrgRhspgZFRCWAcDwyUuvfICeps85fP7Ue+6Bc9lA44jBAwwlvtps1NJoTlAcC
bbPeLXD2MC/pMnypkwbD9L0erdp070NvBVarYqP9NpVIejmYodA6p5g+pieEDBos
FJpaS6cS2YR88CXLcdXGEPZg/62G1FkiKYGunu3khPiBFI8mnFADvefcpdNT4SfL
vtlSpFmknxdfvYjZ+jT0WsiwH3J5ueTdSfVAZrT94bddPLJJqUxh8lk+4yq5GuAW
lh8OYTWPfWvCtDzo44LrEMc0YOCOXMsmb+isNYVZFIATtwcUUb2nOinKCdp+Pght
L93cbRyHYXnEzJqDdAEWEaMa2P01ipn3kHktxff5d0uPULwC5Tbwnx+JUQ82ugNQ
QvUDx3mSVT3cX6YsnCaZhdnHHofVFyQPqhWR2jxyA/Y0qfWIwdWlUW5Ng/zWF9b0
hKAA87EMWayZZOWasDrqs+8HGyR3NSR98gSLurp8//9y2TkvvoAoAKxE2H800PTg
jhwW9lnF6J2/NOAwPaIsx7WFp7NqFwzrZJ97f3j4F44XbSvOB77s0aHFrcM2utii
L8ejEaarjmWOh0teEvMlswpbuUUAJ+YAv+D+8jr2gSxQeIprNIJl2p8RElOu7BGI
GiiUEL1179YsYNSVJtuaH9/aZ6vY4CoCITcFw5xJwtIiuRcFYIQS1K/OadRKAa30
3RblGADatZSZoMivES60LIvT5f9c+Zl45W3k5kMxOY6sf0QDkaQIK8fAVR4W+E4V
ByQseJ7e3O85dGPfZRblDf/GaYNLIOdjerszDKtPUFUHpfG4bn1Ws9Nz4JfLm150
B8nNR/5hXn4ilNCiMb9YCBnAywBXwIVc9hw3rSYRRhriTsg8o+lYTtfN1tV3gUes
xhMi0spfULFc9Hnnd+IU+Uo97fbaQeR7FZMnDcZkXoY+syQ/lR5y0ABpEbnBHnIq
/Fzd02btr68A+ZgKoRe304bPRCycZPItS3UVfbfNtFbVwx1T/pQhiAJxaN+2+CQu
t4xEoFdJ4xjZakItCXyCGtrZRdy/wvsb0iFwWY5/BW4aG6VipfXtrjvjcRI55dzU
Apr0cYxEX9u3hoXpQt2yvmc77GQq0BjnWiMnoDVIy02BHnNN73Iqoowg5oZi3AfR
eBEsiYvfVhOiL2zYby4RUMBzwxTJOR4+1KR6oek8imolxdOI3aFZozbDRIOuiAqO
VOTUH/Ux3usr51f/DthCFvq+wzO59nD4oAW5YvZ/okzaf93oMC2bVlJ/SxKLSS5+
Se7MoeLETMlgVv2HWyJHBSPuhYhgZT1EB5FAdT3cBlezMbuMLR6i+idqHtqC779p
Tu1x6TbB/SSLUA0vqnpdPmETe2bc5BCr/xo288x3p1U/Cgv1Qabx90rRdHykJCes
jOw7YZErBxA7CwnKLN+WhRGot/G3Ff0GFuQdzv4vC+UrfEn4BbAxNddyGTLxua/v
pLTStrNP9hS1QOhQwnfNP4DOJCJBk1bqhF+e5v7Bk4ZnXrT5ky5OS9FffbCK730+
IbCqWjOoQDcJbDzv2nH21Pb99i3z084tvHSwH1JVktQHPnxxxQpRBSCUSeqoKMgz
WXueKDtnaZ5r9dtseUkzDWo+/Gr8yaBV5cpDHi300KIkKge3vIr9WzJ5mlBbDz0D
fdguCb78CNLjJKG+jI3qY8pujj9Ssujyqx8A/wYY4K9w4F9zL/x5NRhsinBfGe2k
DVGc7MJUKZELS/wp4OYpphYlyBCRdP6b+nEnwYT97nGDe9jmN1R9Xa4EuIaJ5P1f
s4I8GOM2ilXCg7YGtDS0A0oHRq6wSowrZPi8eOJf6Yy9YD/rA5LeThLH+o2VZQaU
01SmL0epKvXHuUIy2n0AJkk0VT0DzPiujVTkzLd83RQqKG5AGnf9WisPX7a1hO/l
TSaPNo1KcFl+WTKHfymdb22qJxqo2mGMAXvX1OtB+04eUmbHsVQ7mObIDZx3TTcf
+3GPxkvpGnaIAvwFPUyvgUu1aF5zi+ulLGEfEDsenVyWAebaO3W6MnUbL3Nq9hWR
KaJgiCsISmAT28ekK7QQ/ysvYPTpyloN7KtNQIsbJCwAuiI4uISvIp5iUPdwS6zd
5yj8+WzRtXLUviDgaaBXVJ/89U2lvXHHBT5sV6WTiE/luY/IgiNXjS4ptg+bhV7k
U1ukyg1z6/Otcmk5rNsl6WhzFgLBabLLN5pW/ysUvK1jwiwOyP3ZBAtc9iVUwVBC
XU9MnZj7dMEqWmGyuy8EOp7WifiNit9Jpy+J5uBFexkaOty8jpDm3vZqKU9phSBn
8ms56eQ6BHtCiKvCTLlGCx4YzGRC7RvxsDSm9t366DYwzDRIgYYxQuLjNTueJHNX
TdMUdB2IwMk4Zy5aQTYy3V/BgiofF70JmzaG5ffC/3A2P7VAJbl8kaXg93IPiRrT
skjX5GS7nILxpnNFDhfGdNMdi25dcYFOv+N4Pd6omRLpKIezncobqsKkO5DAgx5t
C8Icaer5wwrj9E1NkQx3/sWLzKuo6HnxOzYu7PErkuYYSklqx40hyyWGQtONjAuN
/j8txt6E7knKxKx/GYZo5q1lFzuqJZpjn+G4BbY7AuPBun7HmAMQvetJUM4UAyd3
0/mg0a/jf5r9w4PoE/FklcBb0XpvpLBZbRNYWgBnOjTKA18SgXderzWkYa0AY1fe
oOQuJMLwU8pEpBAD83djr3EYon6pNKT4CxguVszynzlC4TWRylN9XX5c2qnAzDGC
l0xJLJakEhclLiB97iaYu7uTBGr0WQer/pIHkbMTdG15ky6qZ0qmKwiUL9f/3/Dn
zGLR7wYmoCJIZSUs4REATq8rQy+g9BlhWdWXlyU4tt99W+1kNxpDNcm9tcBwZWKU
UZmxKIUS7kC0C76hDGP8tRBB2Y8FshIXVrCND2y5jEXuSCSR4VTZhQMO1lgrpErs
S2yZZ8p72eXC8o8mgT2ctisjlKToiW9VJ8nR84XwVT1VynRZ8FVgbHsMJnJjO3u8
Hx2TyG7baQGP1UR7COjhPblmsYF5CjJljOg1ziJWCP3/bngs0XDxNkMLsNcfina6
h3qjGNazZCbjXLcjN2TIcFcSvPLWHQ1voMt/DmwPora3xHC3UNAGncDu2+XS0+XV
uJgXptYmR1sKJDE6yOUINl3xtUfhqYi+OZK891VuR1jnd0jlOCG8bTkVqMekH9im
kV39p7aD4IbmeoKOSXz8STNNBpf1/kY+WSLOEm9ZiqOW/ad6cIWB8cCdCwsozs7P
8wjg07PVnOKjJK7zrSXLI3RiGkh+y6gzqg028WLfdM2e/D5G0kYWXZ1xwLsooThH
vfQKyrl6LcSAHkTAfgbbpLJoEmvudqO1YK0hUqezkXJm284Oht++K6AQKaRUmwXf
oCKpkv7MqR2DAs2FC/t7KlDDLjlHKPObRPMnZfNErS/Kb9aHeOAoNc/WlTZK2C68
zbY5SIVxtyBArF7Dg+Httg0ypxvb0zwr6a+DXiCanrnOm6qEzhzFMSulTw6ycV0W
O9LehZ+HxmkyMv90aGUtZW5/33MjpRw8kyLdfajFvxDjOcNVTYg6TjNr5YIve/lF
tYTYNsDj66+iawN2BMP9wp3En2gw886qJJ0W4Q03k/g0nOk7rg4aCxAkziFGVV59
Vc1fJlfuwoBURA4S7PCGtpi7cYLsRjfkFYwg1FYQc8SZJiOyo+8huAYMjTQG1b6i
AEKwUcDVxEm5dLl94gITAF0UVaXk5bmOJWYjmNULw7Yq0f59JQMhTllqXzYuER+K
Pso1RQbpOCVwW5BYeZOtc+piG3G/xxRggoas1jjuO2KWAqjmGkwoJee4psAch4Xs
sDXT5bQbnZHt+TV2Y82NbTslrZCxiykUkxgj30zqZvpR3ZXkzEd5jJy19Qf3GoAf
qOESpbwACn8ndved9aEtoQ1jGMi7VAENf6ixhpZFOIE1dlHQD4sBn3N66cW/C5WB
n3xKLXaZnn7RoBpTjjpUJrofvGIQoyvE6gMKBdWzdoPOHTWvqYf2chs1/JY2t5Ph
d9HdaMrkg04ISpLXu+Nt96DjQ1sKlamMpQDDlA6wZvfCLcPpzF810anelH6A/31r
M/dPG7E3h70AQKwEOuKNk9tTmSGxEGzAzJyAFZbip8zJ+pLIb7mseoOZxYy7O4fQ
p/ODF8mja7Dk2H2gkUz7EwVhYgS2n3Z7vrdlnoMyNqIZNWzVWa5TtSm3tClNSawm
Tq1i7YU5Vqf+SEMVu61nOeK9Jln2aSQagHftvnwpgEh7NX7GdrvcsPlnffRxC3Pj
t1SdYHj1ikFlAmfoIbwsVCHJZnQSnFMSzx5UlZOTDBQc1oRj/T3b8DbHRHbD9GI4
oUb7cImL2/WyaY1l34BjtIgLRVKou0xh1LmAW5yXpao5pxVOmGla9XC2y0sPV2U+
N8DWruM26qvUOO2BvwFni3Mj0pK8G3fRz9WQAGtr4w1MtSMALEBXDd47H0/hCv6S
5SSXZ0izfAmkVSBi1teHvv+/m2T6rWAc/1OGOMMNyRBI9+lGConKNGEscMZmPfbQ
3RRi0HPijUpqrC77TkQoepykUuqsbRcxlvU+BINqyNRs927+jHVq/YMFZQmA7AOh
Y5oIUDstABBrEptVQOQ+3Ko29XerYAzb/TlOf1KTvIlxakzhXc2HIDYlWIpgjtIv
ecJRvCn992vQuk9ROMYR4uzdEfCU1b626EG2sAJQ/C0qaEmAXfHZ1AUSaTV8aKMV
dLA2RSSK432C4S438PhHtMzj5n5aVlfj//l9QY64DHUdafgwEP/c4gEG2zOse5iK
GO0W6MXRlf7q7LhnIaHtbAK+qBY9z82nW1opz2XBUikExiyS03QusjmHN66BMOOx
O7OYpnW3sOoAIUl0r/0CGDCUD2YN+pAIIg3RJaF+ZjEDc+gWlGb5rCBw+42IFsci
BUFuUZupTPeSpaGLLucFIk0PLbHL1mvDNbnY3NE8I4dDB5kRgCuvx7JixUDdDyTH
CRF/4fNswAg5GSzBvRVjDlUjwqUINY0YLeryGh9T/m0yY7U5mLt9WTlhjMSPhQN/
6VCenxPErJwksPedEp15jOzsm7uzzjpct+bTCTP2IRTC3NqISixWy2U2McwrsJ0K
FBme65Ef64MGyxvghO1AG5D6cRNv4qVkjJtHGH+cTmURWL+STz+L/YAGgvpmJy9Y
4n2YCJijZkrMgxH4bgyCcyMy1DyyFOSBA+3r+UaNnZKVyulLIqaQwdCs7wjmocLe
W1wDRG13IBAmMjk4lfyCmijfTaeTFvtrUEOBbwe2mTQ7h8aEgbrqwRJaq25RKfld
PYlGSOHmSiO5wu6om6OF8YPL2gyB73i5ZUFVpwFpcq//885OuBTPtSUd09zupf2G
xULpWaPdtsfPWltZYRvJR2MfMMggQygkgK5Vos0R9NjZ1edgWOKeBGOhX1dyf8B1
n9bK5L7XvG8n3ogebUqAtZLV1yq/nIjJdd7JnOCqHN/N4bKJ/Vra32ZHKwCS6ebF
+FtX89DjPXH8iySzkUUq/U20g4tSl3lXG8/TcwFehxAzva+1DmMRRICWjL0bYi5b
1FF9XfeU5B80fRpWEzCmmQDyAa69eo8kUaUK3wcVt/ZKYYXrzfNMhonAgBXT3Ur1
8FObEMCNDLoxETsp/HUV1qLIe5wi2mQt8Xp2+vaVVNb49XbIWKsMowaYXSC1CV+W
FZ1saDRqlHllmiMtYJ+hObLTyC5bmup/KDRISAYJkj6HijGpAVF+9/7UTL1NOJre
6cv/3hwp6SZMQMHxOwCBO4Wk4Tf0E+eRDs4Z+gxSsIo8frgCyjAFNtC3qDDxWCHH
3HIx1FcO/ZLpi8HHWiEYoTwrgkDXSJED2octY24bs80QeZIddCS13XYarkXuZt7Q
PlRiY3FaCPh6JJ+wj6dATvjEA5MQ2EDOdWEbuTCTP1XKnna2QaqineWqVPqgN93D
PTgOPkTzRrAGPzJPqQ44FkY25GxqoKceTVOnu78rJhZ0C112F4gcuaeGZoyw0oxb
M30GR1x8AwijhvyQ/+6eUEMP0oC/y8pVkohv5O2hKn7C8QFCHk7WNIZnOxTG6LxO
9KqWBNlGoKrmiRBl9L9L3b0VADhd5hsHF6LmjZ6owzuSRP9uZyv36CDrPZz2vnwY
odD9c2JlA9Cq0ZLhmdH2CWJ3l1hV4T4dwVStpZPzSh6okhHZaW7HUVJ2XYnzKH12
DjSpdxfeyesNejE0ecaj3RW7Xc8JGiwgN+6U4KoM2CY1msJv9qjMUIigkMm+WpYx
IapXj4IinJq49dB81rfCzjRR4IQvBnUzXRvn5JUBDSjx1Cc4UIK+3r6pbkpwc8/l
0eLQDaoEZTfvzUO1uKeBxoeZgkE9HAf5RIWyjWxm2hjj6EJ/uoWaRasmiwVoXs7C
LdYtL4B/7XOKLGuaDZ/juYC/BnVfTNC3ZSdCWhgCdOQ/YUIytyZNz8BEGcwCDzot
T/s7sgGbvlxd3UJJY7QdWZomo9wryAfkttecyGLu0YbfyDNfoFIupqZH4vpXVrAY
JNP3g2EdKQedlzzp1dcq1gX1tBcpDfcfYwr+oUPQPvFj1S7TMkSt4yQlvq9QCVRM
HUJTaHYKwMf4xt7frHV85v3IAf1scDaA4PmgjbZp1TjlNSfrVYlInbDWw6FiBtYl
n2H7OM9w4COrXe2cWCG1sbSOE++jqZv+cBdgmy6vXG8J/zP4xazhktNRwcRwcMFL
IeCYmr4t7g7uObfM0YBIiV8mGHAfABY92pxj54B9vnMlBMlMeUF/zFzKg6qEMR9B
xghfemj25rduTwtWU3cQltM5JajpN7LwYzoicESn68RzgSrRffOjEwXNUle/xrY2
ZiKVh43b9H8cpBwvkUH+IbCBSAHtphPqPxntjBArA0Qou9g4Yc8Kx6XGn8gdo6U7
BbeH+jiOq830G7aVvdyLDU57UAiXxKfY0BHjMa4pEwcv2iOytRuHILmWgM2888bS
PWiNu4SDsY5K6NEkJsef1+Kan/gNYRiYuYMEBvthTvobsSqcEMWwvguRfrN1KDVC
RbKkrNoj0u8RYXLd4Px49jZ9CnYcnCcTJfhlLirIbACLj10bs9NK566HBVmQTkkh
hQjOkVxf1EIlqZOaP2TlE32epPpwHWQEtByTBHmBvz9mPkvzE1F+9xwjScVCNJyL
EQxVhpFAeeUuRVDYupWsgoAEH9KZ2hfGCqZOm4wFWpjPImeBIq0ES3G7DIxkgEUt
89ziy8aa5PwX/EOm2EOcP+J+h5eGy19iQbpeHr0ePJQb0CfMwr3jeivBlc6nq9Am
hnpCYHz81IkykoCSZMLosxavu5aofbYA/SzTV7rMrSUzlHAZAd+zqngObhZMcSQy
X4EgM1zHHlKyxTCEYN69dSzcvyvLI/5G6tacM+3OtDplhIApxlgETmeUocxLPvxF
5tdtMcXwOEqxPMFL7sqNbrfahDb5vOl/4h+2hAnJY0a6P/vNahw26ciocZpA+8jx
mqo/WcGd2BarUWZmjRaIkebL1t894FT7q1+/87pN1yUAN5JQ1UOl/iEG0kUWlLck
Ydp9dMQG2hJhW+HtTQRTJQBCPs0Z6DRYU1OFoZqfuzQEMbNrod/xEwIMl0ZG/+I7
VWw6PTWo2WJ3oDuXk4Tk2BGHoADBOL9uoJxNmWYarryQjfu0rbYah3kuSv24bbPP
M7v8nA7px+XJQ0oEg1udzKZTZAuxOMV1iWdG2UczAa7TZ+nyjWsERP9O5m40+WNv
0c5Xa7kViiFd32LGHwIymaqj2PoEWUeiH9DVPa3SOApWYvhHv/TnkHJa/tgMVKWn
UgqNHN64ivtCikHvCurFcm0S33tWaT7KzvAWuvwQTsW3pQ70ArzgJ98EvZFBCkRs
k6yqtN1NMIkzx+lXHafIuLAnxHD/q6qoN4nKwDCW8ssg7vgL19X3IFQf/CvXERQ3
SyhKuG4LlTNIAckYopSW5Hscy1UNOHiLdVfDnI+GgC6LP4N0s5hNLdQgQWNTk6GS
iF6iCxsV/w2G4fjYKpLluwBlFlaiQxv+gOmJy7UO16dJJzXrDzvnC/8ka3XE5S8N
wZ8+350U01vInr0uZGgnbZ/uaqMkRRy2Vib4IKUiqiFjJAUgEDSvffpA/0nH/Xxt
wBWS3Dv8ESDvgG0dcSawgDd6vMduVX1NKNQwiFOYlxWrEVL5ZGpj4IND0AOEwgXr
M+4XIOewcjRMHjdGkGpuAwoFwxxoFrUITqGm6nQeg/dnmLIHnM59UQI5oKdiHPG7
aRXTfVFKuSZkW0gOHCBWAxXBzhe9iHXpcpAWRhjhBP8IlB6LM/czoPOfsB5NUKek
rEwLyjZeSWT+xG9lEzgoN3BjYKHM0+3k59OxXMie3747h7jQhnOaLRblRH7OoGvN
jiWu9IUa3/4qhD28CL5rSgpxIC5ZtWENFZ7oLjXPS8UWX2Ek1p0NQcyXPkiQWSOP
TtPHCSWkCQIGK/2FqVPVOM+03nPyYmdVccPfMpS8RKEMXE5vDn2Hcx0brlynGqy4
F4lC3sxdOL38STp/ciSBfXIkGbm78jMmqqBw/3Vqz5ELZvkK1UTxARunDPNCb7or
yNYKR45MdpKe/hOfgRpAgfb12cjSsOiesraVi1MNLUDsip322ctqdNZTje+sBuZZ
laNkPLkgaxTEeAD4J6ycR1WAczmroGIW7H4nmre2V3qVz14Lb/XbDIpn5pZkLHPg
38OfXpjZNYSwitZzoYtvF6BGwOM+QtkSuDvBHZ3AmFR+I3SuKNKEmZozTxmUVdTP
2fIcG2GYOm9n/Gnr1RRAfZ5ifMvhZqNTG6b0ujc0nu3lXkYp8oLTw7BUt0jrFGwg
+gCRsGo4xFbhpR/HrL0QQGjwxobhopJe7oncGvnFfJUrNMszy6raOzGY5OOFkUA6
WEjSDePsG23FYRH9HmEKthn1JR7tJ3uPDfOSX1suGAlt679p0WRB84pH7v4AV+bd
Z9AhjjoaIquvJVKMTknGlK1FCWq8Pj7eFxbbq9rxIA6OqAn+X2vXTCToraZ4bTgy
LrvYCwt+Z2VA2pBv9uPhavagd/REnV8Lxl5zBSt7G3nzwcIdgnDs002rI5wcjbCd
N6DEMSV/uHPpdNFLtZllpHM2oEvZ/y3GTuYVA4HOrzpGumUIkI156LdjsW+aTjC4
d+G9/TEMiGdiWs1miSch6shmWrVYG1r/6QOb786F9liPy6QpOFiI0aBfRma79TvZ
JxfI5rHvQzaXQq0N7aE+2lH4TKRUTsqkxfGx4A0vDyRb0jwd8YepA29Q39I8K0+y
XxBKGZ5tiAQBlSKli83dfI3gKo4wEV92JXqo8iWRbkLIRjYk5OaScDYTWpqRJcOQ
DR5lyJT8jNIGcvOm8nvP6+5GHz01E1+Q4/GkbQwAL4WWIeJxCZH+3M+LjkTMj0Ca
y+ke8TwTS/MBktR5coSuHCcF0HXe/qlKFfB6+rogvQzsUjus8cONHhzkDy3qKeCx
5enOLSDfifLFA8P3zwMKae4kZHWalJ5mz7vQj9txH8Kb3bAJ3Cm+3lxJdtnFbBYW
qoM6PdSIbFDcFGdP3Cl41nEY/LO+DaNrFLfzBWfYTJLbolRbs1ltfTOh3SPS5oTo
PminptVEfKu1A9SrVUbmKOHtydCOKG+cK99J17qvpIuqqDZ41eMiMyc9DHLIJtIO
naZvuOsPGO3tpFL6KvDMsW0xzpCZmQ4cU4EISIdyhf18cfQQWeb2qGVXlFbIZlao
QnETDtPEplubEqgKfmy0l06kvld3SpNp7h4MMkbgTFvXWsFWEJJ9x2yQxuml02yw
++jfVUpSFOUFAn0BNOTeeiXV5tWdTFMkP3kxXERKG2sGESQ1LY9zEAUpTgRmkL6H
qvdEmnpqoNWJftAIGpc+kEaNjbrq6z/TcyAQCwJDM+YMvCuwFjChBsr4zw9Mwj7V
tclo9GHuav9W48/BVH2dXpDkcAgMgOg106HxF2FSPdlBmt8TAnMcksZsLV6E4Xwi
iDqRP+1qqjkD+2jcisGHxlasq6wRA11+c/0W6uKgErhktNnGQI6bAqrTyXRwr0/F
nJvby8tdx5RviDAysYEg43D90xauImn/PiTdUyQ9qgoaEbIHazf81vf+k3pKbm6L
VMhgciQrIozEFNbM9ykP2X0cgM8Q83FVtzggHKoME4kSJxWwP9q9OmZAAy7cS2gQ
H0j86swhOa30nr07I64WsbrVTbnPyIrcNXT/kCABdzExH99ZxQuUo1cFrCaIobL7
hUh1wJxrH7XktC51PBPz2J6ycvuhpVARMXmokOu6xeD1CrQwIW0Xhnf2Ev7c65gT
dkRWCzvo+DxGh6uDMeh4topQhnLEWxjrLdjUJPZfjfJMhkQijQr+MxG/wrmhkHLA
wuBgaSOUi3ctE8mF6QHUkuLpVnhlYoE/Hs8XeWxhb4EQzUf2ed+7xpHl565Fs0xc
g+L9MyNsEna5c+k0AfZ0KD3fjfh+nCRhpSomCYmw/kNRujOTmgaDUDyzlmfbgYOW
6kPHrtyi65H/N7fWJlHhh5LQqqNOfQC52GujzjuXAzPsAdljX3eej7qUHzgbKVTl
lygzwqOP+M5Hlp6W6pBHT8WuG42/Ey3FztWlKLvNKYN6cWNV9OLx2xeEi19+towg
wBl+kSMKuKk3LMs1jaE4kANqMgLQv3v/Ieb19V2YoB55t/cFU6n5WfEmMA4emsog
TZB+54QPk2SemLWNVVIvrgebwFsvHhkzSMIga+Ag5e0Wbvb+xjb8C35MunlsQldt
z7lGLrIakgQoGeH+90cDJmLtVBedyq+tvnkPKDTA7lvkCXQ8izqtc1P+F/VLfjh9
LuyyJWmXfvlsDAAw8zBz0dLSYbhzCZGnsdl246QINjlPzTJ+b9hH3YyS6ufUdaBI
teARKJQXU4MH4Mwo6BJSLDMPwZ2vdhOtHKAo7R+5y6aqcYhaDQeE+Y5Vl5HwY9t3
lFi42kocPIIfXl2sF9YO/ksAU2vqMyUcqFhdRckO2V8/Yehgb3n64mEmTQutCMf5
6AlahXFSNB0sjjprsGxrCngeYEb8XEZLZyVhkarpcXlKQLDdGhvQ1KH70Ua40YMc
ByC5mXkMzKh83wCKwEtxUFI6oiTKOdipqpW4gX0J3NJgQkaGsoP0gq4Iz2BJhIaI
fB2L/MEyMo0x6/RQ8vzTZCG8fDIOcjfG+j99rGZtRjW7w2JkQhp+cQs/KROt1DKz
K/ueUoEuffct4GRoOpTSg+B+uGpbVDtTMre9X9AD+Jo1LXSwWur79PPAlJnIdXt6
oGjiu6+EibdWgHCJ5G+bK9YNs9CxsgDW4aVqVvtO5NV0P1uxIqpZtGkeD+szC4/g
MmlMUTc7FTzPd2KnR8/ec/df9eib7fBQ70w0uhzK/REA7Dut/wMKlr3xpiQvwiF0
yWgoBhs9q7fKjh7iMp0a6WYa4Zv74iemg/1pJMiIRYn5Ism/cmAxsfOCDeMIqQ6T
vWWK7BlVawFy6YbyyiQnmnpTWLPrsGv4Z0ysimD4IlbFsxGVuEk+n1NbGuar9Ms8
18/yNhkqN6TpGBZgCSozoWgqsoVKwKgzJf1ULmMgi0KAzxyOEl9FuILlAadTdMgF
b2e2pDTX8RiErvzjw5kJzJmC1mqTrR7rQoQrQPJQpJ6OGCAxhnitytbD7+9CnMCg
2HoyH74/UoUQN4dMGnJML7l5yVIHXU2/AkP37AHRTFjU+RPTCUvfkFVRHo8LX/bz
9JvJrHMX88ssuj8qcrSkjoiBEij8GS+VtyiyvG5yNuOM0pnFgku/ZjpMoZqSupQj
B/8elarAVG0RPGDvctPMMFI7os1HLrjnJwGfcNQ/XO1fY77SDxNhG+ufq1ASBSJz
aTEmRa5dISbmcjExIbotIu/X05r7TZs5UuKYhy86XRgQ81/EpLaJCYzpGbQG659t
RVmSy7OI+Qf4WCRCXOeGN1UAOBAnzJKMOuTLgW1YLGKWHNjAuN9xzw6e2pzv/m8Q
FGqvEvkWZsHlu8LTKQP63s3bMlaeotSXokR2x89KUG9nqvrvzR9unBEOM2SGjhOw
iPoCN8PL1A2Bas8cMII4Payqnrr9f04AjkHEjl6tQb7x6yxrHlwPtgw1qp30FEeb
11Bi3E9yBb8n6Z4JtjcJb3HekMmjQncWsjwbgQdgvj2F9b9ho2QFeGPSgRG8S7RR
BmoWkpdSXE6eO8Fpi2UcGLcs+80c/fz5z+N46jE9kVSETyiKFqnZCoZgVjafI3aG
kpoBFhUE5oeQOtrqyspLozuyzt9nRa/+ThKzNsgDMYkkeenFJVUhA7eiODLlL32q
TKZkqXt70KHjhN0mFeHgYDeVteTBLHgjKOQe4WJkogTipQkxRmrICr8vxiOoC/fO
aMGG8GJ7H6uqeTdGHIxLDV6YB5lMAXakHtRdBQLess5haSpzkDOs4EDKtAw9O1FQ
V/QPGVlXgbqXOoqJaoFYUVZojmKSz+e4XedlfDAv+/du5eijRxVQwQ3/v9HDwW60
4VfnLpfcH0kBwQ80D/EQk+CWj/v6aNj8p6ykbc8fJ/ioWH2lId77ntt/wKy5pkJP
S1bjyATi6IDyyjenqYQIT8tL3NHSDSz4Nfx7Pn4RQh/GTUS8mb4xYeG90zNVzScK
xgi2aNJQ/sMO79dwuRrp37R6ih5htuaB7i/4acjVjblCDn1J+USdBwAQUm7nxv0D
lm769raOYw9JKGEKXpvOwfJnikBeKHEX/tUvksfLNrpIaxQWZR9C4koFkDyXib8Z
Wzyc2/U+yQCNsi5KJlnuhV9eL8kvoTeZYnG3t1DDxJlBraUoOXcMEZoVM7XBdr9z
h47XKAph2I3sOSK89zPkolqNHiuiL/ObBdvfobZmEkI8hXCduwqHtYdR71R8GRdB
nPQKluIGAVLhOX22K9RxGiu4HPGNlFxP+1kMV0tdWNLMvE2FQvtFGpwr8A1QQZMW
x+MoS5h22cNALIyTUM0XrCONstJb9/6IxteuVrxdoB0pAtURbKCGGHjdf6Wokob8
JaytYBhjiFk1c0Mvml8bS5D56+0PNVHrmvwcaXkIagghVRVPLpQGq+X+muZgorMV
/m2Y+fvu03eUkf+5+qYgWN8w2u1Q3P4dptmHuAAnCFTIZDCNflx5SrWy14gg3oGq
yU0XoHQMOFMQljS2sLL0TFtfp+yZxx4DStv40wBydI6Xul3LqsKIc8MRsEabTwM0
gHWtEiPNpfZp43uc3gTyNJHLUhEWuvIocmtl7RUDES6I5GBtS7hw4EaHyKjq/X8o
uimT9FI3877Zs5dDzSQV4YRtbuwfTibtOeeDZkK1PHb3Db9eOb4QKKF8rrjJQAbi
Yi1IjAaZanKM9NQAiKALhPJOqa+y8RZfma6WmxkYRP3EYxc3vgs87JELY3zkTfuH
VzX1cFB8jD4OkXkAG9RxSdw3Icb8xD8hsORwEMUZU/P3J5ov29tJEeG+yGGwnq7y
tOwzFm6kQ5FQmUR+AtcjF39w60/yuAR16eHXRAwbqKrJ8TF7laInxI74Ea+me/q+
cnFaEGruSQrKidMtwMGGy0wZOFOpw8DY2X1kx8kUXzGEGR1vUrJzqjxgJBpZZf40
ZPOwjZWLuWbK1m4MpX4+1cnF0jMEQFZA+y5icNrhVKhPFiF6Y+qL21jjeD+S6unm
TEFvvxpFqq1uiKXMY9m8H3cQ+62eWuc24eWfRVzggLVOjFIa9MPydV6ZLNePo4cP
Qql66BmPS3+NwF0wnntDZraJuGBR+UcSEGRHvO39Uk/oyWKakNuvatg5osllfj8l
1rZZP4mqX2dFU9cX2W0LZV+6Ew4YV6zb4LQ2MAtF9+sFUiJGQjpcRbZXvTjSWzxt
8CHWjWq3LmwGQnWuvgKFlFx+rjU4WGcxVQHk/IiCAtt+HVSyxYrOO/i5fB/7CTZl
VAjO+w84eOVPAZOsgZF+ThKHF53t35D0qG2CVxEbsckcn+nPmc0j/XTWg1eAF/jm
XR9WjX0TJkge/g8mKch6jmoHaCQrbYUD8PznD2Yj73DeH7kq6vl3JFu5lwndAF61
AGOdfFv1TwkmOARQhMx/aM9ok2/PzsFHC4hzqn7znCsIwl9yJl0n8U/Q44DPE8HJ
hLginw6WcpdPwVYg+h4HwL5ctsFeUaNRJRYdjkBcBZVeN1gyX3B/yQ3+GX+zGQ6V
hxaNU0pDb3T4j/WQpXgv4RlmBY3IrITWHU8dRozIP3Ny/mf1Re86Wka4VyiFh6UV
8PSPAWsoSAezYJEYOBuaMBxa5LZVHSs4o1yTOuLeDPvar8lkrjxq8I/Lt1z5+JXE
vmyJbZ8wPXTIItGPD1UqPR1/brChvUZSnHEBeea4xoB3dDiFTuWfsWmOSBSXKMPG
99wuJmQgByul5NMmeHSzBSeNEsrX+yu40Y0n8NQOjTE5QH4Bvc7jsZO9i3oaYd39
JFH9cqtf7duP3WIgJid1F3i9u9V644AjulXJxYmEtQP0iBl7ddgS6BWNUnbVOU51
STrSbOVBGKaD5Zd++HJvu6NezrRE8lSL022WZr2XrjAPeNkqhnpfxH2/g5FziJ5T
kPebF00np/Nbj2009cm+xKda6MaB66Sq5UungFstxVhSv6v0bkw5Pz37POkc93lt
2euTBd3w64L8vqlHcmE6FbEKiQ5ZT+nBxIqyl5PjLfLXPkBH1Gf6yXaofD4mKLtz
5kQgqmJAk8xpC+tIxpnmePtAJYAa5aB/j6D1MsEs3EPktGPAM+/Z24oc5wvRHQfO
xhG2uVDxJqeFTMqmZ7tELR1AKroqffT0C8EcE19XEvwTzcvC/j+qs/e0I/nhaWUN
5Te832FowyphURL/jr4z320V1Mi3kEOu7WyyiA3gPymss1edMRCsaoc06+0lqP2e
kvKah5M5+A6bkszaq9imtVHZWMIam3k3KfNqFV8H5HzYmeHpwGpXSoBDJ1AhQDON
tVFNsRgwceZhV9gdRbBRPXiNRhj3xtCwQebOWiaSgetSMeplrrSZysPGdp00xXj5
3ytUU78prTzUG+Y3vQJtejflzmO2bQpnaZNvy8NX01BpHxJmHzMYutGhalrC80/m
MK7FFrVa7X+zX4FEZhnXqw2vLhfMYpPNhg6TzaSFZoGYzpssCHRRxN9341MVN7pE
REuZM//8ds7erWjhVRjx5AmN3v87UaDRfE0aTgBTU6YRwtJeEPmIa6nBQitdFjsf
IygEfexZguAaiemzNM61qURMSMY5gaq7jH3JOmm7rM4CuplUjldjtb5ZrSAL5Oo+
zLQxFdadorqXF7M6GxwMnA9ms0HY72e77NuZ7wxcSW3JnQvCNLnqoi6jBwRC/3HD
ShoSu/JkJ6ouK7u5dpwKpRzFFzbyNoNvSWdr+jCcKR+lmysWsP3poJLtdX0y+3yw
k14oo6dOe86p8/VuoVvLfdmj0ZcyMxLPpuuRrC0Gl+XIj2E+mBToD4sbOVwkrgEH
u75c9sh0ZW9AcpSjnQpGxFYnX6LW+662Gv9bKGbHw2NpdOv8wYCjRBfUiKKU+iM9
Fmt49P9igYeO6Qb4p33K/gWsOJjFEsfBXY+3YYvHrECvWtuugb5oikaXPe0v3Me0
gk7NS/Z//KcRfava9JpcrwXVCF+JwQvhxgMUADev2PpO8QYTr0FLdzIMcHtrGD3h
6bKEoMi9WwExYW3UWMvTDfgRb0IUKVO9lmkIpsI64SHFrmNzZxcahinZ5SfPuTbC
ko7UQ4p4JjERDxAKTu5wnz7wKIaMtjx6Sp/y3T4OvRDCrZkcbXHMTt74pOD7bzpL
Or2AY9ElORNtiG0PwCrxp77Bq0590TK2epSqhY/woErfI1tMlDGxEquisjJwC1Ry
GqD+EnNLAXFxaX/AYxJWyBJkCS118zSaNS2ekDeN9hIUWkzCZZegc7AMyk51WciI
2z98uWhbOgdyzzyFFSuGHgWQVB7Qm+iAGtCKcdIghPHkRt309xD16SupVQtkq1/L
RylnZo+E8BQitSXcZRDi/ms3N6Zotks6iHLPXNR49YtNzJB3jdYB06jbex2Wgbf6
DXPuj/HuHlXKS8wVY0z8Y8ngWqlegaNNYExk3I4jwGxaQ4UxAcHi9e4+WKon5jR1
E05oAjzZIktr5URQJQUwCrlAok/fslMuniBSDx8HFR/nN6sWmgPuIhZIeyNjj6ng
KKHJhMsf/xwrk6IlVj4qSAgIn7LIoOExTPkZpRm0IonfH7XbFOJZdMLMm5bxskQv
E7pGtp7/ZNuBS1zJwS8bsCXGcrHutC/dBHcD494Kw2vDNvb30d4bTQiZhBNAs5Cm
nXJTn8bnJM3wjED0A4kNKxbQWv5zlySqEwXCDziRh77eUNXiY8ycb9nkPQq7viGW
55dKyl6ulZEGWYN3Z+O+/oWI7PTNhtC1tN2R2CSQIta5Hw+FJDYRwR1oxaA07rrr
1HvFagIdHpEF5IS2nfkLZ8FykOlYwx/GPHf0svteyNK7fyBW+HMbrQfspp/QsndG
u1iOALZ/WNXU1eTQ59MBhLuitKPgBbbmNE20h1MiiPV1R0JVOVu8XvqVjcutmRuR
/yB5ulbtpOXSxqRoWjsAbjEr+LOC+tgFnfoArD5DADKzrS6Ja2u4BIlSOze+fabi
3v8RmEGW8iiJoumUmCwhR+NWnHSAVQ+kjIQDtrYtSRphUnv+eU7N0Pz9eUGbF6x/
USY+0GD5MJ2DMzRLKItM108EqTJBmNKI3/uGwwnDgttpv8L07sVHJIx2wGXoOorI
W8O5fVuiDBfdrjNOiIGcRxc4QqlxLazVGY/K6FWMkCQs2QuoP9p3ZhvT3hYgwJP+
ZZV9Jnk9nVNImOyGQ+9Q2HbWov3NHc/0hw6kpnp9H9dGBDlaYt1aPYz2niwCAkbl
H7dTdkRde2l8HtaS5fscLwsv7WOaMYbKxXvpGsKjL5Tlsrl28xe11c7KmEEwxp3L
P0Bi2DotnCbMasWS9EWHWINx/NUrovH2i27zjo7p4/xNx7ySwG5HP3lhSP6zaB9U
6UjnrXTM8ym2mM4ncD/Trkw8Bv64+vd3orzM8PmE7CDPbm3bYdzbg/5AN8Hgl2ae
rBpUMgSWEOck2PyYQi1GcYA7tubsjWEWe+INNzpWtcp39Aea8J5JlLh9L7oHk3QA
yTTcGhnwQyWsUs8hd83IpHhaXKpQu9VWfY5Ws43kyx01ZbN+wIORGGIvnLbtO2xC
FIzL7jf4r+1+Dax1mLe1DRuAl9jyZpHQmJ1ObHeuxILF9D7i1/y4alTaOuyUAl2+
f/XuyiyCoEUaFNYuh9X5FtmoeAHEwpVRZ1DOoEjNaRaNBor1d1kNKuC/WqDOx0x0
mxyhEyozzg3e3g3j7qgCa4Sqjzvu6NLU1Zq8JFAZOOCJ+0tpzSC5xXfj2CR7Z8KD
5wWcttkaYbLptTgNTM7XhQVXx1QMHpzwqja3Y/ykr2zmD0VZNg9jMKtRXpIHaR0/
ScDqYEAWVKWCvjmav8UCJBtu7av0YI1v1hvh7OkRdZg8RL3fQJofJC2fOgYC2y/L
hvQWicSxanycjUjh6spVMB0r+JGL2aoTCwSWyoCTMkoMqlYXvvvNB/rOM55J4Hbv
jP5MDxO/2U/v0+ZnzXNDM0q/dxVQ07rVouq3LEbOjVhgmoYgqaEaWCag596oX5KG
udSWrmm2wdKFmce9Hrpj5C/eJRB3DLv0CRlWg7CI/xWUtysMu2J02JCmiGPZxU1K
sUCKGa6iDdl5CRwYiq/A1p3ABlcsK1n//oL47Sj9N6M5/pkHoWdVkbMtQfZ3rx6v
wRNmlMYiG1YQmwlYPFM/osxsu3aHskrLBnx/AUrSWgxK726IPuUBcqRda4QXddnn
Soa2k9oG77ZTUw2id//eM2L5lGRV3mYVFUQ//t54fKUGAByyIIscotcOwuuq5PqI
2N5eIP9oTYvjEaWQL+UYqwXm709Uoc8PxgOvwnOEc3R1B1s3EqBEfNHhQwI4tQ6g
ncakk0Ruee9nKyod+aAtJ2qka427+i3oXp9n+TTOu+i4wLZf22p05mAVoN+EwKFC
VB2aVXNwL9JhtispoHjNFMGPIQG5kZSBUc5h/+wLdacPiArKiaQOAyNUNtrb+iKA
FvWfOSHxecMBGWE7lsUH9pBi/T99WtF9QRe3TaBptZo0S5hjsJUUQxRlrT/eJfjs
IUGb5r1pxxMcrgACGfcjqOwv/GAWGUBTjIKybnCvmUaXv3sG6YyC+tuTV3UgDCEv
ivCOe+e7ZnOt4yAYFVkyPgB31hzhcNhN/m7P/4xxy05zbfRCLtNsiHj+8v/CcZGq
3R9N1S1x0hhfonTcWyuSFm0JuUwrnsCTf6hfLKu1UllwDHc5RNwzLPF8NQzaW2mG
wewV92rah9/15vf3st+MkqkBckCFt3AaXolrYCnnVG9TAxdJqD/8SJw8skD5rbxI
yUGSiI8Uyuv0B5czUT6yAPhDdsobEJrHylgKSzka/m9u/zWYuhSut0sEAlUHfQGL
qcxy4mg3z1D5ulVhODta3/pHV/FYSGfsntG0NqooOGtMX8zilnoeIqPYYfuJwW42
4MOjZIp0k0A2iIjtXhp0mooWxvOT9c7ZpHeiMGXNthuRJUSRS4HCidDi2X9adYNQ
c9Gbh6s9T7/OJE23R6wS+80R7tIfd84g5CjkqoA2afDkDDT97VdQ7D0WDZVbkzGc
DorDB6YTnSy99tev1RmGOuX2BUlATEp/UY/Faj5sa6qarPdkkjY7omqeTa8jYPKK
0MVtLba33XqRRZ3RSvirMEH5yjk8TVsTvXC8twmKKF7w9+Dlji2/3aY6W5+yCSES
zdXPgzE0PGZBUmlaLpLemgr42vBQ2wXkU7ZohbKpvEsU3HRbibBJiw5SCw6NGPSz
PRcr/1jMKtESiTikpBl8iUFVB9GagXOaaEcnwOHkjXK3zx/4da+LYhd3cREDd4pz
wdXcRCEBPi2DfazzuIMrXsfXzbXP084IaOw/gXaM3nLzqU3PZnnGEMtgd0H/S//3
12k5zuW21/A+Ag1Neoh3VO9bk6VYPzX4OCozrzAJ4j8rXRmXYwu24C/Ln4KZwxmG
/rDNjdTMX12U406eA0lirgQv/1ixQbLiXZo+moucL7t3FokZF7x625Riqd1fqAZy
3EJpwyqJfntpLg2CQNB50zwhlIXTVKJTFphABHd7GrsrP3wWDDNnsj1tYP4ZXhE1
n0m8XqEQYtl1G1Miqk4Q5XlxFDfsFWtudIgfmiWhAQTGeqvkj4Ps64LRjhJgUR+9
txrVkQTbXqSkk9uw7aWrMhc0bQDMCfKVqZVKNDwWyVNJq2BcmKPPusXCYNVMJofh
V3zRJa4xsdnqOfZME5e09O1aBry5TqfyHUMuDGLFbodflOKarlSzn4ukDLvu7ETz
P/nLPp5+0qX6j68YESvOZ+S3q3QFQ7dDmWgoprmWqoSdLmlDlLMrt1sfjer94UEJ
LJ4JynUNi7vi5A4vyBxEvzbZTJcuK85ncNCXLrngmI067WDaXiX9D2jWtIBoEc7D
zuZPSHMJjZulSvNZTvCxldktypVJij3ziOxW4SVcXkvQqEODPajF1iC4yjgNHgQ9
l2EevkX/ZUfiTLgcKeHqd6mcboG1c8+7ntyXt3zRRiTYJfXtHBawnX2+tuvpSkN4
wBCBHNitgy9/VF/vpjhTiaLwKSW2/TW+oQJenNeMY/cSMJUDbXORAj2m2F1acpsB
28xa17IXfQQ1uv3KQRRHiVQ4zKSDJQiIBVaZznlvY2JqZ8dJHIY7PAHED5RDC9xI
InE3EnYY4pxmt1E6tPYQB3jcrPYNWxH+2kzUT11EDI3fDJvXsfT616175sJPrCFC
1uyxoRvQF6+VCUFhuG+4y2y3CZAhCO0rAqm8bWUrtceyAdWgeIEdZ85ulplGtBxK
aYTzk1HJT8TDr/8RmIsQ1kxcOqS8r1rQh9fYt+sSZQI1AZJxW/qeeeG28Y+ETMZl
U+hJUx3NkMePUdqIz8OqUhND2PmT15tbyowWMCig3dbSxmrPk/gsTbiF/4Qnj7iG
rZmJRo/MbTcDrdzXflvsgNYVGFZuSpn98oXJffZ8sudDKBuQZb++NJCgFtuYvScf
/1VxrUPymx7OOldoePHKrAGbaOK5PTkLboM9ONmhH72oqkSoLREeMrD3HKTK2YL6
s5YlHA6+AQBEU1jlMCzywLjO2OULjxeRaJ6iKvEHt6ZwVJaUT3e6/+TQ6rSJ7B1H
6rTeBDtOsAY4ulCihYJn/5BJ5nx5PHMdSYZ9K1V7KhJ8CRzpQXE7AQLL5WkP8e0m
9eUkkpid3Xp4s7ABRl4ZHd1XtUb9JA0HazserWuVyVnmSzuK452ZQNHOTEwOPfwV
Sd8Q2Jvz1EJR65E/RD9ssRDueCbhqPSWglsJe0uhdHbIND0k1DqG2Jl5MYcKLxsT
5eIQTI9UGEQZRPVZ2KRbryZTseE4kXMCHiwcgRwWs9i+PUIhXGxq/nCD23EfBn9f
3m4I+Kzs8F2aOMADXedzKhPFRNMvH68O6RGr1mu77zAGjv+NLITJHREW0qr7u5e5
c4DJ82ddPj0WAjgfUvexhqP8V828V06l/AqO5BHwpPBFPo1DVPFq4DbSpsS/yNoq
AjpUu4/uv/yYESTvmZYR2ybXIi6XHUwwtD3QNr5OiNKrttW9XIKh+4SrjNCPKWBT
gJxRJ6AlnCl3s9ljD/68rCslRlWI9Vvw6WP2eErAIhSI8dlaV6LtGb9h/z5oxglc
6gJB/dj52UaRoIW6iRhQgZ+cfaAdnPcdNnKKz9oajT6MFivy4IfdIg42rKmHquuZ
LHbCTY13LxwpBzAw51VZyFQcZWmbNoH4BWMazYOIv+vGw3/XrZQz7xzoeQvmStMv
G3h3/UpByZn69cAIKdJirGY6cQzE1+VyMQy24IXQRub+1R8hsi2MuR3VOcfgqPur
9QKcbzOT3SU2moAcg4AczRucQbHkqksM5DSmqCkO8sjMhVuDMtVKFB/vhCt6Xm1R
fIX/oW3e7QH1GQVpYd0p/8CoWIvCavdTS+HCYFY/YricbJtho26efyMYAgUYppyR
6AkVn4OoWiZWtZ2d6Ia2bepk1tRX2YBQ3eSggsPwKtJ6fxW8/ImAOAfFDyOGp7Vm
hh2n8B4V6xMt6xCL3zu2frex/wNiNI4M5oGQdQmiOs2oAtqjcunl6Z6Mh4evU77h
/uubU+1nEdwRMCEEhNaJLg3p/+7hfTB7kj9Qpy7vPiML+qxQPkgX+3Au25xUxMUN
+ZqvBeTbcjfhkU3WLuVB4ZSp6gAYcZAiOL9vndARDFWIxbBKFb4lmAkuxvWjfELY
DdwE1gYKtqSKb4GzWJPaLgyf3a17DbCKCHabhz368OPofmSfMVuG8Mz4LirlWGJ7
jxq1qw9CwaPF8WeEmXTolsUBAiUa2ID5fxgUIQWXdtey//UBEAOpzjZgSLWDoDMS
69S4McirIGuC818Oz63yr/ofIPy6yozANNkbCDd5petSKhQ1zvCd+4fCsYITtc1D
9voBiiiCa2A6DrtFELdiP93DcPHZ2cfPoWk98SCx85G9QcU/1NUY4DPLu/RiygMv
7ALA3uk+D56IUsB7o5CH2rzeomUKxL3ugxpR33tCWs2RTSHovxF3veiOxkK2OAmC
VOMY4vr3S6Tjn6BFqss5AiiWM6eZApLwjSMjkun87yxS/O8wUzrogwPYitqcFhFg
IDOmNFO9zGHpUvNP/S369iAgSZgiuLcztxcfk4+ZL6TvbUgUM0UVutmolSrQ1NwS
oAwkG1Sh2U0LxdGz+H9uC4PVQmqmZ7buPZKMOUpDLgEEtPw+wh2ptNxqGbFKzc8W
1n/PAtDZ8fS2ZW7y0bGzcDs+FP8H/r7tG/NwpN+KPd6HOAaVd+urxn6Lx0Vqs82/
W0vZcOvjABgYFZfAVEVbVsNzOCqeQVIOWaFzKp1ieNdJCbK8wHlS8yUQInglWkWD
jkWVajD+zAyxG32KCuLx72nTJA+gmXWlC/bYsgptm79ZCxG8ohjJbkooQ6ESD3fV
H5L+N01pujqu6naNklZctVdty6r++VETMrB8ITpgKyjZsYr88inwMgJ2K8KwkPTw
nLVaeENfLQ3cZyV08vXaaK89y/+IyWEM28v+C5VaS5YoJ4moEchuX9ifTqGYHwCM
6fWLe3ypYGg4A5T8cfaI25lO2lWdhCDAHp/bWELKGw9Mr1xeZgOEHkHMghbF0CiP
4L2XGlPT+Pkjg0t9/1mxcvPfGgvp23qz6/iOuHrt9G0rrLasBGEOBHj6mv06VqU0
2FAME1B2zEkY7GU8qz+ACE2p/qdwR7ECkNnAEfO0/T1l8KUqaA5jZdLC3fCbMgfP
srG52BOnbM7rCfeByXLgfJ3ncD+n2ZeH94jdPbvLKJdkBil5h5tT4iEAwPCtBISO
KEZghqiuNT206abwoWT4pSwsSCd7AQu/Wz/8aWBrhsXZosVH96JbKYkuG/9CzSPZ
uFqqb342MxfgFYsFp+ea8gdQvxpb6Vpe1F1rxfOHVjNsapwX2RuUAQIoq4C5LNRd
KUXhXMvK8ENYHPpEW5BulQMmB9vtDkdfmnr79rtPvrwdRB/zQRzQikvVx9HQMBqp
wEmj2noall4+h8MtSKLYlTl4Oo+rLwFnAuMj3QfceL3Li/0wlu2AFnc1sIHk7z4+
rHXZONGCLBCGS3XxJIkwaVY3Vl0dik0rWMFvVo2qmElMno7ZjsltcvfTpyup6Q4g
7W05nAwxSYfxjl1J0jNKVsl1pqG2yRiW54sAiv4TW6yGGhWMo347tZgfnHLYnrFh
auGQV71hojkLHNDzQEuCcrkJ0700VO8jxCDFa8bN38WXC4efNAPioaP39g+YLsNj
13yl2MjR7qLpbuOqQuW43DCQKHNzq79M5NVTwSMVzzEwKzSanWHyQffoWnjdulJk
TcRPhfOMX/b3/11g7MdDalSx+F+3QEZXlDmRmZR+kaSuFHib/qKDFcqJiGqH4Us9
S/aSFZ5l8ymTYKll8FkbHcz/u1sv7r/Gi04j4/mp3nlhK0iTZ/Gh/q4hseQEGKOo
lvt7HsAHPaDblyV+oNF6xzUGeRoFNYZD2d4tk/+B40Zag7OO4H3JgUex9LB0WS26
6dCdzFSNn3xgEUlfPjTm+1v4664uQaJSNq25lhN3/P1vtDbZI5mlMeDLhoxePD3W
vCdVj6HB3YV+2mvXzB+ODSd/Zra5LuSZQi1x1NVAwRnWjpuSkZRwwtFlrfFFZXzH
zynAf606yi0lfmaN/741VwLGKkCVuXc4jhS00/rL5/4uJWvj20rk08ZY6LHNSI/F
lbowd66d8Tu/n0+jpf2nU27EfpTX75yPtYM34Sp9Lv2nB7++eQi2W1fMl1RjxkL+
zVHMM9o7l/a4ggPX5CVtQGF0g3MzHwAJQN9AacHi3DMrKDrbfHhYVgHB+l032/sI
FwBUJxSd3kGHrRNNCRagyiyConGkWLxX3H9aUHCs0AmivtoDa5T8GMHJgoLwGthw
MmHPpUCdeHPw4CzMeYER3vmH4O4DsmNSvbkNFp1uPFdhKEYErlJnfPhqX9u8YOfg
0FtBA7lQ1NSuRaXUrOHThAI330F7CLFTxTDTBVPqWhkz1QlLv4ifx6Nvhm1fdB5D
06Uro/pyOPvVDoNnHOv52kxbsqcYsL/BanvppWR+ga98/RV+ICM3vtS2hFgVUvZm
nIpshfGn4sIViZxk59a66EebFh9UlbWShpX835SmMRkXTEnt8jc7uaixamJNi+yX
A1BxgN+TN1EC8szMVJroZj/8mRvKDEKevfpLvyfSbhW93XAneIZTGsQih6psmY9u
HATDlIUUUGaIFQXawW/KzPy0aIpRaRh7akh04kpXtEHRpKk9VksWrTiIMnsjfX4I
StHIBk3Z+X4u7xH/IZyaRAbP57w5iJe3d27xk21a8RWrvuM19WmUqOkN/5AkPReN
ly+e41VSO1Om8ARY8/Db0d3BGSJDZsBqL0ttgpzYFp3h0zaulENBK0RWdSpO4//q
Ki5prEa3qW9VAqvSuw5X8vmmZDqRmSQKmEDDfJA5HUQls9wfYXPow8IO6AElTL+2
Uxp5u9DI0kP71ngqcqyaSkBr5NBTX4I0ZCwZWGxIYw1LQB/sD6gUvbUJL6+fzVeb
2UBlwYjb0jker7mqe48FjqPaNpxZF0s5k51pKyFxd+DCwW1uoIDZb3kvOHUUUJQI
/ckvsMfbuaN288ZpAUKcYGeInhxL1+ojd2kVQ2qdXaNP+YUEoq5HnWn/m16L8yLN
yNZailDg0GRUB2OnYpNH1z268cdgpibcEI1xrwjGo7sNyCDHogT6Iy9+hY9RpIzV
27yC3rM5x7tGGZR3/uwIP1fmWC0Vd27rX+uLIMqaBs+s+F/lPHfTyiCMs4Bu5KPz
77hSiijxL8LWqxf4DXcQ76OGStS+sFD9sZnxUgr70jhNVrSb032oqnseIfq9Zf/w
PYAi5t/Eq/ZdcA4TCuN/iFmpx0uO7XVwrPje2jLnwcsoHUGfY/FqwSTqmOWedHak
6yXX4S9E7XSsIdy1L1VBGN0+ikHCF9NQncdIytltHvUFMwzhQA9YYwoC6+iFMRT7
AHcEMr+T84oG5MoAGx/BJmUQNOiWColcLItKd5+Lot+QbtZivZVEEimNMjGlLFCv
2PvJ71zrPZgvw42LrX85JQvDGgmWaTJ5V76SGzWZ53bNtIywhGBfWVsBIQfIzfBP
9cEIGuP7tuepF5d+miBkh0gHJm4leyeGuOj9GBKEz+PGaJYrv1KzEHMFQeCNUylx
/pytANzPLdpgD4Knx2oqVLIoPgz4c4miqM8VSCkPGAzejQkyXclN+O50q/mzxdPK
eVbIBghm5afI8mq3iHfC55y8GMwtaJsneTOLEF4AB0tWGaAuehsV6ILnvmt+bFW8
oqZjZ9pZYMBzyHLrYTsUMHPnkXKpwi3scrmvmmROSil4NrLDlWB4nGD+Qks+OcQF
yJbUwrJu0jwhHdAGiQ+BUstIh0SMDml+f4eoBtpNHpC3ecHvXhO5fJbU7B5w6Yzu
kV/6sX9TwDqy2W6UQStV5YjGNBL0drZUBj5sBThzVz51dC2rjEi9Xda7bvWE5wcD
BcARYfZ96li9cPWir4jIvm+PsUOSeSuy+Fc+fMWiXjRpVwBbmFie0p9MoZNJeRgw
5voYSoBtdJExKEX4D9pIIkL+MJB+m31YntyJGv/V/HmoTNrLN0WqeVOZJLNCROmu
K4vox9yhUZNHt9PzGZ8BlV2n9jyqJKePNB6t0MdRT+9/HSrklNUv1iC/022vJurl
3DeOeoUGmKP8seTECoFyK7/nIQhlQfW5wNaBrqWR+k6OYWFqwlz7+kRaXrCHYMN+
j06gsJUrKbyzeigv7nSBnIiIDD/RTccQOXm2E2ydLFMgCXRs4FgZ5yruW02kQbQD
h/YE0a+iVTHLd0+dVl7jPtBggAJilMOOmK1BlXMepjeeCsP6t5hWZTO8oYeFLE3a
2HNvIypk4tpygB23APD97PJt0AHISiIpLM6Dqj7jfbZ8KBkFUUKJ2lNBkI42WtGw
IefggBDgiJDXKYaV/ii+riIcPMtU0vHF6TEXhlRJHkztm9GgE6ZfVpNvRXlXCM3U
h9hGryeKRZ67tMNE02yaVl77H7OD5wdTn8/qtxl9WVWM+GKd63/BakhVzmv21wAJ
alpPmLAK7kqIgDKtNcCmUSZqbitLaVQlBCIXLTvBQ0vzUehdupQLX8HjbOYm22Jx
cr+dgPnXafaW+tb8nQRK0ss/k9qaIYFEsHBWOGcRYU0dS7TXqQA2CSqSWod7xHmO
ROPrOZDPmtFkK71a+hRtIqPYbxRQvTGvofI2KaYGVQWFN1Hw7ynezWJxddmPSqkK

--pragma protect end_data_block
--pragma protect digest_block
9VgxDW8S58mWAknAgCqNdzGeJI4=
--pragma protect end_digest_block
--pragma protect end_protected
