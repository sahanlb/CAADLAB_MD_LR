`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
G8OrcfpVxEc65IwFWCHdSIp3+S0QrjvLRtGBI5dL56GP6SsrG3UbRK905KQCDjJV
k3Oulq3ZZIFgL7xapM6LVX/J7oRlLphFPrSvwqvM5FIrMT105dO1E/Mvyc7WvwNp
6wr3dzfYNxUePmsy1PO4fdDraclg6Cz7UWiCRBBZf0I=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 11088), data_block
ChWXAOyv4JaiyIUVsXAd7ofuXBLW01pDDm2tfFwUK4HYViCVShLpV0mr1XBq3k0q
UtFAg4uDzRoG3kdPGPdGqD+XBCdZqbjyrY0RDsgheEIpebcMhiLbRl22t/xIt41T
Do+3LQ9XLSYSVmvSagnfzaMdXMIxgnlX8WrtcqFXqC2qnuqyTXyYJ5U+QKuQN4ZN
buJHtu1M+auMzKGWF1jeyqt163TumIwvdcBLe3O8q40lxGTr4Plrtc5UR5GBKgbg
O9LUnKzrdrKrWExvNC3mue0rLOovit8Z+ZQ4GImdrqwFZlXexxFWUqvFigSUm1M8
fryieKbOLzHG+yDYYHM/ZJz1gCD5VGVcucAkrEZH3JmxydP4giC+4/s9ddlZznCZ
f7LbqzLC0lCN57OFB6nWSg3HAbtpoWK+T3GK0+D5KghH/WfiF78rmgE0K5UH9Y9k
L6nzBSgJtxslLsB8OMDPeDODmVzRN0FpjOQTzM3El6fqQev8k/N+yuhG2hT2haGy
xHvC9edUTyxlZ84RvmXdKr37t0jw0P5GW9VzdknL9I1E3wpD9VBvjLApc4mRbO0B
g044mJB1I90w+slv9Y0P/vUId8nsLQKrRkKUKJTPf3NEm5lFg7e9VpzivBE+gD4W
qPxXsbWIoIH68XgSg+QlZ1aRcZFHYO1egk1/ngRT8amduh2RbTHjalM2DmQuZIDH
qqf6SmPr7M76P4z/hzJRJknxJoIj9ZyZsf6zL9sVSsBhzxqRJSPYwvU0LT+UT+6P
7uX5Lsv9r8MobAxpFyo26PeYWtLl5eJDP1ypw6auIRK0yfWCE409i+V5ktPcaa7X
VAtTrcSEE0byJAxy3qZudYwTC/EFHm4q5KSpwRyW7jbaB7EsAPShIDBwICCzB99b
pmICJScsToxOQgLe5HVl5h5voHzauVV+zciHqzqNnMyWXOqeKNYQR6KBPO4mymsI
03xGCYfrEBP9eX+FoF5vAF9BTo4tkoT68TzwLzBHSriV/loMXnhBtQQJEMH6VI+V
F2jMcPikhAEzlgvAnzzCHJ8Tz2PogygXNZmD+w53fagBTj5y9Qo+4bFNbivCwzCS
XYMtDGVVKlJUwuh4zLhixip4RdPqqL92cmgs9jviJdGHxMwH8B9PoyywU2feJRW4
tEcZZsAucb2hWvZJB90+C4suqQtVFNIn10cEgvHE/A+cTXk/KX57RFGx5N0rMlIf
dsrxkojiPeoW56Q3bV0xCDGYgAc/t27U4eC1O/5w1c6GYurosh2uG0+eKR2EF/+4
+ZB00hzGs7ano/bAJkufSD7kJvSTbNvkvKnRW9cM2mDfPMPM3UZRvXtQj4uetMw8
neFzR1i8CZtYCzQTKTEDbv5gSJaAMdPBA9oZyJI8ZhlqcjONhsh/lkXh09KMxx17
dKpNtVPiL5U6BNS8vcJP5rUwqMgKfTsdZg9pUVhDheXZYc6c1eAHXmtIf0K/Jjx5
N+6hixZnM1uLm3Wt28BFXqBCUAMfZ3/pK8Ao8WaClxHBvLhjYjGzeES5JqOZnLhV
8doVVkKFXQ3nQaSseeklfKS+542pi35+F+iLo43JFJshYE5jO5b2LVUtj+Rm93EC
sHOaNeiNFTyVAqIl/jV/yCPXg4DX8Cm3dMhUJe+Q3p8q+fEV+QCSURFERyqvhB/j
WlNIomqcEfT0AUJrG0xWyO0glNiNtyozP7O+JK4aMyILJL+gzX9cN5vZgUTZRcdf
BvPThPpfmQatO05cw3k2zCZCH4Io5GGsGzGAiN3SXd7+liDwNq/pxd09E8MTwYHx
oNQFjeCUIgZWcpr6ZdwIhAIWGfh0eV++V/vC0/9jZP17mBu+E9e9irdJeA7iHU8N
8WKPJCiOha3oupbpmlaH2PJFNrYh1PrggxTvJ1Ml/+TkZD+Bi4XJjAAGlfRP9vXh
fhS9iPavN1BmXqi2s1AGbLhcJ3yJY80V3aDx0/iX7RSMCaL+55t8tNzsqwp5VL7M
3QCXRev59VJS223oDILHpbylH3l4XhJ6y3W9KAzFtOl6FseIHanJKyY2ceKwSPbB
CyoUiKnsOhAjjULb6OVk3fZYl7HHT9McJA2pu4TK4KN6ywlS3nGNWNqOemd/4h7w
eUp6f/b054Qnd7K6wzy0SzfNphg5kRfoS4mp7/OPMKIYy4kkPLEXJ61ryDPR6uZv
Lnmt6HidmXkh6ddKxn5PXop9vzDkR0TTFn9Lqfp8SRuM1kPqIMG01c8TGEIstSEI
87cNfi9epA/ZGTC/0VS2S0Dd+f1QKPaLEpQCxDE47C9Lrm0f5TGiMHy3afeUsM3X
QSdjjGtoRrXdTMWFMvM+/BHW2rHb0ULoX1fkMQXeUlEiOEoKwFvxMJPuWAh+nBOI
rjjwyvB84sc+44L9CLZTkZbwEKLbFvZt07QbKqjN0/e2r/KI2s/3DnWbLjXlxJp/
T3I3m/2zhzJmu22ZCoWDs3wJzBAZLH6+jYQ5tq24JsgijZO+w0KxPPLc1c5zriYo
+TGEaPm0L3jmKwxTsZ+8kgnOyxdOw2nVVNVi/WEv6b+Hla/PWXu+XZf0JJr26fG8
26QIcBQ6FZo7RGo1QoNw6g0fBp/qXdHN67LogDvJXQNDsSD3EGr0MA5GAGIuBsvE
LNdBBP7JgEF1thGs7MteTuLEcDdGBwBioO9JEt+NaaExW2lRbkZMGzsYenSHqBfg
czME3dzYzC9cCqtP2LA6I1lbq8haDGyh29JQt27MH5Cq6JoxX86AmwtWbkPnUiF4
sIyRzJYFB10PH+bpzXsU/6ua6riwT3brG51CqvMjwpo0YPW+SjAoGZkn37XUSV6i
1530gwBv5saToyQdenIfNFGPSdDCZVh8lNQjgkdf10xt3OIQ7ajw86LlNcN9RNWd
IEq62bMj6wyCMkVC6cKQ39o5+zOUFkZ0fPqeHvyLwOMqht4vALyBT0dljYzXAtWy
qtTh+arkI+m6A1pGCKiAKhxMxKufaAUUQ46CvbSHUGHMgPKM4L90USXPgfWIeU0N
CIpFhbg9TtDVQ5LUxUvLnU/b2vNhrx9mG4Y+x0vvHNVGsb2ipYz9Xvj8ZgHgNE9j
sU0k4Gir0px2+SrpK6pZhn6fu2Xj93GOtgYKUgrmK+dwlgyW4JJrr/XHJh3JJNIx
UmHHoJ1Ijearqi00QOdZRjpEPMjUyNAVQc2PO5RPOQOxEW5f0Sam17yiGon45mfq
fSdZj870chqDgroRY5zAgKuVoKyD6JJCSL7khaChd7oXURiZDE4YW7Nr8V1QyNWd
lrihpQnFi0vkTD3NyDu2NDNxf+VZNlSoWl/R6mTGLA2wUSjqVXZsobGHsWJKjl3O
S5nm3VpvkcbbRBar9QPUpiHXbaCw2i8H+GkL8hmvCZ8hu7H1PcszCAYYztY/i1xv
hUjmIt+EoBwFMKS04Vi4agMczZj5PNjmXQSErmciWJSOPIqm6U91g7j92I7BAliu
L6lEVXUE+7lyXr+AHy8rsb9KmpqwN/bFy7FJl+Ms9eIoLLlckE3hmPevE4rcazXw
33hyjrro+1j3cN3DeYup9uCq3STPJHoHntmy8eOxHfidsx3wbnnvu6H32CCnSwds
+BB56Ea224wV2xKCDlMu26lKSn1GLExnEXvuwzAMBr0EKoE2eoHXqfYzv6y5WQ4V
Ot8EnkykcqRKjodm513ghpCjHSNmk3cGFsL23eNHql+SKiteuOqot+5Dip+XZmYk
Rkfo9xRaotuasGr4rSuYfH0BMhUsSDR3mgOSkgrq2DnmW+fHc7otvh+Q/COYpKA/
0kmVQIO9mLnG5T6FU0s+UbB6lBVjxL28vqjwB8Zrw0gQddyJqM1/gThi+f8PRv+0
ECUY80cGZj5bUxA9uS+7idnn0YMsFVELM29BIF/euvcTpkf+OK3XW0QY9CebWGW2
/VZ82SEzxqkI/F2cF4u5KDQO3NuenWfvNU8jCZ/kOMcr+WHo9r2rxxDdTe5/0hTE
eVdJP5w9isDal1N8/EaXgCIUCcRtU8ZWEjhdzVs1n9LBviE7ohDbcBCgPK9tGNu/
ob0rTdbaJR7gqbh2CxhjWOXvi8Wh1ZqlsGU2hVVdPJxQxt4VzA3tNm93LS+O6ouQ
0Pl5ZPvJKvaDdzNcw4Sax92clsBBJ4ALVntczAc8Nd20/1Grvum+1yYgcLCKdEHu
XjHzdK6UaPMEAqn+UnkmBqPaef04r/lEejT0eE31Np+Cj8FUru/GVGNX65v7PW1L
hRmaGqsZSJybPpXjyn2IR4gcHC2p41YaY41hrQLpGp7OdmvXfCr4AIPE3Kpng/n7
prdRYF6fGK5URPPCYJ2uMBjtG2RBHVvwk/PKgRfrQ1zMXQXUKQHcuVZygLB965eI
MF2BKgJLeBef8HHIrn+yw1Jca6UGPP5Wresh2whX9N5GlG+dU3ON5eKLc4xX3RhE
bCqWPxylX1GlHHLK0wecJYt4ZctXocdBj5ICeImyVO93tA2d/ro+MduqRj5MvZfc
QH2I6S/sT9cFeOYhhBCV99u7dz50VvHlR6oZC+IhdjoYQo52PS01j5n7DHTrJxRa
i5AFHQ9fhviltBcBPADUV7YES7a+05Nw+asAHjE+IWHoLf71jzyorP+nPphPZ+wb
5+VYO+IIOlf/qKA28rGxwYSag7ak+KwdtEFS7tDtIXtJeBCY47F5qahX0UrmB5QB
BjI5BQKR4Ags+HaCw+EL9rtIpJW/LEBkBf9iAQIzgK7Aebskck26DyAAmfIEluuz
XBnpqM92ThGij5F8LR9KHTf6q2YgZJanh9zEUlDPXJqmQo9D7jr8+bgl0ZM/DOC4
kEUX8sp3+DoyBLUvAIRXksDSLJRUH870PVvN6dInRo+sB+CJmnSaMb2v4wL4/onS
0IXAEtCtSVyE8d8Y9NY98OgYuC+LyT21GXZmLJXk97l8aX6vbFHtyKgE+KkrzWJf
taUhnpbNIWXueI6VUzeDsOH3XsJxW0aJ/iHr4jY1FPb5oOnXDQyN6LJ5ABQZ8ggw
m09E01fmQrcNB5q2wtWhEgJ5wWb8yy1W43kTeWEbFOiSX0Tiokm8RcTPeojKYPDO
dKEEX6qjBsqBhEZ9SE7KLj543q+gNCkgzuwvTx7ftAxqFqLhKyJYVWOEdV2X6s8+
aJbGRDuiITomzi+Dmq7SAjVUPbaYSzNT6TPQL2BHWinfdLseNz3taZ5GkQUKSlui
5Xz7cJTTjyP2TonVvvTf+tYbfAFs1mCa4NyXA9kde84W420A2sbfJB0aWrGu2Jdw
oDsp0Xwbu2jMquFIlsWOWIQSL1NJzkhdNkvClHWfvPwMsRCYp0LLYCDsuv9x/GAZ
xgGfhhF2y/dq0ahbZy2xh7O033OlTZyXgW9RhGJVDK3irlLkS/uBy9Z64IgAgPnY
jjve7e8XWpIVR/BnTUqT5uWQSQUm/UPOjdBqmCBHt+GFl3VcWHs6omyoVvzDi1NL
jnyfH6mc97GjJty5kT7XsuwwE/BDErfKFP0ZdGt4itw6VBzganU6PB9GLD8j3JwN
sSKOkz02Pfy3HJ+SWLUCu+gsmB9BYZYNmBWqLLuzNN2hUX5z+BDLERefVmeZC7PI
bi7DXjtq7MSJU2L8H91/gbwy6dyYvM5rJK6CVeHAqJdXv9ws2ZtXu4sKBqhM0jju
Y0o0AhVedpBHR1Lo9fg1XDwvzYnktt6397tf3WNUmYsEeBox/FjHMy2ihLJ/pTxj
qT7SFcSkIifRVBINEhu5eu76PKLvcAFyVlKfUaFlaBRbDHzrjG69dpJDAmQJ7D7u
t4uGddEnvmt5a8wpudYuSeLSNIKkUBGHl8Tc9dGBAowFDzQ/dc+jgqTHx3vjyK0p
vKLw1Km5Xrr4hawbU+ZVM0vZJRRE2pWWbvgcSiP+WGvaBqyzuFWt+xc75rydbXJs
/Ba7cta4kqmi2gV6nM7nHH9Ik9AZMKw0zrUE6LACggv1HZ3VtRSuuQNVmk6RjPmc
BqyIiOcayT6jlLOKW25yB7EXPF6qpzvgkHSU0JQcwZH6kIDFg2V56tv4N0W9HEg1
+y/uZ/Se64t+t6Z8NLxeuljaLrzOK2ViGii6kmfMkwsXcRyT+yCaF2/2m8Rl3KW2
+mrfn14Bk3M1pjjfZUjs3BWw+9zgZ5+iAjDvoN5kFPXuM1t65LPDTDDZxQqO+l9Y
/CVYb7aRifcftQhvqwE8FpLktMf3oIyj6HgCJoYeBvyUdVNk4xeU+wbvAseQyYDO
UqKatqftIpIeBG/RUiCcNIDZVk97KFeFJlKeWrrrALEim7KCYY8qIaYFaNZsemWx
gNpC/PWilti8nAGfzpzosP8UG4NjiP2+gXzWZ9EXlRmVaD53cu30bX20n+/Da2Wb
Dc7Wo9NcO1dmO8QElag0UHv6Zs9wt2cYwoXzCtznt4n8vwyUvdRDcNJyxiy6m6Ft
N4JyfRf47DsbEkfbq9/naMFie3Tm3Bvrf1f3i7WXXsQZZmPTIrTVHSUTG5Ei9Yew
bhQmgJwW/DbRE0V/5KfqD9L3gCz37uIElgESYHRB7DKQmlewMI6Qfs6eHw6Zmvli
hASwO1+CyvDwvp+DQ+M5SEPI+ZEmricR6h234fcQR7L7WABuVz4wXIUZwMZbX1g+
icYso/kO8BThZuOfhzBXOMxgCEjYVrtVRRwj+PIke+kW5B7ryrv7Uj63baNUW+nC
4rSBNgKIQ5S748U3naRQ4k6Ods7LSW6vVI2Kv4lJ5JVbgchtaNenQzvrjgk14r+H
y0POCg7cP2zakWB+CabJti9AfiPWmAGKy4QJXRRMU2TFskyscGEqpkqG03uD08K7
sm/Tqy2q0NOHdEV0EtDpPMOaIFW045fFzeqnvwKibpQPxRi3EAeavgmLPltE0y5V
/Bk4HDP98JH8RdIPabN73TXHyJEgop7ZsJigb5wqAOPD7gqPBMQSqkfgQb059+qA
nkIxNmtJx/+f7aiUaSAUpo18q3CxV3VGFCGzEIqyxVlmmaPKZGH+BuMSUbNfcIAG
7g+LfKiYxAXheeyD9fbrZfsHJaK27yIp6LU2Z2n1JJUCmJ3ulFzBm/GBy8vMCI10
WdaoFfpTh0WMcqYL2Ah4mnB+IyAhSTzRuWp6cNGlmDmtr6mc0I1DGgxYLkYIqc5s
mQdBd0HL78y50leHjb17NWHz/JCsKBRPtLwciHhyhiKZX9t6wAxGztkKBTr3BvJ3
hA6FTOgqCU2JOXgqHAY4I9G6MWpijridsPCqNfBjQuMiirHEBrK+h+2VwJGI+VfQ
23rsPvoCn4fUToXEd3WyE2FEb0Song1VCsS02tsUwqtX9/cOYUtZQglQA/K3mCUH
1W2jrcr/n9Jy8xQQjXmc/ANW49a4UbPhLmOsL+Z2R4/s5Tk2bXJwm9HoI3rX3mMt
ZBnAecDWBuTazsGqutPq4NNn5JxwQm9N0r2Bg+Ly/dPwGtzKJ4eRfUBgQuRvlcTj
OE23fnitC9NVQfoNJLAbRjt7gjw2YX3OaJGhnmTkR3g/Z+XGWuQRU1894ezhDj/S
BGi5JljwiJoeHqYIFl7GSsrQLPTYEJx6/uVTy7YYpWqGppU1s9DZ/5/hom7F29Xk
inoZ4B5jrKaFrGxloXHwGcCxaEHVfupkpnlh+eSXIbEnxTDROOz6mkdAVQeyEIIH
K/6iHn7kCegYdRVAFQxOExJyOkecrd6ZrWS0UbUm5QOtmPFFnSfuy5b5e9vE6B9X
HZ23bmGfa9nRS1vJ5KSvmD4jiduuPO7FePDBQM97Uoh91fUJlyf497UUuUnv73Xz
qKzHWVbCyT/RljRVoGzPomH0wNpN5o0bkYqJpOSr46Fqk+aqojOaUpwTUweogi/5
BLHVPRFOV4QSnfAuUtY2nsNnpR7xAo38fKoRi8OTxXhPGDWIBIuzr+RDfA3+SJ/k
5eGc41G0/Z+54rse3wb5ifIMgFtBeYylhdbfG1xQxzYSox9H2og2ZNCl6t+GWo9R
fIfO+qMHnHvKeP3Z7FL23tJ8bWnmvwJrfotFVrbdM0LAc30TwrdNupf/l3G3x2Wq
Wvb04yU6y7WGQGBHPXe4opIbZpPYjrzCahVVX7747qPNwSQkyrSyu2BP5Ko13e3j
hX0OfJxgjgGlF+MK6ijuMGpRbAIT2JAG5YIeiljbjrqHqbDo3bPfLYKCQfJ6bV0g
KgNn+9rftJupy/n2/BkpOZyUNOija04/YL2Hwgbm+597gzYPAmSm3MW/kbhoGeed
1FbyQGIwPbDACtzR2NPQ76z8McM0Om7kdJP8DsqdejaZSuwI2DnQJp2rEAVfNTdk
I+/oECIDQoBolGU5zw8ThJZ0fCmxo35WNqRy+JdVBz+gwvhitGQNcQh1a01xPmGn
xnUBqdcQUvEYnpzYU83DpDzLx9v/wX8l3aJCKc9xKMcAz10fw973lQwGgPcotwi1
ITk57gAGXGGlRljJHh1S2Rmcy1kIrhdM6Bv4Q8R1z3d6rTXUrkboMtkb4o0QwRrO
Q0aTqfo71MfxHmAlA3X2xr0hMPr1ihqBuMdBYmJBIokiJzneOOewJYTwBaZ8gY7Q
Rp3cBjHaIieZCs4rG0pKhC3gMQeIkXnGIkB7TbMSJvu+XtfEKNq+ohZYcm2kQCBL
LiyYbNV/eXol7P3JjQ45k2s4vG2YyDxdjnIH1LSTNZpPz8iLaLKINn/ITMvXwycU
dchnaYD5AxQZlnLE+5RqTxBZcaYoy/Ur2yolpDcIdIDv+ZZN1x7oSxNdwbcc7vN7
UYNi9d6C34DCnGhjQqNmr42Z1JVF7mNUpFpAfns+TnH58eZlnHPcDZM24/Cm7gEp
SuMRvP4fdzXh7SCG276aeuK+223cCQPzk8rDT2dJC3XxiXktCAU6LigspgWAZoJa
iyz4vL5klCI4I1b6m1EfP2QHFifBU9bGbhLSxCeYU4OynPwXddwnWV/XRGzlP2QS
uDNq1M+LFU5ZHLV8ss0OXNkYNr+rio9OMsQaDhJboGMcYwSFL0UnY/kReMOS9xE8
TPtUn17z7qhf8gJddL09rE7LahIh2CPxgVWBFH4MZ0qGgV9OsAZNMCwooseLkmJB
2TdlzOS00yRYjoGj62EFN66PTlO7hfw2tOND1BQxm+FRgPwD2NwlRWKcrRODaMbi
2B4tj1frnzZiAoNaTaUrutFvWXPx8eXishf/IeQPV0sidc3/EMzTlXUZ4yb0LJz3
KbVwXBOs5O2UkKiid2yancLZjP+Zw5yhY101D5TKm3LJFdg/U757y0c5SRp+e+JC
51zYDbMmGpXZCKzwrDE5ZeJxCgWknPIv64rE6sr6PCc8JKjEvyKIrTyBnZCIZlPW
CP8L0KmLMdEAUoq4FKDULDx4k6r66/JRKHn0yzW9N4S9lg/aFYzMiCq+2YH5fqRa
G0tXzpOVDc06vwMXMbQfAbULyWMo3agI5t+dJ/C8FKubpRBbBbcHQND4KKSm4ftq
EMrrmKtdxzNXZ47sW2nEJ9jxejeyJtOt+qRWeyH9MndUi9CA2SkjIS/UiUfQzwM2
58/K5oQVK4Hwrgpwc6KQ8irFYTlmtPdcLp5IwVLT5jDwxChFjLUQ1FwEmFdIUJsb
bdIixgqo2BkD9UctKTylUvP+aGKl4jHPo0LPdAVCokwudtpwSFfMmmFvVWeBz1Vr
hwm/PFjSkoLRFB58olHxnaQTmFPEZcQNTGP6iy0VdkK4gOcwmgdB7vdZIxojrSvp
MlXcBQ2yuhypnXywoGVEQ1lbEykMStyB270cROieo2coSm9ibMGop4DAiSJqhVIZ
qu4PkmI6N8/sAyZDYtC/RNWmToz0ZqXOvFW+Pt7/cobpTBqQT1k3Wucr2IPeJRT1
PtOC9i9vIDA8BAg0u/TugGV1ITlUTpp1yXjvedrIuOwT8H6Uk2sPfghrK+mUl4GC
9yJskWCYKZRWn9HxK+1mpeiQp5toaKWM7STPnTcYQbHN7byGCkwMT97N00m8mIpQ
1Y2ftBO++FNTzvjmxYNb3YH/AQFNzFUMHHzHuYVZDRMVYhHq58zPZjDD5X8atQDb
6tm8P2zC3oeWLr/nuaamhgPZu/zm4VEQK/Ue7WqrexYC2ZGrwdrwEn71TvyhOPNG
kJMxgh39I1QacjLs6I5VyI1B+CcHuJy4dpsRr7nQAGgNODplCcpaOkAg7ONeT2Um
zJjS5sY2kv23DsezfVCqipWnFgksB+3OwgJQZgKEu+iepX0uqTVOxQ/zYldvaVWk
zGT1lVdHnEuMHGzj3jzMo40H8cb24Kak/6tY6NpYeLEuopZaEt9j2NsN6iDfKA70
N4zaHvFaPxPjABdOEJaNH/w/QTpYRqR3j5Y+khG/2/KNEwxfKeO4g+DYxK8DVHh8
LYRXgattNGDZTOp7XNPKWktJcE6vLbvYX91SC0wrrzNBQyXgTZ+vbyfOH4ZLdz6q
zVmIANsEFsdGyw0eIJhyhX8RS6JiB16TAI187wdC1g/lXwd1T3JcVp9oR2cfkHcc
LNz3bI09ykqmOcrTDbU46vsgaSRQhS6jSWYjzYaLCBw3of8ETgRA3sF/G3X0pGAx
9phkVFn53UQMylJQJqBD84gMYJVqlupYC3v46diy6jkhPyUiWJ8gFpCJC3c8fqiB
T8GWhA2fdURmCCeXAHb4Z+02bXyRX1UTwD/BFhT41xz3ywbOyLyiQPOP6tGt6f04
XdD0g4xhSRnjw8nupi3AOskw8b6PCioDjvmRTGbvCcgAVzXq0no+V1aqqnGi6X5s
unr8k5AGsQ8quvU3dZ4x0Et1Skdm5OLCeH+fQ4C5+tgWJMe+a3eO800Slg+eOMQG
NeE7AFVZNhARsi+D7AakMbkXhX74CZhOdIqLT1OGtZBKK3njMdK1tYkmk3DQOlyo
qgJsFWAfVpcuGEut7Z+py7ysF1f9nquxkArN73ixo3GSfAzkRj0Yu+amcJhrjBN2
nqMgP5qx1bQfvpYwJtsXEtdBdbA/+xeEvkA3kUkG/hqxoBaEqvKW9CmNvkaEG/rF
2v+Ty3AqUxNEMh6kWOBGV30jzm+ulHZZcn5LemYnJYCZAP6Uafhv0mK0VJqHhcdC
6eYHr422miThCx/7mz5IqvXicMLcx8YIgYyoKvbkBo+XAPCbRWGhQGVJSmcf0KoH
YU4iQq4/kFEnWdwwjithFRLPZANO2Ws2houmGI9WYd5UBXap7JXNAK8TwYTPfBRc
WPF5lZaAevt/GhN2MN4g0sSALEUe6qb0As4Zq9m2X8vLHDajDMZG0WyXC9g/x9F1
pZ1io7wTGNHPuwpYrqPk2+EMy60tKk4gInfoCdzyJW3gTyxPz2TPlgusDJaIIxlE
YsHIOwO1Rx1m7d56r8jdYjE1yJjOuDSzsmrZcaJ5eonYo+TqGu5cLVC/u3YFCgsu
cY7BRgk9WIVh3wnq6FzGXbcSUclYa+nSJ9Zh7f/OFhnrIKsvTkgXc0wEGoctgN1G
lzXquIKNufVHoCsSCFJY4DSmCnvWeSwyHzVSvAYnJgtRnX1LxNe4x2eJRFcRNCUD
WRAItwKS3V2rELwFiGeazlAt5GHsIgKv82Y32elc5cNQ/o3caYbMH9r8j1MJ4fgy
q5ZxRAKFlUMFmJq8N7uDNKoHo+jPp9wrwIrv8ffct1adsRF3uzFU9DA3ZoQzqM/m
8lT7doHCI8J/gPeHdM8guCzLsgHd5u9LfaU7AzQf3x9gBnLm6pr5oG20PNomfaei
M2+UNjSujyMtUHAQzNCizpbUy87aMPozAYneyXDVLuQGzEaZqb0LDgblJtAE6er8
vhoatYFRQuvn0LSy2SNmPx8fsFENmPqf/jvQY+nCFmYVuyYN7mpV+KD4EGm/LUOv
9BSbhqXbB1C8Q/HeHQkewiHSUw4BAG5Q3QRyUfS/z6OHUUaOSVrZNnelYGF7S/oD
CG4rzgTyEHptnQFBP11qlGsh8N942Ji3YdnHd+yQO9pr1ycJb4sqEszszy4l2fJl
s7ot2TD66sWIqsRYL16QiFn92aC8LAnwm+Z93nMrvb4YCzNYPWDazE5RGsnlxwFd
9iTWlM5/103ygOX+LMPao3jWMTIaJejRz3cmBzRtX50d5z2Yz/beL/Xi3tX45nyv
XCh624BNOqeZC6FX2osTKJT+h26O4WVkypR0xv8Hjsv9x9cCxznLym+8W4g0hvsC
ulCfAX316/j7Fs/8JxsHKX4zMCwmpLFaRq7KPxtfWav1mqii4h+ORTL9ydFPB4No
5QKuWEavkVn9Gs0w+enlAlc51drFBx/sGU87AYFWjWQSul7dh4xS842ylqloZ34s
JW+4OlNDSnrpIzx8qJo/lpw8PQzRAQki/Bdm+FZn+IGuZAdDs41TLGdCYthQ5Rev
y2LvtzUlgdAE/xcSZKjM2jXP38Ta6lJjl2vo7qw2gYAOchiHQL+y8QbZebi40GHH
gCRwRVSEF5Z+mZmfw6soCUGAXXMRtg/G9gQjQV1hIkJk4MF/yYANo0QG1Ubpdf3Z
fFbgVo0CrLncBmdQTb2tbiiQYIMDQioPR9WwoV0tQ3fleIo881mHURaY9m0rS+lz
0qusAx6vrTmKFhy2MD3PObDf/3a74UTpMvcJIfXo4IiAz3GHeDOX4DnVd/1DaC38
0ic/B3S+RbAx3+X1LzTA8+/p6R6+QMkSfPPJ/qNzfWHiSGIwInxc5NOOsZ5Gk7eO
wDC+csk7ZwxIdPWpKOg1Z5CTuZQkM0ZHLuitB+qFDbVoz7Ps3vlpvGj02APtFCPQ
rAc+rtqti+9glBKDCMNJTdxPVvRUkrkLCnEDxaxFLkOzQRm1QE20rzmpy4kyxdUc
GvyYB70VO1HGytDpf+fOknLrCUNJEtTvprEJxWmUP5NNwc19tvtKd1BMtmxwPmxM
YFCSIv/CgaoCCTLW4HeZHSQgAd3HsMD3liiDRNIuXxKrdgLfWW/sv/nORPn39pvf
BpQ2E93EWS8Yxu+p3FYhrupAUAuWscj1tTsef7VayvIX/XRMzyednrehUYcZo+Wy
G5tr8Wvid3DivsvvbueXqClwAON5jQCKkiUlzfh2Q12R+dnuxzYoUmT4uLLAtcPE
ib90nFqqVx3JLlhJbSDr8OVUR2pT/ic89Fo/t8JhedQDXZNWMHdcV650XSmuY/In
D9oc0t/tkwoqgw5GRZltBtQ+gg7oUd/dsraRVCyFoajKne6UtbA7u1/1Z4w2k+CR
Azk1sjWyQJf/gJ1oRhjwuzq6c0xc5BzHL3Wndg9MSBu3/hxD+IOR5KFrrrnkq0Sz
bmBSupfKidnYKW1K52OvgBcy0TqU2L9acjTOSVyPyB1WyUc37C/RXGbjsLnAMOWF
waHQNamSLX7M21cPRZvoMO0VdWFj4nUNKEfAOJsW1Vuf+VHaEJuG37X+EFf9jyI3
siYLA4Gf6gtUgYeiF+MU8pEytIMods0WA376hapN+rN7o9SqS7lVoaI1LaWugWA8
nE3AhzgyXcU8V3J60w8iIoHZe5xOC6ckdTwg3UEUWLqVEjBmntZeRQ/LRdnY7hou
v75pnX4XZriwu4Hgu+bisFRuRKtD6FmfAg7ziYHK9/tcDagFR0AnbGDoEsk80Tdy
dfK6dLDWLeGOvHfpSf+/LZavoCqLLyYWjn3NHLXxGB4RvHPm8C+aCMmSaUNihI1r
wAu5edHscnF/fGCdf5YPmW3q2ELoMMD1vYWI8gz1jfSA/pVslQ7MMFVtvE7rfY8H
Wt44W4SStYWbw49xSwSZSS5rvHyYzNNeThxU6wCXbtEuwDowcIEOwrZexoUivAfW
87T5a2IDjlEushjkW3olrDzebcnljlZPrE5J2fsEBmHUNVAPnvfL6d7R7KHDa+uE
1hv4Xtio4GTiBpdFSfNXui0nAqwa7DTy2r//I32TqUXhglhfuqXg6ja0AGMh/ZVU
4mRTuIFMBn8NEOhBteo9NvQaz+9EBubo5NNm6ajepxhmNq92tLPs2EOD1tX4HUw2
Zho/40D50fc+Ll4Po+XNZJxBldH300zNLrZeltXH99p2gphGHmgXjsfGR1lAewh+
5yl4atV0n/4J6XkaTPwFmRtxTqSOIeZW41tcsAhvC/903QsFb50TOsOr7vbJitHL
BojeYly8oFA52T4uOEkVNLuSGsTxn6RBrpXZOIakbUmwLtVURJy3jyxCddP1JP2Y
rsGnV3bwlgn3No5m/wu7G5ADO0OwKGxvo4haTXrrRpdjvHFv9diCMykzk1Nefjm7
ktag7C0BRoVvSGHgT2W5U2qbKv5Mx7Kgxy+s9wYAmH8uRj1hqFFop7pJZbjI50xh
cPx7hAVqNAy5KmbRxhoe6RDIDJEuIipkHEzaTcUEVNRBx9cCcYAwT+Wr5Qc0Quzu
9ePcGTmLDdhpIBsiQJCgiL88Q0MvTtUuLOgkWyhtCdcvx5h9oLfblWybW/ACLQaZ
A4vUg8zJO5Pn72x1DyJlzTtc4HFHZ56rihPadsFr6gVuFSV97uPxbHLCeSqeO5V5
77ZAXBrTWQonjIYnVdu8hHjY5wWp9FKa6VirTOld3/xooWjcubeTWiSee+C8cJrj
jTvf8ka5DXZnP6Bvh4eJcqS3NbOZJvESdknaprr99W212IvKr5w+5kpxuQ7sc0if
HGtqTrKjzQ3zvGHWP9OQ4a1thEcm09/7DVtToPo0uQY0o3vw1QqfmekqiHpq3jvY
AIbuzlDHlBQgMLG/rcEKUa+seU0u1GR7Qwv/AGKr0mpG+8Mrz9D2NgaiooG+cxy2
UEqCDat8x7xwF+hC2NcrCqcDUH0RyRT9OnO3ffh6ScTQA3J1SUc/M+RoMQObvAUd
K3V22QXVSNCRZqjBkyBuexkkwnIL67u02fhsw6XdQENDyK+4znpxV+530RvbqWMu
`pragma protect end_protected
