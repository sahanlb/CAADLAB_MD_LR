-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Gk5NfgMtrWFaq7s26og8HU2IA8xyP5BwxNIHX5c1K8E3bapDeS2KOd/rJwP/2Vud
7eHlqbb8Ak+A6QuSUnBW0hIPk1vWSM+0JH7DyRkQ5MLtRjz86bYGSawwWNFv3a0n
kAdFT7F8oYnfX7fHaoChFwZ+gJ/mkMqsYhGB/vvH7fI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5712)
`protect data_block
sgJ3+8YKKQr5HHTpHZt61xwCuqAJYTyktMOvsgZ8Uwz7+CI1HSDbL7tRCZm74ae3
W/zmAj9IQGQjn7ZXpLghr56ab39z+H7LNj2LbEQOOTLYa6q1yFEDzLnokr2llt7i
FZg0/TcqdUigfJAAK2oDfFQ2e2+mr8ttF8L1hTAWWoLjDgBnNVkhp0DWU7l0eLBS
XUGmhkNxJmEk/wZ06C+QbXOuFAoA3aJ4/w6PcrwlWYIGH/2/uRB99a5+ty7I9rhN
nRzEnfi6yPU84AiEAwc6weU1DJRNrvY1qgCz0L/11nTY5TYQn4Czfan3U7hiF3AR
LtcTS6EaPEV8iUpApb1Q91KNxWgzVy4V8ttZhMY9uP6AqkEBXkOigJ8mi0rM5Edf
AX5SYruSCy52DODAoIjxSgHSXDLtgIEGokBogoKrsYprR03Olb0zTB73ZEXqhEdh
9O1QFchhwd/tJAm3h+JClfgO66ZtWedVjNjaqe4AabUjYKRa91cU49PbaEwuQz0s
3kF3saACByqh+fgRJDgmu+qtva/zpI+fVdDqbJNRR70pXEwCnSdepOwEuAMXHaRj
SHT0Hl1Pw/QgIrzku2BoyRgY8FB2IQK1pSaEeK/qKeQX06KdWMg7TL/4RdN3U0rJ
SbauX9ZCldx812AMYU+g4wPC74nSa1J3/W3Rn54GFCRzp4Fh67gq4CQ034c0Y2xV
ya3rPgBdKCrY/CkBsuCg5ZnnOVzZ8/bcI44uQVZ7sw7sAkVPgaWrf7TReGNaipBv
vnq8FZwnxfz8liV9wOyapsllhf8j0x/oURSlm78obkWQirp9od8kmTpBDDPkSJ6L
Bf+sxtAgRuhPEARYdsMU/5kQ0X+0+8mygctw0QFmduOfHguAKS159nAVjeFKGsEg
UkEfLaOzYtAWhUiPsCAVMJV8rog0DF40DA1fOOs1R7xmJMo3+2CEawaUmRtG6FYp
B56WAEXUs+45y4mEB4joh0wFpv8O42iuPtJDgW4DwgH7uhHrpimhPAMT8ErcayY4
XyN9MhQyWIeZJQjdChj8ohC59vDE+hTz/Kc9xK9u6qAOim5jmj7j9jz93c7jW4fm
S8EJl1JsbHifQ5iyPPyxyOkuKRW6Pz5IpaR73/mi80QYtOLQFzenGSrySFu3jZMR
y2vLBtBCBrIt34xBhXpxsgtg06JuKsoyaqXft7T2N5fv6HHTdEf8L5T9eTWXU/N2
LNFPaL0Xvg5InMZ9w9JQOv7nieN4mTr9qtoAMaHhHH7LuZF4ViTO3WFT0792Wt8b
om7It+Kt4prWS2yfs5zkjBajyfBrzCv38idtHmwT4LH4X0KXeJhGh4oxy8W9XCMA
Km16QR0sdYeGaXAbDTD25aEXD4CpWjOJKclRtClHsaxkDo1r0MzMGEByl/azvbJL
CdkgrQRkYZ4BisdNwFr+6QNYkmiRI62XLExD5puvr2M/cixQCu2/lxm/unGK3hiK
DrvDgnlwcRrxImTzJg9CGkWTTBKKixlma+BTOgFqX57Pq+OCzmpLDxXht5DXRdBo
7xcpCG03X4gOEd1lcPg2/2R678vquZSmDD7yRSL8pfamx0JGtNwX5gSQYJXLiSPG
I76dAKOgqwnk+9iiRFe6AFY/+YuQIzvOiy9gE/scbkIi31CHJkDEZaRXRvvEADtN
7rGgHgTijWTVdtoyA5tFHccaCLgxr+4isA6mzsIAUy8Tj2afm21Vp/rOwXs2JYOe
4x1qqXAlyqimZTzNpZ7sqp+VTBMY6htaezSJuCvyCRihSENbnEyKwoAnrcuN225n
4ZhyLHGAmUmHLZjMB9nPNTbaq90xLY7o7dQ9Cbea3FphO6eXrV0MsHZFMSL1/G+w
9vSwBbSBlrnmEiTaBPUVVVWwfQ04Z/Vgb2+a5Ufq4NhIoqFFb7eLf6olBTG0oG/2
ylJS+TgtyOOVg2eWKwUneFuCeBJJSBG8muHDmVdpY2B6fv+pQCvUwDQ01L1yB5nY
MDStcd8MkGSx8YVXM57YNBXM7MbDJMkNsltj4xPhFNUpj9Zolg9bPTOEMJH9C5ln
1O785+ZtScDO7c60svP1eCcZxLej2EWkrv/CD97qi6QLk16OfmWfLBFDicJrmmSQ
E2ULD4Qe5Ai/9VJmFWQD1JInxg9gveibh5wgiDvWGDEXeSbdSQZ2APQ+l8jQuywc
Fv9U2BbvOVNWEtu1AXGKBhEv2vpRsZkUiVyk1XJIa2RBXG5uatVO6LRBNEd6a8U3
PTRVJSzNfpDSlj9ziUIlHMLbb6UTlSILY4jKftkZ8z4t/5JjLxs0HzMh5VChId5w
Z+n1VJOmNE3FTrPM90vsnb7JNI7Fjno+Vxhw5vuz8yAKln5EzHxcothTDKZW9vS3
uvj4yUGJk5rgOzF7UvHPOUbqHzf+UMvZyDu/Mqf0sbs3n3R2B38LRcdMptOG7OZd
7VFpizIWlZlr7j7qai4byEdyf8S8FckyP3WqD//yDoNdtBuWNmqRb3D9YnmrSs+T
XJNn+cGoWeGMK2QE3suYF4m5a4/A+aJWPMhkbYZmxw1g4c5PleKZ/z6/CmAMba6w
RE3W+jkQ/4VtYQCWGM0vjMfDq2gdqfwNt5/zykJ/8/nzUIBtOz1X4aTEgM1magvZ
Uv7eThbvJukaxJ1cmVtk/UFMoPnC4RKfohDl8dNy1cQLz2HZf+r4IreAd4F39g5n
udY/3NzJin2bmj5PLRsEMn71TjwAnLvBUKV87SlQF1elMxscymPMezKJp+XC8t6A
W6Sm6R8IwGbgtK3DL22TdRpbEwb3h7e0ZhgDQ6CzXtqv0ctiK/+rrN/DFTRuVjUU
HXzMZpBDKMcMVGFEalYoeNs+tEyo+7PdSGka6hovYahJWpbQfOtn2faHND1YbG5o
vasQSDBW2Kdv/ascuQTjwXA/0bIvCzNnVyF5Qg2MUuP6Y3ZCZZ3d+ELyzhKAT63G
dTcY/KoJLlwf5vhojZxRwJgxT8nDTwwtpYCLxBa9AJo9fa7K96qIGoi8UJEK80/4
sEJ/nNx1mItZ7pKa6NQDYHfHJBjobq0uhzIyCYAK8NNW+EYjkBWHjNmgU3TCwawp
hHLanCYyclsLC6nq12akk38Rp9cbHcJDiNk/MZ6AQccJSwfLuvE6IRJemuiPEILt
9gKLZZOsKiEx9nvCinX/ecAusdFhof8ADfqbtScyGTc7HTrRyZ46VhJZXc79cPhi
gyTSj/ZCpslGTeNWvme0TT2PVyHALT+dZknA26Lja0qJz6Ms6PerSuOHas6QeUE1
zb+BZmYkqlzIY3QgUMX2kZg3YMQWcVJj66+2aI9qrgIsc1F8viVfO/r+3a8Ow1pi
AtaVCjDWfjh8AuA7ze+1D/kteUYhBb/YwD+spYE3f8iXiqlCjKvnnUSjYJY5Z/gB
Hw6joFYv/OoG1W5BE/3a4OBDFePGa2aosj7eekg5PVw9S6YEb1NNFH+ux+5JXaKB
8bT+909sBkUTYGRpcJGc5jIkJZrqsxiry7hNW1d5j9g6124Lc+pzCpd2AzKfApgm
7rtwz40koi5yNWOFXy+BUMtT1EOFXANRtmzbbUSy9YjEdLH3CYMZxjC+ZDbNYqJ8
uLGSzIrrNndPiMxZWnxG4m3NwXYtSxCkAbri20TVLS4w7BA3Vbu1Rd88+7Sui5tA
ClZCwm65FN40qLnEsWGu+vgeOvGuhPgbewfOn5kKMSdYBEgCRs0F1pOVXVo67aKH
AL729Y68jj2AuCYFwsZiBTOSPaEJ2YBgBtRi64s9vJLCLbZmjs0EMkw8l+6WU1/H
Unso6EkwVMAOc5RAsYoQZXF+7qe6g14VS6VOZxTvobm5UpBtefwTFWrp0qmoISY3
ZPgsjRC1AQpIevCG1alXzGylAVUYpUKMpX0X2v+byv5Wbt/CJeJMJY+lbhFibKbw
w3lIWv9WY7VGk4BYmAHo7hJjvHsKtmTG2Ocha2iSKbBlVpKAHafmG2UoiQgfKnEV
hlIvP+pqZzoLLIFHVQp5OfnjmX+vLlPBBunLeMRJ689FQ5uUfXA8rFJEKAgbXm+R
a71DxRRaMyhD0G8BdJk2JmGIeEnhQgHv9yp7vVq+hCqeT08xHnErpCb2olAXK0aO
She8LYvP5tNDk6V7LX6TQkQoXidS5rsjxZnDDfh0obKcESD1wpoJkKzfCNUf+MgS
xKEIPidW8WhEUkFadxevxayZOCBHmzB/ecW60i7P5zUjxCgupy51zCC9VaBrE3RL
AHj17te/2/vKzTAy6DbRYKN0C5BC+ktYiVnZOzDHkbTuNdxBJ3X69M8oljXn3OoP
vttd4Yvu8RXBusuX0b7HkElxXM5APxURzvfsOCs1XdNh2rD94UMtzE3DOEeo9zoJ
qXF90p4nJGOxqUiuDPBwIixg5mddbO8EzK99wF89vaOJnUGMbwjoxFaIOOlkdZFc
fw/dachFJjzlNxiTbnZx+/PMzsxAELuSWqudqQwUkY61R6K7X9gb+++4QNuqQGRO
bnYbO7crq8TXz6q0TtErnLG0ngSpq1vxav++lWdU06Vw4q1KuXqK0p3aZPYsY6um
EzZzK6JpjrHQvEZhztdc+LnzaQlcrIRL/DFdogB3Nbcj1tDEoZMlAUhvaBULu9wj
nziRDPCDpPvE9DNLPrD/l1sAZ/DY2q9VI6JEJWu52JHeN6VXjOGEFDhNpWz0BKuH
eJMA4UOBb+12e6ry4Xiu/SQIjvPUrqwco8pVWnr5mJ+F5mnOt53wQPWLsHzRu4yE
/2NBp4802hkgzYJXhfJ1GJ6zivBbQisMbSkHpJPWkGEPrUiiCjHJutCMPmQZmHHg
7tyRK65shmCviVbDyQm4dbxgIPUrG8JkidBAQyqamQVh9usEgd41MctlRh8RdCWu
y5eS+HhwqQ/umwnEfSd84lymgfV93L1PZqJqSOOakYMuvSm6R2ulAQ/XNtykUe3O
q0WflpqUzXNDAnTmo+q4qBNLtQKfWplUCRehKfCayFx4rw8T96fGSFOZwPASLiy4
hqsLazRLYVsJ9M77MJVnus7TgnlU9vVIDvxz3tCEipya/Q43MV6WR6osCisUTZ8h
XwYIXBNkDLUtuUGbDWWDqXHEo/S3FWTbigjS3QGjxoTBM68rXDpENOuFNlVB3tey
vwtVBfRtRkAlChzd1bdErq0jFDn13r7HrqSOUBlOgPJPKEPMuHjSvC4RUiiWS9QW
rUywy6qaAg96eDu47vd76lAKcZuI3Haut2Fs/QHRmto85OrGISx5S6iTxVYfNPgW
AaZbH5cBjtqsDFFaFQwNmKtk2pADqcqWsqQwXfT50k22S6dZYJkdrMG7RtljL+2M
yi9s4+d9btdvM1g0wId5LBZEpalbvXS3PPLHnCKScykKZISa9t5T1Io+e/nzrRz7
cHsQVxNpx1+P1op11sDT01aZ5YxXi8WWf8I6TNUJo53plsLU1iwQwDwFN1F86MQ5
DVdbj1mhaMgOcUQ/UDQqQ7Qpgq7xKo1KmhZMQuoV1ZJY0b0NvHiNRqNjdU9Ata1N
BEat0KXqregG/RYixk8gBb7aJVAWwx7v36Qfo11zNiBnrDeY2EEhygpMWrfgqDDc
1beUsqZt1STN687I6SOsBxmkuqXAPZHXUXs6q0YUMBKsCaT01nFtKADLD85kEpj6
qBVdUJ6CWtvKUWFYBWMRng4Vjq/BwJY9eRwETaYbZaHtIyvOwXa4M7lhUv7otVgN
bCGLcCJfh8v7eoaya2dDIAH2ncpmmxA4n5VF/UsGqZbbrDGqcwMryi+5Y2+lVl4q
lYKOETSyZw4djPXVhZnI5Xc/2sx+1dGVorYSbZeDns3M9t5xpu6+xQ+VREmky1eT
KTBLc8zraZ+gMH1yvEzEh6V2usv7RAQweH/KHab0QVPg1RevkUNfOz70mCwcBYLJ
+FDCJATzz4ofilmdID9O4SPWw1a9Gbr8o/2o0P/3iOxf1RJCalCif7u56I9ZSRNi
Wxbj3jpZWeHqzAs/fBxeU1Z0YU7oSrV3wXUjc9GmSJaJPITqiWjQCHPiHV1rnrae
LG884blOZ1I0pbhHcAixm+DfzHm/OraOlXrBzalYDF8Q5J4So8Il2uJ+3/mrYHtX
0A8zcgWF9HJoKIWvj77OppqxDX0er+wZg833lK6b32bJOqjj5DIk8qdVHjEPFGk0
TqvyQjMUvC3OltCDUGmXVS1NmsKZwtS1Y/vHFnCifQezr6uvaJal/PBQh7A4hLaU
CaJ1GON+64fFuVSr8INe5yODDVzz/qi8BP3Tuhdj2LsT5IjmfOaN53jULen+HlCo
BOz2aod/wS2/LfHprwZl+RrcU/h1zEzCI/UinNgg1zOlOyryPNmKnYG15xiWkQZu
+Tnkp0ov8um7LFM8wHV3gb9WE2enR9FDgG1P9pmqUvFoSodMylosuwvVYFVDDche
ZZEtue+IXWCJYkFIeu0aFP0M7P0XfwY6SQDyJvWFMMvUNc3W0+MdPbWPau/KzHes
Iwt2AMqlf0gaz76vdSNhU11KIfEipTTeUHf/XBq9MwiQwOyLzqmwPR8Dke5rGtjz
N5+oyeSMVk3Gcs2Jyx23gNNtkpHAcm9G55SsHfze202LUsgt+1hz9m362YrWOY46
OKRnwxEwFBQR5l28ciz1ygUSSdrGia3I+mG62yu+xYrbx11BkzvuG3xUgjAQaoNh
Ap8rkiKCJqsc2jQUBmGmyKt/GoRwnIoQ7jSiLAZ4EVuo6GAzPh8XeEBBifOc6Q3W
DT2no/e4A31cdUyfxDRgILJC3pL4Z5q1dTAIGMsEQiklKRAX/FLcpoBFJp0Xz5ey
5o38LDLSb5L+paXUkJd+gkMFRzszaouIaCVP0xGLycZQofKvOWeGFB7a5Uo0cdzT
rLMVnqE8Rip6L1TIfCACUwAeHf+3RRJVpvT9iu0dWcOp8AmCcPecQfd1WsuETgUp
7lU/DPfHW3xZYciHkLK3ss7xokQyilma3OBPboKgwFiHXGq+aNxv2jg2+/yvPqti
QcpLOXFtUSvI995oULjgW08SkcnP39JxskXnAjRbudNXS0DMHmB3tVNMNuBWnomF
1dJOX5jMEZ9RxTFQt8g3b+E4lp+N/08tDPnSu2Zlvf22QD2CpONjlHC4fbZiTTgH
vX7aha5AT+WSnZgJmxqAsgdTlt5C33efL0Yh9JqUH2WAVLP4ivcmtQXi7I8qVgW4
PMUKsRY8NbiubXQSXWfCIvNfjQuC97mh/YRAQwv+wSFHcutNZpL1xZQu+39anpbS
dhpd7o1aUD8Wq7WHbNniPzEMumJ4ebwUugq1J80Vtbkka95QafKyAtVPxr2yaedR
7NZNqf5Uv0Xj9BZHqYx35cCgL/B7m6AqX8BLr+V+No0Pr4IdwN7cp0b0B4iVbPlt
Bc83JQObLRTqMtdwbgsD+PTfPPS/unqOZAhYU6Jd03zU7wE2LX41t6btWQiz9IDX
Vhmz+o1cvDDHRo67kk2Y8fkFi91r4aGdOpUSp9B2b3+rJxeApYamH8dcVhBT+w0n
Mx23wtbnGkV6JDeNPBcMIwK7R7BlRQ7BgeluWjLIaF6rDc/incYg1hT1sGACPp7J
z8+bIhs3aCrGA+zCLJAeAvU5h9mwVLaOV+W8ruGs2O/MLrXKMEb9XwFTGYuiA7SZ
`protect end_protected
