-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
T3qC0rftmZ6K/N61SQ/oabjMfuPPPGzUTxi88KmJxExWuDss0nQX147QsqVqtERo
tVoRx+sEtk9IcJGBxTMhhlVjOVRmYknvcX8y90d9rrmVbHozXF4W+HGbDfLNfgSl
S4Sap6j/T6K1De2ozLfvb+1+BZKWq1yWj8bM/u9zJZ4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 81678)

`protect DATA_BLOCK
ueCJdG6FXIaD7UTAlp4G9fTsHTJXENeo/8sUYY6HZkx04ncx0D6aGQknzP7imRWH
kGnFivpKWKpZzC8A3I/xofwi23u+6E0bTNF10h7BlBQ3q846LEIjbMqg0Mw53X32
ewZZ5a4ei0+cmfkdkWPv5X8/9eepW6SXvs3W7k9QS9wls1yYqFgCmXL1kd2Plpn3
ZwGqb0WMAPktPxjd5VVrMgWpe/Ypyl46nKuabWm/mLfMlYZaXp97jai+rrpj5iB8
lqncw63auwQMuQevV6es0iiieLE4er6SYCAw4ghXe//iUUHrXdIbl7XE8mV5kk1V
Gk0xDf+TF3ZOiG1qR7cQVIlrXC7HP1GoxMc6Xh1+lUZS06icZJF5ipBWWxUwZ4UI
YP8+4Xz9wGQ3FKMRkglm2VHhdpgQ8Pb+xDkQmqQtz9f8fjpriWEcqofOH8mZJh0H
y6rQhmC3wHg17XrwCUJK0r+84jLfPkb0bHF9b4nBxyaGlxaWSVbmCJpWFIT0j8Q8
gjbqKLCdQix60w+gNAo60p8FdbNuZma4GdljltyZSdxZwWbPM9cKvHMg5KJ2sP6A
PkjmH/ElqGqWQhGnvgOpUCUc7R+w51pun2ZQe9avpCrxZqLNsPJq1dMjzzpsU6kl
u9OeaB2TiCAaA8j4qSasdVBJOpkPlYZHqRzcmnAwj3hSeGKobH7yEp715PoE5/1H
2GcmeO2Z87gDCD8TKanMmkf+/gJ6v80qRvkn8stN18ZwBTzREVxUS4V55v+6gNSk
8zx8HMcFtuNs8QRlQQps309dbG8WgbVjojzv42KZa68Er7zGzi5gp+Id4LK6qU0R
B/hLgx6Y8tHxvO5z9W7vT8M9oRaQOACV9rFuAMHJWqd+JMG6tPFEdukl+dMOV8V5
5VRcSWEvtOXWJQkdJRULqNHZ2DlcpwlskXU2lqXa2SQHTacbK5Clri4DVqx4ISaf
F3fzwNQst95xB+REMTmyy78PbfHtqNfqdpgHy+Zydmy9k4XoXw5wxWwobqRq3UqG
dIaVv416/yno4+xkw/1tNj2xY6uAbNNZWLLZbLogxMUnnYar/YCQGKoAHOvHSQ7R
0Donq+GFIBcNPcAak3RiGkMHkFKgoQqMb867vxj+PgUPp/2YYrvvFDiGYryMV1Nx
hBHpWWiaxHdU9b3shSGeVSI9Z95VPbN+LF8ePnL5mKrAzc9GamZa3c3agNUlSSqI
wVB4cRoywAFueZVVG8JJaHgaK2P/t8yHfQOdnH+uqtAQvuNdNXuYtNd+jIQSrtmn
JQsaEPQi8gw9hCcDWqcvZFzmrzuqa4CLj+ZJrpmZ4OAvbQOV8kxWUbBQn4XvPwov
mGPs5UEW4rxzXhl3ru78CGe7Uyr9L8SqhK+eYZmhbk+G9Z5E+eEWZjqtxbmy0N2O
yHfZ9IH+HAMQOl0xtrRw0CxNTt8Xk2yTV6RrFXu9PRjDioI+/UsMW3oFnRXpRLG+
A3I5Jhj6UOEupnzHy8vt1Ios7F5K+kxauGn2+iBfKdc5YLS91bRdbjJHBCzID+gz
oNXDaFairxL9YiF0r1UCkTRV56zp8RB28edjiIBQFxCScajhDdszwsr5BoDGS0xg
w4hwubPt9F3h7XeYq0NUYIFHSEwuKN/mcHl3NFMwBuTA8ZdzLsdYWbYgUBGMTg/i
l35P2qROkLTA5bG0+wb6+h6bgwczM5MZuE4KeukCENsQIIv7lbbWQYTAsi6JRxx9
8QzLKq9YBzQDD7h3Y5YGlA+0OwQ2aRLYCpBsjpjg2sv979MkBQ6uZU5t5rRNb5vg
wqGFNE+YYxLhS05I4/c5sKPrgy+zcW6jAqitcp6OV1/65bsehV7zZLLCZlt9qYCh
rg0oeJwSNBGLl0tXEeo9rLleMEAym+NsfSMF8n8/QpUQBNhh8VmbOtK6jXBUw3zF
5cC+mN0Q+X1JsKMW4IL/f5h0cgEAu62oqwWTHWiE/x4yo0ucMk+lvOYj2i6bMlCb
4vd6/WKVcTcGcKutcON4yFpB1kQfXlaz8MC33BPZDE7IaQEePqckfjQW48wnsj5V
l9dcN9/O/FNETA0zRGuZLe2AbnICCB7tOcDYdqq+VsI0JuS6PTJScFwfrET/4h/e
6wIhYoCOtPhOAqzr8M6n4Qk25Y67HTIZDsgi9bVHoa7wH5qt5U5HZtr9AmaN1bSK
UnZwVERBYC7mBWXrYSxcie53aMFFDs4HAn7hsLbNium8yi7KfmtjwNYLyo0WMetF
17DUT+SygzLKg37SHMCta5NJVHXeusjCB4H1qodvMjGKISNL0VYkoPjDY6iukf3N
lD5TiGuMgvJUAI297mPKLped220pUNtqnuZQDppmrIVZmp5Uez8O+du0boWWxRGp
efyHI0U0aYy0erQ2FqLIT+kntzEP084dDaVm2u9AjqvMnOaylwn1NgoLkgcY2z2F
nFzOVPa8eIhOgPg+q7qZUqerNsRpiftTKGaTBmySCnXazoc8Oo4c4iJehJ+PzlWW
LS85MPNhQ+sUdAA5vyBOmireRU49zYLcb5s8rSPn0+s7REYESBJ7qnF2JvWNNPCz
gFDbqjJj6RwdZajQwFH4QoWG2D1eZp9KdGJrc1JXj/d63ZXVa+hYyatQOzqxbAzu
EgVdhC8nO8Al2v2toWojoJkbSWG7lD9phBeFEV+ve1v6pYZ8NEdZC/1nXWFjk99Q
DV9izbLP0T13ONMHCp/uqZTMJAum745UIu5cdO4QKg0zFVNx61pRlV0TBm+jcIXz
jlpU8vFuNaJClGrnr/YF+hPmD4R6LRPIfyqicKz7DMdopIqfS4nbh+QIa6Luy5rh
yGcLvyedv96HqVx3wum6RDSdtvbhAEzjqQVq7c5+2JOMmyhEXChMxxpRhwkhwcxf
OlthUZbp+ytyHox4yaejq/Tn+mvQuHBWYKmbPmBN9RPZLcplYRPCzIhqSwpGZJAz
gg7Xx54kEcHmmKnB1FWjjoYcibsJT3Z7AofnwQKHqG+FFUkvTcOwViFPo7+GClLw
3SFI61koIRnX++yuOZa1LpI6NJPK2kZn6GcP5GcMRGnUmVbls61yGzABNgaiA/RA
Up/RiCCbSifGx5z7K8rO1CUX2XRrDKZvuJ7RpH2weGVImuUi40JyxATlCrOzRjck
ygW18K3i4yIym7vLZ0MqwnYKzwFTXVnuNk3lYyod9LLAIvr62o0gGry56HJFO5GO
l4bDTUUQRMDZEWV4Uh+wZGSToagF5aBgAvQ3Xsq051ouZjAZOJXBIpIVOAuGR3LI
JmtGWE0kSaFs2ToT/u5ZIFJjKKpLSMjAtnuqcNq/wLh1RdcfVAYI2ZRdjOqpqhST
XC/i9h2hvaC/JlJWIm0RjSZi4SVjFss76xDHy60zuIYa7JwPivYUnVmxJBofbtTO
3Xk2c2ZmvzWy7UuqBFYrEmGnXmmdLMcL5pL1aA85Wgt+A3lyyKhNqFE3gww4AcEg
t1vy2c4rA9XtloTNIxHksopAHJpGF691bYbKKVWglhaa4surdZCDofmzedWZ+0pg
c9bs8645dQKKzvYB8Qm1VpBynvqLvvKclauC3LUivkagfw5rgof0rcKFtxRVI15l
5Ev/bNeOY8dmNH/nI+tqX34Ez/tDsZVx3lA+DknsEI2/lcZjAn3yc5ekSHker2cM
A52N6FjFFbMH2Vp3O41KbAcCZic/kXYtOfa9sTJMcrrbyEGyFX7PsPG5qf3lfKYD
PoCK5GI2O+eXtAQWAQgEj3pIrJFUAfmI4B0FouhDuF6zlioWCmmnC0BCTUAU0wX/
rkF/ocUYCjVZoAwA9PVutlvYbvlYoy1maPCsAdg+mY9p4pRF2rHcZQKc21IuC+qI
HCvju9UZ8/hgFqeLsYhfwx2vFK5Kiu1tPyC29UKJMoHw8y8cgOikTGQ6yzRaMKwp
MeMMwfK7tKHRiRrmWwDUEfEci889CcxoKlX5Xjulq4xJb5DYRSmoKPd/Ed/0qajy
YAT7lFFh7UF5eBErDs++RIk7L17B3EvH8wyXD3wgqdqTqOuCM/zVyLW2hVna07RU
nEiv8OpKPudpMLM6qZcsDgbInEZtCC1zf+756jcChw0+Y7E6PjMakxu44kSeAjto
HwjJQeC0urJY0RA+kYm9IzC5c/94RFJqTjl4ovZbYS1MnZl3rIOoIJNYAw9lFL6j
MLUY67NL2MazFg/zFCtGD1HSVop+lTLDGFgDoyFUrqu4D4y6O3lgqYVzQPPO15fK
IZ1Vo4r0rGe3Ri8HAMwx4VRT78035xi3fuTD7OHFliNFD8LOY0kZGoQKpTChRel5
yCk49uu7rVb7gr/8psOCmTYWfjEITmKwFSrpPFQoB7m2bBw5OYs60pR18mec4tbK
OPoGLhGmY4OLBicIymxbIKf4/L+p/9MNmdCjQDAqXL8RRzQb/0f3fg8e/JP+gPm+
zeMb6WzB24aIV9UjlCg8qLoryiV7taWiKGtaTWRc00EPBsuXq0E13R8KTqMngJ8W
y/rbDI2xTFp7uJV1KnR27PSjK5LBJUNbFZDz5zr3T+ze6FNUjth5Oh8INSMckj5/
ANNgMkuYDHIpdlFBhwj17YFXdN6KcDYRd3pcFrgxR5qtvPsMLsRMWLTMMTgNfBKJ
23VAXo4F+IDXTVn3NGkc1aGm1vbzt42737gRE4j+SAJxOYLH0BEBE5tG+1ldSCoh
VupqjUPWRsx48ke+rFo1L20mpQAMNRAwf6r8pA3QDSQUWQrBaHAepZ6UJ8sqTpae
X4yIC03prI0KUwtYwGuV5+8EZdrvFFCGeimJuU1fbi251KcSYe+xYv3RngUB9lCZ
RRydf7WTjnKt5OO7vDvobSrVTO1xMq5YAKDTKAhQwbFozJCbh6+TJJxUJvxnNwUM
OJbanjx22MwsrusIDj6QApoCcqF3TniUdH+fhXuKWG0t5wkFsc/oRrWgZc5lzU69
pURq2ZIBNDVnlXpefzlE1/jwk6pXL2fSOjvZ2TULZ6CkXGqdLFnzeGTvJnA7SUfI
1rS2Qw6pDFFciKzF65VypgkKRuMmOLzBzmA/uCOElFUwNt0RX8Z03TbBhiwyBcrf
XKGDAJnWE+ZNNY2nZ11dM5O5uK0HDczEFWg4asW50p1/7Svqo912DEDw6uds56Di
dfl9RLlVZCOIvzjxvNa2XxQs0Z65yobIzUU4RGylNLc39UGI6K4vdngdgnffAhVr
agF+Hd/YW3fR94NbIJXBZfKe85G4ClPcy4qkHyeExhi/xYH2w2Um/9TlqrDHWWOH
Ha1dqq91t53Onr3zPI0MP2inO8AcCxt8QBFNmmBNh9B9kpLdpeMovkd9xfXDF13E
pqwcjBhZuunwGNRRNyKwtLuYK35V/LEoN6WxhTR/i73xgInsR0xna/4JZIHoWpAP
KPDbqFe3XhsJiMQ1D/Gcd5yQmc//DtZqRzQAOS16kkyX0wqDRrNHKU3B9PWsVoz5
g/GZNNyH0Rv67HWMGckpsQUh40/q/vyBuNrRfEzAiF9g9m8WBPGCfBVeK2m9rVlk
5zUfwH4BQUELJJH4xAfqwoukNT3Ll34cYIakJP7RO/4Cbl1LdUrPG5P0VrQrlW6r
zH3xxZNAt+XPwor8SCMvHCIwQ1Oy6PFvKFs7elNF4oH0cIDPsWjo+ykdXeVVbfK4
pxnTvD03W+K4OfT9yd0TgnEPy7fEYE30p2ClNDha3weIj5qxgXZS3/umACd/g3lp
w49ALNlA9hE5TqtZPQp1NA5KPfh/H2y77wUUG3LWL1mb0VeJizLwCUdntGzccjIw
SG892xYARY2osPhpoIxGK55dKhsOMr49dVhqQEQ+vYTbGUcMc2PtLr0mm6sMxnKS
NTLqWFluoQVH+lzpcAVFUbxhgk8c7oHfWe+WRm/UZXE+OoeSqIqtXSNBYmBzk9jW
ZgLSXsxWiL5i8G5f38EXdfyi27MYs5RFjt3IQIz9QQhJ9h+axZP2F903nLHtfeXs
SXhcOa2YdoAJtM9gaZvgzPAJYaPoiZFJ11cpdNjwSWaXvpOGsfOpMX+v3iMSTCzn
TQUd+X5ypTysB6e9MabaTsuVxRDEhNeP5XewMPHLFFqnBfIXzf3YOPTQevN5tHm8
MKQH7xF3MIUYCVpOCGPivwGw7DbAdCgkaS9GfOH8PEFbG0MReqR1ICmKBOVdUuPi
Xf8ORiI7f0IvcCFJAoPXZPksRTz7Fm5zlzjNjwyEZRsAWg8siyct67yHt5VQweF8
CC+gBQYv4tuDu/7wQVQKqlle47e66/oMKVf7XWT5A6s9yWzGmYzyOgkId6gloW+M
e3nAj3+l6oRCmwkYWgy+JGVsDF2emukW2xbMpEaAiuAREpq3wEt3ivmVB8qS14Fa
VKuecc7kjQpCJKNX5Sy2qUHUfn0fmj1OceYPJGG1H8cpcaYtE5eVoHmacSWAJemc
Eb85kWiA152kNZ7vz1EMrKVEkeFa8THDwWQt4K7gAvlfGbeE1+4Qnfdky4n5YxUm
TRK2tjMq4k3Ghce4qMf0XckazMu7PmE6bljdL9yVNb4BZcMgqWBDz5sL3B2Jg4GA
EXvb8DUcAgAx3tlkCau5j3OIV/YGvcEK2Uya/hh62Sg7WudUh77EILPBQzy8NLSb
YLIPxw6nVsuItOZuyP0cDeEle/uPhSdwL+XJUdGU3A+EEoG5LkIjM0gv21B2rb+t
ckCWnzAGXrQRcuN2gu5mVVpC5ZqE7EXcYbbWzsk5eKwF5/Cme1+7H5A8fxg+k03L
tW5Py0zGPaT9FxQGvuZARwPvg6d+eXNonKm3jFNhwcKK2BVsbNnYTP/yKgTVCYDA
q8UD4YhPfvzTq/rRUI5bYgjnwpS4y8W0mHN30fyd7OQ4lS9pp7FzH8vQBU+2RoMg
TOY1K7IQkeO3tmF//CmIZ5uxhyFN9V4RWmpJpfAW8O3/jMkmWdjzvSU4tEaPDelS
ucgiZJnF+hmmN142k9JqZqCGvT3539D8aCnLGjTcT/41x0cWNxU4C41tH2o06OMg
YhUCw1V+hpuZe0UXToy65y/a+1LqNmrpnJgZ2kCo7c5DmXAbMV9PPhZxGibraVQW
hDUkNHebkMwHBKjNhtoJgLwqEdYa0qBi00RekNPzlyXdsQtJgp9GH5LNyrbFlmV1
5iSNKAmQanR9KePuNNxl8efe1N8UIlaO3JyQbarueQoRm0LmTScnyHviTNi0qsSj
msBAW107bzZfThfw0ocaPSIJQb1sHMdO6UY/+iugv0rr6WiAhlbQchRg1eHWftiP
RNT1ep97JRyR0bj2oE4aaoeRN0CdY4gNCWi38fcRG/HqdZOjF3PuHMW0Q8uL3AyM
sahvgMX7lqiuS7W4uZ8OkVcBDYDtknY0OekxQWpU/Ucaykle1L2chJbHzWzdtQKe
JPkyeOd55N0Aneep4AF5a4ZXfP0YezXbE6T0azjjsgjL40QLq8hDohKZsBlUsXS8
cXr0YlWtEtdaqVeTCmzJGyCGfQ+Sv8wt0ZWJAEr+2zE4Ia0IBb8rC0md1k34FA26
qPVlaZLc3m2Ps6Qr/+vtuWSuZIVfAvOxh2E/bPbamKrDyv7hIiXHbxTR2u5+Ans6
Q842/gIAn1rXnzA7RcqRINjYpog1+XSdcKVBxurXFkfwol5yifyQN5UbgNshmmvN
7Aqn7y7wtDX2wPhzymwN2Ni+J0OMYfqHUH+H+FCWlilvMnIShkj60tozhNdnKk65
uk1ny3aQfrbnCnQZAcwnTFTXK3O3hUyDRGcQZLDoOvCROPtiyP4msxgg4DOWln1S
tyJE6u0JcAzY8zEGPBzrvOXWoni9ssF2OHdnDYXvJ2V5PcPVnvNgs/6+v6MM606D
ZIZiLqf54+ENQQ9cb+e6Uo9Rlb63rwzaaYbdxP4sdInRBY8FO2826m/bfsJH0ceP
hoDHj6mDxsiMrUlk+lGomllDgkkBE3o+ALzrMahA+82pfZwPtOLGgJa/BtyYv0u5
q8UjIlJYhJGlZPBlvKsT5P0Su/fiq1/2hiuIUZm7oSUQV9OXxSAz61U7AdAKgxRP
VZEc3aQT4P63QArT+1OkafLAmUhKkA6KHWUz3jWkzpqUAxubzG1x9kT5UbQVE3iH
aFR/+vWQundzNfJFZRJw5nbptwdvkm9XRrUJyl/QyR0TL17r6FFKam6UCjfDUrRy
xEgNRl9HCH7PdteEIT7aYuhS9LpiCHnREhf/27jRrqZQ7+nukVAqxOe85X6h6K8z
lpH/iwMKcN3XJ3MqUq2JMSvem2VXatsmZMQOzPyRxI1OQyb45mbonSyU6RAmxV9w
664JB0iOh9NQQZK0vHi/U8lcNMGFHbPtHkVfy1FSWUGEwp/ZAQMWeIeVv108g+Ho
WYsJuwnmmpCVkRMawAuuKAhER4IxfOyO1nQ9wyHW6OOMAJ+BOe3By2FNdN8Ov/1a
jdltS83p2yEBQCfiMNf4LcsMTjf+lzsU1uNX+NPogefVLwBdouzE/c8zvCKtoLZy
7o/q+qWHG7l9vecSYKGnXwTnERuuoI9g1AbSjvLecgRKbCwg7/DaCNAiyWTsUXw8
8wSIxLu0KORGgHl5mLFzZa+x38N8rc3m86QXJPryWPEl/v4KA5YfJxVTBBL6ndKL
Y3SqL3UdJ50S0tTdsu9dzyVaDJdEDwYjKpzPNTi9fLFlYs+L17ws44JNUHZ3fp9s
LpALizC+jwvGRzW7N1EZEg4acG+MnfCAzRkgY9WwwVZPjWPzslvg7imTMWD1INkf
3jlP7qNrVaVy3DfN6knvh1U/gSreOVPVYr2RNXD0AEAM/umWxRj44Oj75CzjEksY
B98DQWZoQYTUoISXQZrTd/S4ivMi/xTCx+1cplEDVWxGN3k5CzvYQpJFxAzQV/hl
d+CxO/jLB+U6PuDT8gX8TPlSKSLwu+fgMfvDNQ0twM79ErxXr8QYjnuuRtHfr386
+oCCFErUtU+rSWzKmJvKGEU+rX8GY3GEOM0AaB9UgkJeruLsdk1bNw7v19WwPImb
rUQOU/tnVBnMj8GOKlN15MJj7ifDL9uppqGgeJihXJTxx0Fg2myW0PUDAID1we//
ov857kr6juAHhaFF/sWYOQTWCxY1NCpbUCuHm+ZIEyRdd/8cHLKmZK5odg7x6g39
OgEModkRKmcw8Rekw/nG7CV/9GP+uMrwbiXJB+wkXipf2FbchZzBgP10ZkkqOvNY
nV74V/opvsn8ogArfutU5cGZ2nYbSz2p4MgO3DCs409E/q10gblUNWik18t08zGs
39RcVFSPKQHugp1QKOfYxCoeA2TJ8nIuy8bznCvOql993taPcB3l5ipm0U0jklhM
xlopjF0q5QQCa970DjUetgu5OpuBALSp6tcsaTonFs1KDo/JGlQcc/FlNxMuMPRn
MM+9uZyErjZWKqcAaGbo1xYWJMLQkty/4w4sfEyjqbOJKRhMHSkdoX9IZHmnVhbb
3impBV8slF4V/k2QZOBs3RO4z0oUfQqPW0UcruO5rny0Oj/X3fxS70YEj1CSeWQq
Ein26/T/7YygEJWtJiqn3WUrsR2JSad33RQ+l7vQny6FVcFjuDH/kiMAaUIahngy
xCucBl/ql6DmgNnmqbYhTu0OaWr2YOWBeLPyLEKXH01NSLh6Mc6S3F4pSoe7egEm
NgawfOJ26r0CrQzOLniHrEF4NYWOdf3O3yzHzNnY9KLQFhfnnXhghoMR4L6collz
X9WtZXzprto010oadGJJxc4akGUV6lnEiEMfxnUkyJscJ7VI5JDKp8Pr6ndK8Ztq
vvVK+FCWbz2HJdmLRkktHZ3kyQnNdRN9QNsCKPAQAtjRfNv7/lht/dqdhnBqi5IS
JOWJLMrZSkKPGrblrLMXJJWOIfpGE/D08z/Fmw29DVmO/hnlFJBHysB1mjNykBBX
IL9mYB6ufFQ6YZW/dreeDCLfY7KQzk5rzqoslx6+/xThPvt5rAc1OJ/W9IMhbc7L
iJgQul/vZl97IK8q/TejGMWePxLlabJj+k1JBSWBeG9d7m8rKQ+WoqrcLaT96Wob
RzxS4rwAZ6HYe18nD+yuo/Nb64Ld5INxUG2EpxhRY7BkBCbLoiXpJtOtzPRjnpEM
Z2gYE3FRCbP4OdMeVaRtQx09OSwZyyEUJ+MSUJx5RPXVEdfu1IWIZKlbflHBtCI3
ZD9eBWOBeGvYsJu4odKAgj0FArbL+a/IU0X+BPJIYChQk41/ONDulMPjZcsPygZW
MIipwXacWnBG4gV0bSURGeOkPmuuRkqPijLDfEd7ld2NcOJ9tKwXH4dAhDByC/EQ
Fx8wm4C+Ck92EY5Hmz3rFhyQmBK2HjYddeEUxiE0tLOYgqmYbYbeuOCer08iNXsO
itq3R4ubILGN8XrdFgv2leM6cgeIGkZaxtlnCoOFHdRJKOdloIa+0eS5tJZmaoZA
G+s+MkjONbZDH2TcgxtlEetNEDG/BHCTfEquumqC9fwXZox9swkkDO+9+GW+8276
HFenwt7E2Q5CBAGDq1NUd6xYgalAEJ4YveIr2k3ZK6wH0jQdCAWn/bsemZHfNZYv
tIxp9OzMd2V3wNBOjqPJug0MYlVtMwzZyFCrq5J57zUeu4L1L63DsZKZD+q5I5wP
EIPb4i9fhDQGGDCrEPTQPdHeuOS5QDjjGA+gxcVChYVSdF5tNXhc9191WJGO2Du8
lccNH+fTJV2McoCbtmTdlQpM6H+L9QrB7g3f3JEOCiP8JhqylxCls8P+8pwDvyzo
QLXwgHW31sJQ+U6mbxuRhN3TN+dA8RB5MtLpc7lf/yxb/1l66wzKPwPI/qawSWl8
tVgVLl1bp0aCJ3xJI9pyBCYVuUMw9911FVw4NpQuyb9lWNizp5ynj7W0GlJ7RtWo
cbAOoW2bBd3Ie8VXCnlvGGazqEV82g88Pl4A5q4uOVuYThoBdf+s1cyhkeA17MeF
vTXIUFb+DWAaKVCiKmz01inYcIIqtPOep/T6zDRIMeHv8VQ3+HLY3FwGSOIidFU7
36a3X3KRdw7UGbfTWYXykt2fMZmBCMFzBMYLIwynU+mhpbn4sAxiTc6xrU4K3xOP
a0N4w+PPwn2NkwK06v/V1790bgdXP4JPeVDlVZSJ8UNY1LUK6i3pC2/YTl2Ay5R+
+2WKQSxoSbOAm6cTAQU6kPHzK5bZJ3eg3kHLBmnVrSvqNMP5yJotIa+fOgyjajpc
dBF6DbyzLG3lmdehiXO98lZ6cmLldUhY5Gg5yJQiw8LvBwmIEAnugIHFR9ZC9D1v
/HLK2DB3rJBW+XWwyHkzXsl6rso6RHrR+iAOM9mWC4uQKWoHHIMOhQjtop6uGa+t
tHqBECycVrRLjfkCK2ioBhzHO9FCn+VSOyCZG0cfKbFznGA4DjdhReDJYFPAZAYQ
CAUZUgiqRhFAMApustFvsyZaPcOyB99b4IMdL4jntQQzHgsNs3rAvVrRLVY+FFK6
Ay0A0OT9t7u29XMF6M65oV3r6OiKisooN71paMW9DaZPg2CWkVDH23hAq+c4hBxN
H1/bWAKUK9tgc0w5/UUw3F56uEobS2o1ybS4Z6WRPpGSs3yHup5O6q8kZawyeA5d
XYxD/wjXGUJ2akZx9z2o4sP8Ac37yhnNhU4YCXAe3mgD3k+aSU85mbsvBe3ej900
ox23Kx4hAtUWW/3nZboGhJpkyZoM5p/3+T3vH8LTGZVncG2dBJl8HAKi/Qm2ShBa
mlGFTji8lxdx2aPSS0TWktVVwgP4n2ky+pqO3KxRqUIc1OAXnf69lakgClYkfRw+
iK3sv5k1g+L52gvaJASEBsVjeo4CcUo4sU3CT33ZGGMMTs16xUGht7+rnxcyq9yT
8T0l7iBEk1PA0BhUlqPDLslLRAO/J+3xM0ZBqXsWUvqY25NnuNs5Tt8RgxmmZNVn
Xlg+41Ja6QK/kIRQAe/YtwUznLNfozwnkvU4VRs0FTHpyVMi5ku4B2DAo4Jb1GEO
7hAjQxz2N6XrCUrBX3dGdrtwI+jkPd03GHKMYqHrN7s3KBd0RCsqRbmbYk857RR6
CH4IGXp2myopTH9gJ14aYdhSQws88ofXR6bW9xfQoeI1v4TnyyrxffCspOKNELZ0
r7FvIZ6xHVajj19f1aRMAfQpkh0laRRCtUUZIO4iBgiIqqmV/c0aWvvH78Jr20pU
HT933qDWRv1UFpLpFkD9+9E+YvZ0shTXc6NSQDSEgotVlY3f5xijFnfsVjGqZRfV
HHHKDDTY5QuomJBTgYOE9rbbFgeAVPTbRYbzvIuEPuxOp7wVSy/lTVxvRlIdC1fE
6MrKZA3YfFwsbfQlIQ6rBXy0jhl/EP+vtygpB8MVa2s29bdnMGyyMWe6+0wnMI1z
5tFLEiB4DTO+n9lbVKALfusUZhdpP2SrYqr1ShGPTAH7rd7zAkhHIUPnbLchjHKk
g1uO4cNo7nsF34yez4Mnxl8k1t57RJcLs7kSxpnQ8PdJb+qmtWF22V7dzjLtMKYw
M/+t0n1420B/uhyE8mflHs9s3+8/5McEXUsei0wMlB8JyxzmidrjPoCr+2bPvSoF
LI3ZIsuFkUPUvzO/JgrrCZVC3aJBSnN5XMxmBdxSRs159vWRGEzLO18l7nzvMLGt
L0RFz9jltWxdcl9/oCtP6ThUZYfN4k8g03ZcS2WIzq21ukc5uNOqcdAsJI9ruta+
HqX/843c35f2dEWSMpEEz+xU02NLlng9b3x5QvbdY3zNmqQBc1S0mV9ckrHTjhTx
utznMaKsaECym6+JurDcF9INJUelPGGik60DkVlYx5pMrlJEUk3S21gwOChfQRXF
MreybENDZL2q9HMKwOpt3jWycslJCfB5RBpQp87CqjCPuVGPU/tTW78YvXp0FNSz
7dO+pgheQspKGwerJc7e1Pkh0De82aU5le641YSqcLsocdXPr6Ra+U1x8hBrVbyl
82d8/NVNFMryUsa4JK02/4PxmzvZpZxGbUszHuJaKVcXWOHxPMQUkVXjTbl8jWtc
50xlokYSbwVWIbE19wXcaP+xrSxK+zTPi1EkCoEa1mblfT5uFzFsHwh7PZmylXDp
j44Ti3CAQcpcitn4xxT+yfIw3rRASQVOVbLghacPIlqKRwP75bRfNVH7PZmBVGZ5
GULIA9nmH5A/0Px106TE6iU7X3UpU7PhlFfShaHlw1r1a+c6HOzXgGr5o81gv8++
ikpbEG5FnYhgdODn6KjY+pfIfeIKxSyZzWt4jYytnOjvhpCuX5sZprV5ypT24U2w
MKxEfS1qeIR4dK7AnymhydOTmay+vX0LFvSsXEnVR03VdP0uEIAwEb1+JZ3q2ZC+
EpTfpzJD1Nm6Ic8wY1oeu445jU6Pp/AKp5eNyW+q6r+xSwNaODxDiKdlLniFYTI/
R+VEecuJffdH+unHboGnfVnhBvdwHG80hu4Gv+gnfY1x4uXyw8Kv1z7aOl2n/J0a
3/nD1GI/xE7dJr/RdgRXTd9bPEfgH/iylvJlI39IdVBuVce7nC+z4NDQL71/xfca
ZOtNrB8Ng0jR6xAjmJQ/73j4dNMEIrrKyS/9/C2zk35C/yQ1nN6umOx4wVF9xozq
XN27kIIjC9nmQi3M9w6l1PqIZVcXKoTeIUxQZ+xU45Uq7GcqC6TFNHw8++FjhfZi
XCuDsN9GAFQPTAY2nnwxlkqH35BIXKgnHRWbSq9PVdVyPHIzuf9QZHo5hsQ/tvmI
wn89YbrEfDI71FQ2x/zgYVRt3XOq10H7Uzp3cegw8ME5FBHg7xpnz/C8p6cCxdWn
xxAbmropTTxEOB2BUgRQIvY9oEWwBK/Mt0sMGZZGAIV0WIp9i6vOLWybpPqoLjl8
8rQSw8eLT0viOaoIySbYSxSkoarpabnEBymDwrnRET0kXKsX5yz9tINtlENRJlpZ
+Xe7M7Rtx8AfFM/AkSHMxB0irNG9E5/JQM4B9rYlg/MvqVLfsYggB8BHaBR0URY7
ABEFg149iiUg0exMnm5jTyMCOEMWuQjfvfh+9D+tCd+4xIx0wviDgfV7irSXSzOn
jxg/Tm4R/GGNEK69BDn+djjb4r8htiWk16VAj+6RaCRH/O8NmrdUyZzSsWo+J3iM
RX/qMOiJSgJrX1MrTisEc6pBu6K0K7/ciAgZ/T1eV0nkZGn+3pk9N3mx9OVLDJ1K
0qlqULtAo+lxB6BrTE0ykcmW0w3H9SIJAPBjjrdwbkw+WhbDSR/gsDQRhcWJngBN
RUwoukOFMygC0FaFugkE0knmGutwXD4R8xyCnAlHNTr9qu/8aOc46bJZ1kCzEalZ
kPnDsyqO2Qs6ND5ulQ1WFyZ3flVk/rDV8RKkCb4RQdBIsjaVkgM6UPezz9iCf30y
2AGVsGeXJTUZb2DhNTjS/ESCeiDOSJmQ3dxEM0uJxS1XHWSPDJ0L2M98kq2spgRn
d/be9yi9HrEEiUuBR6S7Yj+GRlDq4ONqOLl8ZLiHmlSd49fDojlEIy4NsWv7G+c6
5z7Fvd+5Zya43gQkQiRWu3Bz7uhS6LvL1oV7Wuqt0rqg6XSXjcJF7JJHZIoO/3z1
X6OQdglI3s3nr0XkQi3wOKssPlmjThVhwVft2DnazleVKZT7xfIa/RxLLTd58Alv
ePcFqSZy6DzRSVr/Zi4pynKNFwOu7PY25IpEBw6vb1u95eGeNhRCDPkSfwgJll86
FNLXUuQznxHG7K4pX2oyUEce6qhVeri+smYLssBXwRyh5ngbJqj8L07Vnfhw7Baz
eJdLj1g2ZQiIPMkPxJcPQurrIBeDmheD5E1Fq9PG0g4q4+zs/sqLZvH83cIHSlGw
lJsigjy9QUrWY5sDZ8SwNtaq1+yPqNDOhE1kK6DrJGvmSWJ14GODQxxzLXnmeuIe
a6kXQiF4GbCL7W7Ywt9Uy8yTmg4On6ik/p/Kc0x8nEKByk5M2FIm0v1mKPdc4w/P
FKCzCwWyApcT6PILbeto3Z7GeBX86ktlwXz4v3BOGNQAZXbf0v2TUgT2pagva5GP
FU6+0QmAFRwVBe0SgmQytUJolBy4GuE+obvlXwdVwEupxZ8v7j77XbeC/3dSetrE
HRCb93d5H1nlvvUE2IA8MobM1K7+lWJL+A6vFko7qYnBwhAsTHgBu+qctu7j+8PU
hYk/+ZanaGp12eWUwOtz/t6A9RYFBRM6sGgjz7W6jVvDpbiXoxQ/ybtxBgCbiIrj
U50oe8Pzs271MZCbW/KaGQf+GgRtSkucKaYp+TnyquU664IlIrcEUM7Do2sAik7N
kim1khuZt/48HEk1DK9JbheDGjxz9rNgS3Xdaxf8y30x5sXKrP8q6lKmCdQ7g03u
NQBNm7ExwZYwHDUQzB6GHZP1P+mrCP+N6n68qssYCW2PyzdVYQTEVnuZd/R0SnLF
TMM7Bz2sPmT79qFQ8C+r1mJap/v0UPHs4vd/fw4+7i2lZLVvnOn3os15UFmsKETJ
/8JvvAe4u2ZKyZZuQeWBR6g1+QpEwdH+CTsyl7M1C0yGw/ZjtAgt+A0VT4Pp2zXf
a1CDOBvRfHpZ/e5VbD+aN+7v/vmneRFiX4cThiXDJngT4vJSamMl9j95QOyQpBbq
ywdC1yGjz+c4bj/iDYByEPU0gYkDzhQL2AcoOo2cJSGX5pPJCUE5imAemO6jBA/Y
hAq9cWSffxbtLyH6lRUietp+jj/J9COh3ZT/CSPcr6y/emBfnxsJddTSP19lIBDH
WfTKA0iauGBk6nEcv14bNzVtT+2SKn9IsnX+sEZWsD2pZS92bb0eyRY4rUOPGdGr
nBSm4p9xAZMdWFQ45O0sOaoizU358gTxht86GElYG+Xa1mcpk305c1BTYb7Duq1k
QgqJVlalzeCaqvMZJEkOohpvRibv52P9UwP8Un0GAM1ZXzG5/h3YZCsxZtO+sN3F
rX4xj0B5IsOaKsStw1v2i1LLrAcmx/YzCMp051bJL9aKbP1/SKjFJv4kd+Cc4Utt
RkYkKmNXV9a4pkv082gmJcvy0t/SivhqarPpGMxvqbuAsTUm7R2oMG6LLr9ONtxa
QNVxBJnEsRzfhmfo6E0lkd4rABujQEiJ/krf5ClJG6anobYfRa29Jxhyh1k438ZX
XzIi/+1yLuBMB78XSg9foKmq762BRpUK9YHf/4eDNOH8nGYbhbHWAkwL2a28pwdn
X3CVq2CtW3MgZoUk2UCnOQPB+TLCZ6zvDCXc89aFDD18b0vokbAXLK6OBUe0jqkK
aIPVZVcQkaw0eJYd10CKEr3ow3EHULuHMm+CVhU8rBpMiC7Gefip8RTETYb+t8nq
hvCep6AoBTc1uy0C/GGBRlywRVFKxy1Tu0ql6h2Vw/c0Xuj51c0FW26uC7rtrFNk
eR7f/Di1IokaR2c6I9LCP6GvdQoS+ClyjzY0hlawGD4gbpnwA4PwM58w3JIZ28sr
YWhz5CrTfq96KodRdeUN3Vh0QAKTR6lXHsfjDiSGOCXUpdZwJZ3e1e3O9joJeXat
+8zQueL/ltcjG6WZTBO4fKZp3kFmtvu6mh5l646TL1hYHLV43/vvFBOpwPKaUSiY
sxClLlMtzuRoPgapP4FdmrvGmpH8foxfKGeoNpdIRAL0le7EM+QFuXf1gh+fBvzB
dTky39bkycqqiE46/mTLGZKAbinqxXvVAGPJNu1Zor8JNPqCpYSrLNROQspB0v/Q
1LtXp4yYWpE8B2IJDsFw3HGDCfeB9ISzKcRJ7hs1YnesUI3q2XPTNVM6a3pgCiJF
0RyI5ndjTIEtXRo/VMtkboltXwsJUlUFf+fQW2hbkMtoJiErw+DOjOIwf4ujplmi
ph+QZ3Nort3Da4Y0JD5fpClOpXjBt0C4Bf7/J3JdMhRRkNg9xsi1BvZKpyK3fkqN
+RXjruoSDh7ywaIAcbom6/leFSERrT4Kl87T2qFzH0YnQ0SiwNd3PsemZ5locYq4
o+IlQxH3kOb3s4BI3LZySwA6Ji8zfmrVq8giTFl4eKl1MgWfxDVYTWqhfjxEKf2s
PGVY2DDm2TX6TPG3MZHg9+BZFmmwDyRYNfsVfqHbNVZZZRHcL9VEWiRGZcGA7C0x
DWP5ZxTuF6utojMflaLgIannf42Atp6n2CPZ7bTXgopOdVf6KV/gnu4s0Lvw5DZ4
4qiLhGfb6o2HJet1Bi2kxcMypkescy+vSPqK45DmuPoxa/12QZP6G9/DDAVfoKLo
YfMTed1bwJ+l9tAV97dqNPiu0a0vxuBkf4swXLiyGUVXx2od1+V/swVltqTuWZym
P8dpLreb284XqFjJbyKHksP2+EPJvDigmSj91T/9UYJA8qi/bu5X+eB2kJ3eXdIr
sAtBcIv2qDzpkRnvaEiAMZ5ldXnA0nFE21YJng+xW2EDWhxZDCvtS9d52YOKfKJB
9WemJF6PmxYG1ymRHbS+prLZ2mrXWx3ibrtGqR379DIPb3EKCbNdWKCf7OGEkOoc
fZWOYsi+hON+wSoDTj5SZOG6zzJsTn71cu46FaXZ+5jwpVuqTmPtIysP+rV3aAxJ
UiD/pguzzQkggnj3NcCXxjxDu/OM/S0Gz3Cf047i5eQNEBSwabDWLNqo/ueABMZs
vwlWZ0cmZmRew1Zm8GyJ7UrcHJ+tIZk2wlTb+jeOGj5uI0rcFvK9SJmd+ngTXJsA
HRWGnPGyAdQVCqKl2OTvNJ7CjdXve7T4xThW/wkPdb72kw0fPLPBSc0vMig6H3fD
qMEEFmAlMF9JKpqEUdE8wb1/oIQT7rkWWad0XWLZckio9fNk51KaSBJCPe/ugbdW
dE7+liWkfHBLD4XIEVF2nXPH0xM45O+1mqDZEEZeDPMgAc90l7cH6HzxRkq++wr4
txlEoryYSTnjiQypb0usk/AHEBpw8aF6U7o5xz3Oifj1t35reQrvAbUP/wuGnk98
43f6k4Y1JZKiQNCMdOZaXxZsCTxtJ7KqevGVyHTVDU/kZ0gbAo0jr4v4exYuo6f/
C1/YBgzg913Za7tpohrY7nuo2HyfLR3xElWA1KnLEr20e3htonQ/EMy5db0zUuRb
ak46GVnThOSBLI69AWZjYgQSkJ4eVTugazHoDqRvKpSIQkdXY/TBEnzVgoJk3pYu
ivdqDw9Jr7F9GHL1wGBDO4tiVnoXNCzW44fLRTYDSetH15dTNf03l31BoGHuaS3w
nKTIZKrkmTz2z66DWZdPKjCT6uYrpvHJx0nSUCIgEUfXtDmdYaMpWm7Mxkkr7704
zbjPqAAJEFv7SN59EO40fFoDD8xBvuSbxKTvHS8IZqIgp0TgSVKk10WdgXjYpAEi
0mCK+LSY6yyN94ajNEzp4Rukb3LdAEyKNXEHWVFV9zFWq1F9Zt3P1J5gVndSsg3D
jcxLmyg54wLNfjLxJ9AyAtpdIE7j4J+fqYXo6izHILxe57G7HleEY6ofhfuQzu0h
1/+PyJ8toYPChnH1/Ui6c4BCMfpkMvglzKBs59M4Z+R8H+3yWrdkgy0INIZUXRiV
5trmxW31o1Od7O/eg2MB2xGaPkqXvlb/5BlcwjcaeEICcIOsKfBAqi9FcUVhHN2T
+LzMF7xoZMRHxjI3KKOQcnOCpaILMkzAmc933NBraazX2KifrRYbtXShRM/UlW6I
fPNoPq+kIag+TLVFkyOUe2TcQvTw0oPouVW1pLeweWpJ6sHT0zZfFVErmARjQ8oN
kncCTBbyt55PovDbv96cmUeIJQDmphTwcUozAUSrqsmAFEMiBHMTQDn9Pw74GGuX
jqO+bcKQcw6VmcnLELLE2JswafbiuVqyuYwHGiynlzYgGpxGLtwhBmQ8zBsBQ9/0
a5nH8FwkJNsBtChbO5vP0LDAE9CaG651xreY9YP6Wx4HB2DVNqjUWNo79YspU9Sk
eItck4+zdZl7dlctYt3+L72f9NzFomkKFvLAXICprbEJtDFev0SVS7AU+sr+3v0x
5HyPBXrO+XGplFZoZ0hOZd2tGlVEm2clpU0K8rQh6sOKwNifwIeuZqnbqAE53vZ1
V3aEx3STm+UBlWQoJFUnuhQRp+rSBlSo5kzVU8onlt8jl4UZQHK4wjqXxeCJlqs6
9E3wM26CaIPfG2FMdDDKcOqwdTyZybmnmbVSLlXzg+X2xA/kljm2kCG1ETtQjc92
S4us18PlyLIU6AN+q46JRav4kuL+74HYkhQ104r5a+q6OeCz8pMIxw/uxD14YfjS
iscqNW1IJcCqp1p3YX3YLKoFMyxFYSp+rUp0/OCcQ4LaYDtaon45IeW8fJVEOkYb
89ZVh3t/XcifblQwZpjEJ4rr8XJYdYQIwxktTj/oLkOcbn8QZwBxUBFJkdMm233W
4Hk7KZk0E7bu7FsWt2rG2tBkGGXvBFIpp+P7CrDV4ft02jF2YY/tN70y0I7NA2MS
l3z+poRmJWD1j6SXd5ez16PxWJty1gRuFNLJ4ytjBxDZ007AwY5UUgxpSMNv4kSW
/F7PsV95nmBqhpY9XOQCfJuBKpJ00jBbCt6B9SIk6wvW1VXECxk50YnyfZwaVm6J
8chCG9dRn0Ys4m3SCCz10zazQVtpLjufCb1VakYFG2diR6B6IxNdvWCmfYydHJrP
mM0TPeP6+4kwv+I7MnKH+ueWQc2Y0VmxIiCrVNB79K9Lnes3P9bHDwlXSMfrxsEs
27N6gUbbazVMHJYIJJkWRJhlVJbBua9poCr6Li2rysOpIx5zGCjCjlcykmxSBh8x
fS5gCOTupcPp3kg/8sYS3mPKif4F123eHnD7OEeSqKWda/u13ydxIi+bNK+x+m8H
3EGgk5C7QQDtTEYBV32pwzdZZABsSzsoKZydm8w6nxG2bhsIwFmz/k9R0yd/VKRF
jRrl4vHvfCBHtGvCw+o5YmJ533vB3Nou+TdmcgiVqtJE0HJIZAIol5s9h6tJYQtO
EefAe2SUtwjt215l38MWQhpI10zrQZNyv7XOI+U8r2+Pkg1+82Xv6JJAnBqD47DY
m+aFautmMFAgmXXMDqkyvGfBBCVywUWrGBKRuBailuzpYjccJq/szeOqfQAw1q5t
j//VthBgrf+bXIxlaCsAjKEXrDNsNEA1VBRr3WrRF29AVJo+rQ63z869FG4AyHDD
RINycJ7ipH5yF3Z+xfGAZrWSBs4S9mpECKcufZk1AWW2vrhFQZQs+AdjFm2JmDUb
T/UcBNisTVTGvDULRrcH8UPz0D2ZRroG7FZ5VpQCt71ZUO437WbMUIg50GOKz9yW
NEsIgGa3KgOlxf7bVlOP2pvKQspp3icBd1bRn5JGIAQ7+lmmgYRTZH4uu7I/PYN+
g7ogYjI8kKsQ0JVp+ZJlK05talM6Oi+NnknY6eRTjV5ug1esYMEovqZmtDmuqq4+
RdDV54ksE3W4nsAFbiVuwslkxENZ2A/dNF4sb9KjzWVofMnMA059TiH/PXaMiUAy
u5ffpg/8cN0sA9E3fkB6mF7N2HcRy75YJAM4XjsDGcnbwteb+NA0FyxksaHXdBia
npsk4fz/N7/6Rc6HOaHK1GrzQOohIk8PqMoZ1WUwaQSnVQiDogZNugU0tSckSUuQ
yaM632YfXFS2w7qPqkURKQhNwn4sqr9wYTbLC7HicPI3WsKXLbuXkO1pjVM1R6xo
EdF+alWKjTp5vptKBcwLIyOmZzQOtlKq/qWYuLlC5X8eKjl0zAGJ9lvjnJKX2/to
sCX9EhxMw5qCcEpQhdMI/whoYuLg6kuaBW2v78JA+PqOT294t5KMXlgpTMtQlvba
VshDOgC6ZTpaDrTdD3WbJvL+Nm9DIjqwtJ2IP0mFoJouwQPwEklfo5YBQRYUL8UB
TE8hRlh6nBqglDm6XEMcFN3lR+gKTvuytM8ELfQGuhmf3i1Ic1judyqgW2Exx2vY
tzuYJrf6T+6uKQUXccsR/mHTjKvUGpf3lzUUCMetKa32a5oLBc5g4Ht8awzFs0as
W8Rvw+hAYW2VApKHspd1vJeJCAjgoLql8RCvKKoamZ6ejlNK2S+XC0I0FgsN3UEw
Ewx6vfOuWOhvoq86cgQYaQpYMt3/lLNFdWC//o6j0esrjUdXrxj4O/P5OdZWL6QP
7aTBFcuUNnuiZepg7U8I7FY7w2wpRTHh/7uc/ugMx5Us6rTkmGLXaWRldqv1Ma3b
VadnDGqqUpwD/353ZHu3kaTPZ9euEBgaoEbDxhbIvQFBJJ+4CThklyzubitQHTVb
3dzlSP15RNwd//sq3TPD4mQaA6hkzcX0/JuPD9us/KMgq5O0ccAbh8e9Axao1HGA
dIWblhN2XmpS2/t0xcsbsJx/Uhbep3vz7QwkoQOJiXsTXxqI+5ok1XcWj5Ed4sH9
c78gDs59bGmx6mIcvWKBJVGTMfLqJby/sXrS0USjWAdM6+jQx8TUd0iXQlI4980f
RuOsK4nOHnLaqiWYGYnClU6LyJb6t1wH5EXpGibKQeb1EBQafVW3qU3Lcgvshotk
NINQiPOjetEUI6rjCv/RxmVp/W94kJVIsZinfZEZnHT81Ek0BksxrV4dQa08CqVP
//NeODU63S6n6rwO7DtV/GpwTetaECaPTC7vM38H2YobE5rnVOdr2GnAAkji2r2g
bQyrpkmsXR/XXqtzxfdjGxNs7QdfACgImAE9nsKdfUPVscretKUxAv18VilIujFW
x6IQRbyWyVHOJquImV05N5MlZ1vbdAOIJ9IxzF5I/B3JmfTLB4BRb6rq1V1dsOqD
1TbdMGWKqVsfsBjRJjIxuX186W0EWi/IHc94be0rb/K75SPNjby3NFwJWoYhTEhz
P8I8h2TsyROqhEzdPwYcMbE3a5qOHUpGYK3OpVQAHGtk4Nr7Sa6B0YOzMGilmmfO
OfRYlH2yWkDAasGSshGGrmxwgMDf8k6nYo9MJAksnZ+HeaoYDcOVStB/1tGquOSY
Rgc+6h5Q+HMaK6uijqjlk1G43HScwdWlzbB75U/ycBxaqnoT+etBz6R9vccx9ynQ
ZndiFs7+IWuAd7juHmaS00LtWym+gEdCC7T1DzKvTYb+iTNDP0OkDLOUy/noIPJm
YnVLN7Z8jf0OH27VP23kXmd4+KDXuf8nd8CgtVZi2Z2MbCq8S7H2oRs1v5v+SIeV
vC7rM/GJgz/srZWhiJlIjJRTCdyB2+y/RZNF9eYkJ9iRdVdgSpOKryXyVRWwDQYB
bET70xKboiLvOBeoYQlFpbHMjrZWVNLO0GWpETPC+tm9JUWu4RreTkSxfkUYV58D
QpgT9NsFGFneCz3dMTqEVPqlzcPB+cU9qOvNFW9KeBcQj2xIB0MY7bfP/XNx917N
JSb9fHbZ8UA1JpOXRSugj4D40lNxlT4AhQww/+eGE6dLEFtokxR0Zmq+cLdS2/hL
pjsZXXbMsOXjXXlArIV5hm8Nm766SGrxjel6KclIKB/6TC3+vsEW3EUDSDGZMCq4
G2FixueXc2Iz55f2czu7gdXFXZHzIw0SNVS6kDMO3Qic40Zkh96Fg8EOlvAVUXPd
wxLnc9xXkyQAg5nGQLRGY3u50w5VsX0Q17cgDU/+6yiCh14na2dRjAnVraaaWKtH
oBfWBIzoovYlf4t1bCTKFpKFrTPPhQVSamsbUKyDO78S/kbfcZ6PWrpZHXYB5DO/
WwzCaxq1uvFZa91YKFxrXZxLPbr3eH/xp8NXHbfTv3bJxgDL/FsRQ8enXoUVnaQf
yaE2yCxghPKuWUKA3MvYE6ZNzknq7EjJohaKT8Xl8WuAT9YxPdtDAzn5z42TF2N/
BXMox1uwpdqfJVlJ19CjgzeSLptPizPJfuzsSe2wtGFbU/00jYDmqY4NJcKmrekD
Uiqy8Rse36M6B8PJhFoPw6m+VN64XO5lwVExZnHX8WkP86YbXjG8YqmiI7PVucsJ
a5+du+8UALyeUuK317XbLir4FyADwtuteynxAMAwMvKj0HMTJKk3OfhJonyEemBu
gRCt0pldWlMsxPgznjxyDug7m/QcsltvRETdXWQ7kDdpJlAJNwV7xfUpqWzdoRPa
iOWKXB/yfz2FmaNTQsfxFa2STDNhLOXNFHhv1TMou6oGCpYQ4Z9pptjYATBvPUCp
5+MkL2gBY+n7pSqGvXuxByLPmTK4DKJuiL5dHknEU/3LrGImvlxPTCJ36y1GITg1
bOSsJOf3q3jJYSZQlxBNAWdW5hbZYTmqnc/nNuG2IDsA9jz9Odz0Tc1Wr4yeZ5lJ
tu9QNtDL9Ujc1ukBovbkd+QQxQ408D7q+ko6hXC8F/rxmSSsP3VMxkf7XXyzfhMo
O8aIK9tvNIU42aB0agb1EjUJ+XE6FC5tejFA1SVdqYdnKE5gGbVp04VLbwnwYA5a
LX5dDdg29Cjm9McBAgqBGvf8yysd22K5mQsJnxvwKC924O/B2B8+yA5mRj7Qvfwh
hlT6KekS4gHkjEwuggBOm4+C65JR1QoLMSMuAh2z2cj1QaDX8nN1wHWugu5bsAd0
NDgcBjzJgUQ5AhReJppHvflt/XntT11sE5nZ5Gosl+1M8DhAYf9Y2FJc4bnFd2s8
kRzGFW737NNJAiJYbKWWNbRjV0bqOqhQpjuyFuQcp+j3mbhkYONhKPzBiEbYPNGz
AllipE6oofRuGDD7z2HIIy6IUCe58NjzvsWeVhX4FiNETbbNlcBlsYC5/Ih8zaZ8
WoO8KXtK5iw4ISXQEWLnU0Iq2jp2lBW5KE3LUarirbahFy4D/jZucyYAl+7kI5KA
+/8/UrqitbmqcuFkJXLUbo6OcrmnuqiQfHsQ27utsX+OwUvM9NDBgs2fd6j+Kr5r
Ze1avs/uXVkdzR3vYNKOjcRT9McEDVglnW33H0qtCbFSvR0AD2q6LwyQE7CBJNzg
ieYr0nDj8mfEdiggWysDroyFhSjtKBLUHxBNaeb5eJNZEQYwKA3T6LR1g9MSJw+Y
4bbiUttaQtK/ts5JvGyh79QcCcuiw/92UjYUB7KQeE7w6DAzYT4ZFF39lDs65Mw3
k1y7AdmJP7UPiFChGN7BWM5TXgktODDICt0LTXnV8zpejsO5bWBp0/FM0ZF7s+lJ
VktgB5/m2i+bUFdLIBPC5+AJkk+nVlY3HpNwp1JsG8vib/kct0P+jEdqdm9eOiU9
64/Qf8sHUKq78bnrUch4KzpGVq8ygbGd+Hc2B16SWvTAUBoptFCt0ZBw1CdeXb3F
oxAplvHgJSTO6EVSUgxSJZd4Qqj6hPiJJrMg/wh5EXVHWaiOFtP0lm1Jp1C7PP9f
MGvmANquiKgtoIxe3e+eyCo+siWnC+GGbNZKDZ1yPuX17p/eHvtCpM2jt/mtjimC
yLV9HSHLXhS0fHuND3v+pjlHb8w0wMQbN6Bzlvw6izTnbBl2TuoFSowSgrEhsluu
TSL77BdILW15lg93R9cjyiDz0pvCkM4FRTwchqhfvU/iJEUp1AXDbjlwXKct5r1O
VbX3aRUPLPk130NEum2APmR6GMzzc5cDLks3MQhtBq9o8Cy5toSKAwYE0PzSc3qh
zEdciqRPdzlYEWeiYRCAazEXkA37OUWl9Ig4xJ5Ko7h0TzQ0mmVmmOtrFQAM5R8Q
b+/fyeEgJmD1nph6Wgfswv3bfzzNSjqc2VZHrH9okr7G74Sa8aHXCleKML9ZuHkY
5DshmKASVVWGGzqaN6CdeoVW5ebPJF3Bc8BxFM21vcL5AEKoraAzTx5uIYJUmupD
tLpfCZUjg18QUeUTmIHFj/bR/SdkFYTGhlTiABjaBEKvmbOmSFpMebJ6yiTvz+QJ
5h1lKAVLGqwmBPnN+Z6upNEv/sdJQEx5nRfvQhgOZzIM+0yGiACQ/cemtjR+c6rf
mjt8gncwR4180SZbfEXIVkvAJ3WCH5RGQMqrKkGEr+dh5K/diMu/Cs3zSCpRUDVX
nfcPdaUJaW+CGYIrQKUjOf46840jOU13un+e3PwjK7FFyqndW9EDVoScW+3q3VMJ
/U5Qz0gs2IsvksDtaSVy2t3UpkMB4bFMA0s+T762KPIcgL+0M3p18+j6FIo483Mg
UHu9gbFMktnUO9RxTWojX6QnE247KEhUpEMPrQ/HIRWDq1o0VyIDj6QzXojZxmYs
xtzi6pZQ7NofjfGq2WGby5TLjx8jsfxwrGYf7ILuqtgDRaORf6zik0+9n9WFUW8P
bStfaNsHKykdvxm/+nBuJfKUhsFNJgGmcFLKzGIK5+EfDFZZTnGDin3TA1fGMfzF
KTx1TVxvq75p+qWoNrn0cXgepLcsoagzSOLGZ+8IBy6Drg6DVO9HSzt2RL7FZUqS
7DgTI0Ntg/HvGESQmFDQ409C5J8ntRuUIafFpB421z0A4govZpDPAFv1INusRyqN
lUbDGzwwilAVoL/VOCT1WaSLzfCLdH4zUWPzuyX4wu3nUE/iCPxvXLEy0toCwS3X
phdffgoC6ii/R5b7DEMibHwZ0KYSp8ptG0s+3SysLNuwyMBqzJGEckOtpXtkW+lJ
2gmC0jJW1ZevgC5PZZweQqIe7FvrD07D5Oj0pTxRAeYkXPFqN6e05f3kTSE85euZ
iPNu3Tz8ZfZVFmG0oKKmPD6XpofuSIFNlZZ/fEBwsHbCa/Z4z6FTOtahIPNpS7iy
Uucfsn7DkIIcf+Ho+UC9fl7k3MFTeg+vURWbfaZCt0zHboz2PfME91VsSBFHAMQA
FiRSKX7w2v6LhadNJi+6SMTlA2icCummhv589RTgI7K1u8t7/TMGoND7LVCTD6Zp
/DGocr6N0qT0TSuiPPHSZwhZasR1sjPY9UxlXDjaDSmpMnqK2cD+GAY/U7JbliCs
Gg0RlPz985UHw5OwHRkOXqggv+vnrrxsV0ubzYqS+QqXcdmEXvCDR0nuyY9Hqv3h
giuUS/Qo0BJ0v3bPU5Beg5PTWRi1p3Gs9jRDhY+S+XL2dH9T8/BQYvGwQ9iDfPIc
BLCtskHogjc+1+QgY3hJBv+8Zk57CtE95cigEa6LveiYwuWXuSNALs2mzewWc+t9
Q8tXUM6O7MB8kOfCHwziKDmlmyZ+3Rz84lwJ75YKZ0pKzllV8SZlZK0d17f95I11
vWp8hsJBS9cYbvEbSRlidJcVbfb7K/36xVsix7couWvcfeVg+vWACI4lNFqwhFqT
AzhKKhBHpKb66Yvn/TCmlRtvx2Hz7d8auyOQyW622rD2+r1jtKi6Z0VzOORkjIA/
1981fo4QkIIFw5T9DqJjWm+PRd1qyD1AGZHMvxm4092mpAT9e3ZJGUd330SWGVkq
RcKLz8kjckiyCUb6qSseCwd8PLeQ2KVV6qZkerNb2ZLYVns+dV3hV5cDST72g8xS
bVdgE5XL6vutwCkDsPoWqHR834P8FYdyieCRkFajmaRWCLD7etDii3vQOYFyZ5AW
Q2J01cTdkSn4Mu/Q/MEND0CHahYke7rSc0Agx8nL2xLvgsykVsOv2D7lZKfc2+5L
LE/DwQHl5UK0lmHgbihAtz1HsIYGhxVMTAPpN1HddYNFcRiqpK4Bm6yfdU2uzUbV
RQ6xMjiUE14Rru4hhe8J173RwA2E/WqB7mF1fb9cpbuY/OudDydIMYKKQpWy8TWy
bosA0N079wNgefw7GzP0QQhBjPsRbGv9t3cvdHSQYjHt7hEU+GGeu8exRK+hFCVS
PNndaR9V4fKxaSdRnZVqfXgshMGy9mcXX5ZgXqwAGy+KbvMQdzNf0dATPIWoGxSX
U9sRLGDmwb+JcAWIERRIflU8LjD+fjWgG1vooWcy5ShoXmfnE2esIQEiaDomProu
lmOuj+KZwThZYaczZLz3e9njcjxfJYQ1xuW1ondRGqVkK021WCRazzB5c4RFKhQf
6nCm0iX/uM39LfoM1Qjiu9rCA3GGgJ0HCps4U/sSPNkFlZbiQsr7tIW+EXubqArN
koinJtCB08gZQXwxWC42DIIxa0s3hpfBJA1K+baU5sHQSVzsZMNNdZxC1h5ZHIcu
H0dqbYbvaSaWItfIkZ7ebMv0WGek36elidzkeRSnBpszF/HpVR4EL8hgeYuEJwyc
yWY57s7IdkfGoyRGOMBw8AFJOM3byEwdmjNerM8LmWVzQliUSdPu56rGFbSImzPb
0C/0yO8Vz9wZCvLzXX8uDmp3dicRFhZ9Xk6CXs+5/Md1C4TUudVKcyBAFszjuqsL
nxZeKN5afs9TZQmiJCoTABTiPsLllqaNYP21S0VeEulL90EJGYY37yY3ACEBNKKZ
4GZ8ywiydTeCvBvyXEZr/mbBetfqHNjDDg929dN+k5OuKFDmbWE/4TldwnF49Uqz
lu5xCuFMHfWWbiFUMZx4Y3uMfGxnLGH11zpuDOJ9IHKA1PUFgvmJvK/m8PfJIddE
7ndoJlFVGaqowN05lv9XJqxxM9XO7a5Yl1gMi6onxKtTu0/cAIZhegENGD8shUXf
P1wHoRT6qnWz3M59ghZ3D/BGSRYvfeCd9z7jiuixg29opILAIJ7Eub1Nhx/9bi7j
Iu3W/orA49PS8ia9dzgQQi85M9+dwGQlrlNr0RIO4irldLRr+JC338BF7GsNUs2P
+8R2VntTlYSjNfdjNAUMoPyJyO91dJwBsKkzZrPgezfvrMJdOQZ8ufg/ueclORio
3ItXDb4P+aa5McweWw6rRpVpXtMP2Daa/+Vpp7zkozhHxCGCdwsrjSlim3LbgZoK
Hkt5lPHQBIZlc0Hfvn4FM/oHGAcevpRcT3ADL/6jalE65z8MHxXoFT+VHzPdlHTA
DPnHpXf0eahPNZdBqhHIzo37xW+o+MTDC4yBO6r9rqUeNFRFg9439eZQjrcC+ljy
7dTZRjOYJ4M9HDcDFWrpH6g+IEF9cZoUapxqfAvWCRnqXoRyT9xQUE7gyvSVWnGZ
b34y/UofNclHXWCDxbTy6vecyLV8HYF5Ntxj1Nw+bJTDniuX+3MeVJnPq5/wf+nj
JXr77gU8RCuZwgESRq2+rmfpu2TeexUeHWcA/iTVZJAqinjmJsBN0FwdjtSg5Xyy
pz7gqA028dtBNTc/XS0QFtkK7qp8f/2hL3U0kG0SvHXusjBFpkpK08vogq/yzylf
MA31KKiNsPshqJ33wcYds/NHQi0LU/nhv9WruwpMw8zbSiUZ0DOwQVTVECl251df
EW36Cw3CJY2WODwmSmGG26s55q8Z58GPh/yDTIrrevUVUdbs4JjvChoOicsxqP6S
SdhTTEqdU/vz1N3BEwrauFmq/PlJ9j7+MtXlojsDb17A5w8Xxah70LrHbmob2cr9
nAyPg/ahnMnHDJi28ax7DNYdUF/GeISYwoZC5Jb0K4Li9u3JOVU8zDMSeHuKQS/2
veUkbradvVyo0vttaE1nt2cDc1D+UahkbetyCL478d6QmLWie32+spUtMmduABNp
agXKewfZUFzE+NNhpRdu21n/0hruK99T3XaoC0Ptj8LOiy+GD7TPbHuC9DNZ35fu
UYVRC2/2l+sHhi69e1Cooz/2doSRoYYRg3cr4blYyJx8F66uxtvohsSfPf/L/rAx
NZlrd3v3hSLSoP0ztTMzO7y4uL3KaIOSjbc5oUbNRqX6qXxEO7ybfaTDNJQCh1Eh
NMcm2PAJog9sCwRXoWirp6VcWSkls4/ksPSm56zW67CJA8gviI+DfVzTC3jSoru8
7WhPiab4cBCqzLWPBmVZt7vSo1NVFVPsSKyzwA5e2RU7X9rkcw8B1VrqmgoIsBBu
w3Y31prpfhd6jemhQpelCt5ZYLnvoKjFkKfyWeR1yT/bvqrLaYrpKOMApsJFLnQe
/zTA8/WOzCigNmbC8hPGJTV+3g1X32I7TxM20S9V2pQ1kJUdH13FWDbmde+z4MJz
cwny1weEdPYk8Qfegk3N92qcy/vI2ZOQ5Tf9gPPHDS4qnUfS4VMmVZmtD5m/fPAn
BunS3tDhE1ccU275PXVn2zOZt7e70/z11yWftslo3lB86BQWk+E6KUW4j+Qos1DL
AYGH99ob2tCCkVZ5FFvZtrh985/59wqsRf6YIEriXPKp6+Z8Mfrypr3GE89wWUP9
8p56ndfIODmrl+z4uyHZgx061pFDCc+lrvLtzjOvmOS1jAK78mLIlMo8xvitJe4M
Qbu+M4yYpVC7zmKq7yMtat67JqL5StwkePvnovhjp4PVC5qLCqtFV3FQ0gmqJrMa
Px0WioIv1AHaV0l2ZTSrbSOO+6aQiTZFKCiLoONq2Nz5ksuDoWmD2W9a5eywiPkH
HKQr4Ppuu6XcF98nxhzWGWR9gcZaIrDCGzwrLMIsk7MsOOlK51Zr8zaDhGlni0hO
myF9JdngIO/OeOpk4KWGCwswYu3rYifL9zX9XAItst3K+EPuQdqwwwVo53mRcKHY
24MIxg0w+0t/tRkLDgoThWg2W0alhFeCvCz7sBE4pZNn3tjygDnbZNtw9XAC/qJF
KHLdWQxjs6s2n2mmTQiZ0y4ZzcDPxTuhE792UHyoyIsK1N9mjr9jmyXViE0x7d0r
4S//dBrbmX0nYfbMJEhrTxA1M2Zw6H3JaaaYxuRRtu3Rk5fyVT+8BMcZyz8alLN1
CI3EElngY6uEqwiNoL+4CRtJlm99qEkls6Ogfvb4dzTs/SDPZI8zPoSGzmVKYrn0
24TKiOx+wxI+7oDFlLobDiYvsUQVl/tQxFyIUO/I4qVS3Qc+tDWDx3xhevUXTkz7
4pbozuyPYXONfz+U6OHbT+FWKUj89LbMNJvwQGNvpa3ISRBfmkzcaM2wN5MHsOyp
9Jw/SQ7grBKuEB7VQ6e+rui2eBgnvQxwnshgG21hFPgGZwgxfAP5XDtwi7e4+nqs
VxQBSvG6vmDZGWxaCsgTKpJzhAQqh5cia6lw89WBWu30+Tl/utB27rdoaxFPyfAp
jdIVBvePrY/RRyH/BaaSzrfbVL0YMrTMh2njOw51F0U6tdP7LOwXef50MH8EOwV1
eof/ux2xklKHMG16j2bq5J9P6AUCJJ5SfaemSSZ9wwoGFmlbF3nfW/iGpSKKgJY9
eVkDmPcThESCMY0zwm6VE/+YBdmkJlpuw4U/EiqcOg2YmqIyLeXADpAQ2SRv41ZL
/cnBnIRIXiO4NkCI87FND3rEZzWjKYgm9Q0gUXJ4wADzndFyK/CYb1InmvRMmgWA
PBoShvFDKK4ice5ACcQZv0fjUcM8tIUvuLH1OVhkjb35AN6Onqyu1ZP3zApPTbre
WwiTgR6grN8qYmEEMBwbZe/AJAUtRKkk+F/vCRjDp1DeaKw50xZZFzRWl5p7nV37
lvBQbrG2W3Z87cQXqqhy1XZAUVE/6CHtCz/lDIFomBd4RGIxRXj92GdJcqOyw96V
BgOUKvdrWHMzguaYuWC92N3Xyd2EiyrebiXHhxzZ1XWDKaw/kgX8GCfhlcuhvK7o
5FYdu43X6fIVyZjoWNNqsuyBEj0yx1o8l4ubzYIJsnATO3PEfWYqW27BbOu1plbv
Y6OBdjd8SGKoBpuvYylmdz7nt9wf/UOquAlSID0XnBLWeOzcpCiO/DvSg+/JjZIs
udoXiFlNnznfFVmIdmCzeOsUzD+wHbMgALWBXrjsZFMOjzFrHYFG36/7FozaFFhk
X/b3ri2EWR9NBky7cLHqMAeylhDE0R4D9hezthBRuZ53H9M7rlAprLZGdjnKdmNy
CCkZGSuxCZaXKVhE68PwRL7eS2vGDRiaRg7Rg77pkN4OyOiuYjz7DOBLSBvZIq3f
CZoPlO7y8seDDLKBI5jlJ7R5XBONuHmyg3FLSZnyVZm6DYZT9y89dqx5bWbj72MC
rQ0VVy/n31nitCwG9QNL2a7+R4ny72YjJp3Y3uBpumSDusnCBQwgnDzbJVLZqkT0
EZWOz3TsIHb0urjIvTXfVeFsyT9B2xMjNI96+G7gYp5G1AmcO6NhNRzVron5vhiI
dodxvBlTW5Z1NkDl//cq2GO0jp4V01XN8Oq0RgKWLOFzQll0wR+jqO9/zn9yFQiq
+i9jXNRawHtLkOHRLhqZf9uPIR1/KbPtVSO3vnNA5Qq+AtkNpaChiF+2sFJvj31T
vHLLLJiZ7rCywktuUk0/NwRBDcT6u5S71nVMoIQf3yqmRqoE5ukCJ5Pp3v+T+LH2
SAkSky2+1LYIbAAkjsz41eCEyFx4tyRJz7fjfkq/HSWV7/sRE3Pyg8JqbOBC8AvQ
w+cJAtNnnFtTUjQgJxIEYSVoSOSJkwADXP6BEHPAbWf4cc19p0HIzZecRr4bSNdF
gtZEqD7eO4BZUKs9jM06XMfYoxnsEzrSqmty3gCZq/hp3VDv+dVGkAGrTtvm2lBJ
U86aLqOY6zpJnzxdihEYauWe6iVXIDC46gICuKzz75dAyeP/H8wB68ZIo53FsoiP
I5eAQVbsr4oLw4rRMEojxFASAkGNRG55lVJj/gXxmxwmTuzT0QmIoZvOLne6NYRW
fax47u/VhmY9Bn+ydLh/jEUHGIPX1yd1KCKM3+stUKR4LUglR22bljjwc6ttUfGC
GmATjGWUUXUCGiGZCFoLvaeQ0niNGwh+HALVMFtu2Z2+vKov55YmbHod5mFCWtA8
5Uepn64sDHsqB556QpbnJRXD8HDYEKMHnFv8ZXA6ZpG8K1xT7c3tm++6PnKYUTQ8
JoOP3+F9f1z9NmJMsYBV9CSnXL1SL8N3yUBBoYCtzDwZSFajTfPROJccXbUMAtAk
F+j40MbfR7Pw92rgwHX2NU+d3PMpEWAlb5ABBNnYiRtSwliEmJjdbQ9JDOi+WMhP
kZicI1jSZXmx5mxVzPaSNM2t+ktB2zZOyYMPs4yezXxexyoU2sOp75pVgCmTy8jh
1yBdJhq3I/B5sipuOFi3zixQznxhaap0Z2NrBpXEcSTsHNZmxOHxLFqOKzrT8dAE
2g5a5NLJNSNNTz9j0GjaZYNGbmqlAulfI0vj/IKQ+xtum40HB6W0y6uprb0dZ0FM
+jfft//xfgOc2RSHi0OREemVDmRJdOqBGnYZKftx3kTDGL5MQOybxdvY6Hg8NQqO
Xl/4ufjyTXrzopaXN6tejerx4n1KAql+PDTPoh6ZvjbOClFJZjuXkwQh5jNKZnlJ
gLUQp5OKd3l0MaA6ljlxTLDx8S/Rkxlv4Oq1O1Scv9dbgPdB2qCMGRJrNZ7yE5NX
vZLDmuJSpOtQyWyxwshhXGO1lUuFOZQL7jQrBusX86Ok5UGp3VThu7Hz4f7ivblj
SkNCPhBxiB5ylp+BmZiLgjyrjfk+qJNRoJcIth5dOxmmsAnehKzP73KZN5/RwzDA
vismeI1GKInplYwB2GbNsjSkBfk0VniNpDyzZmfvDmmDEgbrdSNAr7nGIekObGTA
4jx1Em3/LH1OjGUXQiZDXblLuWabNyR5EyOfIEwA1sAsBeYXzdZDqiA9NsUcnwXU
aQZDBeHh01s9tOd4rgRXgcWTuSEwmcs+bWr/02Iq4j8c3Jxki6gjf21fOi/AjBFw
EYV+n7ON9iEeoOp1bhGMvdcxTByuM582lbFOU3vqcvqJHfeiqJ8WGqov+9ojJxrz
ZKVbkqvfX1LcYdfksX/tcKxtQ+5JFfQHNos6D+heous+jUbM1oPp9DwzVvWtN+SC
PLjpVre1k1eqoem88CoSm4ZerH0OPZ6ssEvZ16z+Qy4X1s3HCUeksR9NUDeGIwED
oSCdLCZq/FG47z2x7jhh2fXn8bQD8lUl6ViylQKWGFeq/JQ9uouc5te/5TNDDocF
+pq9Dk4kQTbafsTey0jruug/C/mySDz/0mru2DKsuj4ZRb5yUHIBUhXIKCpxXXMm
F+PM50dCLEHZU3bQpD3Nlmgon8oHr7oc8IkjK0x3lbo5hYAw1OiQAFvskW4F1FqS
TMHN5cd4iUXtWPhnBEUe6Q2W+TlKFSaGdHUGCQ7/Z+cZ0gXlSlP2wQEeViTwu618
VjDYDkdvig2BmbJ1aaoDVCpXwUkfQyZxOASOqx/yXsF3EpuYysfsD3mcPIWgMEHJ
SJA4giwrqh9gaM2xjgeND5fmMJghx74rSBirzelIV5BK3YiESLYqgq3g56xGC67s
ypLtv+XBaCny4542iTl19TzQVyvkjKy5Gx6DPzNoagVdp+cF+lpTWMAOWY5wvJoN
x2SWBBF0XcA1PFV4sriTGdpJVOpbJ/zpke5ohvzJbqJNPEOQVh9LVzH5R4OQJjop
MQgENuCvb9+VeO3QSBO6pZmuSc8vzQH0qJtZNCPHcKOKK9mOzpb4uExTuNbDMI1W
lsHKhtl1hFDP06LHbgABuTjIhf+rRfDwkRIwGa/0mg07S0esptQ/kgMHXTEEQx+g
gX6NNOWz85yrf9EGRwvSUOwoN5XY+aSV7KCHRUv7j+PKg0YVQOlnGp9tkchbXi54
fgThNW+6nFrUFdI3Vn5/P//uUflIAKigCBTOuCkWB6YBfraudv3ZOv7AKWbph6n9
Kpk5aiY3pYmfJuSmpJF04oR9lHkKRcrKPLwaN7+8uYXSBXmtZwwu5MIH3IUesVAS
ZrjmZ5TzUSKsA3KIhGSIXl8nAuSei1k1ffml/GnV6uL3mbiM7FnzDTpxejLaWkcC
AQVSG6mL6vCtUYHRJ4lX6baxfgnmr88sfhMyQZwsjOskDtNk69xAUkx3TptVBlas
zAiELWwMPGY8l9A3Rz7J3yTTckGDNLllXgQrum9kz4LIIv7wPfbFbkyR+wkRPYzx
6NGDyt9MM5Uz2M887xCJzA3/RLaq2TPiqHAVtgX9gY7+HN8eR+1BNGkpgpW0vmLn
3uQ9aJCRXT4P3pR7pcjnAH/EAwIEtwUxs13j5vSIS0543mMLtvnbfvOVM20qGHd+
DJDXKffPbdHrJLMqCt6aMTPCSm3GDfdJfMHHzH3m7cyxGoCGkEb0DBciJO+7+Cmp
Avdur3ndfHUsPUXRC/A3jWPoIx4tU5AXr/W32hNb/F/oDoilXGmyXJZB61posnwu
jVuBKWMoePBeJCW6UY0UAW+SGDWsPUX+kDmpG5fNuOYc0gVaZDUj8D6cHU3S+E0i
pqNnUsS5NSjz95C//XUNFGsC2l5c+3rQsd8yKep/i3FCvAhg+LD+p06pGRDI4ciu
FXyRgBZ3HGlBwLN2rJHx4LHLP3+85H8zSZUQROsV5r8ZUdEVxz5MmrCSUKRIqIN2
7lILz7fg3YCVMNJQlHhn2MNyBlGgoESBzYnpfWnUrgl+EQcVdphOVX0X/xMjXZis
hx+Oglv2iwE3vAN8TculsHwg2f/2vHiJUUAKN9+vQSILsfbBRlHa0NU5QQR1lnDC
s88nlbAjfqqfSQTEr7CQ0FmJ2sqcIq/1Chg8ytBlhy+WrVj/BZ+uCtNWWiYWdxRp
fArtq1MChOfkNbs0OOVUWqjxeSbrctBLeivIIAyJiJCAnBwnhI5MNEv+qMG6F++T
bJiH4G5YBCKj2o4PlDdIG0gh2th0Nbeo1+TBUlRPghp9IiX4idMy5tMZDU1xZbIa
Tzs5l6T+UhY2gz+M6oAyw2lBHK7ipxXRiJ1ZM3k6HOy8PDGbzscj2Ax66+NKUTsD
VDA+RyD4To5JmrtRAP+/Rv2kHF3amQoPDa+innRqZo+lfGSx5FCGP+VsBOwblx2L
41e9RzQOIvfc3TE+wwWjWo6zc1E6059emPBzlBEY5XS2KJIUbpw3kPVIcFHeObEp
fNs3RnM7mxs2kj2UFMVJbKey7TumJwFQwlRJY9YYiPSm3kFuCxQjID7sasAwomWD
aeE4UMBRwIwFjzU8fAXLUJ7BYaQFzGKESxaz+bxBx8wtGnuW33Gi8jQyXktDDlsB
vtIye5FZcarRzNpNJyu4RxO6GY7YQ7NSDNtUs4IEVAxECrKPpkOIOfmqdYZR8+3d
eHoNreMHY6YpGaERmjmRIXlEXL9W3dwtsW910NuQrPc+DeptGs+HYscD9/EkjzVS
gBDfOIbKiF1HXULxwzdmGkR8+cict61Mne4n/i+DHC9t+PTpvSOSsz/1rsEgc50n
pVgoIDX+2KiYMs5YlmGsrL5uJ5VBsU3oppSTbb99Wvu8Tk/XPAL9rg1m8J9Mbj83
HKFXPmaKv2LXSKnLu+CjWQkdanxNwpLt4Ov5cPB0yau5d29CEoQgr+NMC2ff+7Cq
wcT4Qzz1Yuj7wMt52WOyfEpw2rSRiS12CCdy/jc50TdK4LitIAG8IqgonR4gCgkO
DhvSTt8y0FPp1YJKtinqdil6DBGxBQJbrg7RN+L1jK+cj0Ejy9mTQdyZKvhSFBFs
YW1VnqdgG9r2o32dc18cmIO2r999J70eUM0M9FTD3Rb70LUQLYEqgQS4oxgQRvM2
0bvd4R6LFUfhoL6ctvFmczwBu/3ICbkRDKG1+Hvhd1P5A4FfqNZ2Ny1TOwbG+ucH
EI7vp2ipxdByKvTQpdA7fsaV6SKJRajM5W3r2+r+I2LAMH43YZ+n2RCLxcH8HLhZ
kZbnTKbjYeg+xKLmXBbUt0QsyXB4XjHClLFyH0khfOW8vEzWRPjyE+yrtBZ8Vrvk
gmTf5GSlJgza4is0fbBpccyuh62JdfqdYWYsvXgTZ49ex/60I6k7mZV723P/9Q0s
gIideDW/NmiB1XzpO3NRggmqZ1yN9OKwOIevN+0mvZ02/d+iuUvTGxPlDbOyL+5d
Tn987Y7sg2LZr5VIFTqmP1GomdvKvYqjQtKgifMfKKDtLQJKHR8YC+Ra0GHzh7Ib
+cC1DxBDaBmGfb8pKmO8rkeSu9zOxzT5ZOZIZ1YhP7F+Rc1+3qRTZyvIIlW7vGXE
NTV6i6JViLfis5wnptceJM1Y5/azbiNW3WZ7XP4AALJf/X1+WP0eXoNHw4kiLXIN
hGIzhURPYr10gDjX92oWj3lAEbjfflelKptc2X9cly/T5Bf/0Q+v4t/8nUXUUcjN
MvQ+xuf29EH/Sf6giF1Tir/8OWTQAb5eCTLqxEGCvnayoXmB5x+AurFZW1Bn4Rkn
P2cnCHHiBuVJEE+bfyacwri+2MQ9uKPr1M7yLX+jQukLYGfNgOs0uFiwBwmadU8Z
RlCVUnpRcavIsnBcsF4vtnXijG9JleKluRFb7IQL4jtzKg/28UIMaPl8NzFueQ7+
QSueWp3dJ8+uk5oB7RXWC7DoRue8Pa9K0zBJVd8fGaEXun410XleQVhWEOwu7Wfv
iUuzH2R99GLzLFrGwX9hZ51Z67yTGos8T49bb4/rgb7gi2PasYuZWP2OhLZvthkP
WiT2ukd7uuzUeMXS10TjuBcsU8bzMRcacdhetVvAXjtuLvhqUTvZRTTcyMMoZbtz
GDdbVXcpoARmTokfeR/y16zvtM2qeBmyyz21c5hU3qqAGM6Qg+n165kB4HnRc1gB
5T4yE3rKrEDyIYCsboDLSGqUy3nmui6nYBurz7vQdrvKrToXKvCHzp9wqpViipny
2yXik3e4pBA9+/ajfDqJntlphw/2Mv4C69z1aUB4NwSPu04cryICmo/yFNWNuqxX
dvLYVoOJu+6c5n9MqHgPf3UjPd9zGY4jS1hslag8G/XHokdEjgAUk59ht7kf23gD
wg02o+UyU0SA7bJgVmlpAp4NtMMMaiJxF5gN9LLKiIKxiCCNXW2JjGxlpIe2Yhz4
cEa0VXB/NwfhRfuqh5zR5s7R/kbioGEfum9hflU3kbjTaC9js59LBjFJdBOjITMz
7IvLJ3EKnwPM8bVdoZV+3ac27HOEBR/KKiCM8uFC2YUq7O7sq+SkVARn5DAaitzz
m3ocwZ4ET/402gcOVdMU26/4ckrfH5WTxHlJWHBcSDvhBeD2PKi08Mqj2HlsYBxU
d7s/91J3FkraaFu0OWq/yAWysDAV9840nnn9iFwlJuyxEUOIh1eTJVM5kSzSj+r4
kzy3UjfJAxdW7hpuGkuv7kAua2FnQJVdNZuS8uGhaP2iQPDZO1Ms/BK+OzA4sSQW
YDCztl36/XKfmnkBSULp5rhdRYjGVzYoaEdvg3/7Y4sHRT0yaXSc/QVPbwzsv+DT
zlRa6liBEiza5EKKDRTwIZ8Pb3wMQaJT5vCbttW6Hvs28nu5pI9bC0heUJCRSK4H
Fzx6p4MbEVcRVDwWTm3U6pkOtBL9J8yqumrXWeBPjvmFgdo+YZ7LZxzDchW4VJxX
iDloMaRUQCxybUR5fz8PWsY6a3LJo1d27DNTpN/QmXDvFnq1MLLkpw69OC4kLUeX
8P7xr6ejcuNlobw0OTzVzAKZnp0P+cTq6YRJ0oKORWsKupoKar2MfhGKKvTpk9hf
xiYR2z7+lY7HRILOT+W8y1ZBaX675qCNe9Z80YAvVFQSZfHHnaG3mN8E2mC/GcNZ
iz3qQhErBArp80hpyJubaEmTRftKwwGuMCpEXu2WMLreIkqfMO4szFGll+PD6rlz
+09YYUdB8uTxVYfblCYNn86HMFAFjqkpZ02ynsfNpkS9llA/YKi9bK8i4Rd+TZIy
mEwx13Frnl/2ttR86nDFWvGMgJtSLVfkLYza7rWL6cZUmVxjL7Qn7c5Yb9xp9EEn
bAbDnkXXLaFtH2OIKcv0oLhbM9xv9LdmzMurmdvWpI3Nz3MQuNAnh0BoTVlx5SuM
zF0G51skQxVJd8psd0SVPWJm4iwB7BCdG5MTyLzvYbfc4TrADyJgG6ZkuXdUObxi
7HJ/zGZu7ssUMRixYwHkA2GWtA+8K/Vb6wRRQAS1rSqMLQAx7WQIyxjSrYenmE+z
zUIr9XiaubNIYo8gn7dPyW096kcSlxb7uVjSvfwT2RgQmE6/It+0074obtIhm0xW
3NYKLj4oGOWMjYrGqxQrtiMbFvDjJpI91sLtqSZBV/fFCFyV9luG5i5Rvdt44d7i
kAOBRvLDFJOfekQCH/g8r/DWRdQnKyP+APLh0BsAdLiXQ+ABODUsQSk56eJepv9z
zUek3RpxFJ3wM5nZEMCeVFeUj2hAi/Td009tVohCI1qs/DJY/tiRGOznUG0rhBpb
elnaUQ9oqG3apt+bO8QJMl7JjeM040PzRs4gov3D18BVnnw6ZB+ysvSia33wo+uV
O+4OC7+2QKWMCVeDlV454kQ3fpdpZQmDFIotbL4tmFuUn35mZb+q4NJfvwsVJIlX
LjntiWhUP9IFWUiRqYpk9UMjioy8IdMrks0PYbqCnusrYgsH5nJ1ncN7cOCrPhsG
YG8+RMlQZ3HCvk5/8ISS0LFpai83LExOMI6c3064g7FGrDwqZ+OTEgX3PsEhRJ+6
+q1RMO5SqyAzPi489xY/yvXGKqPn5pAhy86ZnfTKFhIDmsT4EIYCAPsJYRJjyq2w
wbhQb4Tb1chY9WmPa1JYc2qqnM02vfiTwIoJrD7xF8cPrc8z2mEW4KpgqY012wuv
bW9Tn0h/xrXSKXlxJ4BgSLyCfLHNPq/CJmdIz0K4lW1LHBlQ8KWoNik6Eaqcj6Io
qvpyXQHBFPvCboyBh8+K2Fip5SHDlot7KjJEHj8ku5dcFTyE0+FuzKsexkhrA+Cn
l4yTG7TVIt1atm2pJ7ym0CLgyRPMfHCUithb4FO+XokNmZnzeJsR4inbrrchVlbo
F/myZIdgFCwYaXodGh3LrI9GQ29KblDGLwtZ6plhWaRWvg6ygF3QJ6JacT6e928V
uNtF9OTVgVrZy1aWamSQ/UR4UoVLOdIOPksVxG7V35ryxX4p1oyoWa9liSM31uk5
CgJIiL4vi+ck/4JTO4s/mIQ2t0zoWk3BU8gDno8TZSkoATnM0xwtvGb15L4PQXDC
wTUhPbsINhnBCxV7ABcbvrYQ44AE2lNMWWKzlSmBNe/Gfoeua7UyA5yR0O4LVI4+
olIMpY1dRWJp/zwg+uX/KdCMUJGDbIXxjf+CIoE/pS1W9hV6fjxunTAHI5CakCNG
fiXanlHuIrTovfjbE53L8p1DxHSnntIzjqK4LJ/H6sWOFZGma9GcTtZrLhRigx33
kSDGIQEWSiGathEsYceR8RIXh2jnknmqFjGXSEg8U12Cvyz9Y5qhbe+mqlPw6TDi
TWXcD9gOQwwBFV/NAt4etAmXnJIZg26TvtULa4zv5EJSqXdPd61wMTW2FxAqMnMR
9l49Ggegl197S5W8IVrFRbsT8FFtY8GEUb16y8iYVinnQUtR/UxUwJWJ31JIfHD0
vN/qxBEggStfTmFUIYS2k4UYDK9ETtvEn8Wx8fwRAQvfEniF9yv0oJyyBV9EjQ8a
h1ojjxlWhVzHhO9fB927J8zCJxwtqEnoN2gVtRUj6Sj9VIZYfV7EJLd5pTZTq0AN
o475jWsQ+wX1Cu+mJyaIEKC9iWQwEsZRLV37Me54CRwJRgtwhvLYl198H4vFXJxE
XGt/xrP0O5IQue5KDwslY4bEwj+xNzyLmNOfgmL2YgVJlnPsTnmTBGzk74nYp2eP
KiTfm1zcRjRRtK8OyM028IuxoToMObiyoG64c6AAB/do0sIEuhIhHp2PZ9iv/r3m
/92S2alI5vfJNVM2Wa7A2URoaYbnhZs47PpeMeeeJRdlkpq2rSottk0eP7uhQA5C
rI6lvgS+DRgC0oK0TC4HTaxOigWC5EJOQzCfTVaUVHLIeZf1B4hvQfGus1Qve4K6
UXnaGhselWJbf6nM0KQMwWRPC5Gemka/qjutqeiDGEf1gh8qveJ7MHa3nfHovnRQ
Mk6n7J4lY1GecqX+gO3Yj9j3iuZGEjQvugi1xvTo/tJor+RzQTKQukoTOh+nc1mG
rFSe6GynON/1tGdTjGj+NGkTB3c9IaUPWKqpK1L7+CcDio+Ft/6L6iCtBwMbs5Sr
R9TcN5d6rfVMu1lb4Q3HJCOq43eVBhsYT5XpssEmwMRU8AbEMAbQHMM/1kJ7M2v/
DZF8fY/Qo6que0EsLzesNeyK6Y1QXbwBLqQV1NoGesBGnwhtvvsXi/N/+deSXfSi
Vd1DJJ4UiUXgnARWUQs99QV4GPHmhNZ6+Q59UY6gtFGEn2T+TgsEG+jCdpGqoj4r
dqxAvh/ETe3SWoqrt7quaxBCLFko9yLqH+/J4YckUeID2aKMZt+tWKjXk9Pmwimh
lw1ZsoPeGXv0rIYiEoBpx8QkklAixxY7gtlUDu9QN9EX1E6BGNc/jT9FGrx5hAK+
2RRap0VV8iGQtdiHkJx7rdkPZR1N1tp452tumO/5zDUVHONIMc2NHJlPO0F/dhbD
ES6vCKAbjQ1J1D+0VwRU1qInabYshCBb17DKKJMl9eWaXO2lVR1Jl4v0L/j/kLtM
3F4F5nUw7T2uw0GptKM26xSFlVj6vxl3n8zF1/y1VnbEb+ddw004Gty45zwzT7c6
/1VATLokt/RDganNXm3ZoQ3hmmiaJVYTEW+GAEzV5sG+7PrQTZns+qkqhSlUhGZ/
VDXNXcTYCpTMQY/29yK7qXH2vms9vUhu1hdnzxN/MB6+47XE5llGH+GvHZYad93n
Y/f8xEfq9JDF09SqUOjH1AuHpwSE/RmwC3ZF6T4tq3GsvPTcFVlj8GEA0UGE2Ouh
TGS2BAU+HxaDYoJhszALuNhvJgo6qzI1gOe4OmNc7MOyYnr5yA8bGy2raIVjSZle
ZmpYC8kyR1WTX+SQg/akzENySnDYXNaazVnTojgSKjDL/jzgruMuiyP31BaYyyyt
gXXg4Cr6zC9mzOyI2TVCIEp0U+NUS96zGe/R9JBkE5X1psblka9sr/cGXYoWcbCz
8W44pkN4e5o2acH1KBF2ps/A2MDP6BfPoeHbSFEK9zZPWg+dngKc1yA10GlslBh/
d+zrh5Uq4UkEMPYQg8EsNzySQY7Z2LmLeFbXfWhyu7ZH3td4R1h+lOWa7zgtCHNn
b13eCppHyA5Q1mD+oVNS09w8fHA5WEgeygST4Goqkacrhi+Tou1j8QVUhLbunygK
gL85oEK9ugN/Ls63CvkOjkbZP9BRUOlqdABI4A4/+MkWbrcWD37eKbVAwz2ohDKU
VmaNXLCWVMaDuMT8m0g/OFubgKk8bzCY1zefMAY9abWI8h99tht4O2RFWBMXH5mB
KXPxBdUxg97t92KQz8TzV5EKpEj37YhsYCacMakKy3OaSpwb/hZK5sB7TPYyK4dX
mAJ/gJ8cUd0rXhBOy4quKddzcNwf0Frov17IMHJtOXgbQAN2cWdBMs5dN3nbasQl
kYjWfEWhvPEvTnnQBWFKyw5AzELd6YKaXFLxm8m8JiRCFd/SZF8yJcBkTJIGeddO
tnjn1A+rgwYF2Sa622heKN5OuxrrFqzgxuS5X+4KgtFRH4Gu0ctjuN/VtwCOhBvh
idtIKUY1f3F4ysBXPfym6dDUAFfsufhrjvvCD7OnlBCgjVeyOpnPJtee20OGNC/Y
ly9sMhSUPojYgE/cahht1vSdx1TD0A8urL+6JuG2wQ7rtIItGK6PQWnNMT/uUIlC
a5vc2dmUNFi2Fw8pbDgHt79Pxu51bXTlC0thcPjo8rmrqfpNIvM+LYQJTzKoMEJe
MnuW5jDWxnkqc5ZeApOiHX8oLandY15s9fXv48oNRKVTRWhw/ZpuYog69+1hseXU
SMJoRWReZR5Pi1HQ8/nMXzdvj4A7pCHPtHJ2y1Az41bGnY+EwUzrfHTGCKgeXRnh
uEUhdiB6lkfqebbwfOkb8YCEP9Ce/E7sjsgldpb+Etzbtiay+jEoCO9PklJMZaGw
pHdAWhGD0ml+y4SfDAq5/R/noIZqoNE0lxOVspqvQx8BSegaGdBNQgJ4qqtVk94P
zK7VPPLyCvck1MXN0titjXGyLr5i4QDTgO9wOYGsodOgzqySGeprzbRmXkmQT99P
wGRFd3i9Widv+yanbpde4bocMDrUa01MubBhpd1WO++OOkT8e+CCgU01q3Lh75pp
PXpz2Oz/awTzLxU8EsscIg/uKqeIaewFwq7tEdUevch8PWqD35z3eqUmCMP/2GuD
+ANI56miwBcMMiZqDG0h5J2eu8hEvm6HDtQ3j3qSik2XGpumknQmcmHkG9CfhNK4
D5FPTUldaiM5+gLPkFSvnvygCPDAg3kWiM7NOJg/UKhnAgXAEIayDO6FF8lO424g
kOMSMuFnTZkiATTpXq2Iq/U1FPMhbjwSVl/URJ1nqW1rZ8ZRg9O0ApD/YEAJ6Pdp
4P8pCE6OAB0mwDnXd9WqvImY5gwdI4RusEBbGr3GgLsJ8/QaKRir77JWNYqQWBn7
fj6P/OM78iWxv0b0/Es0aJw4GH+TeSIYelIdy7M4HgpoIR1CX3ziZt+WnVnJzofN
h0meIiDop4Tywyw8tCuu9kvrs9Ke7/KTnC7Uynw3qbbxUobpZvlf+r3vT+JLxmTM
yQmHDIzayQFb5gmohLExiC/MNkzPeG1PlFYsHYB02quXWsIRx1BoKesKH2y0cvyw
II3fn1cfRmiOkox9GaEu3Qz1ZFcURFqTj1UTvkKCFDh3pyjVwwOUH7ynjeFlnA+g
59Y8oi75Ko/evCiJJ93JNiCErq+sPyleg4CZba7u0fWVdfborl+6W8DmhJIZ6xCk
onU3KrYW1Tfxgrk/hCGehmlBSt8KDRZIMmgoBdnQT3rXkwEPGsV3RriOxzMGtLHu
q032UIuNGVFmU/UwewNDkp4SjQSvGSH5DnlZosk829jMyngVrIUnIFJjMZI5mr2t
+QaCpfj+ScdY1ono0dKAjMy0wIbaxIWHIqtcO/SnDf+PAWsNB5IC75S6xE2MHbSM
aR1VAlWEFot96mIq9u+Dx6xAYL34L6wGGdr6im1At+18avIGTpQTJcprJklLlhOk
jzagXhtHHt+a+jP6KOCZeg4XAfGxAB/Q3REwpfsnHyWAHlx/n0g8qegLeGLZRkhE
DbSDO1tWIzw2/cvJCbDoPR2Pepi4kcQ4ExRLnihGUXNW1+3Iv/bTTwsX6dZQuj3Z
FykqQ4gyYFn4nTkk/h0Wyz0PeGAbDlMSBSfTokAzYc2fWUqV5VZRTvfzfbDqHCog
5Jw5h/znok0TA0GCE7Bkc4A/tlHq/qQ7DcBZb6xYv0qIU2C0xQ3Ec/Bxv8sluNo5
Yub5WOpWROZN90THojk5W/kJJQiy8UJv4o40J5kLh+XWNyOth9UDY68WrYIZuTIn
OBWCFGRDxz3SthoEg5RMieRPKMbwvFPZXeFEY0d2KMfXVYTEpxaI6aF5GToxeeYk
Y2knSVMe1ZUQTrCbJGiY/eQSQSn9HWlHjzAfG93WV2emIQiyWAjnYxW0B7Q8doII
cONNvccbXI0mylUT2xAFZVBxKIS1j701/x2TKkJ5fQmEkbfUfgjGkdu/fN9lyj7v
gH2twHC3z+RRMKFE/M7nnCXXszeOHJYFoaMnsGDgPuatTbsCCkBJ2qRIMz+fK+K8
VpSeWLcQAUJ5sJD44YAYmpyYAJi0oObZPmw10T9bPIortUo8/U79xZvifzZ1A74W
oGgvTbjAHKrC+cVjArT44fT+JY/SxfOPsL6yVAayLsZHwgBY49wjM0SYqEB/Tmbn
HJl3+VAoOK+KPH8IMnXJAvTGMCr5cLDy3Yw5+686LFRysIIFgm9RBCFnxEzyh5jX
zFbxWKq/IVucayUiWVwGrp6mUW8M+IU3nzy0VJLRdU0HSFdL0dLBb5ZOc+XsSm+V
5ySpWS1PglC8Qo92GA5lqTNP6zc9vdwwT3suBXf/7ZAhedbFx6NYVNKwO/ZEgmQI
uzyN1EWsmI6DeBxtwJ4SbFlfQTprKKsR8vUkkAKzRa0ba2Td72lQRf4wgMZd3k/J
YveX8ZOtLTij1iytua4ajDBenvA+LpwT/xjy7obf9qJrFki3xpB2XWrTTmNr/F7O
+YtWSF1t7h6z3VaGOFhhFRZ+3GT0cVuFmN8rOvFUmUc0fMaygQUdO1YZN9cvL27h
o+0flwNHUO+MK1wb2nwy6TaWk3GpTjhuh/apc/Q2dEBVeht9pqXj9ObzeiqSOQcg
Ax8sMHueAodjYdcAzs0Do1nYsJMzZ5TzTIfOvPRqxzVoqYhb57scZ0iaetxIzt2u
gERYsbB2/C+gN7QZJysaS16mY3h6ol+AzH+LCHvXQmcSrEkPkKaIBZKcXzU3YH3h
VIWeXCbHJGRMKpOtfiRUOilanb5CWmF2iHjDmKjRh5cYRJXAjJ6zgDhx7+U2NqD2
D/O0K/sekvwetiqdCYgPMr25pjF2wtvsFXqfJIsp+2eehOPOnE+7E9s+CwlRFcUJ
Lc/kJdqtF7L3jzTDYmSm+8hUtu5pph6zl1CC4CQ8nw9J6trKGJI5W7930WdzdKuI
oOCZNn+hIpmCH/l052sQQ1FnGiHAxMebfz6OZWkwtJSK7FPyId8WDcBo31/1KeFv
9/denmUf3h416JxJFFWKwRhhpGCRXWhCkX5hQY4xHt8/Tv7PpbYfhsNpLTehbhLt
Ekuuv0M6uxjbfQfJyPe3SxFOuAw7UHsB3Mo+IT9U9iL/+8TqYZMq1dagHc2zul49
FUxJE2e6CWfbx2Xp96iDN8mhk9Coa82xkD8/BM3GU3fURcekJ/pv9W/A2ZHM97oE
WDJCd+xITC2+ftdTyQueONGbZ5aELdd9R8eWVq/i2tGKzrYej53KUjiB+wGkaD6g
8ByyWyu/f8OlwRkiXEDqVadcawMlBZnm+7KaTsJMPKBP3GkcRBhD2dFkN4CPc7BH
755icNuB89IqprguQ2nbJjsKCVSDUYSZ5C8WglYUVS1zx6vN3nUxEpLo/9lDLhC9
3m5bKQ9mN2Bu98+YE4lSOyEyysKV88KXipWQXQYgiADW31an7mOJ4uNdHaJn3JSG
/hRGP0WwlMmPWPv5KZSJMvJKR0fjV5VvJChavb7VqWTUvX0/KlqhbZtaWdIm9f1e
Oh4jNJ9YkIY9gkTjx9vrAhY9ii3jGH1IvQS1kxKCH4i+x31RaEFsCES9RbROj5qr
CeGrYdfFkygAa/0myELnjUbgkQYehHDpZjTehpI+f2YIQf6RPujWIf/4beXrgQrV
zMirW+1L/jhHl1PecBuErnf5LM+gbvm61yiFNemZXYQ16Us5hrwFkLBV5JWrhZQm
aYeSrnLlmaPcaN0qs/+aqpHnXcqDRMWb4TVRe9POJPom44llrGa1Rn0seav6tSb/
BAkkpAvQDJRQ6/UVQOxaRezElBOlSVQE/+G0wB6HnexYdST6+bXOaI6CadtK7Qnr
yZgDHbKKyL2b1W/5GXu2PnU5gmEPwyDc1p6XZHJdfawd/+z7fDl4T9ssVtMlZ2nT
t6LPmcueKiBQ+Wq5Mc09qCgPJn4KPpXfFvpjKa8cJUamUbpD1pNbJKCoYEm/ig77
miCMqK8YcdHUcgyWPzYVlvPSm5/OqsHeaVvxlnUvowE4YVJw8Avh6uJNKFEtAIrf
A+8fIqqqhQ8p42JMVPXOhWA69pzQS4+OAkXBK6AyhowITBWgg5Tb49hDXH6dlCUI
VPHlg/7VteZ4ykxPnDu9+LxaWPfDH5MtnjiO6HqPWnc9rxnjSR1qPpfIUd7qTHxT
mg90QDI8//AlEdP1LYB55TUcA0tEnxoq6MSM2p1t1H6i7y+f4MYnwh6+WNAJiwdS
XPOlyZvYIcAR9nP25LJNWBXXv0kape7Npl5aZ0y/CRLxljoVELHh4YFPpePGCNn5
Frm7Nz6dLh5Uz+fdSZsNmQbjGolU1AE+S2iPK7kCwOFMLiAns5M9yL0utCBmOxlj
nz4ajTOVGMygXkVOyC1MhzW8yMeXYRVqkAqSslLXR8jYU28o39+WU+kvnePP13wV
XafBFBac0gKqBJunlkWTRauw/SHew7+4dBT54iFgX82MD6NgyfrXwMUdQIlnwSUr
vdMngrcpMeCBaRrw5Pb4QJ4/2azHn4D+WCO1Dr4RljY3XT1Nwy8cHs9KItbA2jWf
xyjz7n6iKHcPcF+QvxuMtdUMmzpuuuGlMsCmGHrLbCPsFs5eLt6z8ZCVVqRbODNh
3K7DlVzW1o4Ciw/IrnPvzGfRdmhy1LcIwjrxBl9XX7cHfGlMWz/zP/R9qF2W0ifh
bOiY3t8nes8hpxbPfequ4tqCa7VSf9ETS5tmdcw9Okc605tr8cpj+eSOnuLKoWeC
ElMpUrK1PHkPkIDiG+TcCKyPfPDm2mrk8dysyNKQIDGaogQNkA9vwvqe0t0Krqg9
NEC5iv5HNI3xPME/7e/gqaOb0/ZoJxE4y8H/F9ynHSw+sm2UgnQvhKb2az4ps3rl
Vm3nSEKPNzfKSkUjV648OgJKHMpUoej/jFeKxt4UvK2up8+BwXoulD6ds0hfizfv
7yQuaf8kGpevC+ql5vhP8jRtU6aHqWxvqnlejF75R9Bn0Mc3H1sEXCT4QZID77aD
IS76D13uHkVUxLoneO+vmTksxRUWB8G9lKZQ24he0sRlLjefZDfDT978CtUTK+Oy
32jnXURYSkeMHS/FoK5Rsw370QH2cvCyi0eYstqiXknOza5E7xNNVhpbZ3SFqOjo
8+3xRCZrAm/Noh03iHvNiIJ+EWH31Ck+wtFNnr7P7lcDvtQ5N+2gLsKc4Dni/qWz
SMPSgVmmzbIsWlntFM05zz9pfxOrl0ZNrzYqYurLqR6e9YKHBirvBHfBrO66VkoT
lJPbU8Q91N1F2Hl1xxGN7pkSvQjgnut7e2BKKGp985kbDkAlQklE7Jof5bdRMolU
nXZHsl80DI6FYzETZPS3s972e/W39mLYQwukn5jlcfQd/wmRN2QW631vmO0k3ytE
/3l1eV/dr+Cmerchlq5on5gcxUp9EdlIxpUBPvCZrk7WsB+k0QoMSEs7m9i++qOM
0uNQ/+ehasSfmTF14NuCNWqhHnb3w5DrNdCvJ1BUN99Py91b8htQADCgkyRqMLSK
OZQ9NKzfD+eaPZN+ttBVL+ww3xIbj/QVRBbTFWGZ3WIGdeMr31vu5VZeu0CDbsWa
YWVCUw+AzLOtj2QtX8hx/imcOcs+j9vPlviWzBwZA5CH3zUiLTLkjuTNwRvubnBS
j5XNjqnljxgvExDTB7RFwLve7wfiEzHizEFP4MV9tTtng6a+KOY51dQkW3d8psl4
kmiZPBN6waJqTZL7oWSCS696n1ca6E47OTBfIdm4VzsSDVHrRG4VrmuVmSBpvWwa
toskMwmI/RRRlTSWGd0dIUMEqcdTu2Ty5TVHS/d/d3w83VsHe7jwfndjzIMOQhJK
fVcnDgIdjxa3Q3o4/qglsfEHm5Jmg+AnnMsOic+jhdOAAFTgM7OBoM4PTv4R//8J
7dSDeoD3qCvg1eP1ReMVEFXLxbr3N0aInbLKSKVKAS9sOt/1OZ4NyaK3Zm4vz7MG
cQUiPR+daIcsRzRlv/XBK4FyfW/H9a3CbjLVGTTG1qfQC9vdd06aaSb/6wB5de+7
FlK3sduLkNauMmf7UjBsnhKD94bbh1ztOTwv29fSTSnYMLyW8Gzk19CAGeRT6MHH
n3ir9sRD7lW6Vp/uWoXrmgll0gKeBDwZqMxjUMGfTXLYHqdvDP5Vk5+7KRmuGT+e
edE/4LraZuQWBS/So76ezNFsg7aDkBTUVxqHfEhDqt3VwpNwrzyFh8aR/H/rt19D
AIIUDlqCHttriZNtDvcSugIy1Fa26YEL+81bA/DlliL4Bts2/QeycNPX1FM2bA1O
HH1/DCBLmOT4hojxHA2tDJEDffWXnC++MKibVxwNR1GLqB3QKduPmM9PBIu7eMTp
tlbtNzMATCvI05fTOk88hFMdaHXoMbFASRqTuQPtGK4wWbecYgc/6O0+QFYFSbpP
IuMAeXDLARq6KQdbKoRD+Q+AarlqFBla0zcR/x+7nA5VUzOLrJCoHqf7sIyXDEsq
qgOVK5vpF8PnF2ejwPRpIzpKH020nRUO4qS4Jx6bGMu7seIlKg/bpnzo9MBh2NZv
7DAEdLCfSCI9syUjwvGNO28FZyEHOlNtJXimdG6oalSBD7JvtMMvfJOeaSvBTm4m
Yf/ufCLO9aco24rUfF2M5wMpx2dhrI+E/8xDKj/qO9Sk31xI5d3X8eEDMQxHSVUy
8vPmcBDsaWq2QFx8Ib06woT3xAlNM91ehcfBKU6v69iNHtSxVWRTeHy/zKbFSdEh
ICTbaYKREjnXciGnu51G8Zp5WSvMKzfvMX+jyzCWGLASgZOeiU7QhIwMGlhtGzPr
BntOwy1yVc8vp4npS8OmrDnR4luc7kjgAAOnN9XeYToadS3SW/vOQzeSvrYVPj2X
jeZk1IViScE0tVBDnDvi/RLyvsaRXba5NbUunuItpnXhEyWvasXNmEQYi0he4qv1
2o6aVGpEyC5kCfqT0xHUs88fjfr7kALw86NffGG09VZt4z4go42yzFL7eOz2cMnF
sF2tt2wgPAdo4/6esMM9kopSBOvMSN2J8Ba9AGwp8b1+fgIpuV7nvMDIbl/LxPRM
PgMllSrIGmAQtdZrxq46I8VbD7HkClA+jkTl362wjkmddsL81qTj2zEtSBLEPqYs
Gv1h90HqORbuVumf2IJHKOK/3vjUYFmmAwEsy5zzPl3wQ6n79+6LZoBxIlbDP4ay
usyCSy4m3Kt+wLzfNR9DQhxa6XuFk6YVmxBx26LvB3j4azQCjhVjMes9LNVnyp1B
zbnw6+PvJ6b+bO+MLj5zqupgPd03tVJCUK1bBmZjzwZjfC3cHaON3IW9c1m6jyWR
wKnrk673QxUTUABqyU0N3B1JytZx+dKrbvalLy4Go7TjbxzFBTxKSNSsQMQ0DwE2
tP7fbLqRiYwlddMlBCJ3hSjOO0ECDrrkjoBlokrY07NRzdYZA+9TAomCGhQfufWh
rF85hVs+QUaN+XVDT2172gTCrCrmJXYxsegzYjlMoYQ4jLCPzrRK2WbbV+9MQxvI
jszS95umwDRESz1LMCs/mrq0PcK9OEroxXD7TcpJUTYFefy/bhy04EhxOy5KjynW
zoCMGAUwv0RTFHeFaLxlewxZq9iZ3HbQRVbdR10n2pmaI5mzInPOZhGezzkBSDIj
9Q+MBqaJ4dt8ZIC9tiK+DtNfmqvoZloJENnF8nj8U+j82ew6gUO22b7EVMhKW+nA
7t5XOqsC2lNflT8lMxabr+/+rA+2P7p2o+cm1B+HxjuImI9aSKpwhnxZFUJccHVN
C2FaMVhg5w8Kj5GObuceSXNKtDKZRegoORHc6oG/lmX/WVDR7PfVma+Ej0qkZ6dG
gfS0POBMwfldSVTCpEXsngpD4INKHOC1r860g6Dx8zKDaVc2a7xMUlpPRYpXgdq6
jSocgliArMoCR8u4T5rr0/Ys40dSoF1bGDMx4yHGHy9sJA2q+brN7d4FUJdWxr0Q
pAX6GN4pcAuyWMWRhkry8elFKA779wYRC5VIDB+WKKBYmGf7HA9DAep34xrkB/l+
FY7FcqAlcoybVwgqRwvhqE05yx5K73l10OAJXYxr6LPYjQcoxaiEf5u0wXvzzua+
0bSwvQsY1g5I2XVzfZiQ4Ezl8z6EjwH+c3UJNcfH+zgJdLDbmToWSUsuHumTQ6CY
okW8haLjZrFsvY8qUMi6qy1/MiVvVYDrow7/EZP9M10vWWYEYMIaUTw9KvPjIR/y
+3tWE4rvN//lhCICtWHozayZ0zxEyBRh3vlslJ3fN+NNGki3Zw+uq4mPrm3O96tZ
GK5E32f4weM8pR9jE1UpdEruSQVHEjd82W/yb4E4rS9xz+2NfiUNQ3zty+jndOnx
h3bxHgDm0AOD7xEsbz9r3H1sD8zP7YOM00SBgf7gF4Af6ZveAAj/iPpMi9q8aNDp
+3gef+j3RMncSoRp0oVO1PqB7J8zDrnnlNhG3Pge5ZionLJ4tj/1O/6R3a2pYp/e
LZwzqhepuZCEdohEwARdTKi1K5X+Uuo6lWXAlrq6V8kwZYiifA5t3s4j3s0C5gOy
Tm4xhP7/O9DBSB69AnZOmAWHnKRnELr3JuwS4MIwAcLiWhOvle149Z/9VN5eV/NU
QeJSmtztxK6by6yj4Zkq3QJiYUNlLDfT9q/R4dIQ2Q+lbWgT367Ak2O+nUtFh+Ej
NVZw27p85sm5FkUnKAGafiVUo2uoKj49qOH5hh8xGUdGoU2PQaIobIJfJlGfA8AJ
3QaC+DKe3lVkD0QCYTg1EJgNK50dVilz23zTC4zDi6AkbuSmnFJde6OKq+xjpP3m
IIKxokVpBx2lwdrIvQifc5E2/p4xVfPhKMFWYbRCEwKXEQ8oSZJkssGPZ8omy+Cs
ic4GVc7a7EH7Cs+KUmpz16/KvBodXscYrgj34TffVmaz0s4H0Bj78GRVjPSrQ+TW
qd1BLWBs5j4qN8MTdqc7Evrg7vGoXojyxMsbyZZ7Ctps8YIa95VAklAFFeU54spu
avz+pKW0IAuxULABmLd/3e2verBE+UUZjFzbexOPrnan7eIzzIge7jti9SzRy3wX
3SIUWV5/OHHfKW7eCAecbe2TO+IcvO1FN4PUP3NqfoTE+i/TjPUd7J6xaITjfoM+
c2HijEV/g1DlJA9knoKh29/ZG7daCiUffPSNOSaF/280zGcYRETWRJCouVzVj0yi
A89l/E/FlYGqvNQ5s/MJ2eD6PbIBuJTriyV/5CfjnKX6mCFnCYWq1gxeRP84jsJ/
Yz5Pgs7UK/E4LxFRYW69NFHTeLfBippsDcu+KPvQrxBJWer2CvdBZXswudnSOmPv
iN2lLGBa3JDiNUWhqD+nqIHH4//UZDegFP6n3ME35ZohEnxMaNy1jWNswxH+fjt3
kRqaggsXFdj0ZRPftvmkA1H5WolXSAw75EDu0TB+p/RFVLknklDNx0xXWyMxxx61
yptc/d155Tv9Cs3HFf/XKqkgjlFWsTVRpns+3pAnU/LhpqCHE+QZjienHN3IsK5Q
vLxi2NJn6Kc965YlvgOha9SOtngdfZNLOxKgCy91JTkjHeAq5XJjpNOyRpVhdNK8
MD1krKrvdDWk2E3dh13pDH6Ok0RKSyo/8fpigjPRYUqqHSCf/oX318ZKEf8T2ByB
XIJQlzGKNG/HrQ93wzy+TgEli07/uJXE5c3jYUOLCjqxYLxO8ZUKGQSgDRNNgCT4
n/kxVKjFp27/JZcot+botMm/5YhAGWO9XiIucbpDKCOXJINFKS0DXtvbhEF19BsD
YRbaHWuNOCqv95iaxIwwg/Rfd+iWAx+eDJfm22S1mKjfBC1caSLT/xK7IfMtB1k5
K/6uyc+LJSh1h2sqagc2KHm92eoB1ykmsiFr0hEo5mrhFjfvW+b0JZEOfYIeRoUq
smAOiXcJprMDaQoCuuOQL8Fz1wbE4D1LDqmsg7Rb7K1fL/QvkKpjFG+ts+J/b2VX
ZcMLeqtInMTCIRoBoL0Fuvdf6bwAskowskhCHV8OJvdHftsO7e4caHI8c8HsDVNn
Aa4gKxNmCCZKcnyAUtwAQzF4oYhsaxSz293d/g4BYTKjckPrWlT6ldAvVVZ3KV3Z
bybnvcznm3GyJvauLYasehGeerdgWg+20gjqgxxAXKBp8YTicFCuqkE7zmPh9DTc
3FktZI5HHD5W+SDr8ylJsgYTXa9Q0AMjoiR6V8NqBWyKelo3VD3N3UxgGM7BVOMU
OMAWhYUrU9KYO6mY+gmAqHmeGmj6xDHMrWRW5ipyimeQ9/Q9r8caGZ3R9EawxQAr
p6ms1Lv2YolhBQ6of2P87/L4rs0ts3J6qr8xVIeOQkP8DwdnoygWPWncwx+tbm8A
AxKY0E27BtcB4/PF92sCsh7Ne60ZYDXsOzSuk9tvHMdKglpHzBtY7auHnMmf7qPT
bKD1MILnggMA527Fbj8BjsnJculmTTmIlaqOJAV/LR1USmzmeq5ziLWy4W+vD51f
/IKRiSzY/Bi4zyFwdYrim51RkZkbK25nXR6g5gp+3SwQBbKq82iUlpRHDcXz3UJh
VPND+xjm167wT/ApPWM0VM4dOjsk8/sT1Zut/N4lg7LiXfwNIn0kfysKuXdKoVeG
8nXIVH+VIbLL83D0SyXUDrWqxFEPX4BlIqwpdLXrns7F7+wyhhRk5zd3ipAJN9nF
yuog3oUvAZWOOrrVeTGIpw4DfMjf7NDHTx4QaGBlKwiiuG4UCUSjNxLYUmUqhPbi
HT5dp8e4ar3uHlK+SyJldUuS0RbdvGKop5iCSq4JaM5waRJT7YSqvaSyCOpYJSyT
liQbv9OjgAUDyvXMMB3BmyQmQB/PV5o4b5em28MdCaqVwiLx82gX6OP61yEJxLoq
kuXHOwZQsqUpWXj+7w5BRGhobzNYrHPMos0U5Ad1o4BU7yboghzfBF7xqBY7Yq74
SzVmg4xLHDWclfcMmsBF43r+tzTKJPgILI/3qj178UUxVfJSBzqal9V0YcWrCN4D
lsGz4pxCyvl2ewRXGiBR8hrxpm76QlYIz0YzO8pXKhgNdUPKXMPkVO8LTgWhVG4P
IaBX9IiKv4hPA7GQ3R4SvYQwgqgANdDq1oIWaqIXXLA5AnBN43FTZvYiHXL7kCp0
xjmdmiYcus12lYcI2T+xWPmOIdlbzOLffzU/8ywX74lkmcTsdASZRxAXOX5Gcajw
F6m8bC8y1EMTu+xS2R3n8cBQ8/eM2km+SE7WMfMKMXjnITCWHOFAnoIwpuB5kwPH
QC+wLtUAQpeUDftqApkJSM53N4YL7/9vzL/I+W3TqJOnge6rfVgDj+P26kCvhD3n
IhoOyUemW9LD1yC2u7yNrY6Tyyf86cRp9RQ1dy8hxOdOb7IIs3+cCISqQ+CaG7hc
xBvw9zgdZp2vge2MOrmZOoM7idLZmfrtbPoQ0oWevv5kmGKgGxjuLGqz4g2tjhcf
qyDImH4nzXurmTt31Xfcym78sZEzn8I/xzQdvfdtNAclbncqjAiIMPaOvZqjJFVT
NiRGorT52H24kuhR67d2jbO8x3NlBryGD78QdQxeZoCOmq1/5U2a1QVFSJTHODLs
BSMKfydZVoxQYbExDNaPw2aCw/IfmaMRBXX7jk8pnzbsvNmchtX2umRLrL52Ye7i
L/uv9c+Gkj690igq5gBGlZ61X2CRlekP6pgvZCVwjfVzI4gSPiL0OEv5vnjHn9lW
KzHrFV9v/TBrDrwtuk2g6OL6SDwWcYUt/73hgaq9ZftiIpnmpeGFSsAqkbCaaIHd
ZUrf2eo7gaBhO30GHkAdbHy8uomo2rvgrR+n+8alpEEq7CIKGEbNZGwCHlPutzW0
MDVuNnH/IO2yxFZX3HPDA3fxxXExB6ylDpHhDkhTpH9w0grvXl6r40hM4xD8ZU9Z
mfsifSKE4ZlPktoVcCAXhHhVMEK4dSPtAxAeChwZUVTdh47nK2V3Aghkh28k1Nce
WH3M2l+aVWOnHvLdpQYVmh/TgeiJDnRudjEFgmcl3xSKdQMuz+TMm30rmPFcKZz0
5cWlT6Tsjz6Y69JUePO6pVWFCGVU7DfXXUlf1wz8JmSwHz3DWzJNIzhWKZQLn6HB
2neUzh8dWvRNKyf0701R2T41/5e2OndRq/4qUQ38Zgh04zyW1ZY/xf197IIcC4uO
HKdCndfZVRVxG/gYBThKpI4OBROg4B+o+RuVGM1KFA6iSXHv41+LWpO5iF+JjATs
zSMk6retVUrr9hd20/8jMxvKLKyOFLRdS5cLUSO9FzEL7EIjXXFPQgPNq2VJB/uC
RYgH0unL22R+5Hfq6IAEmnAPKUyYwYuh6Y8QtGQefq9aTjZRrwvC6LGqeTn865qa
wCc2Glg2g0r67ziZm77ALs52JiOxMxES37HEtCsNMumRSFbJr2XY/UX5cmgABUFa
H6EEoX7ELWUTDCNbjci1MaUiLHQJhJeDnhjorptWpZyoTneGkCBQqMI9Q1jE/NAG
EJOLroTGD6yOt0QQF0sWjOMLNzd1sqbNkpkiNxfxOH1Ii4R3VvBQXZDdvcOdrV7S
AF39FYS6lA1Y9GMs7LiPBv2GVYZ2DOkI0i+YFjcwmP9uJc35sr37Gk7AYEycL9rV
exE4IV5GsSCmUm0YbyBesSO/+UTzYZPCMtkqvIOLRj9T4E/dcyXvQlIiBzOsCeXx
eBT7oUiv5wpsk+19TRfg95g4sQbgDBWAiyHG7758zP9fLoxBOyut+5ooEBw7k3UB
TOxB6oZ/PK4DzVFDf5iSL0ZH3nuJUr+sisrtx74dRceJnIocgDzTUjwGxOKlr31D
swg4Jwg9EsCvBjCC0snLrMWVyt58cH7Ae70KTy+Y2fEWFuoX/J0po+cJcaTRD7ZK
p5CQ77nUrEVoj9fL7gzvypUhhJRiCUjE02FhD6qIiaoYxUwwntxyFonf8ihTpZ/f
f9CI7bEZOyyYK1eK2iAc2WQR3jcy6P1BLGvDKJqh8FapZLPLaqjGl6Q8A23yVGw6
83WZcolDyz3ZxIQSr2xC3W35Y1RY9cChLTauxs/dwLq+2U9761LDlM5qlYuyV+IS
SRcLY24Zi65TD25MR5VS4zEFv2bh9ccuE89d47Upf989kUPCrmtVtnaxY328yBF1
p0yZZKl3fULqUJLdoa5ZcafZy566u0GW7fftmDdPCe9mIJznPj+2rcUrUn/HDBm3
xb2ZJhdaee68bumn4s96ZsdNWvk0jPuR6qKYRLrRRXWwAmwYKcQDU3v4kXdudHQb
pzYMJjbfzGCEhlofpBWDLlVnUfTvgyLtd5Oe0NEmuvxP3TfyapwssF1fbDXsoSlG
9OMlMaXI/jNhxn27W+4tMFTXWFIQ5/9PHG95yWoM9xW4Qdj/YSCHoP6ggB84agyc
V8OGjU0+88EAcatc4aTFw8S0G5fph/RoWwCx8aJ5dnWOUwIFtWf3BIIAmReZio2v
BTgmLFviZwPkhGDw1vZW+BZOOZ/LLj2krbGAEMhwsU4C77mkiPos7yFBLb/a9jKN
ZotukbwVo9FUquqTaiMZWntYYla9ioygsj5RHL+eKNZ1NklXfAhIcxgkD7RDCezz
V5x5bU6euFDTE8Wz8DWOyE7Y8ya+De74fi19WvcmFJt2pMxK8VpSYUBt4m1OmLCc
yDcRsRt9eYBCFUEh1nFJBAdL3Pc6K9ZeFUD2FjHj92ij8FDvLih4tbauNvnsXCly
CxnIo4x9SpQibk95OS5xxNm2AwI7PsIdXJ9hv7Vof4e7Azes7vssRbzxg4pD5DhQ
+iqpFFPXd4PnIlA0kE8hoaQhKptrOfq95+UStz7S3ws2/mRoJziOvupahu8z6YR0
1MQzKApDvzl3UhEhJguUwwWwhAM4v9kstAaADd+VbuBF6jy4OrdCLL7yvSFqcsNX
64SioiMueBSg4IsB6OEhbOnAvjUdU4A25TebAPpnjxITLaJ8TR3iWEwwx1jskCXy
Leg7FtP5YHGA1A46PwxIPlJMSiORBlyUcaivWMnn2SZ2sIZeqDoVnZpgLwJM0hBx
fqGSG/SjVjfyumycrAZC06x6D1GsJcpT5B1PKx4popIsEqn2Ra0lYGSVCNsp5g7r
C9o/K7KLc2j8x0xQn99tyA7n/3XMlWUvMI9vARDzy8O4sQD26qzanO6OdRBZvoIF
kyur9khTBFkYQneA7SXYRMraBG8ZVf0bykX/g9h0ASJCUl109jznOf9RZJpFospu
ML2nP6/R0cGb9bjmWtgXXFF5kHpmSqq9v1Ig/tEJ2HBE5pY9moDfqvqFL+l3QGez
+DcLH90A/U5D4pEUOS4G4E7+UF9SjHNBAapbqOhy1/xriKxMnXFTWQ5KyvPxPZqI
1XP9VSwnG06C3lvOFnhEgjyaPCKR3IOO3qKFf2QaosKBO8WTlrdhw0Uk1VnypvSm
nzRE1cpMEfrCdUjSip+Ig1Q4CdSGNG0SOyJY9y1KcS0KtKvjNCobS96SRHlFoh7R
eLqBH1dMX9oEVfe3vdyNxlUgavmA9SQaHDFGYS6QFugOoTSH9fz7wIBT+HGZsD5E
A2AZInGQIi6KmdhVoRgqGRcDOqRjHwiseHtvDvhLA2mOP03PNY/ffX0q+BTfXWRI
vlfxeUFuWlyOjHrZCtYJCAJ6uQEOIydNeux0/NFiMIGKRdYKRXeV8EKlrsmzDBl7
3gMpo6fiig/cTtT+73/5eqtCM40YCyYetiGMWqd/PEDScvA2sriz5J93+RNxDBm/
6theCWuOcGIALIlj7IqWPQrEa+NQpvardR8gwuQwWk0hIXPtziowj/SCbT+DAODw
G6t641Gx4HJuNAiupK+XOpPjL/iPOK0Cuv5fRu9zkuC+ZAicm2iG4iDKBxwZGnA6
6DpaU+Di2D1cn5ddAUaaBc8UKXMKLspY3U0PdSgVsGhZ3d8hiczb03nPt3U2FYDV
D1U5ZRbg1sHyIDnhKxZb04KrS1VEBASHjge2O7+QWTaZSNP57k0kxLTWC7sinVNI
A7vh9uwwaoMxXOFpdxj3Uy23sQQVCe4u9GWTeR0LJT7p9sjwmI+I+RkW7p6zkcQ/
1KK204VCBAPbP6VLPyLChiUf2+ZEXiKD8xhJ/pSQlKlYMAog6r0QuAkjIGIeQZ/b
EXTosXG4r5rzZW2nHa7EajkskUYQOo2Z0ynObHLsiQHukliB2FBVx/LLo6aow9qs
yv0SK5VQNvvonB5ajAOsxvaVNpKEngx0OIUXhe4MJb1ubRYAXtNKOlTyS0VsZaTS
8udhcgcACa9UR4aZv5zUB2Ntw6wxh9UdhQqaTDHxj7dCtGkjrQwqKVDbTqSiQlqe
0xIy+g8YSxubCuY2U2rvKQF7lNKWwkGUWqj9B0bNIkqObsWZQwifDqZRjETP0pk9
QG+Sz/fNR7+WEF1K/+qt7UDDnaz2l13PyRjNPCyLhf034uvoSF0GtQBKK5hGXtLq
cHQ7q1ZiZmkxa1JjHYwCC6TpODLy4Ug3AxHfzjQVnke/IRrFTqxATE4a836vUm9G
wdTRpKJk4gUn6OSQwzfEOwm8URspra9MRfcMJgCT+X5Sly18aaKhqSCMcQ+3W6H+
ft/Ggy3JMlIZq4ley+CEHwCwsxMQ3vHqxumqy8weKHHW5x8NQOUfS949xK5EozLL
1Q1S7ZYOqD9lKK4zIcKU6FqE/28Fdqg80UqgETfxe83x+xDQ5svzTHb7KOWHQ/yt
IjB8X/qPYCW24YaOXd/Nk/AoEUthiFquf/Y8LmXAWCr9TaKcp9z3OKQ8sC/NKE/9
7njjBpgtlrQYHqDo19EjBkaKfDOFGw6cAqksXk8NJbDUarCXs5FmjwIgqIrkaRU1
WmQl/MyAaTeXuZiR1Of/kp35vwYOUBwfKg0atdaHh/UrJOh8DtyOV59P45zaW4f8
HgldOz6Aw1s7rDJKZIeSMTRHW69bBh5cZG2tZ7/Epexnq+rK57VvAm6mIv86UyqW
b2IEcO6rGchuV/1eTuFHzBmYu0GDUnnzuWGJYipTudHBm20AC3EVFWh4JkQ3vOZr
r7CX0DDeXupfTvrlD6mfK5KLcMUlVzh5r2VuhO73H0zPkmTHvDWkff443oFFDJ7D
4Rh7M1aJJ8UUfI8lxVWBbbDJ7cQMipfZWWSJa9atK6asJ9Qwyu1LzZKpaC4V7A0I
7bSrNGp6CK6WmCfWBfMJJwVlKXYE3ejWqA23yic9iKw5htOiTWuY318x3wGFEI6t
IXjDFaraI6JLXtD0EWgRU6iGHA04monSMsEZMxHcovTQqZjuQI5IvEUjMPwTik95
9avX59MjX2EGfn0o8hhZ0zNQe9U6trHYfIYCb32RKA5U65AM5DxfIH7MAITwu+Zd
l3awtc0aOp2I53jOZakmI3Zz9ndoHGZ5/12srvNIsxg3zwbUJl2r29U3dwfngtrt
1QsxvL/OgBxXkP35bq2kztJBpDb7HhlUe/zTdYStj78w/fDiudmnJZtsTU0vpwfI
9k88HN8W9wEQXvBNxyWi6PAn6R9ykiLQqQRSA962bk4D+Gl45yWEmLkNNHtvAO9Y
48Y1QBTNBXcUl/SdhwxeL6ToAsFQNMxBO8vLlMZ3YeOanZBSPYVMW0keiOMiEl32
/ioTUMcPRzdMI+WzSHFP7lxUsw4Si25/UjaysboW/OHLTqlGkqUFwmuak15k5RXT
CK0TbuxCTO1tWRMDJYeRyporZey003KS2a6Sxpu9bk8M0QrCeW9g2TApeCMTgIFa
4qofI+6dHPkUxeObN74TkYBgp4mDgJHjiChNbXjoCVPicY7ekLo51n0bNIxzEylK
VUtp7XMu5vO/a0xWAHI0Om1krOQKEei+W2AYOLKi+tsyCyK53TIRp7X6V1dhTWHC
48+8nCGCvGSEpPoTeFNgkGqOxZyiruuIenF7kz5VlGKwsPBVdAIhKcma2sY0tisF
hc7BCSVzpzvY06BWXUicDm9dXlXKK0VotA9mJpPYhgB/ZhrG3UALb5AONmhALVgN
DHFfL1efzvPfqeJWrxo2fV8n5As7tjvMD27Te2dwYE5L913Y5zxu6NvPWrcrnz+r
8K39jzeMtXvqltF0px6nmmOTSO27yOkldtr7wweCRj5111lzTIlQ6t0GWsRpk4m4
5h5pBOx2QmalWlCyiHnUsdw4XiAby8XD+dEsuNz1Pskr5D2xEpu5TcyOh+gIq5xJ
WX8VsqOPpWYf3GzGyOn0FAyHJEHf/zkeEfkSd3dc78fALQiZJMU5qdyzuyD+gDwV
yg5uUJZw23beP9SLG1FlcOGF4wbE/lPfvlPtGY7NzgmTUsW7ui08pKdZAEon5LlE
YZydvmqMFpDU80ZQ63vpVL3v+Mc03i5nhq2BvxrJMnHfPfLKwNaMY0IUv/JMlipT
j284HbkUwfHE/cqqOZRF27j9SAmDKxNWzHJlhOxX8LuyM7RMgHMqJzQwj7fcJoLb
a18Q3UZH9Q/H5gs4JsBcurA15IyfatuSGcIjEB7fNq+ci+K19D+8flvN5D/S1T4H
Kxh6H3K+5cj/5RQB2iEhtI+9PzAwqT4iqv9USb9mDBqPSXWZoz6zfVdRZTNDTqfc
3jg+Snm/u0hE0W70DH10gnijVtiBeFg97kBl0pDqmSXe3NyjvWlnip0b7dRIiCkW
ETz6MviergO59ITuHK5dxBASauiaviB8XWzJZBwLgCU+EdEHBhifAQgw8mows3l8
78STp1EvFSzTpWgXeG0QXENWf7ktxCZZZPCWjuo1uJmQlJMlsoEyoWRTDiQz0OJ+
u1Zb3cHy2Yaeasr7gEqyv0aF2vn+FyDL3lDlwFmq9C3bFRBKUjdHTLsOh9qt+Ixd
Y1CVq4qBFn8xS/KdTWm+7OZFzttkjUxg9qklEC1fz+9JRffB7/HRH/xmFI1St+2P
dpDIlMyR53YriwPfMBpZxXz2wGYycK5xUUvNC/1Y0YkREzvMoJ0QvhAXprcNt4Ag
SlHoNPmGxv9t/7/UU7u4NezJK5CP7bRAHKiMwfhiWehzGHeISvo7OR6//XLIJ2mN
lJXKsw7oHqDphuIUVcru6FkI6mVr5RLEofmjMLhtoIHOhTlNVeWaesnnURiLbToI
srEdYlZRv43/JsgrSm6Zoodca2ZtzAnYbUQH/7Frmvc8AQhRlesbWA5PUnojMTR2
2I7GAqOWGoMiXYLVj/DmNNt6Sxq96IL5/0XDZQ+tQocWqhSzuAFN6JtXMTFUt3hV
1WhphlEt00m5rC5juSWWTXrYKnL2LgHi8KLYi07xX1K5V/ppdaBsxzTdxdOMk3Ai
1EINARcnmL/gtcMdN6VgJa0+1nttSS6m2O7dy5pwVVFp+gVRITUCKRiaCmeWSuml
A0q/Makl0xZyBlFXh/zDH1IA9obQB2uCxSj7Z0cS3mgbPE9jZpFA1/4nAM3rvbhp
Xpe5MqEWd9tZteIqLPRnReFBU6Nmr7yEEExHPQjambbBcqdRllyfipt1AiRYO0iy
SgUGEY4MeaJaFllT8rUN+rgqaOzZXgAWM/AsXeK5mcnvmYbdAtxag3QZjDRj2JUA
etVV+sqxAl/EDaxyb/3xZ7OxTJrtOn9SmlL/+OI+TtqXwlrcqMdk+kZKYNSx+dfy
cjZXIRshRX/0grqeENIwfoei7UR2l56Ul1fNkTN/uS4rFZkx7BrTVMa832yIN9eW
q4rc9WCzZd1Hu2asHNUr9/GmZK0Qwhz8VuTzkCsI++CkJyUGAwKt4JuT1F+XmrGa
YGPG3W/GZG4XII0s1JodM+2E5reb/zALstfDYWQ2UKzJCtG8dkRxOHqQq22zSRzY
2KVaEdcIPDK+QVIJkU/U24gDRtFw2J2ib21KFlBlR28nPD5qHHj1kMLhmxVxmgsI
ANeG+08iIiyl2qiZMRI2UokDsohMiREQ5yglzh8C0sOGWiJVZpYh6XoD93+oSiZO
+dqLh0fGJG+Cf/1BjqFShIc6iVsLoV3Cdjdyf47asvQUHlw25GQVEuZjjruDWbLF
OUmq8OG84e8OoiZ2c5AGWZ7nzbvBogOSkx7F0y2nkwDrZbsSW89zDM7iW3AF7Z/R
wDjTatG1KAmnezzQw1R+faVoYncQYJB/uURPRngytOCYC/B+KrFXt9DIaqe3TxAL
2G1kRE015b74Gtxnf7Z9/MZlF67kp5EAcVXnfZqlq2mcOl6JvBlertHuRwaoPFuw
9OyWfT7UUXpCstn1C22/GAZwzXoBVVnbWJP80kplMXOLDiu8Vp/abqMgiWjy7lGS
oR+Hrcvx71+AVL1F/7NzMMPSryxuYlSNeKX4wquN2OHPSU0/SHQPKx2FXMFYJBsL
a7D/5Z8tW+vEPwTepojnVhZU3IYYJR2sZlONcy95Q53lVB99s6qCe2dfGtShpg9t
oOuh2PeSq7dD9XuHiuze0eRoDBB1tjGFDdiTgtE+i4j2CBwqThdU7QNLPicFQBA3
mWzp3lK5leXh6LdHa6n9bVb5E8R6kw63/XmFND+IScx3h2K8p/JF53m4xrWjSfWD
raYinFn9igPRPFd3BNoaZkoDAeQvyw5G05+G2NkhIgJ1Nn7zGhTclAamT2CWg83I
V/KQbIQsPCyjHmtmRNYnriNxpPub6LWeRA6HYL5VXmleT7yXoNGvh5SPVubs2ThI
pjgLfu0YdZQ6Rw0mXHhlsA6xrigiAI3xyjrW8G/ozxBghkOs7Zs3JQnigm8KoAA0
5aFk2hwDWM748+etb2hvnKYrtCm8kPW/l0ugjmNn0RtQgBKlppEdWo/U3NMwXzKm
W/qaxoa0xQUmDYFTqZsd+HgfkRM3DuMhRMrI0cg7PN5EwYxwgK2KAbQZ1Z+U+N+f
iNTmvchdN301hsFMwnDdIAbjrW84Myo6IzxD61DRk0+WdaMqWrTin/X3sPm2OwSf
696ppL3EjJe2zq/ir0yYfZhHXSfREViLLPGkLRdH33ZV/iWccxbJQWdzosoEVPHJ
lsHaPsSpJZN0tkRWeACc3l5KOobtmdzrzIdpR3DkFrhGsqWkUJeXrWwhzmOQa/Eg
1NZL5dbvdLwTXH+DVotsmtIRDs/mx/vez6lKSC04jpOCKKwrjyQ1hUv+ka05dUls
jj4eesQCcQWTxdSFA/U5iP/FnX7Gha8gw4k2hJUKEnOcs27fI9hVqktF7siQRJdD
W6+HTbeMJEQSVyJ9q903vE7ekusyl2uBpZfly7VFuTk7NGwcQvdtc3LjNmtyf77Y
94nzIOIV6T4P3NWZsK5nnuClPazvEeqUSBaV0nAbwSZSAg2No2jfeixdoxxm9egy
LFyH1v2RcjG3EazZi/aRBHSBOUu/WhyqION6HLBMySF1TtDmfAI2H2n9Jeq3lDcL
ECFR6ZqAPHm0UThrF3ArHK4YBThiHU6AF2Pp6svbzEK7hSP2Axs1UHT15baAPJ6k
AEoPhIXbh5vb104AZQcmc9eM8FtlZyfitjCoyPeW0BuBlLpD5WWh4faKPyG/oJaC
hxERXAYNmh8k2LFEYyZhIounaS//Y+nliemufrrrDprCzyyJk9x12DD1epo7ZJ/r
9D/moyRruLKpqwIiHVFgRSmnVfFCZXl1d8Yo2oEs2HgtMG60Uii07MA8OWGk7dD8
24wnL0X71gettnYu3RL1h75wj5SnaicO0IQJI0Rusl7mUCJi6hikOS8b12kmB7A3
cshYu0Akc5KZqGzhIKzq2Efn3vH455aQBSs331IRz1fogyd1xA9sDUAZWR27Z75+
j5iA8yPUsBsjpIZ/UPKVE+0SjWt/YalPIgQBag34Ukv6UTwNrc5LuIqDtrQ6SWZP
1Xxuh5KPetCFEKenpAZfpbVwMEoJssjUOYKOoR/c8b5nuYp/Wv5Kob7uP07wKgr7
N5owT8i6i8ZE7M1ziIXIkFIENG20lTuhM4BvBzzpK5Uk0Q0z/9idoXhNWs18FZQ7
y4KhOLRXOd7VXuIFQNm3bGPOA5wBfs4RFSKKuCWZPBgPrgiyT01Afjh5k2PKGc36
zBr6dfrUVizVcIrXWLLfMlhgMq/45PabP66v7pMZ3i6HIR27X1ERvY1QsG36OvLu
SBgmgxLNfCMeJYLEYg0J2nIzmjsy//9i643y6FUTLzr6ReUz43VeCe2mizHl6JTI
dvjJbAfDFyIcTHTPqMgvcc6Kml8xpXNlhneoO7TLcldfIFkRTkWDdZimnm6lhtZc
ClD6ck13Kenq65B2qq+qvv+35P5Rx81YJvkJuqrLzCAqiyoGzHR2n7o/64i78oAf
hsiavOvW8Fa8XFk4kje8fsgshv7CHyb5eMxTx/+03hBAUVgxkrg0cTh0Px9rcnBJ
OH3yCRR+xNSG4RyAXn/qtsD1Vln4jrtNrydSgZAw7jOFKMzERe8Otsi9MIU7a5o4
bVrfIPPMgOxhxbl5NzlwVQRwAaJgrI9tv1PHxFr1cIpZ+9dARFKZyO6dXauUwIJz
JRQlSkvxOixuAdcE4rfrMPkrLzUoHM0XBLPrGL7SIofwNtBygucXKfEQhWQ2PmJl
mQ7wM73rqTA12CFpr+NlkMgFnztA0DniziybSbOzZPakiXjeFuyuA7TRbeCnmlso
NI+pV4IsaAinZi8RTiGRd8A0H0JvS1KC4aWUMK7tAkRajCUh4dcSwa5+ucyOoMol
HHHTMGn4Vkwi50O8JbBfF29YBqJV5tu3HcldTHVmmPmnonoVFNOWdWQeSAnQ+fOt
XJfEFh0TlF83JhnTEasiOXxSC0YzFou67jvtgYMIv3oTdnSaXp+GZHR7H2N55duy
/mBPlQvmayDkdNeEDx7lcMn/b/VCbC4mnJNRutltxX7GiZlG+uYFclNnA3VgzIFi
IViTMCgKDJ0GVn94phxcm0WT+8U1FywolMHG705Xiddr3ggtYvfKNhaSU5vhVkQM
f91zMa9Nz2QGDc8qxRYOJKlzmKv2t0pi62OEM1hdF5oXjWl8XcvvzjR6ke/cP87M
VB17ks2I2z0CO/HJe70QxwpPT5dwFM6pizdgCD6NjOcsFEBFtVdRSp246bcxAZkx
zK3pSL2tAEvjVk/CleQftYfU0zVwC8srXD9p/hOzL/HEOTagHOhVFTRxSFdLdvd5
T9BJw14/ijlrBJNdRuATpTkrQvgLF00Tk4FZIzMsnulD13NP298FzW7znNary22P
0NgrohwejjkiQTgeD6A9CXaBdVk1fCZbqsOfTiLX9dGnxkzNlNM5Ty1dlIjdGQF+
KHkDA0CbqLtEohdN2BGw1xy+wS4S17tD0STt5M6FsyU1Dla/nKwVeWPEBiNbU8jY
6IrakIBpzd92+qT67IHpJ5E+joQpROr7kiRDiwZkK4nHhDi4ESpAw8vxcjWtSdnU
ib0Bx7VyjDYQ2bmQsUtmrfVmFWK3U/nHEvX0KiMZRwXtpWragXe+vdDbXov5HJsE
DyaCCn7PC8MyqN/r9AzAgYVhMc1wNsdn0bg4xdcjp3mGnC/cHMh001aVXjO8NIzj
Kth2NNpYytduF4bhIL2b+tUvlkirzmYlv5X2ohRWTkHmwAlbwEndAC2ftDcM7suO
aHD5WWz5fvwAJhsnzpPyfOCW69c5zMx8ooU3SXRj5RvWUBILHIeM9254m+Bj5Sc7
U4nEO2yeaTAsZ+Ou1neNm+NAT2aHsFwmLJbqEQmBZNTB0LMaRgGYAexpIRIKcu3e
KN3oUgpKuy3Qoeu0chZPn60ZheGArAR6u24oBkmDESeO3aIZHJ/GkJgx/bWq3Y6G
q6rexO5RPmUXq6hmkG3B+ghJD3ACXCkGBr0vA89DJADerrKwYsZl48NQOx0bfFVL
UMClSacmpR2f8B/cc+BxyPctq/JO2kKPZWHLyutGcmOVvgNrYlYtLaG5ZAqTLyv+
E+1B/G0bxrpa719JYyVN4yAjSh1MeEcz2FZ+USsTBNOupBXXSybQFLXAJHYAd0OI
AFeNmKQOmtSrWZOHMvV2p50MXUrsuEDTd1dNEnw6mS+7A50aJ1KEHTWTHNm5C/J/
qaH9M6lnFR4cnyhFHVlZXDQ5kVrBwTNUW5F8WldFtjk9RjCdo4kmLr0vec3FPP/i
qGw9b7XohKBBB0A0eYhU5a9rw+ZJf6E+1XmubP+tSko+5LdVMwIW5cByNRoeMRCy
s9J52OdNk+VvUEF1dyOj22hs0F+yN+cTMcC6rUOScOcsVW+W2BSrHB1T5ptu0yNH
TsSF6yDx0xkVjimNqH72C54Cx+JEpyODm/0QyssqF0oY6F5tGYyUp5PbDqBs2PxB
TvkoNjLSOgYhNnC7/dQNKIjH5bllL5zgclIuVph0xWrSLeXgu5GXvW1RtoqqEb58
NQ0M1CWo0pjsCDH2g2aH1brMXn1AqvWzEQ744LXOdFiunRlo9x9ol170hEnnBHHl
yjNf2UHl/x6AMiODhJv15Qe1k8zS7lXZw9sa8TkZWre4By9+LKdIHqWqWRXDPrr+
fXGnn8CVZVXU/2MCz//obZBFAXSyMXZaP5et5ZVrYk+CUxHeg/6ZbUbpoVIJfgiG
/Gp1btR8ynXK5W0h3+vhRYosGHvIbMA7HBTfbOrJZkpKS77BRF8KuEbXCowmRI41
/8VO6EAts6UNgI7rDpAy1t1t84qFotFp7UcPOFEd8XbVXhl5zpWjEeGX6hMaidVt
AIyhK/sU5o34MtDQqpX5uQVACHtYkSnJYyMAz0KJBco3Xw7Y7m8arLsaFN9hXdw/
/bA+pHM8+uylEyHzzxuxxCNnQ2TOPZaahW7khIVGUSsMThlYUXlLKckJeSIc2vwX
R0crSe81j4S7eW2vDUQ1tmWk7EfIQWSWnRXQXy0RY10UWYPaZNpUDlkX7fuI85xu
V4wnlHCEEAx4u8FlN9okwYhiqTTjA9Q6ilEKqXTpsDhiQy42lAp8fLPCIHaESdja
ECTKb1XUpOQjTqse5BVaav4K9d4njp/r5ZTydSfB3t0StaVsap2qgs4P1xKY6QDO
gl5vJjddpL3SQPerGMQokVKFuLkYpnOwB2SxtbohVYoi+8JBW8oWt8pQc+P965Lq
LnvEXU1mhUWG47NK3ddrnx7PvrJJHX77VjO9ADrYlPOaIxKgRk1Khx1Bpv5euvN8
DvqA0cC0IzdEKLFvG94nHYLCiS+DlxKToZctseQlOSEnFnyKlKzNCGugERtUYmjE
LXs26TsjXzh0c+ItGtKAVyqGV4M6OSMaH9PWvK0fcrL+mBYjTfO/FuZgxv4cw9Cv
2cYX44a9E+E5we/HCbxfQnP81nRmms+HQ8lWaoj7ABeSHXm28Dm1gBVZA0CJ2iwe
HEA6MsFWRLNAErdqMrNnp0OwwzGjot96CdtWZLgTq7+6gNACXeF+GWVQb1oKXPh8
LaMNkUKecEmj9ME+I3guaqGaKbNE14skpejIPhYLrJUurxiaa2+wjW/33WcU/mVn
gFk53XuBecQXqY1xz1lVej+rVjCihqVcNZmYqmD53uFHbvGhq71pQNEOp6qmqVNJ
v0hnfniEGBHdJu/KvblMe+UvHtCG9OvOtoze+prIpQI2bcl/l4NPCr9ydehjb6Ev
eJ2n8n672d1mT/iMDNsbUsJ2zS27gmZbkDg1lwJy4obGeBnXYC2rL181+opvLChn
dcGapaJOu7WrbmXtbF6DUAznjZDQfXv5rntGka4/jIHJ9ldg9PBhOn55dLbZT7De
AsrlVvjvyyU1/0s9CKcfKLIvXZWbzpXerwsXu44NKwEzsjgMBvUaQdvufq4GezXI
34KnYG5Akdz8znkZnKipcHDrq9T69rkLYRnyJePPIQuElesxPq1W6+gkxTuMu8qF
BEdicu2faVwR8uesIwVdAc2MuhZZnYNvGz7/M3Xv/Qm1jJIq5wwLUgD3uxWsD3EU
uS7om1bOsfwwxfq6mjvZoWv6OQ06RXiMQzO4Sx1wKAuzId6X28e79GE9W5D0dacU
WJcnpPFsLzGQvaIkBZ1Bsxz3nhcHfHkK9p7CzM8AvvXoV4Xen85TECWfN1LHd1s/
tC4hCGRw5epff4KRt+YdZ9piTj45RWDJgJnz7oUWJsDQ/RnsWUiXtSbtCgq1lcPE
0y3p77htckq07cGlNAtLS+CV6gYLuHbnsEkfJAUJLH3eER/CiYVJSJmGuRA983G+
WSu+5zFZLM9iQmg60is9pDsjCG7zBC7+rJF3aSUPw+0E1qJZCYqtyzDsodHCC/T3
aO6TnSiPzHKMF0mZZZ5e4nBQ4P14dUHXVtDG6+kB6+A4qs6WaRTyEaTRgwc+78Q3
Huq3fbJtc90NF6W8ji6lYGsYssfX+2jE2BXtbhHMQXNH7xAeE0lNO2T/2xXrC2NO
Rdg0HZ33Z/en3z/5UA1HtcblSpj0JbbjG4eAcfYGlBqVIrcJ2LE+KFXHTgG51n/k
iDf07899hJlqF/RF8FQqFggYSoMpedORFaTybEitnj1SIcmi2rDQKxl5WjNWME6A
YGQyznoZgGvpIXNv3DzGSwpij3tati+unMvgzr+zeGeaO7fo5z4ddn6yjmXnfWUu
PqpyZgxw1Wh3xOIeg37eVGxy5fY6bf+piShuIk1SSanO6KdKIw6Bxs+46pDxdRgn
wRM1qGM7HVAYxmYpmbDkQjAPLolA1LqdJbOBOlPZ/AlT1UYG9aaMrSI7EgZdFom/
Aljz8gXOaDk0YhKmogBO6FvfH9UjJv/Q/zW158D8MoNCNpjiXJXsRzR9KiXhbP7T
bjoB93bM2jEjCb91mReryVk3QO3eV9sg6lvmqSclvz7AvPn4JrC1PDDNwyeoFUtN
WIgvjnOr17GN6Nj02ab/PbjGB1CNHkWPzeuCdOvRcwGFN/o/dRTo8B+xwoFaHlKl
XX1DUDgOHUV10qq9SXru34DwvxAw2BeHIu1i7tqzRxNBCseYdCZFHDWAZtphnKSI
ETEp6hAb8fkQlzCvrKHOuC1YmSrSKWmPgMuBPREIsar1EchH7i/+LN2vZM+bGA7P
Dp/fkD8iw2Ok04tJMr1+978ACnaQ0xV0qHPqf5LYxPHFwOo/HROi1um+t/v3PEaJ
sP64xZtDZMeQ/RGDwUWHekOkJcTEqYwJgYnEMiWPnlfq3Lqf6kK8pJZLKRpU0iYC
JgBWOfEgvBTNeRaV5E5fkudw+Zf0+mldV1oH7Fk6+l6OBwX/fEdN0ABID3maIp3A
a2GLjifCx47+SCTwEZfdaaE9JYzOwfclOLPQ8mSPAf7xrcoZkCU8Z/hHYNwnIJYk
Ut8brkyDVfVVJaLkAf1W4JBiiJOrrAA7TPCzjMx9Vk6XhenYaxXP/AFp7T2MriBo
5ks3sFAJflL+IP0A4700t8Zrc6dQKNsNx3xjAaHwzOZJ700zZsLz4XSS6zuD41WO
KY0tVsEoyIF/BQbXP+7ZuW+N8cBEgyl9WELXxDiEvEDTqo0GZrBHi+EE9KudvH2v
79ViuBtdiFDF6I/IO7JJEPlOJlFRCnSpv+utu77kmr1bCrxnDQoMr8jwnb4FTWg+
SEDk62OZy70L3Z2KL4p64O5jCRsG3Tl1U2gQaBDiJNWjBXcW5kq2LY7B7xHC6iWZ
2MoJUPZ7gIMb59q28MyLXfs+JLfkHQJpQy3TwHHaBOm/kk46uqSEB6i7I1jwaJg+
iQVe2Ce1jOxgHslrZVos9AUMkvY4NYS2c1gw8xpxHxvVDt09JTyiOjpwKfVA3mtK
skatAGo2lHSzAYLDlQkvyLWJcJ9oxtO2eOOjQcXCBMhRW3CJWDDmL70fSvpvXCqI
NDdZgr8hjOea/XZWXLs/X3R9b+BHgolklxj9PFsHs0SJwxrIE9KRqeXYBj9fd1/s
Qjm8ALWkJQU759ohMkCrPiYHehskAX8Iwxh1oUSElwF7KbxpkeHMMWbhaMROK4Tc
PLumQ9QZefXf6dlITwAa052eyFq8oJfoDhaMPVvotU+0XPr4GdjsKhFHkilpM3tU
uKjUqTx8bh8zlzjiTu7gGhaF/fl4BeelAxanY0Awosfg9ymv9mIKRogn1FfFvFLf
WtHPIAyLe93p1iGdLrhAoXEaUCqcwUq9bMYRc1WleKSGdf1twN/WU3LIL21ID8IP
MJ0DR9ZwTL4y3gPROZorYO2aOWXOrTSvB26Mvv9GAeJERqdUcS654mjXvEcKUm7I
pxMIfByq6zBuKqmWoTJf+Sxzlr52FnuHojjpkFA9ftQWzVq9tY/1Hv5NWncnh+sx
hsgLCuh036F246M5CE2I92xhxdx+U70XzFf6mtmecjTJt4wjTpleSjk1O1Cemx9V
5ko2fkCcQI25NznlM3EqP83X1Xwvu8D45DLYvS/8ijZbHsDqHiisJWVVulrcG8c7
oRWrWChadnll46dO6AUXD2RdGr9jSgtEXZXdGA9klnDJvrpLd4Wu9gWyOHH0BrA1
pdjgDhcUGtBe7l3PezK5HNvxrlfODsLT84Kjy6fqZUd1PXlkeyAZCV1gN7FU5l1X
/5y3m0zM/id0MpA/4BWf70UdP+Bwley+PpNgHPV86aJWfer2E+1FGpCYiFva4AWy
sEMrzH2NUh1afsxyfpV6b621P91CtBqX3pnrSV0xUiyija6YI7Nl20jhJw9fM4YI
Ffk6+5HB2gCKS6dDtPfI1dxKATVEDyAAaI0H99oWNMCQIGNubDVgb1u08p7TqwQ6
GOsE3fppN4HPQnEnHoTs/YDveocflD1d7mJLuof/p13VLoLW6YmQOEb7JxWtfwB/
dhf0xX1KEatprtxKy43v+/FkI+tCCwY+QUNteOji6R9nABZhnh7Lyf8BnaVFCqpS
kWKFPZqS6UDmCNnVdt5cjZz6jBnjFNZtU4hdBC5mYKfJb7CnuTs+sUWw7v3KFAbf
F6MVaZV8tTSkkYrfrzb0yOp0WEJmC+P+jG+JFh+KjyIUhz/skb0ODZZ26PwiveYo
1EDZTgP32vQMXjxgfKITIY66l3yK0P2fduEmFA/zfl75yXel7/mzWW3xsilh5EOo
fvp3rWm2Cpg74IygADSHl7zYYVV8awZsAp+JCwkhC4su88MRuK0GDLvrDBtqeoUb
lWGO4oq6DQRxpIbudXIb9cbU8+hFUsNHWrzR6M6bWs5s24mzMdZnnCjeNFOQOygG
YRyqMOPFauweOxLm1XgdV+RDj6U+V1HcAADrE0OMgQUcXuorFf8V8Bz/C9SJv4iN
qMAsSNCuPx6HqmyovfYBjpDA6MoZLvsgBhDWK94V0vG1RAqIIZBdilnx6LBsgIjo
rDym/VGOu/uhNZlmFI6P+jSqCQV3JTZg3SfcRZ+naA0xMSB4bxAKpf8/ixUOPr62
9fzmSDmVpNkm5hxEuokHNw/DFMIHLrpwFbK0Ml5S/vwddDWE0+0xOQ0rOTTkC1rr
lYBesMfg4UfaXIIPWi2HXyHvpzMDMk1jqwLws58XPiG7LgyGZsuqqOestv9dmvki
c3Cay2mNMzIZJ6J2enwPT0kuy7+9DpkIufVcu25YEkz4BAt3U6J2tlkqFhbPejdE
deicVk1WosqRho3yElDyzrcfsogDIov2rNUxjCzH7pJe55Jaun5r1nSUS5sM4uN3
ojMswT6H+Kmo9NQ+UcyN7H+IIKG+lZnkHeIk1ezkB/P3KufMkfOC2Ox/VMEyybHP
TjqRmKoV/R8cegEN3tlhkBtITjg3xPT5NC91K5xT60Cfo2zobY5F5SnS5NmELJSw
U9yXUl9mazD/207EvsYwxo/28BFS+XvcBcFX3NWeux8eoxV688/JST1o0A8RmOjk
UObQlk6ICx/rfLPOXaWBex9o8BbCuSWtM2v1pzfEKvzsAS5cXUrxr7tWIJtpHdzm
ZOmsTVd9UmPqRRNdEOwzIN3MbZ7YUzZ25Jk3UaWA3SXr4dZh91YYmsOnln07vj+B
HdkQ6fupJFN4RzWh+nL++GII7VmElckrOT8y/c2yjdhoEUtX/jPEnxaem0rsD2ny
zR37lwRJcWl8i/3M46562N+tgM0iIizY23opk2nvs0GIIkTYWQ0r3BLJxNDTSQAC
De07LOY/+F8c9hDw3JtjwkYMgBIbB/TM7C7lav1IEyDkv+Vy+TfF3y2g4cgA6IIz
fmd94WDcJK3o5humdoMUGkO6Rx2uTfwJQ+RVlTAOxyCvMWjDUmRKo7SODnBIK29R
DtsptoBHIO0gQ3+bCF+JQqbGLJS7HwtY7ennKXfu8FeoNZ+JYKVs1omfpiMfbCvh
gwhQUzwHPXCBs1tTksjKfBKGN0lVsrkaAzyES94Mg36s/I709HTSLIqYV9A6F6ru
C/gevH0i8PVT1CS/rftsQX/ufN2w0fca/uCvMderB48orSFLuqIDq3PBNjg2BE9O
ew+2m2aO7tgzUPTHVRDWlFqdxNun3DMbp39Wl87o8b65QlG6SRx0FIDSKFk6LU8n
R1u3F+0oRsLGeax3+waNBNlR+v+dhW38TBpTWySEsCBfyqUbgh/xr0FkyTtNE6Ii
ajbYpsow7ewVO1cFhDZ8xNxwr7q/w21fw0Ye0AJ1sPIT3wUsqyC8TsTW1DCI2nDd
ivH+B8D14osPq/bS3sU98zej9zUPyX1uYqAuV2Qr/ax4BLSWEIHzRG8vjr/eRMs5
0GOO+4mrmPFBkP2g3cqzB2WL8WeiuEFaDKVH0QrQk76EUHzRUxb4nkCP79qLC9r5
IM2u21M0cCJGEOdRAyWnuxs4/ZW/3QGTYSDucdDy4PfeUZWqpqgvKdHscdkVKpi4
A3vyKV6eSXQMopr6zNL/78QxysKNb99zpzRE8JYbcyVg4xVvLchB/kLn5pPykd6R
cIUiQQCx/yOxgU3P9I8fj9ku0uBTi3e8ThQAAk8cMUjjYZIYeC1lqOxDNJyIHxrQ
bn9mt/Vr6NKmTVE1JZdCcR8PRmBsrSq7lFAqAlqbUY5hU8DNpejMqhtO03EvbLAc
aioFnZAgQX9VFNi7vLtAgK0KXwO2yYYruXI0IH2LvFvN1oTIwWlILMOO3XIARn+Q
iahgXPp0SI28anacY2QY/SyReVnZqztVuPKi86Ifd73Mc7oDn5EzOMPmkeWfc3zl
nuHjtn1fMlW8Uy8Dn9tx7v4stYFB4VNHQM4GJ1GCyhNQ44c8iNvazqzSVO5zJYxD
tZ9acBrsdwkcm3jCykpyMgMfw0/NQn00IRI2TkdyE6Reptf9+tfHQReAuE8EVGB5
xgeiS6Iw2GpOVv2rvxnKW6/iVo9bqBvTQli/jewMXNfJ/STk+xJQwB2RGTCrOrp5
wWa5U8FtB3+uQ5/lEZbR0mX8FO7aDB+kueQ9jnD0XZM3s12YTRCr0n6jopevwDMh
Y4zcSDKdYpqUPCcBL8oHNFavYFvLTsB4BdJUTRLGA44x6svcuD878e1dOQgFsr9t
9uWEzF2mG7juzJFHLKWRoc96FA3XCooxi3a1iKmVwW53nMvx3pUdbmAi9i2xQUkR
FTh/sV/RFsLAqsS0z7rNFYQQtOHkkxBHnKRPNrt+IGNp4fvFK9IasIjbzN0smJiu
hLxZNvU/oPXT2WPMFkqhVX1x8pcndnUrysAc0wq4TX4rJ1OjvWkuO26gTHbbTDF5
T0rc1R3zPtIScJAlyVoIEo2ntlXA0Sd3cyXyi4Jkh2NmeN6WrHWSVk4SHGzLTL4Y
3VrosQU7HH8TlmZmaq7XHua8mIW+v2Tp8AWWKBUJYr/RUz+DC3uKNRT7/BNCzLDI
5rmJFfFXkmgQUrxR2F3oVTlWM5U43efMqNFqdHaY1wiNjBrUYrz1SSvJ1tdZHVoE
9NG0gxEyEt1sIPX7cdPNoDbwJ71aFk2BzYAvCAP8RrnrMqYyjE/WzZO+TSHfMVKS
rexXr1o5JQDC5tBZUUypU/Lb0NvhThfa7PjTiALE/oFQ9g5IITsWNTVrRReF08AP
3GWzodjcp4Zlz6d9g7Wt9g51vEstSgiE/lvbPWHWb1AY1GqS94gwV1kNJ55u/mRC
zhHSAAWVAawwImd+2XTu0AIvw1IyWUfiUBmeG7lqmERPj2MELCAoeIm+NQ26m992
/rkWjVRYmOmNrq3TtcZgizltbBPB7HFMBsa+WwXtNgtkJWsO6YNzaW4B0Ue7ctw5
T4QipzFaGkkhpemnCoz3q9Fau5NUMWi5H+lBV7rVLvdHb27UE2GfOR9/69BknR31
KMTt461MQn/xWLVDhVxEJ1pktAtrZAEKgsNGJTFLtw2SRAlvcGkiedcg4stJMj2h
JZ+P7N5CirgoLdaZayNZAyqgnsw8tDleRYGvUmgPJH0OLeLeMnVl59N5/csDEqAv
s/5dgFI3YVnugq0gQ7PRF9E0ujadggG5GLe8SdcIO5hueyOtPbQOCqhxbLDIhjBv
aWy1izCbVc70Or3r5/5ExrvQcGdm6HHv2o+SL0kN3NgR5PDKTlbNCbmjFmkMQoUP
4Jig3ZgrPe5kbmZuT6BFjL+mw8AKIekzPbdojMLHqJ+uPOdK6GheLoCtGeLbJ+5K
ZH5Vas8ILMWdWD/j1w+oUvMYsnGNaQUgPyc2zSqxDvNzLojeRziZl6Rs0dwEhvms
i63g6fhR+ACewkeHLlKhZCuVDPIdNpjEam5hLDuZbrpSYjgVuh26agm9oQfD5iBN
AVUOwj2w3ZPhOXTcChxXTK6CBbovPRjaVnoWdxkueuDAqXOrQQiGZs2JtXTv2w8H
1Yb6A5VRdiWneRUsQDX0c7ut0QZsWpCvbrAbYc/lwvYz5frJQ6p+6ij+wXe68lQs
kTqDmYuCqObcu+vcWj7S0SnLA3hB6dl77f957fjUiiBaqBGTebMrlngM9jUNzusd
XVLxY953hoHBb7Hn9o3VylMohqAscvz+bztZknaSW6A999CsGN6M9FjDiDnSFgKA
8rbpPRPwxsaVEZJGj3kZ3I7LwBVmarG9CwY2K2FHsDgTcq5AwvwwY7Zzp57C5Y+v
Z0N7WMfNqSOuyKKlTfx3xWGVvsyGODyhBmn8xe8nB+3g9jGUIJ6qNg8q1vFbqMV2
lyiiqDc2krVkqFzEhC1dz0pAN6lX+zDcD1tl1QteBaIyIJkFaowjrLcT2rAxm4uM
EyeVDf1B93k2xRE64IQdLmBLpxN4wjPlZ5ozPnR5PMcmBHx78vAEX3QHRaEsEKHl
ul1tM5C/w0eYFEt2hFHapyVHwjskZ4Yt9fcd8xQKmW0D7eLgXWTW89N4WJXTsCX1
v05JX9ILhOuOSl5+lW8AB9QahnaGnmmEIbh2eCf8TrmRMJXZe4AZ9JXCKnXJILMv
DotUPtL+AzUbqbqF8gNPw9jouzpMVKxYEHEXppQPKhKsC1CIwcgbT/+pDj7xQPCZ
Fugn1pKEhGKyCCSGBUif1OfRoNixUkh5vCUoPsydxoBBhfVgtLkMlsolbNt9cnXy
/VtVFcuYTZUQNc1b6rHrcpc4AJOHpUj6p6nLBvWk89Ij+hs8W+xLT/vyXCRPgXYd
OH/PFbMJjrIGrqeXH3LOPw4Vv1POhzaLvfbW0KVntkv6/h7tb3QECnaOlWB7h8P3
lC79Hf4vv/wATWK2+/le0SsELoS2+XUJRuH17LFJXBNVJb9rkc4fzZOGdb7WNRE3
WAJoi/aRHgKf1s3Y+jvahmGdpdz9KxeydCPRXPdn2v5uBHhX1IF0htfU/Y1/W987
5DFtShflkhoK9j+fKacEO3Zv/LXANZBkaaA0kTwiudZL269ii5xWWpYNbkxelv/s
sb3GP7ok+gB2l4QGAbeWQLoKNZWtNkQ4/Eoirq3QXD5FyG93GEBz312x59oyjk9n
6NeiHh/NMt+Xj3bTVrDdcsFdEoJn91CAIXAsjrM5CJXS/3dUPQIecTqtuIHTn82g
+AOUFGHpHS6OxCZPDQmL4ufw3NiMvytUWKIaKkJYLt56+0kOkZtEUIdehbd5lqUd
s0JbEjHORjP5rWqKUIgtQrB/mbZNZcwQFGV9RJaOs4z9d4BCM9va7CT49a9Wdn6M
ZKeBONHlscjXBYMiwmciuHHgF6WfdcWj0StEmoR72S3HNq5QsAMchJ8K05N2Y8OQ
d/TL4EFqJiqttsbaY5XynS7r3XfiElPJO+ZFCmP+mPrRoEz7r8ZFt1LD7ZKovssQ
4pfFZquGVeW4a1goUD0kcHZqKBjH93El7EilmOHK4Dmyoq75v0UWL4e6QB3+VMY7
2jo269gbKz/z5ChsesWyJmAlPv2AD4yb9LwrsJ4sfuSvmNsmdpN+iybv7oov8bLd
YIS2BDf3juFUrCp4SI7x/5NWGcoALLXuG+5UuEeApUzjrYBL/i/W03QZFLbO6lqw
I+jtDbAzg4sbGWc4AANUL73TZmXvMX59HT2U9/6VNwebrdm0x6Z2k0TagxZTFDMc
gI2QhaD7owVbSEDhSPoDtHtEcxItjSFUrYKNoglp3fQx8s1nIvaNHq7xve2MYZMp
2NWrvLDjRTO+yO5oBacTYevVLeELCfK3uH5fhGr/cuRmK38WsPI3xY4uKt0o3BuU
BQylRRdmA+47LxHZ9ei+7C4Wi2tXHUNUC5H3L2jAmh1Vf/xXVr5S+rU7Yok2dXAZ
xPWG/OT7DyQs5rMX6WdH3fCti0ZWTjO6LR4o+1ZqmVdKPwFU+CBiadEBmPnOExTb
RZjcXHpQQv7urytRynFWPrL7wdzH0zbGVaCVyiE3sJwRHbrljhYV3zVA6sCMYmfS
zDkI+A52fKh6e/WfvOZW2k6j4xq1R/Hqb9CYSlRO6EqZZV6VdW3tcrLi5w9ZhRQZ
62Aodc2ZDHJk5K73dvx/QfMnB6AncO169DevWoXDBXf9UK83vQWyfTe4PNFgNZc7
gRYU+bV9CLszqJnBRXpwYWQqcemeui7bvintxo05lezSnqKLAqfxe5GmNZsiRQpz
waD3oS3N1OEtAWlirxUZspTriAkeg8PZjFvlfLruzwuKkfNM7fsNckOpeLTtFeKs
osPqoYyr+EKobw4JKJfr4d17+NF66RIDdOQ5Nv8Jb23/NEC53HVUKq94AS2gei/f
Qjxm49iE+Xs8DTEOY5k+AM3CK9Nbplcc+775EB1qChoAuSqmdr7ABPlvno7ac4f8
wvFA3cChmcM3zAfsAhnjwzjWRY1Dt7x9H5/JFqG0hEsv6SZHvobekWAKTa6Mfhwc
ka3AnJ0O5P0l+xQIJF/boDBsKJKDj0KLMQkx33o4TiGFHnsw50cMtkBVnCiB5f7X
kqKwJdSNPL/sx42i0ZbKI+aMFgVFuq3nEbeBcUKVaMNDL+fF9MMHD2F9V18jaNur
CjRb1tqeSpAIOguOvOnx7MlQJlUNg/+WriTTyscUrQSotKFrmTbZFArlj81kdY7L
3Lm5M98QqEqkeKQsZ9Tdw44rotqDtolUDlLLbzbNETErquEmcDYdGLqea5o5ASS2
OFk4R9DcVtLcqeG9jdh9pMqbzfpqJ01g7sN6zeNuHq9CQJM9w3NznokmWe8BVJzO
ZEnuwwwJBwc/gaVCYVIclDqX6/cFRyL9Ll9n2/1Y38PnjVR4zbyK0M627ryLoJYy
R+jn1jZy6nRmL653WLEnq011DjvxdyY6PA8bvy6zgp7RVMBm8yzxYKz81Md6X6sW
v2IsoBtNqM2UOVXScYwgHSzZdNALxD/wIvLwAOupOIiXTTp8aJZgcW2Q05AcGy67
5+moCKMPC4oamGgtvVwe7u+fZUqPcvnWyISo4SFM5jdPAlM++UMbwk+Bwr5qOBxo
9JOVudihUP8JZxLRoAgcA1WjyIuhQp9/AnM4DgjPoVKGquVfqbYZMi4mqRmst0dm
H/2ZQPTAL1TfQlDQ1/v4nZADrP9FHBKhL/b4pqfXqGimIsQDX6fpTfgnq+HaJoXe
/FOnEhl3ffx0ONKM1+HaAXv2u+oYjaNSH1OXXd6zcu5LsYsjE7eTW6bFzHkNgIGh
pw3ukIIUuQJ32SV3kIlEarzSl7Uq1iPQkXcyZxiIuFAjxDMqN0GT96majOCuODjH
BfZzFcXaoT9/6umTp3M7CowjANHU2lMX68cwjJ2zybPksabYbGHKuBaYB0dEbF1c
iXfYjooQFsodABq4EV11/7lAeiA4GeuXyOBQkWDlpuiHMpBrhvWwEUsvy6YO6w8D
wK+o4BGm682YQraH71HASiakwuzLSZwAzunth3EV9tLg7JrjzSiojkvNSXlh31/M
qMhi6M8phZzSeI6EsdYNKTygAU0HnTqZfSa7gLEIU/EwRc/WCv+7UKsvyMxolGAj
eTH8KBC+YE+7OaYdHwR1UQZaM3gTHeZjdnrU8ffQB/ZiDkWV84svz+YVevwBXon+
s8dURAEcja/ECZgWWhHwImP93CHgSw3LGJyWvjnFX/s8ZAL6hqOniYLx0hNprBgG
CMZ6Hfogha9299GNsXgtIu0qljpAObiF6+mI1ncIofHtXtD7N5ftww+hthEaFRpN
m4hYacj0bHsAwr97Lbfv+bNJ9JUZ8aJe+swhZhIA4MNLVk6uzO80Ujn0Gfku2j4M
09wF2ml04qdJDpBym2iJf9Kwxsv1CZUs3ZtLWp2d/VQikqmwzYW1QyoFvFBW1Jt7
b5IRMHjQSZteN4sxY296lORj42PwViPHXjoSnsXYXS22Z+WUCcWZ1INIMiMOkKHj
WQR7vxB38VGzM3YtBENML/Di9vvxkP5BsM1wv5CsyvMwgIgTIIU+fz+BOpfOCJv6
FdgJBDcDNBLmGv+VT98NC/ELQA0kxinYVXA1WFxJMd5UhPeEjzRJ2uTxJhJxnblc
/0ebjKxi/zHM75NBYrm62b/u3xf76RqQ0fLcoEyVizdl8YQ+ZsEGXj3grwwvJNhK
WsH7nw++FaEiiW6u2xz0FiC4vDBADvWo0gAcADzIhWlGr49Wo5aylONZwyRKC0Wd
aHoFMu6KAhPhLddT128Kkre42CQz3dacPNrJtA7yPS12Q2bDITx/z3TG99rqJE1s
em3aGBqWYkaZoa0e5YdWSccsZL4EPXMwCzcSmH3iJ3kL5rY3F0bPbt3RS2PNAGA0
JzLe6hF1ncIGwwBBlhNQcoznDEoNnN+EzbooPODnONh3ssIDC7ddTnq8BaRx6J+c
x4Ysqj+OHHx+kdCJeTSZC5kJDUfPZESYuKp0KzCBrQR+J4kse6i0zTLL4Grb2e2V
Uj6vTUWj8bPTN824lJJRC935Iaq80RbZ4Ivt2GQCJ8ozYz+pfL8E9LfsntoaCa1E
JpxVSqfnYF0AUyIEzpIM6R/8UD2MkvRSyN4et9HU0EzJH2BahprK5PDhVZU1dWPh
C9ZI7FkGdImTMgf/rHa6t2R2Sxm5lP0RM1gOCRP/9t2MAWOyE3x7bZ0O3c/rVAt4
Vpc1cyuxRujWOkTkR/caXMmiFgr2mYH7tB6JkBCHVHAQbw+xNzAVW9ELxPcqGHNE
pi8AneUg125lm7XIJTQFV02gmaa0v9Qm9mTHEcEc5fjfuuw/MKM4wMfd0TMEGm9v
jvWXY63N79ihjhpqydc1NpH2rSR6BwCJ/us13wewFRlir/uXu7vwTqqOlqZYoYTt
En1t2Fac97wOfFmZj6FHi8dT50V8/C1pMxiUuMZN7WITdsCrD1I1jDLC12ViixCh
OzfdDmdhRMFNpbn32k0s2vt8HbKe14b2iaC0cjOzidMN3xbebjjtpN6IsTh0wkVh
oZH3Nga97hmOVAT2xAMdQr+8bGBuqai/CWjMDCYEjL64gS/+f48lh42mqZPbwVzb
rxpMVGlkdVZUwEwndkPjpndWaLkcvzF/f235ndNOpVhp4WbI3ByqbQ4rXsWf5M1M
hPNtz/50n4adhBVd9y3SinBvsG4aX/7gXdXDz8DR9XA+fNo42ydpeppR2o+ClMyI
SP1KYSPw7WMRanjkIyEXybqzXV6bYHt+tmEVr+AGNtxANPlcB3+Nl3IFAWoY4kOh
7AhhpY+ZO4NTR0muclvnY+vvRQjfhKYXaRXHK6mFvZoJplgBqxl7lRgV4q9niBn4
Kw8ZqRAnfaFyBxWgsfB/RcYmYxnj+92GheFEPfybL3JTSjNrVmfq2rxvpdNaQrjq
wVUDPQFIlk/KUh5dbyxZyd9bekXGJEyiFk+1oesx4tv6WTYU8dQT27pKd9oWGE+P
Cu9UdEbVOSFgfC6e+UqcPM05PemjcXojutvp6bNDrdT6OKnCLzpg4CtaMSeJtBTO
lVZkcK/7FM4E9D7Z5yhYADOOku7OaKJR+Oq7sf0oVK46igOGx+3CFAsgb+C2iHPD
3MuxtMarpAHlySIevFT6Jrz3AIBUonbhibI0jmeIFGhhYJMmnX8bjADZVsXSuRka
IHidVciHumH8B/MPXKgLB5O0Df/GXKOhJtQHRwCYsWtfcFKyel39NTOLZA1/52u1
fTn8Xsql37koVEwX7crwVUvXjpXEXBhrF0YV/7kmYZZYy6/Vv1uytRmBD1EE5L8t
cc6Od3a6BgXIzY7xv77RzUnJf9Nbg06mCqkrVGIUjr+x0BGh4/Vx9bFTTGlofgYM
qhFluXeUaKNYLPP5T8EbuawOrhbLDW9vYCEibD4k5NRnz5IldK0WO8+QEHSEAYY0
7QTWAFxz8o8faxWJymVXBXB4tv63zR82cG5dXgovViF62dyeFOyp42ePSOBNqyyc
O4vyVtwMk50gHZUbNrW6c4A1oxEeZppD/G9CIwTSS7supj7ZUwnlDDEBTK32wAz0
odY/GloqWjDbIamyF+BmtNMMoPVGzxHiGe0xkBVlThMHZnQK/DO+ak/9az+2MrZo
4h0+n+LVMnnZa5acZvqy4fjBCVQw+f4/TYj5u3uj+6uVJthehtgJifSxQzDNyYZz
8lo69Uo/dJxnFBWKYf8knRAUVGdaETWhujIVFeaGlXutjgVzUeAEGu8fhl+HleM3
G3cUIT2NORTTEkiDi3aDrLaIhdQbTYwZcVPf/UZMjEt3eVsveCK3A/Ym57xV3oWz
KtbXS2sLh3OGlAFu5z9pGm6UcyyiStwxKyJdTmeN4ZWQw7FIZMEHzNkqBiaYKQBp
iqu6OF4zKYwWd+Ao2Id1N29iYf2b8I5+63n+eN8qxkbR/+tjKWaOuzhYFvbsLMBw
MiWbl10dsWPOuj4lQQGvK+eCNyHvSN9UCPnJYqJAPuBSTeHIlCJidw+UXgEtlLvR
VHSH5AnBUicZK2M+Az53Q2I48cz5+dg2emi8yjEmSydQmW8TjZCcL5pQ8IgJ/zZh
sYEhd1hyJ/fq2jpkWdMCbVyBsEQk1OeFZdPZHiNQHpz8CNE3W69XHiOO9SSotJBA
SK52+VqgSGe4UtBDXdrtRAvAw45q4MchGao3dARGiCQUsZYIkNYnwViQI8bzGhj7
z82B8U3gNo4F/9r0fVhcqGIrZaJVLZzKwtDvo2+JhvlNvRa08NTdJrPYNv8OYw+t
frhQvdXrhBFdshE8mW/IKwPQITGHSxo9CIbkDmeaIhBt21/UAByDmIOJmB/QVa0i
9qb01DxdZkBwUL2/6A5CWgwBOBfYO2IFWlXwtDRb7JKLOamfyNFz6kcmLonATYbs
5KzDOzhCBUyMeFd6vuR/6wc3s/kAzCOinTPqrTOS/T/vBjGTJWKaVQbxhLlTkUUw
Ywt7bj0iSA7fWPw8/71J0ML1ZEXk29tVcPFhqLdC2zCYjnt59RyVIIfSVhI4cyeH
CDvDqnZStDvDzS3X2LxP9gDaWlsmVtis1w9y+4LJkGZXcRRyKaYpSiVi7ceDtK+U
FwEIoym22RGZqqoXdTO+F5fwvEDnhYfHtKA847rZxgSUKmk6eZN+dr8eH/cebIHK
Ke9i9Thrskq+sNpgc5Am2nHt0ZOF2ubc1p++794bjayFB0cXYFnCtpWKcPIX+wB/
xa9DIkLxrZq/FQye1l+B4SXJtiotr3AuuHiXJlz5HeBqc2ne1UDZY25tC9adftax
0+vIyCh1q+mO23FUrEtF476X/+ytcewRhQHyYCX6Tsaeq4cokrgd4aeUekJxSvrA
u9+RJvETJuJt2biOyQn9mRzz++/ve4lhpsH4dilYMMnKeTr1a2yljGHw8jCWzrvU
5bd3FsjsX6s2zRNuucxorx0YT+sxNsyGCJsduLcCdH4J4VdSLpLF2V7V/sbcWCVE
VmN/YGO/wTs7EP8I+EVCP/xnwEdqwOM3Cdz5gfQ81ufPnXLSDdgSgRpFtxYntUG4
MTfdLBrGuefjhu5Bs9vG9rGk72VrV7kZ8HjfW9HBqq1MPj1QGoJ0DKI0RuIp18vI
mhUOXS0oZahANtKDAMO3zA+b1PNAYaHn5E3q87yXtkZbXsejIFqSmUqzkeizYaZ3
8JMvnCtUFnym37khuSb0scy+fZw+rAYVYAom4IGbKtkb8v81dRz6ds4vYHfQK9WE
sQbTtCMBbrgLupmwgXurnKT6QNF9qsRSFP0GVD0eQRIWbhQlKMVsVNJq/HyrD8Lm
X1qw/VHmG2NFxJU+gk8uUc6WRMMcScBbvc0SsW2x41Vm2JIJC438tXBnzOQCtJn4
XFmeHrTvzVD7/ZG8jVicDzUMKggbFfqL9jK3i8uUSfP8nN8r+FaFEQ3nlvWXF4mw
I+y59ZJFVrpyeF7aP6ZabWdlueLHf+175WXdGE6QcxigF7OGDF5tMJdkHzn7hdg4
kqq3gbw02lNvE0HaavqUgkCEf9XsYhmA6SQA2G0lLEBxqibHAxFx+tv/o/F56SGk
Ax+5LDetuYsybEwtKpVrScWZgmYbbk8/R0NEw21VggctFBzcXT1JR2fwX74MHdWi
F1QAAMjMuu3zd8SAdpZZLwDY8GoxjFlbsZH0niamZjrgbMBtMvyUyPVgJRNeDVpb
Pef8QJ77CgcLxmsxx23rPxj+n23a/CqHgWdYeC6FCQVZFVffYzfpxLF5hfLPZZPK
Jc53QmnOhkWo0R+oAO4giSniJ5ouXCUaOHNnUgifD8/2OJMmKcGH7ElI7103H3o8
14ADRbbxq+kY1yWAGj8z1wUNflqFe8AMq13y5moxdw4C0q4mIi0eNHCaDNZ9FLmC
hsWa01SpyKRNQREvdiUri34+SXDjPJy3U8FEzP1woUU/awXcLKePmD3/QO+Lix8x
3vRvp81b55tGK7WS1pfkFrA0F3ynkClsRaS2jXfau58JR7fTUnMmk5rPAQuMEzNQ
l08a5WmHgZoo3tj3vfHFMIraOwXoYB2L5dOZyOI1tgYstZoSVqZcGOc3uICH7xXs
Ss34GimFxF1SQMb0OZLkS3ooMXYaQUFlMVpGhAzrWbZcnzRanC2q0B4i4zWHyCdr
GnT87MheMXm4PitbwU1TLLWKTaAMqG00fv0IdPQAzh2kNmZCmGcpua/c6BbyuZO6
FGs2ILQVuUtUJbGLKzA9GHcw4SNS9HdxeFOaPsMiweDSbIJRU85YwCQ6uEZwIFw2
kHviR4pCyKVqkvXvnhtKz7f1E2BLz5xNuiYqjQ3bezmzOKyMbBGPApQV1ArgrKls
X24nUt8qrA/p4AjUwDTKZhvReMk3G9hjloXomRpes+csS/Oc1eLH34HodOiJYys0
Vo0W9A7Ye3nvbLB+PRMuyw/e3myaoUEQs0/9GDgCYV6m/p9KKhPzksBSyAc5w0/r
6QErLnQthp2dM7Vn9VUzVzHPuGmOWOKiN1gsscAKvsectM5JZyG1+1ZLuhjBar2f
DJjXGN4GpR7mJD6Qixl8oavzvZFV1W43YUbjWAX5G6mhLOPwskl1oz1G9B75XVK6
gsz12b5ldyUDvlzVwwEhK+aiPP0h4FghkuIv6v1N5eldbv9GnetYxt7NgboEsZE6
LclleTWqsRSfCK4/ohlIDeaSqU0rdDpliaNN00gIx1c75o4qMLX+jg95eRYo1FeL
R9mcIa2TymleX3O5LPpEYf6ppF6bRd83OM5KslphvkKGPhn1x02aw4AeIxddhSt0
F2kefZNo0PMJMAoPkdQdeeNSEcUnRPDAiAghHWwA2W+wWGJ1LKTpGe7n9eCGpq9D
lhRLw0HPEGdOMrM1x4Ki3W4gxQNspAAVucJutSB160ynbc4YMyjc3kDLU5QqHRax
oEaxWeEjgUCXWPr8t5d0F31MSlmgNJOEyzzuJnWpjajULtOWWkmNakV4JAyMMMbf
G4BpX5s80BNBQU69lNtNOzozBvpob7lSWvoywrkxFY42aA8H5wsM8TvB2UTCDYKC
b8Bi3E4RuovJE4/DkGg8fZDwM1LuIQmUDEpO4DGJtTkt2mUX39/K0g9Y3V4vtloB
zX8jE5ISI06FOsqi9lZ18rYfqaQwu8ym3LGRQ+ru/Xn1gF3/+/b0e3meT4LnbQR8
uD91s9LuiZohs6YUcUgeWT83V54oBoThXhaQHd8cRshm/ea6qX1wGbOgod+tJAU9
02fW2UPqzUVDCubcBOIBAmNp8R1GapoU8X4hqa/rVAo0pemwkOn7sNhSRHmWKoSH
0TX+lZxBjtgOK+UPh64i0wLOB03nfJyuD+kKGiR4sbFTs9qm4GRYMlTUQ0KOuOFl
NP4Sq3J31mnGCqknikljz+d7L9SsNldhte3TudWiArgrJq0mHxKnXXKcB4Kg2Y0e
MfxyNRH0A/vSxBQO1y47Jcuapn/2rpyfvHBXJR+lZ2KOwH807kb2qOd3w9cxd9+y
onqJg8S3oIMF0mG+xDUbPvNxjypwKOSF2wXV3qnKHppwUwNeyHBE71PPcOooKOdK
nXnOtUHNbort+g7u7v2sIVS6HzKvVgvidQwMCtBgbO/selAW7ni+X+3RMosqu/pN
eMDUZ2vi+cF9u9vOIsk4D+yZkN4NzlEyYWvUhNUJx7Qcd+vJRjZyFnaTfyMoJEDD
jdScnKixsANZi1p29V1m+eqLfKbDpQXifYbipf6QwiuIH6KNFOrvUQUzW8XtN1px
A1/L/zxUn0P9ZV1zwvP+uP04IjyLAVDE+MqQrFELTbEKPctlGJFo24a7BG0pcfnb
28uwaAxIXSjCyuDzFuUO5u+XUXbxxshfHwJM+BlgaG8LOcA0qlHVvP/8GzPs9zXn
ii49/AtMVzUrAqPk9WJgJrlEXriHILZV0Ku0r7Azl4oGNrpeqUv2c1JORBm0sVf+
jmC44bkjGb736XVqFJy/7ZsakYQx92pqYaWdlGnAS7WZ/WNQ52+8J0VN2F++5jGb
Yjz9lsrVuvyJrwQZyw5I4u1xjWJbuvH9sbPBoXKc1y229AM8YVi2xVkTfN+MQvdt
Yz2maMaTYZRdLlrN1JXSU8NdwtDSnBU6b325NeJ7VmfJ9AKWLo7LYsdAW9F3Zhlm
gZJDGxUgNY6VkntmVD5+wHv9sK4vk6beL6uXa8F4xA1vgL26YnUXCppiqWu0CBst
hmfqoC+1Wq+1lXJ9OyQm3BlOvPe1f7M1rNwU34aK/UmZsnqh6Th3NCo3+l5n1DG8
thKpAzNHfFOMlPpvpaT58K9vFqyehxtgio9NztfuDVDtg3/2hUiyx5/nu0agolX/
PTXkpbfTcNOGhLwYmUHJczRt7jiH0ggD1y0/80PdPthRkhIUEFz4trAXGfMb4qjE
UXi76aGqIHvQhJza+p7O+wqyrGk8vlbOuji658XGFAopqia0Lz/AsDYIXqJ2wG0c
JVn+kp1fCkvH10YYwJnzf66VjPn9CCMiC3W01YJXSMCHP37cvW783KJy9DHHvpzH
iHao2WaWDS59sMD/L0uWLeevjiy4CjsmKz9WB2dcJHOfAt9vsgo6gqYDBhRFsNZZ
kOTa0SNibdLY/caBJAyW0HP+LgvIWUfdNzuMIIxJW9eiMmDyAtpYhe3rqPAparWy
bF6nEm9RhEbIIaolefq3RHjGDsaloq4sQyALAclfWXNCB+gj7jVmtKVFMF1lx+8e
hN/qfjZOD7GBR6bYzaa2vuMaEOYUbLfX8HZgH+q+SpSNDodEKrdLs+EGPt0KjBqA
crFI1U0OrI43bMmCEK9SY/PDws4C7Xj6VVqt8B4ZZMnrYYtXL342q8p+i1WoxHFp
Xq0AwzRXnqBxtftjRMww8QvDzy31r5aQ6StiU+7wHztOdkHUA2T7SrPMjChnKU6g
TdOPtV8CQPLh0i7Edyi+iu24UQL/ZP4HXVaEmHAgPsuCNE69+t8792DzpPxweQHy
mYgsaQmWx+DHOqvvjYFNPYa217I5NtXD30OkyKtiVM+u0gK+CbwFCJvVNzNrZ1XH
BNv6O9pzSKwX/u2ZQ2ailBbXOb9TMQjZhl19Yz/mbL5SMVZrlieZpY3AKIT7OoO+
E+KC3Cj7idsIN6mlMG0+kaAo8R97ne4ZkAFxA1OYv2OA7JQOnAaiHUe2/P30l6gk
uzwA5BbNG0t3YNz9kkJghnXgGjPXAMnLTyHeUdBeDXY21La9AAmKCwnZaeDOsvnL
kQ2A4vEgi4cyAu5Vl+ku0q0EaEeweSzCk+KRaIPsQlDSiZhiXSyBdiwxtdtTK0P6
0/z8NaV4VuwEsfLS9vs6vl0YJF7FmtArxlfJH854TbVAJZuf3uN307+LAZNllUJi
e89hXynsKcylZeFj8uCsKQjezSSney7HR+CGLcc+rp/Fbd0+q83LKwg8jApSSrPj
doklqYluEJKioq7AEZJ2btQQlb4BAx5f+Rvhtx0Q2Nh/XXN6kMBnqgWjLsfttM59
4kyjbw1LJWKhI0tv982f/jSbdOA/DOGDTerEpSh4MI5BFaT7rWVvZyL0HJ2ioQn7
H35tl8q9xc123xUWlvBnXIc2NvkBIY1ETYudGUyclq6L6vp5KXb9bJ7XlZUzyMpi
HNtwahcH6uaPKslmWYN8R6wc29pbKsV1YGdGHovO2xQMT7UoiASg1RzzREwKB61H
3YGHWfKhlnmp1BV1lh63wZuM6DrIjU0LIYaRVRHdJ1137aXVjiQtEPt2jUG8eizm
y5j7corpNBFNrln1GXFQbGwhIizjnm00Xq+puibZj+oIjc8CY7ebh0LzB9SRtAAd
N3yWV2B8mi1sKuMlaf/uDlQRDW0Xc6X9T+ifAjd+td//qtZxvxmgnBSOZmfdlslL
N75ddDSdYl3a0vvqSW4e7wivA/jqJqh5EFtpHCq62YS3XjQeZOEncd8yVIEPBWZG
2iJpHZ66bKwPnqhMnN4l5qp6YcXn8HnkcIdF3M9/A4DWidsDbKz5QdftBvaMF+md
4jgfQi1k9hwr4sqnhcIMF2Uek/BQlnh5QWhUz01X4pYuZNMZEchSFfAeAzrsYbPL
+MALdfCinu9+4gKj6zz3Btsnp2kWh+uXYNlkFqpYyGhngYHB2vBo2Voo0mi2E1fD
4fLA8zEW8RxFPlrHlOo5RAVoQgRbgwCdtMd5yTaPsdXVXaM0onSZQEEQ/2P6Cm3U
VHZ9JvTGzd/FXvnDe5lm04Mjk16QPXTDa4KRkPX7m/sTzIIQmNht1Dhymeltj0gX
UPi1I54hTYL01r9pdem2eL5yKACTynhJeUMB9LH3K5N/fbbkhrf/Z4tZ2fLiwvxa
nm6F3bQsPKkxQFsc6AS2lCk0RfhwPXNZX5oLetag9DM+2mRZOyR/17XsaC+VW2uT
ae330oMlKqFf+bnrLLltJbxqA6q/vg1NJEB0IQ9irnhS+XBCAoNfHq7WUDcN2ISM
AQWpHM7cHhenV0zixsOcOXrgDR8O/VnzVrD0y+a2UAwHAHeg4d5PSv6xqN7ELqq0
7Ug4LudO5eDJk0lyNZGtFGOjUPI8SHl5IfawGIRWCbLKFPeB8jfIXZNlD3xNlNZJ
NEr1ErsPvTbBCqtctMeH9RG6ifj6MKXJ58CR6DVsllqbAOecTYhWEdL8DLyLOqCh
+ByGt49+44faVs6tgV4ugq48Gcc+5KuHznVPjqODN5kBqZMTluoIRRcN49HGhK62
LaDCMlaSUXv0cjxrruHhV9ZElU1IoZu77CnkKAZzvpo3RSx/spPFJv1hk3pXY+oT
w4c92P0O/h9xEspq2YkFScD15DjlFG7ADtJy3psGnQeo9Y5LpF7sfSkwKAyGhYev
kb0bdRI9IYhPb8VJC1ctfLVURmYOt51lUpc0B9gAl49X9I1rY0DBnLoBTAxv+Ecq
NGva7Fe+BAt8FLE6xVxHBBAUQSmyInN+Ag92JMafnNJjmNZKwRUK2usBd2ihhYht
h5L9Y/pAXCc65oVNkDHONMksRz1k6V/eogVEQBsap4JOvMl+JH/RNOjrgr/A2S4s
lsvpmnf6epap32QGH+rlWsHaJDY8ziOgLvttojmNPTekZJf5jtFAh4mcHJDGFdMZ
QVP1O0OYChmU9THjCGJKzazuGurqRz4JXo5+l43jrjjh6brtytgAcUUE4gncVu5F
D5VKnsiOmuFlC1skaN6Q5xgOMX3t6ZxM7S+hmpAnjXS0oMoT4kZXDbVSowBBz2FZ
MthyoCzYO6DoEW+o19tUuXzF4glZaA6JSpFcWKc+lvXKcD0BqVUU2te3XaHpOKBa
M3hjZyeaJjrwzDTkNd0kXw/yOpjmaWz7PcQmQW/6Mv4caqqg/dsskEVjUxVEHy1T
AnwuSnbe9V9FJbNMaBtLvrImAr6B70Sidc33zLf9pcailfQBmurh69YMpEoxufOm
IZcN1XeXiJeSV0HVinNaqmbo8wMqCCmRt3jSqTxqpxCLAOgBDCZmWvOHHiySN4jp
U92o5cxydTLhnR53Dxu3WWG5l86Od7pyvftzsrnblgUJ4NxbC/0PUZjo4gKaWnSu
+nHwefyF4EENVYlzqqt5Wxr/30RPQVgGVQYRhfve9RaM3ngbfGEemQ02Tew384pz
xzJQZHQ4giOswjHe3JXYNTnJw0ZBi0e5yIBg7nS4wHfcjkR33EDNthC6i0xVoEGI
K9bCMbN3xIE0ulzD9o9I3/BfSDmpht7jz2mtvlwLA42QvT35YdmwruOddYjSgrhd
xekbPcVfmIhp/4GGAuBBhriQCBjFRG5NCVDT9XtwE4TVAjg2x2yrxCjg6V34FdnI
s/C7kiV/RSoYp4ivk2JnE7kIDIbv+3vLJy2QV2uU/s2Rh/87mQV1bwi3aVO9uXcQ
qJ110urAry8lFAEl39/efGvn9zCXiBQKb89qIQ3jotSwEUOVWTEsqHFkah/p9X2V
oDZQMVm602E2bIcd9tq0k/9ROEncdx8zoI8voyxLkPxE1KG5I/O7hd7Hd6+8ZuLo
fTYpmXuonKzfwHI36CMbV7CgWChod8UzrXkNrl3XwAMF1WCs9s3xR7UEeOfar+0Q
HANIDL++rKAVBkuBmOTfWHnA1wgaek4MeSgSZg9rcvi+weg2jG1nqOUIyMmplRr5
NZKN/x0nYeaMuzkbxC+OBCeRUf3ZyQINSdelfRe/fPBfcq7YaspqIIHy+wFZJXZw
8B02BTMesMO2VwJrr7R7SmEG1QQM/hx/vsKAs6LjKvRO2ivQ4AbUzAH1DuyVzAqq
nSr1uI+5qryyadYWcfL6Ua361urVeFDqto/vXTfRiTHz5F/eSQf8knKSXesIsTLA
MZKpnDdGWGLKMMXox+peOz/c63ZTDadPMUqaFErRziwGZCspXRCpdaVmgrmxPgHF
5ID3UyOTT2bD7EVOpG3xCekS8ZpW9umAHuBIk1YvZ3ggCFcWSECja38nH5pZgynX
TDSOmLpwIy61yYaTPe7Ov2clh9mkav6TYZ+jkERx+QwABmsO1nVnIg0q8p9LRW++
bgn6RLATvQIEnS6TqYXxCuhAh8QGoBs5MTuAsKEUxvoukZpErCbVrSE/OyeE8yqU
Sx+gMJv1TW2GpMZGHla5D0uRXRTG/bjQka8BjNyVriMP3peMW6IA1BwLnwtpYfzh
sWxqkK7nw5rPg3C1sS6fDv1zgg2Za4AmjAYikg5sARI+vaAWfwxlEleKs/a5J0nn
cJf9GX2uj9H5v9t3tEOdBU/vX7IRs7zI3e6tuU7WjhXYyYUn9k2MylcxCmFQA/cP
dsnMFOKSuBDQPTFPTQ79Bb1xHid+Tb5fZ1u3nkzNomnr/gAKFfvTirvJMA6fky86
eg7MIKGLpKL4NqIaWe/l8azM54LW2hZ4ApM7HEQ0H7UYqaDS1eyN9FeHkcPuhRLw
JVOsRUjnOXrYKbBG1zrUL4ZtcgrlpALihCLJDK73XleZa2E9SPel7AEWIQqn0ADp
bhPsYwskU+emUKDrGEtpIOnljAAlbipyTboIxfA/+nyisdD7FeAO33NhEfR4HzjJ
j8G/IMxdEyDtfcx3jzusBqtmSo39/yx81quUltpBAB8RkXaFqliGZrkCgC3Q/ZHR
5NHT8v7RBooIsP5McfMWmV6lKqRY2JlXFEawk368SjFYNRyswxhe2kMUiOwMJ65E
pz2QEDQDZeQcjjgkZcZnZ3UAJPBh2fBvvTq4bdfQFtHEgq4ff3o7/LAnLBcgzJXY
A+H4MnsNQS/2G27Mws9t7Sredwwl3jvQ17qh6/ZPLCoqI/6lRnyWj8sozd+25dkM
dcriyYPN6aCrp5Dge623jJqdfqmPw8s+HXiAkeYVMZwPZ2QqjTDcUulUM4Rxi1P2
uaZ0bOUAEtsv59/epTxIEsFztR6oCHQ1c58dPwZnoDCl+LRLxjWPh9oJvKLAgG9y
YOX7Vhd8O08XqDtbjRGrTbeX/CztVU+qTYD+V/ODdmOXZee3PtuIx6LjK31Mqnus
Jc17+BlDrJ4Z5qgrv+7pUq37ULMikQMs+GL6nrku3DIt3yXq4NYgwYxJUlhx9QRz
QBxcAR63m737e1bszB+3SOl4VAwAiV9nbOLwzuAGGOneEqtnfCeO/GdXR8dWzJ/p
gVKlvyGQ3k2xDMjrnDWsfsrnTmAvuqj+kKwnCgLbxKRXOOpV2qA5mmY5PUlY0utg
YuWwtmBbbQSeaU9wRzrHriVNpyKJvzZoRrNU0ZLx85a6nyIISb04i7dIr8pntbYf
COYgSN6KEvIZihYMb0dgUWamfTjTJXUilxg1+1egV4xwqoCb45J5Cr0o6DWoL74q
UlE7T3+uOXBNXdxZfhKpfH4CRLhOftkN9+gDQi2NCBGPiMC/Z8+tCCE+V2ZiS/HD
hCAhwHiLwtBPFMUwHWVsfYozcB5ucQJgdQ6KOQbM0wdit/4uY7j4tymX76o9+Eo5
LYjV/sOOv0T8Mw0pjytPgZN8FpQB0u/69CoeYAWHtbz+NxPsGaEiYr0B7IAKRReY
xltPE8YjcfZ0LmvI0umPC7oQTsgogVd2UzAuRc9dA4xV/mzk9hlmsgzMqs8ct2fd
xO092PORS3eJiYLfvIDjf9W36aYplpVG0rFeFlELZzxqGmz/j84sdhQ7U2kA3gyD
hfQ1xNqtDKrY2cTXCJSHQXociHtH5EMot7RhaMLl3d7h/Z7Hz/4s6oSgpYimsIhu
9Qdeoe03BOyfqTydmISsTLL29hoCx1OFhg3s249uPukiy6jm5DqG6QCpNT5PU4C0
6fn33TdVeG9/ZfaV01v8m+kwCns0YufvVWacYlj6wqfJOFy6gJdCSj1USPqfaWHT
47NxwrYcDzRcmN1wW9D7ggLeoka8tPF4ZvWjIIIr06biQPfHOWab8ZJ1g2hA6Tey
YghxLSdcU5Tv0ZZ+06ozEx8gkIiPcj9WhQ6LSK7YdWwSW6woxI/3a5w03AYPeVU8
kWlf/VqzIEYIR2VzhPSoyAVMIl1VF9jncs4nCnfZuYqr1kLOVaxYS8sMwibPDqMI
p9GMoFqdhpmoOW48Y4yFx5jwz3ujybQdneJn/QAiY14GCHN/PfnWiJ138Hk51Kw+
Fn7CAA1EaH6zAU25z+d990Q/7xiG8oNMEINO4spx95lM3jXFWwtgHNLfK9x/WdgB
bR3+IQSAUaO1REDlLxk2gH+eZ0H+6I+oDMEKYTVMxRDUV4vw/hx5Sv3+QomWtdCi
xcR3iXvlhtEP4CA5vtnt2dcPDICIa54vDJXwqkJkrVvzEDvDfm0prsR3he04i5M6
0a2D4kn1vK5Oo3Eokzw36Cb3TpiUEY9Ifl4AxvVjBwst3gs+42SnztCZ6ofpvv+h
rndX+uSbFS8peMfEG67ye8Izu/YYzPcjtTM+OPc4DIVl5x/vZZe0LKhmcTvDNskw
GWqRFAnZF5EkBvRmj8xAY/tzCauD4297BOWhveDXNIMP+3YDsxjK1ZQZh60I1JQn
Xi/RIWWditrcIDjYz1t/GUnBBdTA3D9SgjEhBtaWUbVzSqoenbufYKYUUM4aOKz/
uEqTClxC+wl0VD/eyfa9S7mJd15OAR1RDh1I/fvBKB8s34tpOhDWtLvBp+5/zGbA
r8fY18GTesbMeLFsEnSKco9kIv697sfsTzkn3vKnlkNgn2jSyeuT/HMd8CZAuymo
KBPjfubS3BNqxqI+W8BDGyGVI/J++w7WSDMBXX126K8zLV2TeJqf3hPrOBBXDVna
xvaYbBs/D1Sh6I8mkqcrDYDWO/pqqTPldr96GlkCol9dJjdiPXYcidsmG6PRdgqz
GjnRwOdpyK/0RA1Zm0wztCN1OrJGXBQk5Cx2J0vlEOMxj1aD5Vr8ZW2eGoEgnnBf
xWmTH/bNtLhY9E8peQm7sOmyoSkeDF9ZbNex1edabgTvZc2p2EAl1PCmc0Rqc/Y4
uHYNIZ9R1c1LpFitDNA2njV+TZ45kW5Ec+4p24eOGGo0FQdn9NgE6RB9RhBcBg5i
FuVNxVbawo4VDBL27s9q1CrGSCI9FOYOZ3DiGl9H4+003i9IYoOXWi4qSndg1tvw
3Vbv98vmlmeWUPrw+U+8b95AuGP5KpisXAf6oqEbHkDnwvsRZ8AJHNb8D4vLSTH4
vSHgB6e6xYPJXrcD6HzvsFTTn1uGttbkLeCAD1NkB+99/ZqKWS6be8KqT4/nRXfe
JgtGpoajDrfoeymaQg0RTS5QBjNGssgJ0zv0p6qPdJsyluZe6fiQX/RMclXIUj1x
2uNfnyXlzoCFkl0mSipFSx7UZy5lbXpG5p34IQj2m1UvBtYvieVnoozayMo9Qw0E
KcJuT9reownzjMoZa0FjqQpYXxhqZ+2mh+z5CP0mdfLtJDHUbZOKki1GGDMCSdUW
2wED9RwFinbWUDnIm676Sqs5Tpuwrn2OA3IpKbk0Q5yhQojZB9Aum6kf5MBRFiIE
erNGvYtH2NI1Sh6ycdtDwX1xDfeVe0OMJlw23dKxSr1seZX4vVn/S5kP3mRwKRbp
LiqHECwfRVzNjBZprfjzh7qcmp5E9aSgEjJX6wX6oE67hQ0QFySgxjK41ZbGpYrW
7Ml/RRTj9hbPBh7Svmh9+myc3A2IliyAM6biFCfBHpd+wla3dx6fMGMXCBNzkxYt
Rn4zcyCk7ttVsKbm7tQplWJYfqZH/lwWvkTvZq+Mmkc8g+SuOW2EX+a/OzG2v2lb
LU3opmLBv5tPutMXgHz5d/Mzd7SJdwXiiqshjKk5faAYzwcMfk1XqlOaZoK4Ui5f
nAkpmeZGt5jk0HqcnckCiwSypYo8ELfuyqM7PVq89wesWl/frl4l0qu1IIS1qSs9
QBo0GiT1p7KKp4dfOi3+VfK2cm3GdCh3qxIX0E/Nt05sp8EmMzVyzGTo8keIm1xw
AheR0pD3kfvl2mgQ3jmOSoESf323FBZJXWJyJ8rujck8nS8EVqETlP52mXtHinE7
aNlxdG4iC0+K+ecoWzckcluPJnbwuR35hEq0IQ59TMBsBkMvc0FNaTh0gnnrn5Gq
RkgbaCyJUGfHDl5FPqOIivNjXd+deFR29Wrx1PCaaVR8+LPPE7XX4lrW7H/m7Z1W
Y2BcMZy9qGMfnzwsKzLAVZecHFc2wLXUuu1FXrq7mYhXtKYDSckqe9zHMwQO4hU5
oenVeROBeJLOza0GHhG7KA/kxkXBMHh0qbQBrwJ0e/59tRD0+qXKA54hv1imvK5k
tt3FyaiNEmdSCl55IT/NhmsQj2QUXZ3GXU9GAo6rsnebOp2yy7sVeS7chnJ2j8mN
U6ZBqKzYyZV4tvhdvDMN0397pJ0DrzJPIBxXqloUfrz969ACQ7Cy/KmznwRv6GST
3veazysuMeNkb8tGlLFpU1ntU16fkn+shnv4SL0qDf/ofcV/NQISFOGa5cQzvwYx
9PVACMcDU16JXiwXp1gIbBA7ArI/UK51fzZznFBHzcyLwLpDKiCDfO2WJ6p1IOZw
oY3MWiB27TfvDtG672EPwl7Q4Lad90/xbXgrT3VEGETbtgPKxUE9luwQ4kzcDrnY
s+lQBEFb9XBVF1rmto7mQ9P50uagJaJBCDoqbcVpEKueVHx0QweBga/vyCvp13jD
hoOoqSYu3kt+33pV5dNsab51bVDlE40PYXqQCQlhlHZIbvTpccPrNZ3qfCHQz3SS
21ffTbXLnSlwCHLp6Bq7uK6gEBJWn8f/D/dZlAHwgM9BQe7GeIMILCClXNHxkm6F
dHQ05/e5ySG+q8lzF2Lu4RKUizUVLFL2vFEH/y6sCtsNmPdTtubJFiK9iE9baXQ6
1Li3C769wQ/xPa913TH/IyEMf3/kf4/p/Yxeda13UYVpQsYMc+7SGVy3Ecnqfe5m
7xD1Ft71+m97R9pS2J+sXEIilbB0hvddp+JqgPmP+Mj822059wuA6JJD1mv1ZOrZ
UVJmv6yJLhkMiu8855ZGbPeewl4SCLChpaO/tlNONYbOluSVV02Z7kcjlcohImja
IbrNNzy2SFAJ6dynZOW/RbCA2KcL1L2IkwS3YEcPxnvkPR/vwG1T3mwzrUyBT8Li
Ei0qq4p65SN3k25xI65WZFe1DV3F3vyggbrTH3X+EpUUPn82+tBz4Emf9DBMRN6y
GsR0IW0Aru2VnUs8tIJgKvekMsgYZQvb+mpmCpoSgjRv3YhehXO/LPvF83Ety0sJ
NaFiPi8MPzXmcCJPTd/0P7j/+ToHkCi7xU8ZxjZEnXBNMACrCnyZBQuzUUEO/9hs
qzi84dnzU2FxiZ6WmgVtm3B/NWtHMs4G5eb2bh0w8rse0FQVXM4HoGhnz8Y+kZ9A
LBACe9W8mQpLoP1lURGk5ohGWIHfac1EgP936quah9whCSK2IAzqlXRqqhvImbfS
Sv71afbbitkuUBHuyyS4pHfzaUOakMImfwA52FXO5CXbuuEDSXXMDUwQyWcCN0at
0m+z+hLuhM6hIQEwysjzDmmna//WwBMXg6gL8ZgQAZfk7Oy9Ey2L/WgoOTr2KpsI
hKm36910eNj3E3xVZaou48ywAoHCa+nnQyu5Z5eq32WDScm9Gc3B37XehbP7BZIs
WWIug29jXk3abW90U1F9gLV7OtOj+lSmKYbRFAN7WKJ+1sg2Ems++BJnoOnfR9c4
W2SG0O3hw3sGn2NpZxhOUcSj9b/qftyhGQxJQUpFbpWiBODQN6yrwkCaiQDjMlk5
2r7SUjD/oyGpMw0g2M9U47k8m0teCq4qy8UaYuANaJ8oIdjyTYDXmLsz4YqB5IOD
+PkdnvXAhevhvYznckyLAXzsDV5wPN6QBFD2nZZZpvSHeNxdk47pAjMzyhch7fL0
MCPqqy1FB2RBdKjQ40h6vF1KyGw7W7goA/H7aHHKnhfiNjQyTjoVoLUGKBwG0HGB
sVuneA3/hJFxwKJF1WyETcErN1Xg1a8WdWq0YjqCa2HRiDKcYm45Gb8el43pz2Pf
j/dBUZB9PVoMi1vcR78EysguHu0Z8QT14E57WX288HJNuRfsgttT6KFkutHGtXXm
Hg2QM7iYFar+EVzgBWU2FPFJGzTL7T1EtZWWy63QZyv9I3tDKiz3MjEYvBBEDBfA
DePMyhZm7ukBJTZAszGOCSXSr3cX6NkfIyqWsqpg00/8i5znk9Hp8LudX9eu3cnI
W+493YhlyEegC3ViMdfIKEc1wBPq0MmseX8Mq8R5y2Bg/jK5ptCNYv+57XVwjeu8
l3Ik2SLSeNqAuaXoaQRl9ExbCqzQat1dW4wZHMI8RjAdW61xyZB6zyY2ogWD3zC7
lTcftOeD0v3a34d2liLLZCNVaDpJIdjWFcl//swQTpnUtBmQYxFtc45XpGaytguP
wr0JbS+Ytt9Nx6m3DmVTGUmoVrUqjcc5cCXb78rtnupgjyxvbmeHdiqZYTbAj/S4
0uA/sgPv4Y6PitJ1Yfv0KdybsTLpDN/H5mscj+meLhuHnAKSOg8mZ7zLiBeeqRpk
MTxsmYx65faZPhcfjPPty24zxsaiQt1TpiC6F72dGkUeMJ67I4AdJJorkN5V9DS2
P62bvF6CuCRRvWXDYPBXiOGXsgtOskxHsRGlcURSk8rnaPOlzI/GqEzPqbiQiXle
LRYr+EHwhhyE4Gw7HHB0BEB1sK80zvFK2xIvbXUkUwSWWeBGqQoPv4EpFxWyNVYM
qWI0armhwotHV6XRVub5E2mTzFkaCqKAKl7Q3XB5rAqiYAQ1i9XOEqVzJBNYl14e
ioSPgB9AfnnNz4AywnuChA/skMFkdOXkifYfENml2c1xF4n9fyqHYMyxd+Mbriph
dk78ITvM6cqjFrOgI+o4XHwcnVHKpBpH9GLf5I9OaPG5IJmBpAE8D+6N/wHENyiS
xt2Hj+MZCLQadN0dWxIL3/9eXJEzBSSzRsCTJTHCCXv3VlGtn6L/bBaczua/8KzX
CeeY8+bLHyhXzktvwonTGHbEmdsmTDO5rleYnLuq0hx5qAfTnggQbk/JNa8VMVdb
z9TfHCxApOupmaux4IlqZdMaIs4cYJ+HuKocwn2ZlLeKAaUu7sDe3K/vl0QMeGI5
ktuHf/yH7DDDd2nuGl4vTaQEUFqmA87mlWRM5YaNAYQI3wtiSX7GK+V/KwCnt0xr
U6PX8r9Q419qA/a6+UCanO9z16NX866E38RMHQZq35gXNx3/xn9La/OuzhEYfjp4
P0i8Kn05Z7Ad6XIUkpgZFN6xL8738E/6zihf61GO3zgOYcR93xAF5oCKYndIBinW
zemlOTqLmQSkZC1FIhFX19ZYyPfJmtMMYmaS64UZ+XoGHdEpKH4sL/by84LM/FC/
V9+vnCsyIOXGviuayKbXmhJnZIUCSjmDb5/Tj7yO59YoE8CHa+u1fQQONKZsCYJt
zBvDFcFcZvsQGCN7afQoK1twAuzNnejMTweI95c47RstD/zQ90PDt1UHiCBu9uJ7
epfto9AED7AVjMfzmYxmqRcYec8c7rukMBsWI636mUg07nL/pKJNVOrc5pKs/RUi
0zH2i+5LykxXqIsDoYwwi3Nx3AKiV4W1XAyLLKI5CsN4tIXQYjpVV4NcKUeR5+lm
j9KlZjF0rteF36eNWdVFS1McAXQuXlYAyByQNoLAqld9nCXsAOGOGAGiMAEo7+1X
VwVHj2vEQ/xUHobrN2MkjcOhBbytxKttXSlYbLK9/bt1LsU0iEI/sT+018vRFdHX
sgoeiD5h+Y1GpY0zuzF0YPCGM9EKZEnQ9EDc3quuKRfkVA6PE1G9WHdfZzO+HS12
x2km7uTEBZw+rP8y5mdnn02AZ5mdvCYhOdemTvB0EGtKoxMHUVX2efd44v2YUeKb
kBaxkEVXUJzWBvaEU7zf0YfdwzAySs0Wx5NUeBi++i1aPJ1szflEYK9bksgwmFKE
U8Z3/IgxsTjxuZaj+3OpcBShGiQBHtioPxllXnjNdVRVMIfmUgCZRpl+KRlUp+tH
cl7X4jeK4eGjwwfgeB5NtaAG/HD3f3OacJQWZhld7KJ/y5FfNx/U26FIgrlQd4y3
h8LjYmA6GpTtBM8v22nHiJoDm001C3s95OPuF1W+FWmqyHtO6wSSJPDQz0t5tFBg
NJEU1BYa5z8IWNwMPob+Gf2qOec6hPO1KygTMrwmjVo8BhKgX3NZhoY+Xu9nc0kn
Uq5XqiYu1fcdGHo2ZsBNwwKomZoDpuxnv/1yTg6ByzvDdFzNk+WS4DHy+IbhDdiT
TK3wBYvadE5wZhfGIF5r8X3Xe6G24C4OWolFYeOSLqGB2HOwgELlgUoRStx1oJ60
rd1lsiCzSwAiztOm5xAJt5gZCDovhjuwWbb6cVOhUPKdyPq4Sz9OFjbT75qNR+cU
8zACmmNnne5kniII5PHgQ5IvpVIOL1Azj3Th3UFT14aAy1A/Q3wpXi3FrQOvCK8V
l17cXGdz0QNAbnEJd5WJ+b3FY5/5q41SiZ2vK07eDVSmnsLTR4cOQ/T3Ih/uyoLr
QnJBgGmcNzezAdiv1H1LkWMoccWHS3uSS3nbiPpaJzKVqBD52v4QLu6dEg+F23Kz
uBQvtKyjDMAiT+j/B0a55Q05xnUR4oCbcTJmFRXgXpgtnGOXKWlNe+LdfPKdJciY
1qjadIVRg0mxgSzAc/6oHspb1ywLex8VamQqQG+x4vwR35lBlnWX1/j9YR8Hd3KL
btNDVdaMqWtPqEJcOEmlyGTcUPxZFtCz6fl0mDK0uIYgz9EDUqNg9e23nrGLOFG0
8SpNCVPC8ZxGLmZfkTuLulZy2J03d/3JakBDHkzkxcIat0X/PQR/UdiWHFFYqsi0
vFLsZ5mZOzECKN9kc6F58qMU5gvKyJ3FwNg8n7iRrcstNio34o99q3m7qE4yEYe3
3rAYvX2hvSTH7RvT5Zq1dsgGJaptXYmqrBuWW+KuYcCX2ps9ZiDb9G6C3u4jaCCV
fj1nQrTC2ubLRBrX+qOvN5LWKKWmmo+OhrVsBqhV0JCX5ft9mzPkll75XpO2mt/4
5p/KTTJps/oYuTHIerj6enNHJoh4uBWTOPHngwqIcjt5e3fgW7ivnrhI4YhvwEc8
lI6WtrSBeEJkVi19B+RTEfqi1TGUqFPQElhxMvnyRYvo9/uvVRpNQLrCYhg3uutn
S9pZ4I9oAvbii+1TRcdFZ6GiZopNXB4+tJby2w6D5cpYjuIgnkOzNaLlTh0HeIia
sXxATe/Peo+K73jr2nfvH4wDj2jtyZM5NfZhkMvgzDHeBomW+jUmn4m+ouwsjP3B
U2uRctdoSb30lt8O+Ou7PHtY+VEKNeWgdixhbdLBCwLZ5Y03WJwvg6Z4NbxWd2I8
BhKUkvkmCp1hc0RRbgeaMQmPSwY6RiKCNCcxnhVaBqTv+10jRwsSwRRb0vcZw801
8Fj2tJffODjJ0zDi5FKMxtNGZH3HtTWT5c4M/AgK6+RWGH0aQTYG/i1U0bobfoHz
+btklUkkuxBPosyuqFcW2xQ3tV2QuprY63rOGJrQ+v3dlNZoct5qOI7ZqEW3Lgkk
1OnMKApRzwNdJ6qbAQt1BpNbv4ggWiRVkxMZ27VHutNYXFUFtf7NBlvQA7YdV8Hr
YbDZtG+lGXlYe+bufUJqdAMKZooJylNggG4pJGFbyBKdgpbHvBbWVsEKSN17A9mz
dMD1S600o6hgZeO72M/xl7625jB519fdxoFqsiX/I4E3syoN0Dy+VwLvorvNW5xq
mbq9WLjqcG08GyzMA7Fi9FWLXtPaQqI6pbaIDqB4yB+LCqu+JEMOGaz8G7dBwjxE
2q/XN9C5TxDj2wtRlalrio9IzvsQ2BAYNW1IUt5DQzR6V5L0y1I/1UUfV9G6vO55
744D5/0y6u7/L9VGjY6fxMqwYyWveqbgHF55kTWtz/jWqNuL2rvMF36NdcGc8AIM
xvj0vdkv2HVL5SCc28DNUkV5JRjbK465o8fX/vwcxHKY/5hg6Mp1FsDxFWHCEcvz
UluTDBMS/vAbwhZUyWuxyKADgQ14coyCBNqFBR+phUsQANr8DmCGX2Lfffiocgyw
GhpNnS48mDFeuc271weQVW7Qf5XLnXcCSSU+ZZl5l7JVSHGPvGy7S4AXiv/8MJgI
Xn9aQgDTXnRcAau2BN6IcaqUGsHRpPY8l4Ik6Gh5W57sELDTYU2saGw1dj47/iqy
UXDf2ytPLt548kO0s2ltzVEEWpCWGeYkhfaC9k9pf8ypS1QzIXUPvb6vYcNm+41l
iOMEYD/fV0JznC+KI4PPgEYLlYN1lLOxoZlVWddz5I8D02m1ceR4qMYPp+dKVlmZ
pRzOz8evXe81wpG9alaFlvJo0i1NvSfn2aRWtCDbNiPc7SmbZQ2ZHfnpYlmo0Jxa
2g6dKcD1b2uD3ofCHcEZAwR011e1JheDwfTgnDATz+9FOT0EENi1EuGajSxkGwWE
bu+h9P11wij4+j+OAoH7TMVKM37H1+NFA+R8FwzrPVCzCoCP+YVXEqKN5ZEuWjUW
oxiNxpblrurlQj7x20m3J+G/Ty/K5wGNmBipzuZH+SNMTJ6uRtTIXMb4mgO65gbe
1N+IUmtNYZoTTKsOI2+o5btqY63qfkkLX6Ct2ICSnLvSYdMLv6IhlysOKQ/yd4wf
hQbWos1idWYrRmuDuJ6j3b7/1Zvk4/ikMYxKRMHnVsGeajWCq3XKmBgWZ+AotjQK
l+D04Cj1cAoPCaep/Mwo0LXyP75VFwmhh8uQVcYtzWi0CF+hnpb0MZ360w6strP2
GVAabccOsjCJKeo5yNkdW8kP63mUb1QVGYO80nlUQBQ5q2zBgWBOuCGT2ko9AzZC
S5YsCqMAYJh/dZdKG+JtDniIbRqmIteruNaTeHoqBqTqANzrjN1LcwDKv8uSxOvK
op+pne7zS5KDPopgfclYEqg16ISOTdE2LUwOlx+aLkVJQNR1B1iNaL2tfkrG4OPz
9whpFYloL1aGF7UvwF3bmC0rOYhcDdlwVF8shRg+E3bj7F/t/CELS6FAIs4CfMkR
ZTgYm3uAl3ywyZ+BSVS8OeDwD/kIyZG7KupW5aEF0UL1Od3DlwmEduFy5nYie4dt
WEk5rZK4G4qig7RbCpxogfDGlHYFgX1jnNddtj1ACHvieAwShhDW3j5a9xZrzX4L
1AlP2vGZyzXexvCbpOYKMjANHPAlBsqYc0Wcb5s5ICXuHktCESTatSU4GiMJB4l4
760p9iXDiT32+GE3tynwJkW6uFod8h5cwKlFWpNAVuAmUZiH8LIY9fK26wRH2rnq
IxtF/6BsVsi2QVXc8mB1NFsD+mhHRNzfQr0Llc0r5wI8vqZ3iULclgG2LgZXyMiG
dwNVIdF8KSJBYJmLuDrjbXa+ITjCD8F2dTH0LY0lTRpGBue/c2JHKEauZbmUA8IR
9xjcZG2lSE/R9WKpzri1cZHIpx9q5sAy/9iWhc25qc1Vba7ApkBcUqrnlfshHYuH
jqyx4tamoi+tkx15wagTNH8NVripz2EDDEDwegW30xd2k+evHN/sPUnD4y3qLxzG
nIx2ekU0PX6RCdBb5nEovrKTphbuW+verv32yX/UmeJdNWXz0lgU9YJLP/zhJY7P
y6+vRWO8r4yeO7Za0m/unsp7JfKouBP7J3DsYDflECg0ai3UjKSQeQk3R3NdZGkK
Lpc+zJg8o+0n//raj2Ux7SlRzqgPtP4TXDjFQ0AQnAawca1nOT6j4gktbxg+QxZH
bx2lYklDrSKyE+N21urYnW2fMD9vNQ0bArt2e7d6GvzD/69XGX08QEnZrTIAYrcw
lCbhRnpqZadzvk7JQ4hjUjoMB9ws3bbtPBbxq+NYksaJnZ8BqBbjQ62gAafaJ6QK
iPWN4g+4C5I8H27LDc4E4c/1NQLL0A8aw2IdvyA+63vS1MzhRfMOUCAytbwW3ZsT
D0pdcrlta0t2VTS9/urNgHocC2hG3kcsbNoTuE+ZtZxNpgxdi38wiFc96aHJEV2e
RF8r+PliIhn/smgcmErHsFryEqPqQGdYE492O2rhPG597K6+sovYXu1fx7fxrFIy
0+5Q6H5gG58h1nOzp/co/oM0Uwi2wPs3pXWlCTx4ABAIf9z9swzDQ8fAQQTr0AVP
XcfHQzgmqKguK1LBKshAGSxytfXIrdz9qlV8QF9wg/GsYNEU9HRByH96bZMbOupi
+S6/BCKA9aXiqYU/rWTK7YTTdsdxh3tVETkZJuSHPldgP45fDaPA9a8YdAGt5qQo
LeWLOxvqP4l22c95A0/Lb9foMxjXaHezA7zX+VjOirwZwCIIDuBhSsKMxV18zZuf
f7gXoOFFJDiU7bKLsLAva1aAqPlegn5IQPRpmpZKj7TwCxTXCweVO+bmAxCbDuOu
+m1mWCiIb/mGAYXtkLXTmuOFrQ6F4v2Kn91ek4vKyBTAEdNvY+WK/p2pXGC4DkKB
YNron/FaAWn1EbEKwU++joqRSyCS1FBrbIGpNJzd/RiKwNJ03abE+kEE5yDHp8v0
7jsVBS/7loXOIvYNSIrLfT5/lfzBY+bp3JoXNMD+6j30IYox953S5vuQ22vqhc7E
ozRXpeEgXYpWzCDoULgkPoKHuEKq52JXuEmD939LbJxvOyDSCFLX5RtjTCAkZg7b
iLJi5r1oSnFVV61XHuUXtJTyMBqn6mipyt9MhVImrx3pW3OCXxi/r/zzhHq2QY6i
9FXuQ1KOelxQb1U1/odAO7p9HIEROGHDx9miJ62hb5UqRPwWSDzOc8dhY5ZRtKrN
JwgiC9Z6HUFM5RYhOUzADJ1H44s2EQRFEn0+LTT+5Y7DL6vMDLAtKqDyugRFZG2l
AcuapO0UBERkVgb4WB7I2CrYXMuFcmpQze7O84hx5hLvvGVSYeeuanaS3FMkEi+3
IX+zFID2YP1jtv2voP1NPfvHerqogxcOir8cG9f8XgOCahYXI4wdRP/IQ8fQhtPO
5MEJCIcQ85z99naOYdrhmljWdC9URPGs9uLSmcUTWzA3JqsJXRxMlej+jpa09ZZc
nz/eHad6oCfYqRJ+fOV9KFPUPAfMuio3e0ifCX4PAiH3k5graKS0387m0gJOO0i8
qRtFHB7i+0lrQDTmrtT509fSnDqO8GUqys7N5vQ6aBDOqtlGgtcKfYp4WPz+4k5M
8s6cLpK7uPUQ7jebxa5giYVt/MXUMNfMcohUCG+YFCHyF89EUnnGGL9BjlgbBzMS
YaLM/jxqo1uLM1tIxX3JDdcX6m0fcn64C1PywOjKxH/+Az1VBm1clRmEaDCaU79o
O2FbG4Fb0C4reFK5UM5S8ghG6GllYHRYbnDO6VSiCo7hritK+8NqntQy8t9NjC4q
qBAkl8Cs2QorBIaKFLz73AZnTuDLH63dYRQeC6VoNNqlod50ImuGz68OXtzTMcFt
Jmp+70pxkQ284ZW/ancH3x8OHCdnT6oPbtnjvbbeM46k+1zMPJclqYd+CFr3d8dT
EdF24y8JUMJyBwzvqPHzPrtZWbCPQQii6izbaBbN4w0xaeOrEgQI2hI0i0VnykML
KARhtyFLTDgMUGSS4YhiyKpPjgRBoBTQJk8KD9i6B+1MbGg59jbsVZ6Bjq+Ynuj4
9ZAJJnX/c74vmSiwLaXLj8bVtyY0fIGkw94h4J8NOJjdE3f1qtA5aSeahVV7woay
79C1z1rkYfOT1xFch5cH5quOkAbO8LoEzGcpwYvw4JznEdBEo1wMSuWtfquH8MtX
6vHP3v49is4Xebr12aWMvATWjPu9LEFpbervdS2LBJDnx9ubpaULEg30rerUEIwm
HnYG6MBRoYoEgFxdngslOwvprZL2G7Z8w9ZjbI1gBkOvl8ThnGpYc/vpMWrWVQvk
Pi4pFdmigVhjd4IR2Fq6GvBXrbDMc2VtJVY05RT5ZVke6emN5HKhG6cSQ8VbAr/C
KB5acXGkVW8qJX4S/AN4KU9JmU+6lk7PI84yYhpcZ7hJyMtGacQxzEK3JFNKMQh2
QcZS8dKZN201zSE/T5q8XD47N2bJqFn/QgdTE9IMDolvXLGJOxHUrkXLg0vyJNjf
VKSVMVFkR5ui8xgCaXBmtVr8pyXGIDJWGVhvTBlp1rNKbh4MAf8kBC0zX+skqHYh
tMZQbOMMy5z+AZJJS4+aoZimyuUMmknRXL2gkgDJ1/TwZq3GEablZ3WsSPBseFTv
K+7tNJK93hvOQEQIqCbaaWX2GkNergVOZsO6Y8JwF1Zv0rcRNsn4Tsd3Gd5IoI61
kWUeewoemA5v2ZRAVcaXGKLAs/jQGKESGvltpVHJcxbdon8tT547iFhvuMIeZST+
vdVN99xnmf+UBA66rOzONT7f0De0YP7P4KXuyj7T9HyHQKJagrPNS88SYoIkxsTV
65D8bZH4zbN8FpP2DyzqOeo5I/NKg4NgI501mm6a2Jvq44q5yypPmDfY8DlEmLix
Xr96501K/ZWcRuZJCF+jb9SGu+ICy8CysNAC/ZJF6DIHWb3jpkEe5tNgk73lyNqh
sZ78E+s3afbXaBs5nW00B68vPiBBagkxcUgB/+zYBige7B6BiaLHkkojdV0muaMv
9GqHnRW727cs5vUpYzagMBDjTq8/PCfq+nIgi8slY0wJaYgJY9WpFS7grNJEvlA0
lZgvADTpDpv5NIuZ9evOS27FodYkZ/MbTNNd0n2MRpXfo9A8W9TZ76q2wsd2bsqT
PDZpWD8ZxPcXVd+MjugM1GmXyE/H3KXEPW4WUywf2Sd98NEs5ctm4DxuHfJKGaMQ
KWXUJFQhzVyi5C94qZD59cyhYbHWIzVRPxawQkgXEj/Na5AtaKRmhWQaR4hanT0D
mh9FI858IGwGXeNzbSS0zTzHI1UKs2g1DJhONOPUUEeOA6fnKxHxGKvaslqdsOTO
xDTvnvEBT15/vBpPnD3rl+67ehBTKIFNqh3/fAzCgnOFF21bYHohblH2R0ndn6py
CyTCT+yPB2tlJTG4PfqjtqGOFtdAiL1W4HFnNl8XB2LlqPUYNIJGWVD7q80hjncs
cUrXwb3zd+LDcuSn9gT4IqteBXlN9n8YD6JC5rlaWDB9ziqHe/EVGs77t4a6anUb
llP4HF7ICpUoPvaTPQQBarJRzhSKQr/+rTJRWM6sDX5lUs98jhZhcKB5LHQmNgpi
k+aOcnZJHNTU5KLcZobpKBBK20rzgsXott3fr0BFYWX7FcX69YhWZSzgemQglhI0
xnQ0cRLGZPLcdhJyHbPzXRYZbVfCnYtFdeyf/rhbLLmSi2OQtn9M3vT0Xdpo3MaR
4zg/Nchy2gOvtbmKmc9UtvrxT3BmhExz7U4SJ1KPuak7+1lBxafuWZa5L4QFtuxu
g3i5jZLVXaaN6/oyMUHb2Wry/+jykfDo27FZ4YpPDS9dcn/2CuXwEKGiS1FeepeX
Cf0M3YrH2FdDJFJrwuzaKVEMo54EL1H/0rUEWtP2QXfxdPMvhJBRMxRQ3fNLg9hq
hAa5VIJDuD3HSjeY+Xzlg94ib/59do1FEbHF5++/bYqKb4iGpnuMZwYw0PlMvZAx
Jw2rYqoJZUsrtdRZ1k0+VrQ0yyRdD6QGCuTpPlU9WbkxTqfqmmAdFs/ccjuYW0Xs
sMR72Di2Or1AsANgKReSUtwsAVQSZbJouQG7ZGgJ08x5Xydnypmus6tIyhr6XIL5
l06+QC1L0/M8Nh0lRYDwoV0pKyylT0zxwEtmhkUn4HdnOHJhCkkUBBQEtEmd0kg9
90uj/s0m67L4Sw5a4O5X84ln0d1P7Wx8kTnOzmrvXznX+4ghsg2xnQUlmws7XfLa
8wQg1TX9Xql6rt+kUUmO2kUs2SdhKZSMyOjD51el4fiT54IzxMVxDHoB9fWoXEhe
zFLF8VimehMBhimWlOO7U4Fi1gIyZB6DmVuf+tje6Xe7IFSUx+AlCgCN8YRZwQBZ
ZDjj0hQ4ALZNf4GZNyZsTSLiaqGRA70kFAhGH385Ev4KBNW4kLmLfK5RirkxOYAn
1ZXf9DX1SIl66Syjsww8bxRYGSFaiqArFX5tHEjt9Yh0rCtQZiCw4aGCTDUXiZtG
N+6ZEsZH8zS6s3os8t4CycPgNL2X/5NHqproqx6MaXPPDOt2HWeb5BEkzXT0Ecfi
RvEDC9jn4oaX7LRVtosF2n67HjZxd0soVYbpvltLUwH/A/yyl4YnnJqo/VmyM2Sl
/+QIYuxOg96MApYHKtP5LbB+gsOMBqNZ3PCDh77V2UFNeDrGNJgGZXmuJFi8fcH9
6KzmEWU5xcnMNHGkXO7JvWY5WA+ZctK4IKEsD2HD7MvKqqXEbcbTZY6ncRvrsQCt
SMTjpgAlMj4UTRZuLZAiI9feJ8XlrgEXR5t5pxwnfT7PVgZR+Yg/f44l8kOXKjj/
pIol/OZk7jryNunpsA9JkJSGWObf6XHxlDWhM1UJhfgE4K0jbUZhPqZp8/vtWJBQ
ycA0vUdABDmRrx/+5rRqFT/OgyRHKzz+iLQT335AzMrQ4O4kqPshJGCGRr3nbIcF
Kp0kc6PNIqqn9FapQwdAxppl62/oUN6khVz4ztCCTxT2Ex3IvATpA3FVkjiCVf2N
tg4vu42E4VNWip+qP7+bV5Z3M33NnvolPsoCslBCt1uybtK3niC087hBp7C8ksDe
aZlp1TMMaP3xWIhcrBelKjdTyKpj60Hsw/c+mCtZoz9kxMDIgpMd6p47Hsficp/q
jvBTERN/ba1u/R4iNBJoDd4ouYZ4JKDku35ODBDeMMX604beyurgh7z5Z2gRAWAg
G/tuyaNaCyLhvikm7YMFGup+vYHLNLOt7eikuzRukN64jvmd5vZ2dkkU8zd/WJ2o
A+ZYz7jik8SEsaFHIpUl4iXMdR9l+LHzg+m2oVYWcLG3tAsPTImPHx4T2NrNC6C2
xUe//JVUPbRmxQFEHEkUW9KhE2uk/7NRdXpmtSXcoRRTmk2KrrFy2ABq+XYWT5zy
QK028YRVn9K8gmrJqRZbn4+nTL9v059wkXsJcO20uZRscLLmsyr/RsJ7YkFCRuK+
Tt49H0UXmKh9j5TdY4cEtyN1u25UWeKCUa6F3g/16pucZcOlB1r8JR3FCFDmNz5w
u/mJaas321OS2VS65dgaF4PidVi43O5c1r61MKGN/jp26Tz9EXuKxmfCsj9yEvrs
Vb1N7lOe72G7zmIOspxF1MpEizKA1t9Nh5yIj0QcIRHReD5RPITD3Zx4t3C7Ws07
sjeGumVOQSzzcCd8U0KAhNQAWoQ5Mdls+zum23rUcwE+Br3H6TXUeDPK+yBGvlTQ
mRspzsWVNr7TquX7KMUex05W1qePRfXveJKyCwtItCQmGy0oq5toy4o3kFcJpr2K
7CDWEC8lFWut+8aR3Qgfpy6w+2HzNec8oZtfLjGgW1B8lI5CGLPvcfZzyp6jrRMU
yCw2XQ9BdWXklkPbU1C/uYeV2qXH+bJ+9e+IiYWyBt98tDRwh2B8talgjjrTZa9m
VHroAwLsjhdkyby/kT/cJHnijDQ9wa7ODTaBHS0jSoUhukx9QOSMXtcvfeMslffi
tRpNhkz/P6ieDd+J81hRuZ+fRuFoUSG8xzCZGPyygD9v1odXSQK7KsacFe/bOgSR
P/62EA56abVIUMaCRQpTo95ZxNHIBt7SF7o0PifpBnN5sDd34riQaPw8xBuQ3wcB
I7KWkL+chpkVbOdy67nwxvAFckcnhiok2KLv9bWyMOHwFJDgGFMEE/N1Hw3Jl75o
4RSd5hSnET4vtcJZA3aVc1ri1a4DiDe2S5lsfnhfnkrW6t5tHZ2xANx9jPHBzrTo
y8g23ABDIpOFqQNDoZD+HmVl4toQBx5K9d+bMPb8wEnPdeGBg8gMv8OLxEMh3w7U
QIT/pq8FGvS4xkrDewYc8rwFuXwbO7urmek72q0s5+mZF51DaaxkpGTbeur/LMqs
+9EIz/qz+bUkIrScbc6EsO1ObgI9Lhblen8CdnXrTNCgJ5NeKeBcur/ac5foozf4
PsXgjbaSDrpJ4SVwBspEpOF/VqG7CXdI/rFomLy/zjTSYKsHmkcrDzOYi0M7o34S
AyiJf1iAoE5agySB9UNxDiNCbFXyV1P384qB/TiE6gdDQVnNYffpbOPqvrZjT6bg
VNqBIapVQ0auvnUBu8gbHTo8troehkJvuVjxepNzzCQEIbksjP3qmakQOHvqCFVa
P4V3IyC+b2FHR69yVOd+2scWUliMH3r9I7Vo5ui8ryBLeAAKJkaBSH2dNh3aH7de
XvtmWeMczdq5YwEkwABJIl96v7+B7bkvzs3ZLg+YfXY7IE64iyQg1X+DXXZN6uJz
aaMKzNfFhyq4XjAWIFk8gM8+4iu/CnEd1Uka0Q6JhDv0dQrZI8bL0JnxbreQDI1H
yiEgWyaPbaNVpgOvC13URUU42exwd4NVJXAIpD0QWW+2h/F4RFNqHoina3v5q6OI
fkElk3GheRZhQgFkaNDIyxsVOVjeBCaztwmr+sS8t1oRiyuWunjYwoPzKIcWsrd/
sw+VekhusowqcV5f9/R+HpxA5CoiveR29G5abx7eo0bCMfWRugUz+XA2eORJQRRx
+WS1Njhk+wFzxF6NI8t6agdpGEhgmd/RIbDbuWkF88BhJBycRRb6HKdSGV+VFSm2
IAxAHNiLTkM/SVnA954ZU6dydXxfVSkNeU0RKQ9dxBSyxN2c2Mm9RuOgkn9lNpvD
at23SxU1yEkBa/YfBXYeDInWsQ7r/p0IXdQHRObvvoXI/yOzYuaNgP3Cdnx5Rmjz
qin+gXsZnRdBOSZEFBfodzVovTwFe1PlPBeV3aUyljpm+B1aA1evC/iqKgAaYLnW
j6C+/EihCijX/bJX3D+ntgwKZyoe2Zj+M7vJkrnSrKXqSvPc9CbWntms/Ktp4Irf
vQtGpjQ9NTHrWtooHjakfd6CVOXOcmPm9YtsTgREM0OPt7d3MTtVGY5CJVdzvT3C
lXEl1HJjrJau36H0g9vAf8goRXX2AmoAQvX0BxyazlqQLzvGMCdzhuM1fha/hChq
PcU8zbMUyBfg5HfCg3vZD/+fALDXG1bgejOQo4EgxrF4bQmR0kWNIelgkMyLPy2T
Skk4/NJloUTnfE7SPqwOCqI0nffBpN9XaVyDQO3aPAOqqOzOYfSvzpaRtvioMOBf
XK/Sciu93tgARy22W+Fk1mGeu46Z9Te2f8eUmoywAC5fGezm+pfQ0FQW2pOWxxJB
/BiwY9nUOyyXfkPpyZOMEBv/KSVcTt7JmvKX92MXuSuj9RSIa9tH9SL5iIoMekR9
sJ3e2ePzVb9ITs3cLVIpXVH+3SQikqM/7JpsUnWXo61QaNasVSWyabD6lcsWj8xh
uhNE9kvfJAuT1qe49ZiXCy47IojywltBczbt+28Nwrsa/jnhIhKFdKFRShkLqvgZ
8idOWT3unbdw4RLf/irnFtop9T6JSdGBX3sR5x5Xi0iTzh7wYmmvwhrGsZ6pxkEW
5Yx1SOPz/5FlhPN/3TupwsnGhCzx/S1pqi0Y9RkMWCqxooJ+SyI7mgpqN9o3PtdZ
sqHcbZiP88hMzcjlDbYcVByaN8/FZFbW4Jifs0G1iKCZ243HUbDF8C57YDaWd+XU
VeGsNaXzVgFAiW6mvCnuayh9SHjcGwzp6osQV6Eeo3+dtGW3elD8bI0VUDdQYyms
W5yfNwcyHuwYmnjkkLEXqwSpnpval6y3i7fCFaR9yfIHPXCToJFgvLktrADs1XzZ
kCAWLwAnwwlYtc8OvrpOr6FON4b0XRgc1WeCdLJ0b3yxOCD9+KSkv5VwPFUAJM9H
Ez6GEIjIfXIKhCSQYc+Jih1t1XvJ8DbQDCrCGpPtabEDhgDZhzGZ6V0P5yFJ94Oe
jnPgqWoLJrx/FhBucca8AfC/msWrXVg0ZyoHA6qf025wmlR3a/CBEL31jX+eyXN7
ZxHbQoBMOeveaIjkAd4vhrjTNdwVsTJk0/y5rtBCbTUgNpOqOnUOu4Gp6CflkP+t
ijyrHbp2HM+ef6SPW3Dg7NaDTK1hHiMq1ML/LSi09NkZ+mUg41qwapj+Oty1VJR8
qDz4xj/AqMbch08YJAQSH7E0ckHWnOEFwLgPsuOG/8fsNvAd+gtWO+0+ks33Ye8e
do+a245GD7Z8DGerIr9jU+JBw+J2ZcRX1/sA4ki70pOE08OnN3BFkpNCxQoGlKJo
yjAXvbnAYgf7rjNMsGe4DoJXBTkhAOYShjM5IzOAcKDFm97tT6WVtw3wFU8C4WoU
K9WaQu6w4WzUUwdgJDuD469/GJ7jBY8QYhUM0GR2bzQerjHDz7+TnTzV/3Grg0oe
6Qv0zixpdx+En63xSxTpEkcVGYy0dtOv4KkmVjETSDIxYEdsNqYN5ZLywCLuoxQp
I9+hpQR1Lqa/KY2DOD4kKOAySYYI6OmfkIBQr8mOTQcGDFf/VTOimApW0cS4dADG
bAa1yq7O0herZOiUIxQwH6uCCyjFRJ8u4I5PU6ski6Lmvz8P6Z30BmRA8K+G77U2
+wTpHgZRFdfSn/cN1ShYzWAEkJM98XIcl8iCBcdrejndxRLPgGZNdnXITM2v2KCo
ZKF3qtnF7jEJwN+7MPoWPOBl9EEzW5z+c8j3JzuRpp1SFH1nwKFake5pOcysbd1+
i17AuBCM7T6ehxrlH9HVs5NDJ/dlVlMzCtM1RNdEEVT78LV6r05HuphmKjn7cPDV
9OkMA9nsx8q1M3jHLAfeqsHEC0intCge15FN46J2Az0ebetoldRN3ZatFqQ2Dgk1
6KxfzbHo+RkW6vaWNXpsmRonc1ZY23XXGZlAZ3WMvF6m5jGzrGTjuJN6Z5lKcjOG
brI/DE8JTNDjxvKxAqhdTxTJbLUCicHnJVygvfdltZmYIM4qGsddv1BA2sO1o4nk
Fz/AE9IgL51SsFy6l85e1pOXWeqt8W/hPOJ7TAIYOUC8GJn/yXs9VCspqXS8myDG
4dm+SRuui7InQmQsfyhl6BUadV9llCdjtVMLUAUnlFPwygg3/4kD3Vr4iAyuPa3J
XbB0AVZ54gUPvnUQrwjbEe5zqH9iN/fYJsaoH9hcuXJ4BELPpJDC1dF4OHCAKkMp
xYTxDalTNKy23xj5JteQygV1SWBXkoTbXGPjrLoi0g2WyshGDBBSlNLRMEs/Jya8
eUpnH9QUk8RD0xpDb8G+Orh6CPGE1CySEY47Fm9ZX1igB6AC/yJJllA71thpnMHs
HD/NHXMjJMbjljKKtly2GFv1s4H/jwi+BzFy1pyGuVHJ3T/WmCp7cOmOBZndKS9h
2zC68G4S01DjD89z0yEWaMb1eijCGfm4M4vGllnmRs2z8hfdAkwFKLAHDlyqzKeJ
9NXy2T0GyiyVuMRJkyoZGH+B+LhhMi3y1w5+mzZ5GSptkD0HyjTAId+vvyyFUcyl
a3cwLwWAEly4pcOiQkCyiHg27AN6DGWydtra9FxlSrlE/OwCBKPat1mTjrs44ik6
SKShzj0h2mgXK42D68o/tkGzDq99EwLq/KGyNKbTs+W+OVea20fyZpRXfdaBMtqj
/dH60Ig5gmE5VztLGj0G6OWWPJCoN09NtiHuUbFrsSBStj0jNShvX9DqsQonMDTl
MR6/Qry+abJrIBd3bcx6ZVf4wPlfpWJFddc/bGsqFzGtBEpTp+UM8lOuYFtUle2L
d/4Nq+SK+EpvZ6b7fWt1kHTVtArekzGQeOUk1wkc5lau6Yc8e4iBSvYhEo1Mwk4o
1pTkrpre+/CvxQqpI6tc/QmXI5U3sHR/Vnxrm0VBXIRcsC1bD11xeHgqJpunOamE
us/fVMdq6YoCCi7xV+vBnCnx9y2IGai+J+pXu8lETEhFE6e3gII25S7jRu2NqLaz
ZWtWJ5ysyzTzTBkFLRFF7OkyD0CNmIPQrD8kZ24jkxWlmDQRfdSSXD1e3+FFl+lT
sLjQZQg2jvzyyzyUxdtEn1RUsVKLqO6OlMLoUoaNK/g15ofC7fYKpJSlB1GaPgcT
`protect END_PROTECTED