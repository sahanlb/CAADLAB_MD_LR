-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
KxvL1fLdVfqm0/zCzGs/g/86qHNcLH5PvIolfUzpWbyQdCiMvShWzkoXGev8sVGO
k1sEFBdaBDx5VsNrNF3J1VokUWGoNe77egNOz8p9VGfWRcP8y9Nwz5jReuMOoLA8
+qHZGXBW8jIRPE7/kEMejqp67kzuYqrwM24HTEGdtkzam6AeHJCMMw==
--pragma protect end_key_block
--pragma protect digest_block
5YQK2wCfC5Lw4cEq/Bwoup/p8z4=
--pragma protect end_digest_block
--pragma protect data_block
N2VfIvMaJPBSERneYQmBbg/otA54EkTK8rUuLAsgTrnHMvQ/0eXMv2awCinKnUAK
fHQTO0reruiboVbvg66yRa2a+0Sd8cKqj5L0ZLXxJYkZNfdxi2Nyd5WsvLTlQ1FK
Mta2T0V+YIk7hVCDB1QGJLUcfX/u4zPVVmhk/8B6ypvMVKulYPXWtrQ8AiWvK2Dv
jKaHjjSNx4TYhkVlsfoP946QqjmKAL2fRo50HxtCl0iGlQ6fW7OafA3AEuWAEHWD
g2xokTZMPVxRSJ7/hEuS0x5s9JdMMKLf7xcvzfLo1gS3PfSY/KIWVTByKI5u2pZ7
td8DMZhQ7/CAcVvntFrON7VA9NWQm3zGSqOGC8m8+aL88q9PIfQWXsVJ9wRkf+Al
u9nXuBvETq7PTd6dNRLBkJnjDgrzoR3RAyGM7USlm+OdXGYwUssULzuh8YA1nWBX
CDeAlBlArZwhMZIdFzRtacLspqmlOe6jox76Ha1eBhskMKRkMACFbEWA6MBW+gl2
MLjcrqub7BCrYdyk6HiaTNLkXP/d9O1XMBIi2WstJcO707vsxT9sdMtdYuPcLJoB
IAdAd+fvJlzQZt5v5FVB25frFZjhsnIKJXNEQ7lpFjPLo2PRCrdsIPqXuxz6FiY1
Ue19W8HoPpb627tInObPYLtPEu3pMywlNPMh3Iq0TbOAy1nnZK9nmEFzOPCPnmwh
OcRCuY0Ff3Y9kJv2NrmkAkdf2hs/xv7UeSIpScwaNWmpZLWSCxXxiY7g3HL91tkZ
rcuLiLhFadLxPscRj7hWHblXuqtSzjiLiZBu2jlLAts0GGvd7q39B57NyEPHLlrC
nO8r1PpTA588+IYNgxVwQtfpOKuLz2Wj4cUdg2qmdEbDb/zzhCgl0tWUuWWKIuLW
Q2ge9xlQXI/kTFWRrwkjzDVif+6HHLM2EFxcRa2HdGTthYKUVfTAVZRVKmocaiqW
xZJAZFFMc1Onli+JL3ocph0DyGOP7HeKtlhPi4ONrF1vHDDadPKmwa56oBUVO1C1
BBBIw0fVFK3R2s+iHWh8zSbDJ9fnZZocqtTLi7IPaft8oREJjIsc7sQpX8w3AukY
WLtoAOZrRhent2LWeJvOGyxZ/GNNgonZCGS6oWFjJNvv8icNaIWUPBHZInJWC5QT
HZcMQpT6IgdJBoDoAHrlLYhzSqrhKfzWTwJLo/vgtbTWqAD8PcP8pm3lCvS9rs6i
YyxwApKw+Gy42bX8WDODE8JaMbZpqnhH+ZDxlIu57Op8du6KAJ6he5kJTqSUgE82
2xVcJpyCq4mulEXhSjXarNaVKANRyVdeujfEFuDgClP0YZvyG8CdkaL4mRKYt8Zj
Mgtx93uVHYn9h1dzjCKnCvAsAe1YZzxnzRYkBrbeGgi41WiTdZoJDaDjAAvDLSkg
y3bHI0SzYqu8b7HfWPU+S2Ulei3iCT1C6jLYar/oH7TiNIKUPf1VaR9z8QwhZEIt
ubUszjcV1DWXu1IXaOr4GiSTvCNUja+hCjeFm7+UQj/NIDtl5wFLnypSUepu7Rd4
MbAPfcwlHMgOVcRfylwllGOU4tyN0tXf1NHA+rAbuKNKJc9dN/0nZg0isAoPPVGj
h9q5BZC1/RQkM38IkwkCAwWAyp1Peasx0vc1/VKF61wTZ/MmQ1X8VzMcKoi2hXdH
KoYVwrak97oNlqT5QIJ2BhryxhxKIVV1THSWURa2fJEZfRnrHWiq14cLlGdl5FB9
1M09twMz0C/8toZ2v4lwW7vzmGvtb8ZCEofMIaX6CZ0p4DEmNal9TdUayPctN+05
me/hYyit8jj3xrYA0b4C4ce8JVDQdrJ36xvt+mMidvHM6hppvWCrULQYSFfcQsQJ
c9U0CZaFkP7Il3NVwotUT7U29Z5KWkxN0Vu/NoywQpRfSx+HXMPzVBLxX6ulopL7
G7JmiodXHk/mXmAnSw24Gtxe8o2lXXBnWO2Tg0wMW+6bkQYrVNVQGYWLlpUH/2bT
jVNEUH9gyXky42oNHlWUizbisnFzx6dI7p7qs0ZWDVyvWWy3S7zsveGJNsCUrwHd
ajJRk+zL1JqFsWLFUeQvradlGYo3ZdtLcd6xBisECR7PUymri5BguL8/iHwtjW3j
5Kj988hgr4T5B7P/za8F1Iq00/QF2X4B1Oj90iZnt3naNKRdKCJg/5fVnoFoPUyg
+jKYSu5J7scT4Yu+BR5V74gkRcdlAskggAtm242thYUGNAFk/GVYMvSLsx6DRXkc
ciRWKfPFLeyxmuc4L3nLFBxjymt0ueXsIXF3c8yNEERRtUkBHaI5/eQnSbEVnz0e
acG0pc4ObtWqxTI2SzPIbOkZahGheFSyD/6461nVuVD43MRFcVr4lfX0etQZ2qaj
f6Z0OC1XOYRXH4PyLAkvs09nJuZ+1S6Kc4XeR7MDYlJiRi1SnSNcnO7omgfblbMa
Q3Ytc55oBVDUXi9V6N/h4m8ZK7dtGujdvegPetiOk5JOPvrhqk0k/YQCt0+Gf6E7
6Qk5oX93eereUtNMyBFhQhw6qr72+ravCXDdWq3HHmaj7bhq4VNHMTVQy4vjr5Or
ZlhP1QsHbFKW1mX4cgA7Z5ROtUFCvHtIdRuLflG81lGdWl5SldKQazxlCCsfkfD6
D+R522FXmJY3jSo9YudcpXTc+oXC2T+xZR6GC/DXymACJ8jwQB4v/GodcLNsvfrY
j5/23HZNb3BkKoT+Fp88tM/XMdMr+oafqyHkFgqcgrgEOieavxdoLSx5aRD5O8/O
PDxUDEOGl5WzktGKGqqLFDCfGL5Qikblcrctbn6Nl+4Pk1ITGSqDNuVZXtZyLWLE
o3B6BTiC4JOzGI0Q3Djtk9TB7I0gjUxegiTy3rpfJOKwc/E++kL+18TadS6CJ881
MH7ftX5C5Nl0ScoTUFxel60dUoX4WzXPF7UmizoVWkOwt2snxEOwM7XpDpkmbL4x
N7MqFtACiHciWOHTO80nqCuZrFz3Eg6bLsNeIJNq9tbYa8LkbwjYvvTaLqqRkX3L
JC6Hkc2dDmG+tIV5hEwZFPA5tRTmT8nKKA6X4GPxmydqXmXMSsiAHuyRxM3tUyqd
hkg2vmVHM15Qem1uUnHU98cVQCLRqIW9WQIkn2ATS1AjqJidpGM9bdvtV4u+i56p
r/Uz9cENrp3t6nSH7MP5tocUpbj3X6rChooFkJmcceprczqAQW9+pD9jm2z7b3mz
L/6ZM1GbfPHvXMImUop8Aqq4w3fV/GHAMJQ0RT++RU+QuJLB4EDw55BlUoRmsP6l
g748vvWN3noFfKtEoW4nnrVWQJSAjK1nQWciA5y/8LRRPCzwdE24XwXSETDlk6tQ
XU+W+FKIBWvcfmKepA8ecbwYgu5dUAc3ISUn5gUX5gMKMadejD7F01Mhlnm3XPVu
NbjkSFV92JlSOMYAQMQ4yUtAA+TUWWOsZrN2P3mQCtpReoxZl0jgik8iny95V4bU
z1seWVFlUjpFCuT6Xmzb8uYKFI1gEV44JDJzaKHytOJs6/jfahmfrJbv95Tkcpic
CBwjRqLBRDcv2VV5MpvYxrvf56uhfi1VGPjhCrXhbwSwMQr5NY0Sqd5w6qlpMyBF
stbNl8a5eyfSTfujcjABI6UAxt1e+lv9KteEZfc048gkrmlAZATYfWJP/HkTMc7/
fwwKDEM33xMYi2i4E2yX5qEDluCzbRKXS6vLAbvadP0LTOrP5JXJqREwc20QvtR8
neA8cC9gcw8qlbva4DX50OMKhrTXVM4t2uxLo40BtK0KW2ULMCv9vnSvg/99vPuE
z0bVtKy18MifJkL5s6/zAU9pYxac+aaSsHmA1Djt4eJ+QPoqWrQNYTCKlvxhQCyx
aZ5tSdKNCMdiPDqMeko7Q7piqDfXK6SnFNLjDzWTRQy4V4ErodA09veEIRFk+jIU
aJpc2HbczJRrMBBfBHLhxNUbNPnc7PWGftgLr1XgI6D+aAVRuxZCy9RMTUYnC4Qt
d7A4QW4GWDtVDSWVG/sW+UwMqLxZt+fgdPp4G6ZE59P2C0vhKfxXKIzy7IVk90SH
Xhquwm1uQuLp8eJQTQ10sqGFSwWSFJyYNk2qlZtGXo+GDQahXMSA/lzBAwjhN9Kj
XmKNGTcRgWmRWTZsFtA4UCriPv/0bolzyauMJEcZYd8c8+yyqNlLJ5Z4sUpagTE3
KBdMqyJ7E7jkQujmAITeZZToVw0X883Yp+myO7jrX5jHmeTEdtd7cOhSnveXySQ8
PGK9RhyCeRPGgZmSuJIrkXv/UYqVhtl4Y9rmBMSTC+4bFtonsTNq8znQJHe3iZTu
zugx78RygzNF4R8BaNxaHm0ZWm95JMLfXCt+dOjO53I0kVINNpNIqfrlbVz3y1ij
U5e4F3SEAsA7m84CUhasWvrhNj0zuLbGge7JABjgLrnPZCRuERMMp9JewD6zd1Lo
Q67q8wDuhJ/fARSrUis12qVKdrrj/0PAampR/LdDfZ9VP9nWRTP1RTe9GCDpLIkd
soZn7mWSyopg4Bd2QYW1JKnUh9mn41UKgit68YrAHn9LI4zUxGqsYLUQ8rQRFZRM
ArRDEC1TNS2A0wBF74LG9y5oJn2vvhX6j0HJYdI5e+BqzMz0cMfkZkoqalX2XT/s
z8qofJRlbJlc4FQr4xOVCFypWubFBIpz7TDIgo3qE3sustQX8dyUFPhhXsgr8GgT
7Fg+sLbMPzkdECF0Os0h83Q/HAcgpN/JmT9MK5Lu8fjjZ3ZqIQJicg1kcs6UHdaK
3+oSYE4SfJiv0vVaKAJUzKnBQuBTY8hwmNmbfe1IymE4jffXoE0Omg5KQyP3U3rF
hup+LYXQVuTFdGNW7J6y0+vzcbjPJJ5G1pcZldsd9DKyefKs+H74DrGcYEHyz2DE
MKJDb5aVMS7+deRV5YS8828GfuB/Xsj4dweo88KH3WiwUJX9YKZz09Qpb8l9znm6
8QvxFg9xx9XN+N4cNBsRmiueU2F2G/uMljje5Aeu/1cJ+zuFy1iDAlRMnUSNVM44
R9u3ZQ6BgkoxO/agsk19bu5szafoe4aGBeIFEzx9NMMZPI68ccNM+505FCrNre5C
Rfhu3wuaH/YFvpmsqgjLL3FvI1+W17lmkU5VfvFcZcK7e1UFZ1GiprHnYOPePlbu
kFBVyeLjwuRpoI6dm8WF9ZNe+0JS8ezgkFSI8kRhXHMKO4VpwftnMyMb5n5sK3qd
AzalQLATVE2+FaWuV8YtH4AT0wjLtniY/77ygfN3IPwZyu8qrvVY3ZpE0bd1xoEO
tq0mjm403YtN1UtPAeyX9AeI7/v91hHHm2D3cSqp2dbcRhI4LlVj/jHIiH0dPmaB
reScFXQjLHsJN6Ri3qI4W3mSOkkrVN5iuUWhogLIQAJqBBWbq2I9TtSij9zcDmxT
BeAvFG43i+rlybYY0PAB8LMU6E1IgqgJYlVfluBD3bk16eRZrxMjMrQv7E3fzCUG
IGUOV+Wmauk7mh2AwbchosdV+YrAdmaeqMip46fR9KoBo61dZU/Te3wk1KW1QcG2
PQKNQDTMa5UT+PpJHyKLJtuiMgVO8WRGyoOKIaXT7QO0D9UOWaFAsjUDgRwR6VQO
VFw6vme1tqW3Ri8L7TvNDlsDgm0490mYKDuM6qmZocataE0Jxzhy03LMUXSF/efR
uCgx+Vls2wti6gpvYAOWdcysTlpQrJfBS3+Jq6aNi6WzgISKH0UR8qjzJzE9eRb+
vlcPS3ozalUj7AjHoA0NO8HzPPRpPFGq/87BTRXQjAWEa8k09xyPY63Q5gst+uRN
pBc+8IO2rOXePmZMGRimIbwWux9TlAdztuPqFhnnUfpeyWM3PZg/TwzNS/MTpNPe
Zjdrfnps46MxqmTffzWVlP73rxmmF9B8v2G1ad42KwF59YVX+KKSkGarNDXpW/nx
VDiNXx8ZwNQoEY94Nk5mAJ8RwvGYQd2BpgGWgxJxFFBAurpj4UkI+z2zuJIi5zvu
F3yF1lB5JgIzcxyHSUYlqR+tJEwmEsHwFj3IpSUkT5RCx82jhGsgIt5aB/FTeJk5
sZcVHbKs3IRUzOTtt7rL+83sN2renk4Dobt9nSyTosUsKWutG15cHxIdw3kdY8Cg
k0Qlsu3nJ9x+FLswkBRt1Wop6xIwsLeFFFSE/tw2ENndeN/RQTw+/G3FEJyDTqxF
ZVNN9T90wCOocTFd1NGdQpcO2lijlLAED+iev1y9hggN/ZbNjddTs6QFXb0SqMXN
6aEgw5nVdB/MyF1kMV/Oj7paDyzjOUk22if7vQ7VAno8zJyicRfL4Rynt+KsHiq5
8rgPB6miBhB7rdHnvtNSoK8izpzQF8d7ZZUBTyhQHJHaSWYwb7GGEs5uM89HaEsm
BDzHZgVFPuV3JB93aoaQPWrggzrtXDq5MDX+FvjqfRk8tf3bJZb8VMgmRg7cl+kM
MhVruj6soY5/2yduZufSDxhqP6aXcRMzOJAYkRvl8C4q5abfFSJ45pQtmtvlBnpt
UcqUOcJ1Dsnpq7r4CyrL4gJ6+Mo9XLqsnIQciNuOIUM+J+Lt+hhmn90Z7wZ9WSKA
sFmo4xHL4+xa6dGF01NvVjf+uCTOWLnPyhSp6n+DeNnMLvFMqh6IcK+d4odf/XxH
EeED/lpfZEyItQn4rpTtD1qfC1uEGjd+q/qOYiqEePrSbAjvufeRsPXueh2jBy6m
dwKcLEeiRfF5FoAtSzwjZ664UkoOwud3pbiuj7Py1y09K2V9IvSyBI6Paw+8h1ni
pJH60ZcFzej9Wcjxk8yln6OadLKFu7D+7vU7ceMR5FG6rI1yn/vpy0/BpRAjflu2
OftlTbcyo6YtGge7tIqGghdgPaxKpwIJU8l36hBVL8f0Ii86iNrbykfCU59Zf7ae
RyOnH4W6VkAiTAbGPNpslqKaCUcpXs3lUyfOoCgK1uD8uvTDc8XbMbNeytZ4lH0u
hqW1ll0RWzsD1crgGdr9KqwJMS0e12LHV05bBueTAWRjjrZK0LMcqESY1Ti+FTju
0D2eulE2Q45j1GLqat0oWMAezFxhC3Z3DgyKmvkY49MTh32OwsIbXHKn3vmtcQIe
vxh7de0knV6XDoK2UZcxWdWYdhkLbgvqE0U+XgaSi07KDbQv1TsolJ8OUST+hygi
YK4o00YitxSAnlTWABO3liBf87XMDJ7Jvji/3fym/bWx/0nMOm4/HbygqvxUJh6b
SEaKU/4E9Uam8wGLbwyAl9sSKGEOmVsPV0uifPJevH/vdNnuSb+xPmQeN1lNvlRG
WNneeXZEwNDvxnMvw3ecSUWNOY5iXOKhhlMuaBpKIICTAi8uPxCgP4GBfoWfiusb
KvrUevjmAdsV16+44jX4q5BYTdKuJHCHmQsVAC30n7uYiom1LznGcK70cFDE52J3
Tr4p1juJztL8LrYAxacsUOLCE5lduQEQcnQmurBB2gNCAY5b5nYVjKUV/zDqjCOE
xLtYOXNttl8TlMhuZrpyybzy05rPuUFKkpkyeCUps5lz2L+Ad9bMVyO2IOeaPwJm
Fr8Ta4Og8bRfCVdH1/KF2vhh4w85a5LdrCim5ln3SZhfH39mtNZXDmU4JYvwbLiS
gJTVPNfO2UvT/bieNprDq9JyEbMRBKek40Oo45XRGkw8ldCpCfJHJJEB3jK2kyTa
xnH4iD71HOtMnz5S4brgofbrpIrnDaZuQxCTUAQWEa+8UfevPJtAR10RTJG7D10w
6hOCIB1sSchDBosJNXVDhmdry9SAkBJbGDpxYQiJOhrGQeX6NSnNBGHVotagMgkO
D+3vIXkr6Y/VK4EfExVpJIEFacXbmSyOkefRUf0sEtnNwOJxOXC8QLjd6tAQLiuI
MAYLTyxRL/w9romSB0bBfygefms395FVDj8wQtpYisiUawa0UCXgCskN3F9epnl7
f1VrkQzinOQzNht2DJkpD5J2KRlhSmkh+nEl1ya1y8bJOI9hmUg88iIo6WWMEQ33
rmAP1KC9o73WDK9Xsm0fCeUu4SoZgiRtQ4qY57LgxrQ86yKTqZQW6l4tWlXd08Qc
n530Go2G0NahNMx3nwc0yq6xX6puvs4cBClv7RoFBJPRiJHUhrmQSGl6gKeUXJHu
IKzF4FVOwzeU6U8lKMK2wbEd5krp77qvg/B+ml5wb3oe5aZzMdz3PObptPEEy2Hx
3z059npp55AMnlS8aNKluFcwJr0sMadd886aDYdzCLtOnUV7Gckp2QtVRGJvwfdW
B9kHTPq0p+ZXS0K+SsCdmwt9FPrjEEB5H27j28ldpTNvgzRQT0eH1nXeTLv7gKVS
8h3Iq7YHJwb2foKUDtV9SEXfWU1S7roBXw7VikPxu+RHckgS4YJonqNvQWghepoM
6q8CuyPN7N+TRe/YBXwhI93nrubCUMTogM1e4OlKNpZPo93RSiyM3m64Ewat8t0Z
8QiJNOgJfFxuNTvOXgcHgqRfdTr+l40w7O1FgScRTz67PhJE9jThzyJ6J4Cg+V8M
i//h6ZRzrI0+tBeFlAe96R0qTQanghlQGOqs7yF+wKy2MAolp6cycLcFlax5aVt0
vCJXCpOQcMhVi0aVAYdDUh0c1gIoouD2e9euBznyugdFJx7iVTymBiwOMofZktr1
ak0Su2wnOkpPmQOk0wFJpvmaTEZLaqDpSZbS0vh8lRg+SdLUs7nkt0o5GbNfDxJ6
faAzSJ4WEj0pBkxzRuQp4kXvZ0oJrozAsK6Y5Z35MrI83NltrGR+ahgy/edkMTXS
GTtmqOnrW9xESwc0CdKnf/6E8+oZ84leBXRnnS4wCMtnIfzYaXto/VyWytTt8Twb
Ndn9im5C7DnNYxG5WhgwdBhv9VKWOXTPfE1MQaRQenuQ19HXaHIC0xP3VFfswglD
XkKXn/o6ehxc5hLRymGYpDm43YAlg611U1lxHYEa8elNCbO8C4Nm6YmlocNPsjL+
CsF3ni2YyuFAk7j451VUQ1BAwFC5ZRbxQje8cHLykB0ZkrwHEsNkxzGBojBovGoo
IBbakoVP53xNRpdu9R4jv0id8s7L2+baMbDDWJMj1yUQnwEJwGffV5uVEMkHAe+e
wEVpmV19Ct9TL//okQqsaPnRpne/U54fv3ii8CH8FqoZ02q0laV4A08aNHjqChQz
PJIuiiM0MA3wBRdljpVNCFxKgK3lqpb/4O7wPvOkB4wu//MqluCwaX5DmXp9Ox0H
Q9SD8t5qpYXcuzebx8tFrdRUhFGBuAUSSL3NY5Wjm4G/wwnzzMLqjUmp0qp2OkAH
UVbDwf02IXNJbFuCMSPZUntzKI2Fr6yn/7VncwpzbBekAQ2XplboCvqz4LVNhyV3
h641SxqIdo+9JxQdwev3Sq6j+x6sv3HWW3uPjDFqi6Qe4m/RkKTOivyJpdBIBvL9
+fVixpJkjTfP3u3VoJQAVbz7+2KjzzW+rIs8xJVC3QlpfmxlPfVVX8tfjh4r6HDe
fkKVubi7BT9UP2do1sHlW48bmDZ0ypnCG8AWS9nBq5hgUv6G2ctuTgYX6nj7cjJO
g8ba4fBdK+YLheAT6uMjAY+24h0Ve9qTKtO38VD4EHOSDuri9AMneQmVr4TwI3NM
70ZDZna2qWLe638bZwU7NYdif4PVXeh4eJebd5gD+jdRD9ca9dBrPZWc1h4fg9PW
VZg97n9sDTEnjkXsEL74XojiIZZHS8p6HpLKquiu+ZmXT1pttPMwKPhhGjWquyDK
mvM6Tr3LTlN/6Eff7mGrneQXn5szzh+K41Uxn6f6bzCPRnfabRvdTKF7lhse5Vor
jX+bgraFl4wEASUOzHvyU+7sln9UfNiQH/gDULyHIRhr2NXwbYuhc9rWZu5IHFK+
EBoz89JkJYQ6WvlUhajfL/rr7U+14dtLvZEICAgsYZ0Pn62HPDYnAX521yIs1+BK
Z055QpXNQFV0Mw0ADlhEWrF9WX23dxRdlvtTGXRF+qvNd8aJPajvg9UCSMmAymLL
F4ZUgcPDk++cO1P0kxkXezQEpZKQ27zekJygfEWnsS36jEV7q5jBOjix03DJuSj+
D2AAFsEXu7Cxa80NI1HJV2AXKUkFZ/e+Vzjvc13oBYkXom2vASu9LuyVIDbtGarK
6FDXu0ZTGmY9UxbI5HbKlFEVUf8k5ar5A1WedqrmhLmYdgmiWhcwNWC/bIO94Gqu
hSJw/X4TMo3TzN8z/0U1ifWpfgAT1ptEtIRxq2eGsA5KId2cTdV3J752DdSKxWUw
UJN+3zDXNg/1mE8DGOWLHqajGFZMxsCJBr3gRBLPB2SharF8EVGSm9EPbPpJO7Fi
TNMxP2Y6s+xXEKq04wKEylS6W0kEjjEw1DxgZxD4XRX2DBCtB9AttbaneH4OG+7X
a3VxpBPHEATws9YgIQl9NHR4wRZ1+Uiz2y43XOgnDI33OgnlKRLOR2mwDO1xEKtw
Ja0LkFWgJTRK8tqh2AW5DMgqfUyoAN8uAo1ntB2u4/R1tcGDTZErywLOV5Pp7UM/
mPnfHz6tbEbQb/Ll653tO4qUXCQmN2Q38Zyk6pNr4H6aHXrcmgshcTuEhG17s2vg
R7X9vmzBSj3WI+O7bX4jWjumpXykhI80PjAauSKYSN769WbQl8dlwhf0LgVoLlHi
QEuQPCiOZj+QaCxkECevtftcGwLBMmnqNLFq98k+En22n+xqv8Gv6BXjsHMI3OFg
xoaXEhtPPHy+cH7WnjFgbmEA7RULzZTJxPKgC4rsrPzRJbgAW3SQXm1e+Ghg/beS
Lk4rC9hkYApheQ0JNmKnVaM6PCrh+bo5nXr5YKwZyqKcguPHX22nX7neobka0y/K
H+O/mV9fY6ehEoo+hHgfw0SLCmx/XoxH+eLLpu/x3ZIVdbijSy5Y0Ad1u0JCjFuN
tHiJ3ZnyBE2YzUf2nqdDl6/jVUHPf3/A9Rl+k9b/a2a/R+j9wI6LKj6CJ2nkhZzT
1VY5CqEw3hF3xgb8e6Zs+aLGPoDzg5BSXRdiJxus2BNWc834k11oTCn98HghD1E7
2ElhFp0uT6cUvLHwDFdzAebmG0sjuIRVsWUxd/F8/S8JYqNMw9K0plxRJ/aWWmcz
EIe6UEGGhblQdMICABG/Ep09wzFbmddUPWb18gEy0yLjeWYFDjmJtj9bs3na3gLJ
wl4ve/i/CrGOUTjRYxIR3bV+RILeTM8sjjTy6rAfaUee0YH+tSMBkV7AnBztoUJN
9kM726X5fESJFIvZneCuI37zuFCkOiAa61CJzgz8pmfeKZ4L0TpI2A/eF6QXLezZ
FQRDycBEr8BXJ7vubd7NB6Gs+4otVDynbH+Nbu5rYiaiEmzNqDAqLL2yIfDDhxOG
ltj568EWK2vpgKxxWO5Yarkw3xHQ/1W7wqU3cFc4nyeEo5i3H9QBa0Fx6yvTntSl
d08JDnWtJUR77x+gSZfJTg3RryYK5VpKkbOpgPDv4MTSQF3dUKCztlMHKTXsZdjY
vNVeeoDkTawz0wyFAPMQU6yVm7Un6eUfzsjFyfzKSXFgPJAPjyWS+x2wgXLb/P7/
IlvakP33LFkZW9NF72Xw3aOcrhRBoM3zDq8zFDGUnOXPZJiAoYEw91xIto2kkyw9
LyIl8sWAJQ74U11OPbBajDbbO9DN2dFN9TwDj/QtmypgLM/k2+uN5sw/NJOiEJuy
F7V8B2ozOTgvfqGgwXAEVkk/zloy4qxYWKKFKZ/HFHuZCWIx7Udl7ZwKJ+SY90Mj
0eB+Ci6Bry0thyDCG+/ZBiDwW2M5/RKoo4h7xwxZji9ayK7nWpBCNkMKba/Tbgeo
yBWYT7gXm4htjUGQ1EvNNSE6iSLdTIGQyHYpqur4pxmR9I4M+8rN846tAbVcoRdE
McRv3Xd3gJ6Ueahj56etuQBzv+pdAS+SA6nWsuxuSt7ICeMoj6nJiNLqREcFwMNJ
rPywOoqQKXFO7GM40X8PJn2xRIaanHFq8kH5sZ8viYt3YRB+aJU4B+cYz8oZUgvu
Y+neaFb2RDUZJneDW78erYfzW6JRrjcREV4qzATYMDNskZsR0/8KE42jUJZ7GTm6
P7HwPrJD9+tod5MjTc4HlMf4Sv1yjb6wX9Kbws+C4/g/ONHA6Y76eBssUKhSOBzQ
2OjL1g6hJ6UdfWcC4RXCKJ6eN41fbM+TmHVF2a9qjTVZUTt5q6maF/qG/pMmgU+G
gfWi5J2o0gwIn7LSrkkckw/wqJCTJq/XWg2I9LUtetTEc0yd624T7InVCqGAf0vi
ZaYDRtNQxLfUI2I36kSar3YG0sSrQhLb6KnUVl7PC3RI/V6YVoGNTaRJPP0qfJdy
9SrtpH6FxxlF/aDFxZhBCDkboh92nzOFehsFHjv+G0UluPu665vPjj87vZvM8ifj
4vMiVA6EUwkTBWks6QffbApQAMK3SUTLUWfYJygQLM9yZImczqREt9/eZJEzT6Tj
LpJUXk4H1M83cpHZ2pApevFu5Kp3OzpBhDGiMTvADouTN97IuLrd1Bqpxw3Cuxpz
c2o4TkZZsX3Ry0ql8e7bGpL+EPMN4HuGE6wGpYsB8rt8NhRLsWKNi3xjLT/8JpPa
5rxIrW+Lx9GUJ+YTFWOzenf/Ur89Qp6F7tUn4h5fVfJOwJG6LjruYmzvjkAsYiBX
W+aAxswZP3UZcmfsTSDW6qjJhkX6U43tMvfy7a7lADzkIwic8TlISXaKX8t6c4dU
ebIt7gsMw2QP5S7UnedmFDnHYLq2Gh45v6kmuzxpFaXN2tKtHfmasNcSOpPoNiQR
5rt2Ju1CpUIINolIbzih+L5wjSGBCvaxcua3aA0XNpRSXIgd0PBdSN9OBH6FKlAt
hdh/Xp7h8c+Wr8v283EqI+jWlMQSpQUAYYHp7mJPkS51g2d77QLxC1f0W/H6iB7q
McUyn60QIkju6o6e2aC+emTmQgZ7vCrl9v4/WyjdFhtN5BoMJHpbf2WZGEqzDbSB
h7wSeICAEkmarBeDVD2Fg3D/XscigF5Fiyyhl69dD67QNSe6mFDuyqIc0G4L2l+e
mbY98cZHoYJ1A55FBEnRt882Ht8MQFq4G2sADgz/PX64Zt//PV0YOWXL1hZusL8M
VubDVrabg9tSZgQslWDkCOsdhzj8RD8omhtH9U/9T7h2U/s3EY2CeMKHznYkZZOH
/TET5AJkwTdRBW1nvqxTc/yI6GvBe3so0B7KxnQ9r3RPUwrvRYhQapTRPnXqG2ey
nXUdV6HEnUYwzX4LwjAolYTuFI6x1nstVP4OXmpdl2JhiKz4AESmo/Eq60ir2kuo
tr6AnTY7smoulZt3BUKRBYLIUiRj//KArNfeK8VBTiW4MEs//PfdsAvKmf+wTTff
bt1ybgMMj9MCDdoDkivkRl8lvImNXBCgbGllc5waKkZY52IzvU9RGCizWJP3JQUf
B08gCNwV5Y2muBzPRxvLmkh8S8uv9ccNMXCKxpKPKBV2N2yZ079R9/r6t7CL7wj3
cxOFi9yfyeq229U5k1A0PW7S1OZfNwFBYsPHsh05wfgsc7TkdH2bEDx4feV9DZWd
c8tuHW45OWHst+1z2kg+APk6NiqTvsiW2c/VGi/XRpbChyNzR1QPry9QmvKWuGy6
L+gWS+gmQQUf/AfAyPfKV52hmsgJOhqTal23DlcPEEnijwRSyNPLHjUyiZ1stfkf
22/zWpz8kHn14EnGNelDEOglwBi/MbfFRVj9i9ER171c6SqeSOpXrWFCrQorGLSC
7haUNbAXuU+EWy0B/fa2HYzFa7JxKuoXX+ZGVqvvx0jGVUJ9uOHfGnwkJx9NvuTj
cWDFxnmV544bTSM4i5x6C2qF9QWt9RpVhwQzl1gGRKOTZVrUVYEofO/IZpEKZg9W
2FIq0Lx++CVsQJaB6DEbwA7oqS27rzbbuxuMGYPSXQh+yFHow+Jtd9Aqg1XtT8+W
O+4MH2/5LjE8S1JQn9/ujRuZbliiQkNeOGt9lLc4jV89vIo/B7MQwlzGknVVDhAU
daobilasjoE99Lmm5gacZHHCz6oBInITHQ7JsXOVNR+wEHogtJewoQDyjNBZKiHh
3wCE6nv9+D0JMF6G8uvsKROrtPUd0Pcs7prtonnzsjGNr5b3PfcSgkrH+LtwaXoN
8Z0tLxUzc088TP1UUdKk5f58fjVwWcIfK9IlgTPGi6jP0i3Rq2CODAD9I0fIMV35
UeqZFeRuIf0ozfEv8Km3ONcY0wPlzYTxSq9zKOBR8aFRyWXpRu2j1tDRSiVhKURn
NGp/c1aiWh64KHd3l2CFUQ1E/dEmdGaHqHuDsJVXzDfwLs3MfHJamqUBYGzbxaMR
iCJ6rOzTKeziXsmQ4h7RQLa9JWXxjIpI72iRlAn7CIvATOX2PYcanpLcENmLho8P
M2h7Ow4y0qGHG6iDA/TF2W38q63wEA7mWWpMbR1odAs/NxtXOiV5nKp260glNix7
/0OpNf3SOd6wlitvaUJqIH69ToAPoa3lOc3fcZ0vjMdRxOf49LQ8WghgCq+O2p+R
fr8IeKlQNKp4s7cJMEAsxJX3DHVB9WELetgOTSpk98AlUfiw5Nja3in50qokmCta
m/hnK1sDUtJJT2+5beDyp5ZH4dhIqnkN/J+5cz2mpSfCBx+pRfvnjzbOgfXXqyiD
9CWaQ42y0fiUYIRYnU50V1TSYJsQBYmWp1fwWvtTJPwXzaoy6pTEHjDS4qFSZ6K1
gjOfvBuA62L2CLkWit5ywcvxxmbwP3ToGWDrwtzsULDsTqV8uRUvUhUcK8LEBXLd
wxit8ya1skd4/p64F7ozM/a/FlfJMbq6Glf2j71t2nW7VqhmNmpIaG6vnyQukgrH
2O2pU0IrrfiWDACUjsCzvvDw0thDIFSiPnteMmPFGLEoiN5uHCmLQZ3OjIybGrlm
MpJqvSniX3KJfgfdSbEEDMm9AsjpC2KgOI11Z2rPov3xu1a3HCDNMSf9ngQarJjt
qvdMXFTcMDH62H6tYbuKBRw8vhyptZf8/maFTJU5pVYymVLJr9S+R3mvKU1aGhyX
VN7YJuaoMuDlBKRnNjAYVv8PCFY3xjPn4KyxGx0KNFMftodt43PQP5RtOs5O67J7
E9vOMRd5cwp24d26zY52li4lmd+6Xe9ppIColzQUzdrclTylwfvZ24D7ZVbeSivR
wTC1WlMRHepsN7umjUG83xIJcfyhp9Nf1XyhmvDuBWJfCX9IT1wfLtS0/PipqcmR
t3vLZxCJzP62Uhz1MKjD0sMu/GzUi/lITpqB6aoOrjZNzqp/9bGh1jFBqR2LWz/c
37UE31P1PI4A14MxxdRaSKQIRCqWmXYp+hPFxPFtYAwmgO2e8r346n+G31cDmgFo
skfckJeirKdPEs0ZmyutcVe1o31Wxpr0mR+CouX+uNGxWXYulgqwzCDMXo0HIgxT
yFkMvmY44srXzI6TJQknjElzz1UlH15Wi9ew70iXVyqpePdzp5CfUJVXemxEEIi7
4D/F386lezx0ynYKW7UXea0eaNU4jJrw3aSLVBcbrp/VNsM/DQomO+sLqkDWWh8C
WxI0nzkF+YYlppzp2XKguYARJz2xWRLMWU8kIpUoPtRcv/TCzM0jGLzLYZRU+8UP
UB0EsgCN35YlTjoS6mRXF0SfFFkr5dFKCTpiLmsQc+gDPhlB8FLoCMgyhdcdnb0O
wkZhy1nq1PhLCGX49yJOJ7WuJCK6hdCr+FnMLaY0CD8z2zLq0QuNapshAtkva2GR
8D9ix4cPBtgDpIgCF/uD5F0IQHu2UySAsM4yYVE0nDQQL0XHfyeuMcWrCJa9pRi7
xho4qBKBn1NwyzTt9jajWhe9tLIr/rdP8ebK8RhBGVSq+2HYv3EtjoPNuKyoZc8s
mQyTIUgN02+p3+yv5vk66ZCt0S/OtZ1DYVLI/qjaGSa2eMbvmaZ4nIcktkZQSSJR
EF/3AhoAlQg2MTAaGkACXn1AwBzQ4Zm2PG/64QD70PQVaRv0PZkwwLAGyoZHZYjN
XKMtlwUHxJTVv7hLwx1OIA4XoZbvtWPQznhhVFfhx+n+y/Qdx8vVCUeS+mv4sVIR
sOupZuNM3afrtWfjEdhcFkvQuv0Ib4eIfkSD2gqK2ycTlii7t74LpI8SanSbQk08
EhiK1BJxiQPgpoxryDmpkwo7jm4lkmr7UHFTLbA/dovaQHGt4YO7zC9vaVF6k5Et
5zlFLeeyMOiYDNIMrX5eguvwPx7k927EeRvfiQrxiRACJ/J8Qozd2lmPwlmHf0CQ
rgQkFmH9L0ayWxdYyHTwaPW9pJ+6KmtJ8+5R4YKBx5oppuXc1yeSNx1E/Fwq/goG
/EgGWN+yWsWEXKj6pAlpdyx6Yqh5UrU6aGsh0uwJMvlm3iqaPTLa4jTBJncL7vyt
D3LEylfyJOXeoiL+mkOiCMuvoN5qUBUDStSBnZPkJknFTg6wf5Nt/hfA8xJG09HU
LNIAkvFOw8Isno2ARFtt8QCnER8WEwJkF8yiHwQ0cjKBTBUvcaEgj9PBkBINPNM7
FKa7UwPRA+G0FgNvZ+MK13XfMWfJA8p4EEeAZx6D0U+v06uR++xU2sA0/HN+/PLG
B3EB56zKmO5l5h7I/K3o6hf/P1ZESLKDZB+Vi1huLRgXeE4McVTpguMf1hUx9/71
I7YSff/e6MxS0duaM7UK5XeRCVnrN1uJF7KxxalUGW0EdprACWLddvJG1cfBsbdR
203I15lbV2UaeZ6tDG2to7C3xIF/+CJyehldf0Pj7uZbNqzRDWJ2tnAkCzV7Pbsy
5+M6XhyqU1hXKXwfd/PLun5Hun06cBhci9VgyF1covcZRH5aJ8Ux3M/gxRpuDOfE
qfE6FR+Nr8DIC2/9YvAU6amNGBnUChVokOdIMqbDQOUuMYRz3CIAv5rZixRL3qJY
WZwGNoxcxJZeKh5ZuXYRSz91xLUNTSlBg64rMRJ9OYqLN8mfhO3wttLA9vUAp4LX
2aUQR8XaH7y+1EHtWz3pMhtM2Gpxir+WFrx0VbSu8dxoNvGkzAnwEgdlyVAJLvg4
I6Nid67thUYls4opX3cefboz3alCZytIcmhV5Je4/aGX9brhPVPS6L7p3/g1WWEn
psZZ03ZiKiY4Sux0mjFc9mwQ3dULMdDTCxWBCxmtJ3y0OUYb57nvkXLmX7DL9EWu
aqI8zwVVe/ZZcfjJoCq/YDfJwS8wafBgRtC0ibq47IexbBNuUAQY5OoTDAdBpsir
9p248Ts9z8U6yipEGV8oVPJFtGIp/oBjnKeoATmAiz6w8S72aONdarVJtG9XZXv9
lz6z7ZB7cfGWEMxVbFiBaSKkmUfktitSsObSoH8K21cFQmncE3LEZWRM23zpgpwl
EOB5tVS8QxApNsyQ2wEVjB2XR67sEH2ttU51H6N8/koGZHAwkyHccw6ING4Y0Ej0
1aIQtbpWbDbpwaFRtAZGR0kfQxhERHOB/34FZvGSOvvsH272icaSo5oZLxB/pbjz
iK1EEfgkf5/0vDniBrwcaWrPPQsymoNTBv/24+0YOO3rdfn1Us9xmFYwxwLQK3r1
5AAhAgy80gTp9XzsHkfXOTXD8pzAkqgOPd9nxa8+45NCSfFKMWlGMPZo80P3ymlP
2jP7zbaeoFRj00fp6iDO9Ajju4tdelx9sE+Ir4DNb9scvghPVaFoqZL3SFQjpUHu
3wk/WG0R7ZAAplVmi3YYDxDGeN1XBWMry6/ZL3WZw1H6DGTcf3f6dnc4osrw/EpV
D28H6d07Jr8ynj3Y9rxH/AOpseEPJ//Q6t5uZqzTlIN8Um4srAYfq21Q6cZxJmDx
sNgK8dTHVzSOF1KW/H6gDNIB56PPRGGw3Fjyb+dWZJWR0mwQ08CVRea7Dwoj+7y4
x37WNoGO/B+mdR3cT9QzMtpF0ZGSsvJr5tVhUf1DM+viLPZr9LZFN9sLLK+1pPh3
BNrqzNlasWVfMvJrRrpuoOQpG/URNjpzBnDo76u1hskYVNO63GJfnkEA6UGbkUqQ
FMclNwQS3gqaBztBAH+DcRsbGRgBX0lKVU/QqozLEHPq/mIFlQuC4zHbgB5z22sk
wL2YI6p0FZFbjunR1lmQeEvX6E4CqB0ZOuPK7Q/fTifULQbyfzz/7mEMKKVmbVvT
lFsW4qqaGfHoU8DLMVoguzK5SklGZU/4Xq/NDUPooln/mmk9I6bNFbtsoSKTjowl
HXlbd0wrMiGY7XkI1RyA4qhtsX+FLg4syiSqGC3rMTTtk1+HzqxJXmrJlIucZeBi
gQSw2Fv4cbUqBcoBBvVkbiYeKAa9D9pE/QHSaLuM5TXU8T1WqfCfzFy24uTJd80S
kAkE56bIq9xhUuSrZL5GXCP7b43yzGLwHOPYYwKw3EJBCQQRUvEZZx/qwvvtvchd
lEL9EH3znwhIIbh1TZBF2d16J+hsIDUEGTHXHUiuCanYVScGwXIoI6r8PvXKdpN0
F2nDU0wDSvcsc5t3udhLUNAlKZnqDQRaBl4m20xnuDd0f1x+gv4g/fxT/dNufbS4
ZAR1ZoJ6iawKNkA5wXTdXYQFlVb18Aqlt+irzOvC5nvMo9Ik8vfr9oF3TNdRjV9H
U/aVngyIV9DM0d3aB9scN8B+whdOK38fawzUPZusSmIEjnYJQSzK+X1BbUhhURCl
M9ECkjcpl8/xzCZ0FxPHAdfw5QyClfrjhjzIWfUgm0Y6/yiRrkCVImaoaziLDJW1
v6iBvbQFANUhnJTFewpHi9okQ+YMxE3NuMRQL66GJpGEwwhDir64HIpWioh9Rf1n
aFsr7exhceYbcbGA1PTV+AJbEi5FbgwYXuj8eY0I4IGJ4WXsEAGeXPUZwzZ8k3Qy
NwiEra5c5rkS2KTV+tY0/hgiTduTxD72nUPZgk4azciCDX6gq3U2uMn2SGgtLIhL
1ENRMST91AEQhNVLfluEZFPQu1j/z6grgbWymE72yrE4f5IEnMULcdaT0rqVeHRJ
AAYzYnZ7wEIyUyuAfQQjJnLuo/6smoBIxgAX0Nb6MX1R40jPhjFc1QZyqSZEIPVg
YcGbRGNuJZ6OPWSnQShNB/NbKXFIJ84G9Qev0Ej+kEnDJRwp+2l+E2lnZtP8azKe
7PPhId0g7P8Z02yx5FR9ojTnwlMp7jbM8zpYIQKMNX+Jgsn9VTuawn03y9fem+Hl
oAV0TIH95dC3Zu5ePEsebhkW8O0tXIz/apuP0jM77kfjP6EpnIysOgSuyD721ObH
bKoZyt08zRF0olQIaCR/9gdEXMgJdMGoB0EIb23BVDWPVZvGvs5c+WozPs8m1gKt
XbEjcyTXAfZMC863kgdlMzAUaTByjp4t4jOWgSfr/RybZP0An5HPuShthqDLLYH9
Hln0r9+FY3OsRJG9nC7f5ps3ayLyojwFnk5OFimEEqnD9oOW6UTEw0XyAXDkWVDf
BksJRCGAc5tCy5VkYcq1POyntqslMM5jVj7Wyb4a4E4PuU8no5so4xk0juiBeiR/
PuYVaCVzDdCS2ucW+ntu5FEH9kk9iAZGWK+8CKI0WcKV2z/JOrSceAOQoqB8SH8z
y9GzlwY0KULIbAEE8QxdA80s2kTcfvHo8DTvEIlz8pbSx8K6zkPVTdPZlJbrR+NG
nyFwW64J6f3g5QTnLpe+QjhtD8twdV5n6URyE0tRN7rZczf1tGnR7bqrJNF6RE49
NVhS0g5F7nk7pPgjqMerM/qfL8O8jbzDFd6Wd9WG1gCISbJUA+7ndnlxkcdRTuYV
dMXVzqAZFz1dajfYTftMvnHNeriuZfc4HlZJzxrpWemWBWC4jzrzHvteE/URWvXV
wf6bGwLRDrqoFQvXCcYlsStwwwkm20IJielNnKkZE0pO5GRHp1yIa38/7dmHHBHQ
6aRBkgVZ2CfW4MCNo7gNw5wvfrAS8KLBW6Xj2+mwXZbK1GnAAqv9tizyzNn5Fwvh
vpewSBB9gO3PJIQ/Wnzn4WzFd/XZhsl3TeRD0vLybZhPSXmgNtCi5KSV0ZtPJlmv
QmJxyDOhiXs8FF5NtHbEl8DVDLqH/yWg6K9HCpVgNKn72K1ytwDr4zvjebIsJYdr
IFdweuV4dLz1237dxMuz3Y5CG0yWk985uoIP8IUqZDzaWhMF0/iDefkoKWeS15mT
jVmuQAJ5tBGUnWR7ggLwgUmH4fjk5u0gnZiQ3rULJZBixoZm3MRhi332zOQkB5KX
xwCx5/yZT9t0tyl0AwGPucREHDHn7HK/XQ70uJUtdApCwass61oOg/fGtmau2vrU
xdEQetR0qQ4iuwiFuhQ+VaQjPjZQ1qqfeFlnwzyjDGmO2Ju2NWLuiJPh1/bebBgT
Kbv81GOVKu+GmZsmGtNBYBE+CbOvCEBNC17LO5bsaTEUoFRExxNtld6hZn6iKMIy
Id9ek/WdHP5xkgKh7awazpYzSQK8lJpoRHbU0wJ6I7SE5/VTfMXROYr9BAXLqVUK
VJPnQDxAGSuo5PA9iOq0P2h2a427mf8UHycPSAGlxPk+rzndXyzBSJL/d74PtEc2
ryXrrH56U1dkD41YEF8vcu1dv1FpUtbQiDxOnRUm7Df1bJnN+Nc5qpWDo26KTKU/
tmdcqCcKM1AoFsHfGmlyDUOe6u2HhKebi0E7m7F6FCJOhziX3dxzURjhzPfD8bQ9
ecNjCjtS4Y2ThHBS47JwtlMaLRA9NjsVRyGm0v+jU9yXcOQ0DsQyQkhN5EzfZ2Rh
c9XWlYveDcHggaPBJwrFYLIgATK7u76qP7xSRpeWYaGSldFtlgCLM4XnEQrv92au
4WWlnXWS+rlXCUw7htRLd85a8LUY4SFOYI5XP+d/3KpqDQ/dlsg0/y4FxCcCk/Sk
YXHQXAKJrxnerryEOJ+Ms9tSg2l3gpay3ZicBpBK5oG5+OmtMuDeil5SUqkqhG1J
DZuxqCHMZbOFQRTJ9nlc7UXiZGaD5jaHxkgwNHKU36WDVnEKnXZ+C5a/NLkgQHnC
KJVR7qI2ltOMjR9J+y27SH2IauryHZ7KmPm1r+l2D2qEQmoFr+GM5alba+nDINbT
OlU3dLPOIeEvfFT1V2Oid57vOdogcrOhs4minHhkcgZOKsMjxLe3RVyOAisSCUwk
S68YHQR4U4LbuhMG1jW1HyUKQ39FxUbeAGcbNEVSQAcZy9QrFS6IMhZ/oeGn1zbQ
oi1AtTvkpz2HbdFotQjQy3fcW0r3+ml/DfYsrtyjANr0ixGT4Kopne4VSlmvhx7u
b2U9PlCJAMtHIJtITb2J6ipU15zye9JIVm46PfC9gBHGTye1D6u0+GFPj+idmMS3
nz4/a9fzvhdAA9W/leJb7grwjqpIgZnSZ40/nk9Lpe4IcRaqoZjHTrvCFUh5OHtC
OrKyweh8GJSZqpsLy87N9VstSgIXvhij+14he8PnKLnZegfY6mD5arylVRO5iRjV
BW6CZ6fLABBAKB4mZDVBqp/obFhAXvRaWIJ/OFzbSSsXgcQ0MWl8MliHNT0qUshV
kaMA++vLNGHGLMmbIXULCRjujyHEznrI2xbATbq0GnJ/VSCCpGr6hRyjNxBKJstB
EJMaKZSRKJC/+rlsI7vCS5Ywbt9ixY1mp8sPdTLrWKxtpOUC6//t3pEWYAGkcLKn
cXr5pTEqJR8lJAyHu+8gdfFiXzBfi60SbsvsD2j7tusfTdkj4/GX1RjeKaH12NTt
Fyim6fTmBqBRc2A1V7c+Ybp+yuO1o3tDzOAkBc+zfLfb2bX5ikXGr6RJjvJs1IGN
f4jXnYoDBegZ7+FZuBlB7FFhBKeIWRbT0uTlP2q+uw6+fiUGWbvHkrcnHIf034an
cFJraHNr3l9i/jCyAB4bSB8a6FjKQP24W/IQYES2O9Nkbapfm6Z34Y60UQ0wY1QX
gcM7iX+HWWeGrW1ed/277dutTWl8//5flxGNOOqOVedAn49kmTOkcCsBmFk1XSkd
b895Ftcw29UI1daSxdWRnjbtyvzBzMTLk0LXFCnojhgx4x7lWtrRCkEOdrOIXA4A
3uc80wE3EqBwvaxJDE1AgSkQKpH5Q3w0z6A/iYjdaQ6D8y9gYCNMbHrsiJbKCFK6
YwH1eqRYc1xIui9ugz6REJI5dU2FSlAc26O/5CTx3i/sRqodjEUwHSqXt8T3Urtd
jy6XyAaOS+sU4muekuVn53V9G3AMs7ZHM+KogpcBT9Nck0Rss23xZDhn8kzUs/2C
iIF+lW+esUoGO/UU/kToiUeM/h8EULCQdWxWt5Zjyp9xVOk/olXbVak3qCLoQI6q
t3l5WX61YMJhHsX/0RSjBMIQ2sTrET4WwCXKb7jrCtWwKNpKazzuAowlVDgQGKor
v67VrNgGrLIynQigAzTvcXJd0qOvhJoovVmLkE13hR3jKMfLDzHHL380Y3OlAkbD
kQickl+lqrtyA8zepTtBJmxxnbuj8B9ywelinwKGNYYcP+ZgN/f6Rc6PQbFEOsCl
IfppQbMDX+uLv6QD5pgFfpIm3ylOBhSy+NfGHgxkmbIGZzMvjSe4/eXw5EFqs6v4
PSNACgZY388rr1FfPwb+/9aIyNdqWrks6pn07zDjAcgad7SPtIK7Pf0KsCCrqJ2x
XmnJlqSewGOsCka/6O1pipWYV/oOY1/TcAx5rJKXW/3Ij/ux2hNegFcIp0tuyVJR
3LKQd/5sB+QYw8eMwFQTkKtJHdrmEynv/VcdAPSTQYilzUvx7drvzS3JgpYmMg9C
r4SBuRI2Cp6HI0WPgviRCfcMdm/zAQrrjGR7iVAxtS1AcDh+FLIqKOyFZybNp3Z0
GnPWBWmQLsGReg77niJKToypNkxjnCwYlr1vcLPtWRaS/60i2RqPkuDOCpeuoh6o
RSkhEw2qW5j6DP4a5fSvlIjdkVLB4hxkFATz3MX6TBJqf7+pp8xqdZ6gFVuARdHI
Q01G1gOsIxJBlYMo7uU6uGfaZBfrlDRyyiLLHdXb/4SdsTNHgMlaZzoB6RXhx1WL
bWQ8zvQmkPBoxG9o8d4WAt0ZX1omGeMKmnMTrSFlWn95R8GUl+LYe8CTlA7tv9YG
Valo155OL59H13qDnX3+aHupYgmWf1sE89LKEQVjUY3a99rFj+iyXdnPBEhCiavd
X56JQy3UgB6xWj+1tJca5KA3RLcNJUrXorlERsHotyNOAsoF474XfE0rmG06Ri8K
zrW0gDsUhOy8AHsJdyPtyFSdSlG8oJUujpi5+0Z5iaR3CZOO7ub8C7pjOS5AmtOn
mAijdzC+ll+xZWQx+WBKhDHGwfzXI4/YEFbTfQ4cm/vnIklZGsn5J/dj84BxTbN+
pU48hUZg/KaTcbO47k7KrjVm30q3GerYw6xutSFDvA1fsCjMVk8iSWB8sHqOiBZp
6mqrodTiYl3red/jUTH3o5wr3KVL/SsUgZueGRgri9CGY1dw5HJCuTXZj+Z0B23C
Nn7MqSfiypWikM2Hk3387jTpmrFCvoouMnkT1a+SM6LYvXee8jKZ+ZlQGd/8tdqU
YLkCeHe8BgrGTVX+Kia6UmRyCsvRBonlHv3ixzYxKrsZIkgReFG+fI6MagUu2Z/c
4bD4mpm4lBG3eECJLSFv/i+U7QdBQWVtxkOdgI6pmp8Q93qS9ZP7OgLzFnwC9EUO
Mx8apVrut+ZxUgoWVMX3tXPxHGTlGrsClt7kuUpHjF89Pywun5r3JyWhF/jG9znU
l6p41T2TvC4gaiCm5pDHlmjC/Q+WzO7Pd1pPvNniP+7EcPwobWiil4it9kmfI24C
U47eU5KL4RScNKyY6JNu8riZ8qTKK486y5LbbDKEiJc2vI+vC9YCIfo17WNftlK7
IwFYBxMpRu1T9Yvl24VCtS/aZf1n+fJ4A0ZUBKAmUe9e5rsizxvvpy9YNWOqhHOv
D3h9Li8c9VRjc9eaiEabW7K53QncUAy1qaE7bcM9W3x8KEOgpqHNcuLqc7H9U0+6
XpaXgLhm3TO4/6sfgo6gaM1nFKu1DWCXXihsdcN9Mv/9h82u8lpK2k0r5QmX/k4h
yxnFMYfMaE3tx1N3uBNs411yoHjS+OY5bG27YOpZb5/zyF5T1gSJvcL/J9oqmlP+
AjnpKTAra/V9u9pQ/lPZi7w/8rmli0JOiU7RxIT9EK3TlkwNj/mOPA7Zc3p4qGe1
alCZdyUwormzSBcvyHdiIvGOtL+xOI0H9ydyViS8Oknj94dSXPNuRCcBh+uycRgr
kFY2UqHTl7rxiO4QoopMDqmRC4tgsIrK5WUYzXEfGUAsbcOTUX63njGxSrn8AuOd
Mg3IwNXKDKmJg+MclH6vLmtDF3ANSngFKHoPvQO547fnGbP09fAzsNrieUJ3lUaD
XoIiGC1Bhs+T4WUT464L0lA8lJU6aI0zOfSiIPzWaRyTMsjFVEUbl2ZHbCkqbvDb
tlG4dJxwG/Jmm+I2L1PILxLnQOyL4Jt1b3e5OI/AxQyh6K0+bgQCm5Y/K/rx2qJ5
ln1CF3hSorJ1yJ7K5iQ413pSiHCNl0AXoin11HNjidtiiU4WsKuF+hC3QYLyT2LV
eNZ7ka81xCw2lVH9ssjGP6XuWEgpCDq9jAECI8reOyIliNwGaPjSO0lLOt+EaXrU
oKVt3F4V+djjLgr66d1F5v6teIHjEyCyUnrIlLsANKKEu3k10XtvAcya5by7QniN
dqfyyUhsgFsC7cEJmLKjOJMKZ91GKzbmhcRb3j1Mj+mVhKUeEz4HlwvX/qGfcX7l
gyVPUax/JMONLyYqCeemJGL+9ynuYQi+OLy6KWr8fx2h2c4FsMtBleC6Q9ByiY2P
TgZUzE4Zevj82nuewKp1NF3j9fumVd9L23jReaSvUYLGVbK+tX4i3YtS8vO26p8V
a9Il3K0mmB/A9rcWCR7MbaHmo3p+gZ86XBLGVL7iPPLZBoOq7ExPvI7fdwiNaEkC
f2s8Ndzqp1TmB/Mf15kWtkzZYcuHiQXXOsNzBpBEanWI0uXXU8zl1KcQktnQeIzR
+2NbW4mYU/KDvSMf+v5JDqyOwVM2MkGxk55RWbAfHE7qXDOt7jokTwpLDPfwoJKz
EIUWOaeX43/A4qXDUFPYqZTqR+DhhPrrCdinFI8b1FD7/38CF2HIYZxukTd0Ri/D
iyjvLJ2G3l54C3zW+91c4bhRmpGjz3qfK0Cwnsrxrgq3RScwn5BSiNG9NusLV8ni
gA/Pg/sVCOxDTvKoMKPYkgu2MQpdKGL5yYkbpPjM3u1twF4RtNZOjGskqybQLwTH
LEckdvm5hWKzUNRvuinSxlICDrG86yHs1sC6pPzqOELMUAROiNl663ZZYFHlEuxM
5QT015ylv8KbuyBYQo/Z3VSHSTVFIzlRusWRIlPHxdwFPwLetCrOPi8njZHN4Eg+
hBxu734Ln1pV9A8pB4XaCz9VAFv3mzOz8fuwEtc0BrMNbFbQRM2Xz5G6tuSIclhV
P8O3fu0BWVUdw0wZW0ylvQ2pIETjQVEmr92CU4szq6IKANiYb0kSI568KwwikyRn
g8myz2c8DnRd/BtPdWr0MgoztiiV8yPaRZt1z8d9DVvhAK6xPhgzMQ3g5QHHeYBP
GUD8fgFhJaO987VFy3rMneJqN7jv3YD/XfyB1LUJcj/3A7ZYe1SmSQpEwsj9vYzm
D/7MqMCA9st6GEFvF7wYm3V2KuCnaZRSLiwzp6FLEVU9n2KK5CyvZEFfsVz684kP
jhfCjWUtxKqS6frqc2rkfzKEWTfz62NmFNdtCI+EFG9mrzLGPKNaChJ8KXRzaMT3
vknO/hWo7c8joA6ucK24/Gw4N0DDzUgycGAbjXu0oJY6CG8ZmmkyX1KInwgKInWC
A3fUoq43sVyZIGAd1j+GF7eJxagG9SQw9MoXBgXgaG0bVVdr0Zf3Y9/gDNJkgRI3
e/u+3B2imoajdC5hYddE49zIurbcuz4CVNs92Eg+NxFkSXgxVxplzJx7khaHPD4I
sXxQXLh1swhOwSlfRaKvhaXNJireS4giaggFVjcCuEi0Cb/D95UvehX74UAKt90E
SbYORmrNXsgBRYJ7ezCngpLbPaCfHo/n3EZmGDQmQK7JvpCeXo69H2U4O/ghado0
89EHjUTFsSF9fvTNHfLAPsBLcRyCTCDzv+EG+6XAiJL3Z8+chbMxlMK50EVF3cmq
/7RZl1CqogY3KiwTogNVVjDNW0rXEglB2ZtKb3oBmEIj5197bWrMD6ZX4fc0ZqNz
VZY4qcSRL21aHE14u9wUh9PPBLH/TBahNDmEkGUrVR67XvU6DV/mTVqIObMwxE2h
pO53CF1anIIAPekk7DfA5Ivf8nvY6Fua4YYMgetteSYsh4g6YryULNOcYTJMNMfX
J1SA4yYrCfixX3OE2Kek9rtl/JnswoUUh2eqnRtjXoTEbN24hxg3c1xK5w1ovjNx
Bcje5UvmfWijyul4lfIeTuDqbyD4m7y29fGuLQvK0nBNrsEhfZZ13lUMcJgJfMI/
O1Lxg7C416pF1gk793FrJAzKKQbL6CFavsMsaREuEQQ+tAs9QRcoVU4HQwuAFOTu
KR6YHJXPyjLr3yiqOGjM/DZHXBlXoosYRcMe6HKomog2tVust3HtCRlHYHbPj6P/
pnDPZBb40Fe9j5qu2bmd2xIcC44Z1gr2iP96UjVWrsZbXf2gEJuBgBOVsUmrXHRd
ZAHkggm/rlVKWsw7LSvT44iU/ewCPhTXPwcP1bef6mmjMg5Y/1rr1DIdfaQkdV0B
hLM8RCEncF5iZZ7xGNf5DwPwGaOrSWvUGzKUOQKZmxlLnNTTbHEZ61s0Giz2LqlY
Lkt6e7Wr4t/4FGwfLeCV7W616F6/qEM4WM7VwDSWDIDRjn9BLCGsL8k+4CXbrqVO
pBWJOHiacHqW0v3FWICCks0A3V3NRP+S88GnB3+OvDalBl8m5xaPhsUFvkbuY38B
E2R+Y9pvdwlCWVLreepOueXpvfiuSMl6bt800l7nsFrYqG9GCWyDUOX2ufFAugsn
85WkFfXRuIeRrnJ8wNP8UVgugbmY7DKVYjcFUNhEYacdxjARIFEie5nxOkwImCk+
FcmC8h6MzpRGcpEGEDm0PK50CngoPIw6+Kn4qEjLtSDpOHwicFZoVtczmcktHPw8
q5IKQsRdF0xOJ4/wY1YbqrhhAuDl9GpTIaiiXoh/opwB+Qx9rX9o6E3CsWLUtMPk
auxifbyPEpdgxoVP+41LkPRJG1VwG33SxCqr9xEmiUE98IDi00ESctG3xP9n4sxC
gCdIubLBRlBmmblXARrEivQhmQMEyvnskketOgCp1jion+9dlSf5rYx5mZHDmlfq
oSL29ZRX3O0+ps29/jXj218T5cl4RVDwAhsnlm1sYA692C92rginHczYLu/oq4WB

--pragma protect end_data_block
--pragma protect digest_block
LNMTofFDwknPqi1lNBaWvvch9eg=
--pragma protect end_digest_block
--pragma protect end_protected
