-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Bl7Rq/S6IBlYGfzaSdPl2txmFPnT2Aa/gwCU2dbtD3+o583R5nYW2Sfzij+kT+cb
W7S/EGkezxTwdH8SDZQXpo4MXMvSp57FY4YA2OCUyn4yFYlvi1iR9KR4c68j6Y63
7BLPzcpelz421GxsXEvqtWAC44Phy95h4WKmB+t2X7Mlu2EOS+2R2Q==
--pragma protect end_key_block
--pragma protect digest_block
aVZU1A6cgrnJlmWYSO5zYA3AwPA=
--pragma protect end_digest_block
--pragma protect data_block
lxsiypXP/1Obd8Uc1/c5V/Xl/s3YlnSZESbHOdP9gTiH3dzNqZxLD8/vcODE6MG2
qeg3vmHV2Fm7LyUPAvzUuiyeWxCBm+hUgdQGyPgOOlqiguW8hKXXAtFxKSspghX8
enDbMj9K4vRsgkLQzpzp9In8uhUaMRy7EXd0/31S6MWLOEBW8nwwgjIEHwKzCv/e
ysPl3P2YoC0lyMAEO35urDlmY6urMiYGnwxYjidxv/85qlRRjz96OSnaOfHgvRfq
bWTpPCky5DT8ePQrDIPARDctf6kEQYsuMWIzuERMiscga/LbA7QdUcWKo+vX0uSm
V13cVMYnvRW/qeL3NnHJ+z5QZSDEOEy9kfJT3IaF60iJeN87tDxqXmZK16jFbNg7
NPavfs6gUBAX9UxvGTE3IMkiRk1OQ/C5MsUWcroxgSxj7lh3Xlj2Rf0oOq8C/SKR
Rq5pcvgTeBcR6kfqbVrZAC0zm7HXvGHkARhjhx+weW91bxjPTk/FAHS/d62tzOtS
r01HrWmfhMAaMPIVl6rd2A5YdDTnFqOkm93Ty4xiQhU0Q41Bq7zfG+Dm28LKMzeL
oztyE1WrwNpPoSTUcDwihmPoIId74HNC3AdsmrKnqFli/UIY+m46bYxECEcrKtD4
5CO5krBEym9RiliRW85v3AJXWH9uQ6NcmQMs1JwKMJ4eCe8E+kph8LKC704DAG4x
b9qW7Xj7LyIYb785bUim1fx6G0YgbAU31e2kcqbHTFrJeMR4isRoPolR1Nn9XgO9
XyVBlCBEsLkp3Wa9vvOkLYNyjIOXMEBUToOdrsGt1jxQSlTd059Zi8Z1hXD/qLeI
v5+HReOtmQn2kmnM2DdER9a/FWJWuoOgWJVf+ID54dmZlZUEWs5s7ATuvVQKtzWq
4T3PCl1j8i0x7b/swuHyqmdZylFOPo0AdjueZgjeMIGfa4RQgzKL9SOx9lN8fhoW
oyKhQ8ChIoFntDmIwMq35M1p9qy1sXn7o07eCTApZzSMb0wxrZx0kq3SD7e3oW1g
jDVSvVdM1qU8zJE5GdlRe2hdTmRGBnosbp54F4w7km0v6zxz/XmztxgOVMW41vRp
i9HlV18isYYnp9khe7ANI+2rs15lYwbaFc8Haw6AwA9KQLZr8Kedg6mnToY4HRLt
0ornG+EO3RopSnBSR4pXL81QjWnXOGcCLtusp1fFrTdZO6UvaV8OwFSFBK917gBA
5dEMn+3hCKsvoFCSz/oB2EUiL5cspPvtcCflDWTFjWR3BaPVbqvhrnK95ufpw2Q9
V0kFOsT3bhQLr7BcgDLPd7mvJf1I35L2AhW3dlgMtWgTLo/xF0XFcVpGzpR8QL53
gbd3NP4lDvcd+vKCHL+TVqALSnC3n/eaKOvPL/nRsAX7pM/wax0aNV0dco9JilTZ
MZqGEvH+Obc/6W06fVtiCB1vhiL4lheu9dKqe+fzGYVa2aeS8K4DqSkzgb9cCB7u
2Dx7J12YQo5+97iNRr1Gn4Y6ATBIw/qJnriLWeGchFRyhbTe+F9hN0TLfDAig6WQ
nx3zzJArPrfg3cHv+20C3vlgp/KXvUdYYK5r+waheLdhMU0KDi2snUqTtMAAIBXN
B7KwMS9HQtQIIXeYyCJb/F5I/0WvdnAzzRUEy/2PTPvlH5QQvzIM5NTzPk36TWyI
rb7pM6pMpm9TcxYohnb2uA==
--pragma protect end_data_block
--pragma protect digest_block
NTuc4jSDi0Era7HtynEz4KLD7es=
--pragma protect end_digest_block
--pragma protect end_protected
