-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Hc4j53QQ2sn0WuqcIGitOWmOe4bzhgAJ7pLCB1+SzTy7p4TnMQJcJqmcsz14nldl
a4F5QwhbifolriIoYW9Pm9E3DNL+j5oOxdtwWhZOgmr5ef9NUmxzrKgOy1v9Favq
llTpduSXsHjEJhFYvBe0GiN9Z1VA7ouidkqJf7yXw/Q=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7574)

`protect DATA_BLOCK
H6VY/GwDgI2O2m5yWntmVvh/3U6NjHKJXuteAgtprWa6VYXtnOADLNkN+5u1JHsy
KnVj3/9Ew0pjZx5AbfHxyTVlP/TO4yM+a3swzrp5Q4pP/eQRqsZqIeUIuKIqHo4u
P9RD0BA53GXRX5wjR53uTwYRPfVZZCejho4bg8wq1/6K+ZQcsYA5MUgabGdH74Pl
lCs5Jufw54uxHrTrJLP1+Qte4TqRUYObg2UixCAY0ox+ol3djgT7FVimZxqto7Zf
EDcznVL9Hrjm4mGENcpo5e0OcXecTIsoc1c+KueRtR43XJibCRNdY6ZObachyJjH
CEGN85lz0kvmh5OMTVul7V5/1y4yO7bN9zF9bfQiUNoce7bKuYKCSo3BGjF23h0Z
Ypn+7VuSHxjF61n6o+uv3pF8SNPSZYSRgA6kr7Z+NI7EcL5flNq6AIJO/j6CeVzp
aPcR+Aid0RpUnLoaBvH9Loc+x7bHysXblpQhj2ZbzI7BKXI352ZRsdTnVTuR35zG
AsHcGEQU1JUywPUu753uZKQK5hR7qyB8yF7YQvc6mHQ9s28OSGdJEJKFhSktNaU0
+eTu8/OH8H63WJD7mJaxWNq5rGNLiGErius7QCSayMYhMyiX/a4Ti8rh7c0y3O2y
dkFDdEBJM7OuMm8E/uSJkpVE1tSQHHkjpD0ytWj+Oh1TOwKqXwl9V12C8zWPhiR8
57KE1e3jXNbnkKsuSecGsY4DWod/apK+Y6TEEqnxRXQBRsLhxB4FdgDWpmUEtMc9
8+Q6gzqFj1YF/v20KX/eqKiR/6GQC//6ynL2pnZmpH67eYSJ8r7TEaEFXkkfyq1h
4F2EomMT3q1ALWmEsEJ2WR/OgHAGTXNdi+FLDNmMVpuKTw/SosJDx+CL65WyPgj9
nb2bYoi0EM2qiPdj3Av1AMqcS+eYvUoo7StCzIwuKra7QH9Fbmw1d9aOUm2YuIpo
GpYChNEa7mLk3J/T9dObbgiaNGhOBzycQgW1E1PhmqNeNN3Ubj9P2f9cVUa8uExV
Rf+b7TV/DouuEcSrWONXVwDrWfuUIYwSgWb5isrWqZH/Q11LWLaMTRS0qKR4sOxK
Swn1R2Jv2GGc+2MSOz4/aOnhcgW1bUWWnsnyIQaYzfUJnly5EmlKWuGhOZ3Jf6Rl
Q6XOcM4puH9b1+JWvKZHVWxvoorQ7cASBvxk/i3ySBDtDkv9MRqjFrBOhQ5HfpYf
VSe/hGCvz7/Y2wTX7eTbivYdNHra+XzO5SaxivGOX6Eb5qBUPopsZZMDMiqKRP08
gEO8fsqh3btJ6Ql6M1SMWBLkbdQ4CQ9cJsGqhcv1EzBF89H7ithdwiSvwUL3nZgz
0Xz9xgmHuWS6yVq9nbMgd2TQYp8C97QPdriVifwTgFsZJAEIb9HOOcmIHlHa34FN
9BdX7qT8vFFxszVh+sKUxNb2twNrgXksTca9zRAcSQLY31SrT/RyV2c/X+PPxiyp
XkFxy0mdbmemlglLEKJB3512/7NbfrIqn+vVHXB/34x4XqlBnmchnbe/nrg8OnBP
DLgUIiP2pvpIgxDpSV7WZcRoucInKNxC5zUz1Pm8ZtC6KH7kkOBflA/DO6/xd514
4YKOoK0n0oIp9LeS49ZQeIduDtoSzPqq846r11nyyIz411V99jyI2+1BHWohbflT
Eu2FAc7tmSi83IMKkyyTyuA7sdskELpN8fFbAPCbsYMovwmYimgg/jZ6dtDU5V2i
Fu8AgMu+MbiG3FQpp4PMA2IKqFb92/+zZAiIyP8l/s34dpvpIUK3zVdS9Astt9AK
ejCBAHLeshCZsuitmll6Vot2hnnNVMNxzr4645F1lojihxKQy4Lx6+KibjYqG0g4
Uaq0/K/ilwLKxhDyVW5nYt0Cg9OEZSQvDsjKPQp+7ANDXBedlbGb4yIOQBjBkiG2
fhSluGFY//Dv5PypX3dEnAC4hY73R5jBzu4ez83OU6PUXhxxK1BQXhjKpOLOkCGH
k0SmJB+n1+5s3AFiEI6fEnLxd4q1WknohFcWSf+ePNpHEdrmAJXV8wQ2nDIIQuet
6ntsrQR8Nm2nE7bnrOwHDE34Tx2phXMuHzLg3+TMpbxsVmFI8gtaw9iVALXH6aw3
7DZC8N/s1tSWbaCjELSjD6k5ABIAnsUJPE30WVbpCRQAzwIjOAVy61cqAj8FaRyL
f8Q8FIYE3KUw/OIOH0pS0AvLxAz7aHsJubNfd+iqOboRM+pXlT+O8gCFmoiPpQDs
76MoKSfzMJPP84pMSCg3uZXzSHfA0+vPiFKaZ70YHdRdoFEHBoQNX4TtmBFK0+pF
Abp6MvuzckL67vsBo6PSLTEWLtQSZA+Aodi3xA6/XBdyQs/i6egHOINcMVGBZLi8
u9p+v6TphoNTFrL4uPhpR4PzmLSl7u4z/yUG1Z/yuNFgqJYhV3cJW1T9yJjyPCWu
m+/zun/ndYNk0WK+ulfwEsxVQ0X1TKzz7XAM87IB8wNur6kbQ5/nLm9ojhY3tKm6
nuQH8qvn9HJz+vlHBhYyypOh5GkucDtLK+o4hX/HXax1SIlAMVqgmq1fv5ZvJucc
EOrJ/H0IgU9hJDRr34CkhHOFko8wcvgUi/lTfr3stzcRsZ+JSRNbbFPOvQ2FZUKz
BZbsRYgJENs7ZqKypnSzfQWxejqOiT+yv9jq7JNHVuuGnNkTGrk0ZWSV4kyrmlOw
yu1kUxKeGqH1DNdaV4KJhVdLvpw6nDVDOAXoSYE47hGxfs1Ea6F0t7GHwwkjLmMU
FHigeD9HfORfnlkvF4nFlAFBfnwqmchk4IgJVevrxgxLsZcUPrYLUsuGz1DWBqlK
EC/NDdm9VKLy619Fj8z7S6HDIaAliMkFk5fRS2dS8aM5HBJH859JxVB3FI2Wivpj
njdVcbw25NVZxv5a3oPIveJWttWsXs2lWJC8LEBetIsYCsTQY3MdElh9uyVDhJeu
RrF8kqtAga8gHj8WwlF8DCaXOJhDMcHFqNZoKAdQfMxbp3ICsRffHfayGPkCFNyu
5ya0VkCTA2+m6x4xEnqH04L8AewDabHG7yR1WKTG/v13+JHJtr05VCakeGcqUHmq
I21ENP7sm2CFDupZ1YhG45gpRmq1udZ9GqaDmMrHbGwgVt3mKznjIj/OgyJHiAaE
RzLLBjPBA+ygDGkHy6z/1Zwr0+6EnT0NcQ1g/pbLf9X3I38p5s7RnycnslHUQp85
qjynUXmg15Wc9UyQ+f90fCVcY2N28JHSz5jTBRUpqxCZXSgkA9Yfy3Aq9GBXK3YL
BxfUz4vUb2ZOOMqH5dwpYLJLixt3OjT+lAnUc9iIe6BkWy4klPva+t5CmjyVgeia
KlXU0OX3/j2SWLI9JHQC1gk8VCztfBGMWNLSXyPVxd7UESNoT8mrFxFiEUzrnh4Y
Ue4f8+lxidwTDXppMO52nxEoKc/zDX+b5rOCaNLIxBaAEuY35RdRKTvjjRODrc7D
nTkWHHI/UNaqyYmRqnCwNna/f8qnjOZSvGBG/BVZOcMascAncRVRKzYIH77sP5nT
CCAlHxR4eQYR5QA8u6e2+yOZvSdypwWr67SOgYuMZKETrYtgG6+0L+3XjrOzeQew
VewNUhaE0zXoPB+vHVObha7+K60SyJ/Zz9i81MwxMcIix4+aSrTgKA9LpDga6EcZ
nSj9sg5WxL/0jg0hGti9xqaYikH52TUJ4iZtnTC1kxzDC3CBaq8CE9UQN3xStwMV
51+W+PvLdx+DsIfEOoJGhgylEa7ZIwujCBg2XlCyl3eN3yRTgSye5/6XA/WYWSu9
vyzK8J8j4Maz5zK7x1sfUgdRzCvwUZTG8ThSpoGsPShzEeA6+7iKWVTzdK93gBWU
sDVjwCwq/4xsvuP+gqDCzw/SRF0bIIWTr6bFJX68zf05g6hTZ4mukmTqsMUGVoV3
Rq71GiZVc57YQ/0xBuGM1qaoL1Mv2hfHcHkWKamDCkkiEHrJYKB8BurMPUrz+qIC
wIz3Njh+YHt2l8HlN1f3z3o+OgnAGfXTIRCgLfgab701vW2aTEURKlv1KVrgG/MA
UgwJjibiY//Y81GYh8EwuWwcqSclwBVZyUBdjdGZn1u25gPzQ3ydIXqUBxt08TrK
m1zMknPExryjV2ewl7mENjL7vYouFyCMqy7htpiAlnwXZCz6HCt7gI9MWQ7IhDwi
npBDDFe7wjFKKUNTR7anCKuvFHz/fTOFaAr7d+pQcy5Yu7k1Hzfy7teYr8hqk5lw
/9/nrSitDJo8ZIQsGig+tkTfTAasRZitScdYhcWVOPAPIzegpd0jx7GYh8bKhIKA
e0Y0QSDWAAsdz6HEMrApJ8cqnQJRI0OyfUHRizcuQ7Qk79WOXqDce2DvDdaj/xtZ
KfafVpBhCnSsIdiyBB8Ob3nUatvQUAICL0HPwDLTTID506tmrPqBOC/+8NH2wXWZ
uKZTOnOAvoIXyJWO/XYDrf2lh6h9OPaq+2wPSMTEHOo4XS2AWYYTmbQxmKnRU36I
nwI4/rgddX5+UHhH+LJl3f+NmOR0XfDXXDl+kNz0fuTvW9wiV+wfXYqErQ5HC1qA
Ot/zNihn5YB8QPp0GnzDOpzMTmQG41R3hlDvb6wZ9KPspz2Vt8+aTUyl+c2TG7Fs
+/XHkL7hWxdcuKts1guyBbnleQhzSq8LBzXftHrkpMP143bU6tAcoKaw6zVLe6mI
c2Iiz0qm09aqdKYt73gRwP3emPFmdK/iIbt4NK5O+Iy2ZoB1IQLfsrMsesExTqD5
f0ugZeDHmbtaWcI8a+lIX1oYa3S15Ajf5KSwavZ5QMguifUxw8lvA4tiVoa/ZnVI
UUewFcCwUD7Og4y58fOrD2lECnptYNUU4/wVHPOSZl+KH5+pj03iY3QGCKOIseYb
ePJjyEDl0AcTQ+kHfoqmO5fXQJ/pmX9T3r8ebqJGdGAqS3MHfFCZACVM/XpNIrZ9
vlPjjPESYWK/WTGEJZ/XqU+p1VVQ+o1f4iDZ04dTghRosFtQCvIj8PnQ3Tb8q5L8
CdI9xKYCf24n/acZDEl9yDWU7OxFmrUZWB6qxQEcAe2rvrmqXTrjhSwLJVoifUKa
iGQwva9r4f7cFgvsJz51i3eCM5X60XFUTSueb26JnI0zWPMBt7S5sumn9u1ITe6f
rxb/FiMsYw/l18/kJaj3p4Q8+73wV6krxvXupKVi97gGpspFI2BKhl+N8iHlIROn
1RAe8RhlpzCspO0zzyeGMimKRpRU1YH6y1uUsiEzGOBTIKQRJndYpG6oai044djh
sSkXCc6U1ffxC/QwmIVTotIdj1ulEEKIGBpcNzYxEPJFbl54QZOno34lOUjX9QW8
1A852oXbFxyqTvNgF4iMLTB0wSD5Tlhga6AzFVGiOyr3sVtUT+rU74LuJK0m1EDg
hPwfxzQ+Lgt6N07LVEPXVlObu0YRxngfLdAOvj4XcrIKJd7S2tL5iqJJ36IPYx8U
WvFSTXkvbom5jqVARVyPTnBkZcEKlNxtodSD8wSZxF7xE/fUqqXpFhTr6kg/vz3p
tYSJCvNCL+OyeTXSSNKXe1Yb84VtJK6y29CI8CPV4RgqhAxB6EV9KuUwOQPXjZLu
Cy/8VkPju8zzMKBOurEKGo4mjWohWeYwiB7GqJtERxvfat4uAb+HAOFAgJqZ0Rhf
mBVLg61sLxK53XzUP+QYAG9Mm1hGUmHmx2avqFtipRfBB1YCFVT7acqBAOfjLkgT
L8XkczrGGjnmJ2qTCV2H1ayXWbwGiQqXuadj5gUZMPhd6bli1bFEDgpUs4X+NYIq
iW6p5W5Qg1UJ/610xo878D/z5bfwgCIkYUSxZ4qVueV7wQnhrjgJmVEY5R/L9kdL
Xyyb5bFCCl9htkd1jfHyKIx7kQua5a66d2RBl+unzlQF3rSHiNkCFx0fPFfoWVtW
G5Wtn7YZygJmtBEHVjN1740yQb5QUfkofHCV+Y2ekUwqbfgHyTwk2p6hAGVw/XwI
2xqGdp9CkR6NFYOXX8yARatwhTVni6hRFH+sVV4ytpRWsV4Pdbdbu4K+YUCUX6tM
QF995TaOw+APCayg5PqrkyBPg9RYDDmN8Cw0GAx6lLXL2sMdeQjM/pYhuWTeZjvt
qWcFwIQFl9AcyfUz65c8PCcLXLKuI+qS8n01uTYisCYLSRDJBRZp0lbMtqZ8eAgB
6i6c0Ja7TyZJxzzyrHcEp58NpziieBBerQlMgWolN/5nU+B6BucCL1ZNrUHis+Zs
PTIuXnCdAwF1qp5Zy+Pk0qAZn1zeMbXtMk5o9C/NqfQzFHkL/X9XLuZWEKyKpEjq
YmB/FwXFB+FaY1Y8q2M4UZ/15zLjsYbWewmMKUafPmuVKGXeymxtdytxbXqJtngc
m9u5GjgkLzT56DMt4kBHbynHKsDEJ5gRXGjc8+ZQoe9MmyYfv6vjrQPi1d7MuJ2Y
K4Oo4nHTYFgtRoAlPkMgiiSt7QpyvKrafzw63CmAXoJ0X3q9tZrJZ8yIDTsblmlD
5guYreAAT1O+FA7NaAKuWZ77M7wO6reUN31zBzaAW2r9xrRgGqZj8CCIYPyo7tY3
nTToDxKSnev2BYo+lAttmOW8PCJsFvg7WHqBFgAhk6xD++KmmiQ/8xOMFQbBj7EX
q5s7YcQE/d9NTvspeoyWXqrHaV+LhswCJ/qm4PlwsoDsW1aSlvwRzD9SfLSt1/E3
GFTEgZyLItQFpTK/vnswrC/wiZDrCZxd/SkOHEFASQx0HEW2I6H29Syn2986uew3
9VHAVKLV6sr87O407q1NTmKFEHoGyet7t4JDSLlY//wIv7M72WiF9NN/lM7M190o
9gcWwCywnBktY3vF3e9eYtiSJuIMCFQOeCjaLvbIo3eAWOWrkZrcAUe8/19tBKJ9
n1pjBGhIYUuDkst3a9uPSgDP166SVeQNybe6hFvxjiLkvoIcn1+meGTXjFw7YJB9
74lm0NNL+l34JAtz+neeyB3zY2lRdHpZliEPu2RCrSLkpZsUO50u/oK+U5PVv2mP
mw/nXpIMUIy6VuHQny5MJtxoc8pX9L2CI5pj9HgHyo2avaeoEHC32qEF9jBmYuyb
aNelI0XjVRs9K+QrcLqWXFacKYzvDPfgHBSCwlOFUMD1LmcmdY3NYAnVN91B0fAg
jSAVjK4xXIN4tVuqn15B5Gzrv0azjaUC5dDbzBP0tF83v6hsciEkYfB3NfJKkT6w
yDU+NgtgNAR2ODnGKU0ECSLy8+csFnGmNc+/VXaaNepOeAmk7XSkKlFVhq8nHE+f
jIdT6VLn99WvjauZ1DLHukPTyqBwQw/8zoVcmKTRL6fnvQceMicKvhZCjZ0YXLqw
SExigrRKP5LElrQuLKN5akjUwM6zqbnQO/VpqkdhpD3D2nW8GCGPUpd7JFgbQgt3
mJ7neTL+dq117JDdYe8xyjHhBn9CZuVCx5sSNscTVVW4aOa0nykUS2+O1e5glgpF
9H3mgD58JDFpN+w2QBsBc1ohfsIotFY8edr7+0anwADOQ38wmR4J6efGMuRhwhLB
7u6U+3bfLjWoMeflrfKSy2KTm2MGPHolCcLXRnLrkDS/RjOiGWOJ8MbuQYfnrpFh
O1BKxs84cNLlxGDkr54p7GYOPT9zgBXQHvPOKMA4NBY5bLlPJo/PNcmF2nXz5OgE
Qe4SSRFvo9vKNXKIa2ISg5s/N+nsmYIH13Zymj1jzOAac/2lH8pt7GZM2qzZfXBZ
iA5sDV/JcWdP2/r1h5MH8L5x6FW0wT5PueYpkDRsygRGjl7BzZ0uv+hW2df8OAg9
RfMmFrTUhpjQ/oGkpHBvsoPM/vRYdHuW0oywcneH7PjdrqqXKnnp0KEkGErZim9r
adxegZk8ms6mjjajrPsFfFmvXzFi3AiRM+MdDRgGWQlIr8MFujAeQYtTrNlW6OD+
T3JFyeQ+D5Gy/NJOV4M53WTHCQ6iiG0Fx8qNPzc9x8yXWdQolkdnxNVq1qhsrY1o
KEV4kwg571UEp/iReiD0DxBQPOTzXXFn5j5ij/StARsiw+0NPB9TsAneZgMVky2f
s3bCI/DvsgLmMw3mloNw2ZLoJoLI0+nhFkOAavwfZDsye2xDaNTpVZ5FMFXB3iiG
waAZxRS8gZfQEJF7TsPk9fSgOP1PiKZ9m/HGmMdq5KRiH1h8duzyo+vbnXx6YOvc
E0mo2AfA5Vu5EntLWqDZOwQbcC96p5o/aee/1fFsJ+wPJf5e3QM9jwbAzf9XtP/J
jjnCuGOVN1Jokewb307wvlIsjVgZoVBPrfXNjlRl53VVtj6njmk7L/JEH5a2MVxj
inrtqGH4mGFVaB/da+SWhhNO2aXDrhqJaNW/5zzEjyYRds8bnAv+dd7ElXWkYd0w
ZVzwFVF+UTR9f7/UI4Xf8rDXvuzPaLDYwTAgfxIUOUXSvrLEqHRqF/giMeIhytDH
/xfvEuf/iEDXginHoPNeIV4rGZtbF2A+hsQDDW9y6ZH0w6C9n5nay36HRLCQnDv/
vL9BFpUrbt/WDevjTSH4wRQQHlx6RhUVE6Frb4hyVqI1auPKIEO0H9aoYgOSWmJ2
/aZDVDc2S3orik3LWRlorIXj8ACok9LJbMdqDNgERk2oto7eI4AntoDpB/CByrvk
ser03eGgwHt04w5Z68JsKhh74s+L+nXXjb/NVVxAqwVikM13A07fDw/FmflO9I7U
c+TrwxCAywUKtRMAbtYBEyeGNbV3R3Bm6GdIQQeB+z/CGvWUHCUgXQ9anWT0fpbh
lA4nQ2StC+2T1krsFAsmMo1jmtjrShxZH/wha/4SjxPFCr2gm8PZy0mSTBooVPZG
ZtsXqUZ+B5XbA9trs1GlIRMVZvXXtQEL9BjOS/Os6ODH0EoZFrQmrwYYvh9KxoGg
Dby+evp/tvYchDUr/zUrLYqIVpRVEA+NBQ1iZRoscSeRVfpIJNtLu6izIPV4aWLS
FS5PNaQSqB8iSzemgUCXv99e2K7T7nY5nE+hZYpn3+uPliIpXg1E7qxWw8Z0zx3/
5L7TDnMog5+WUvR216WjeihgtQc3eLHW1SZFq2XfAtzecioRqZwyJ9osyaesXZqq
QW2akUuC1aT2ZzVEUw/38YxEDpJSJXPxl+bZJm1a8fb59HdwDkwNVIPhX/bvT1Ox
2KLoTJWym7E8NJOTdNjHJdFU+T5FcFfiDr44CKL1ArMW7IPt84/Fkwf9MHZ4pn85
sUl5iMi3oHj11+EqR5mP8WGWcTDq5jIcMhmJ0GZcHPji0UTf3fIeo5P9ODAzcRLp
9X5EQE5S4DCTp+IQBentQ2fldCYxX1m7SwPft0C8ybOfcVi3dPtnPbZosHH3HraF
7sNEtgcc+6kYJCPQsB6bdyaWOiJobRv/thlrCK+YYb2K4w7U/iKmSGcklA0PKpGO
Us/BArYCSM2rVXjm7/kFsqqmZxzNnrCIkjIb6lPkBD3a0ILyHdKo3HEmA4A+XDSp
2uJayBEMLtycDPbKTC6RWkBe0K+u3dF7EedJCEhqOv5lTYM4Ym0M+x6cno188hkW
dCRYBBusWMocXLqkqaDXGV8Zh0VWPUJgyUz80/eXzzfDqBCp+SqCAWIod1wF0+Ry
J+tqpJM/uMkPFb7R/kQ/o61uL5g0Chu2JEun/uwETOppAFZvdipf6vklJd/fqh7U
GCo8xOVfu8KG/tqyh1Qj6n8XEAUUMEPt1HVBbzgQrqDqT+BACvd+/1mob4G3GRaf
vZl9pc6Va9xmIna9N0XO7scMI6PoaaOCX/DCTUUdMi+fSI80r0gprVQuMBkOIbBS
RCPs1gJJFm1WQYk3qn2jWPOng1P/lhsC4jAKo58vu5W1bQkSRVlRugfSuoRU929s
XqCpv2oP17C3nnHlE777n5XmOl4/ydoCX4FUZPckCstlLLXMfcTGzvbQguZ/FlaD
L2LFSVbRmSBKLgCgF00SUS3cVoxxxWR5hn8EyVnlKdp+ubY/RMsx0aLX+wnmAUu4
y1zLXofM/oTKR5a+oFhEvAD7FiWKE3ZBcNtyC4NDwvsZcbc+5cFv9fk2gRY/lh7L
qifgLgmarTPUA3SlRRsTrj3std3EnPj9bbklDfuj/Z4UNvFOZUfBDFgTAOqEq7E/
UeccuynpPGfoyHAz3UP9Mcy9kBTccL1n+sagLi3aLam59lNHOaB5RQKOosSboTZj
COUTAUxzQ1izVZUirmnlOA==
`protect END_PROTECTED