-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
K0ScUozbnf9Rv7sb4v7fygqZDMU1HbZrV5txpbdVnG+HIFhXJsQXWQHZfxS09yKI
9NeWuV5/2IHOnYK0H5oGEvbavBPf0q13opUGGa41OvaKzH0oDXq0Kb+QdHOmWIwR
t6Z+SQa7+m3eWU/pyLwYXLyF36vnA9xR1ItEh0/dfZFUtQI0R93RFQ==
--pragma protect end_key_block
--pragma protect digest_block
NOesvd/IdV40Gw+TOdeAdOjDYxc=
--pragma protect end_digest_block
--pragma protect data_block
++c3abkoEuezUEU9nJul6qyE9pJtFQudWUJg90okcsHbK07kqk5hAwcz7eLgJ9Pi
AQCgaRpc8oYMr8wvr1nbMfS9O3zmTraDdklZHvW7JYBa03u8kruWBwnmjfb45nuT
imFKkUQpQCgN/18+I8TLLbtwo+11/SxVw75S5RN62eIqfxnaBXsuuvnts/hTenD5
E47jSwb5J7pxq2apRhGS2e7eag4AoYAIXgGVXWBh72Fqi4E1mruUKFWrNDDfF86b
4T6YvHtL6J2wzqMemgSDr+4q8Q+HB76G1WTL8sV3akOrlnWpRuOALoaJPmJc9Rhp
1IWi+QNjOgvxwUBqCM77TupXDLYNbIHeiN2iy8omvoHbyAaGFub6wOULGyyMsY7I
HpZEtejsWjTWRqVOUvVaRgXK6syj2RlQl73DSptCLLFuAS/7mprcF9plCPhlYa9T
kUjvSkK0Se69AWm0khzakXMUfw6k3yGpXpByZdJGUxk/JZhnuYlvxXdmm1hxMbN5
d1oOYv8QjmmQeYZ8+pa4cyFh0hjSJmSPtpMCXiPz3n16HSILw1T0I71Ut+fpUhen
rAfCcBnupplbHzXsNa52y+a4wzB+XaRjtS4BcXCx3XuM74AZJwaRS1b4pOSqpoHz
siTiBW2kBhmBTiY3XOdZ0n+47y+g/gNh3vLUM3b0i1zrwUb8/CBAW6nFNS9iuxjH
IBueCe3QizwPvF30baSQ3vTQiUWDwaH/NyO2xGIo319ilmZxuYmgNwUlJhlZmcp5
SwW2+Xe6G1QA3sj3cGeYa+z/U91bzLj2Wbl2up4MkqNM+xbNM9PJaw/QbXwBwDGz
Kp68sBXisz8oCuIupeV/dgjVfuuSyML75pegTG5op0dY5GY9HI7euf2pJERxB+TJ
POjq3DUTNayG/+nFSyqMfRs8o99mqgwbdGA9hsU08kXvC625stptx4lfArKR+ilf
nUw6NfT6kCmalSd3I8UyK1NxX9w8JGbX9ZQXvSjrhQViBA8BCO/toI3NP+aVJd30
FcfNtjxCLCIu87bPvgESAVRBIGsGGsf6pyQAQSm2atdM7w8TkhmJnh0lIK38WVI8
FXwoGLZqmhSoPYRY/0lqpeG/bnpUursNpFZJuQ28m0MZUsd2yr4tpx3W3GHburjG
SX/E8V7+yd0QgnohO7eIBBMG/V38jmV7uXBN6RmL0VMnlM1SYrlPzwvl32CYAOPs
XFS4so7Z5BqSmFiDjwMKwiRewouLdHrT1Mdtv0ezi78vO85B0W+xY1FWWzqJkCWB
SBJKMy7USbCfNLQLjG4biOfEzsyRVhJqay4mMK4O3qYQhl2NEmV+hWDhuoJfxBF+
E68EXVRmc5XqbxGGYVW531joU7uw796BKFTnRSzYCuzQimFS/MTRGA/ch6XtrFud
tymlFF0rA/bOy5Povs+90cJMvmxbwv6q+PXxxOUfbd8+AKwioo8jxNfEkFhr1nz5
g8IaGUttexAWYpNxjGxNmer1Hi+S/S6tY5V59/awoyGrKRtiNT91bKSacy7oVj7Y
lP+ISljpGOy3QxcKGqkmNJfomakJOKU4lCgn8ybEAk3mdV9CstZMInFGIRmgUCHa
ySdh2cvUY8F/s81o5wysR97ZrW53qBBx3ad4szlwZm/1V6iLQzhL7Qvgzt6ApVq1
2cQacCSEfs6DxRv8LWyHWeMnq89nNVqwDyzTbf0D0vEteYlZtJrM8VoPX9hYncRv
DoVE9ZCMLLcDTthRn2oiixSmZnh+yi27AW19r8H/rKZxpBmRX1WaIEK3HvUkIiYh
sKqAlqEZEn3jQ30vrecOrkaFwHNW3c+uEUFwmWZlewCgJvoHh77iXvJRo56yF/pn
NCffG5T1mgnmNpRRUYr6OAiINLbZDdnNpua4X6If8elW8OadfkxMIttUxIP//O1y
nPHyYSd4tEDYQ9uXYcfY+IHiqTwcPMaWsYHRDRnBZdqtXKE8elyHDkZCoX4U4eqh
YUrDzwCcGGdRCn3uM+AHulsB6gyD80ZeBH/m2MhmsEtH2zoI425se2VbxUhsnbXo
YM9ymNCBu965xkC/495oN+eqTNu+PDB0llt3Ho8Fsffrs956LIfFtAu9ZNxqZHqr
bI+Of8vEPiEBryBACEH3YxW5QSGO+u6n45e6fgoluxCPGcIrX3kx6oYTPbAI5cDy
JX1iLGdkdJoIo0Bxc14n++t1kGzU78Epl3IRDlQruy7n4NtI3D6mg4oaWl6KmDQn
uXCx65ZTdT/H+2xUyj/qBGlM4BIFfs10V/uaw1mspiPIrRy6n52wSS5YGcKeVUiI
JGzFY6kBYAC3owxi5ASzJcgZiL0Bfqu41WJ/cScQoVyAv4FO3F8tyogwezj1I8uC
ErWMxgD6j/hI6gotvrOlhIFnPajTwAl0NxFUpR/nfzM2AGYxyWwEztY2oTICFpan
XwuFa+e/T5PgiwX/nHVA5VGY5CUyjuSFB4fbzZn+/krVZs1yG6zXOeRc/GcphCQt
6Z7OLALbYRbh3rkqf9rL6ZRgNfBoSa/4+WLVsPPv/J1rvruWOT3AIk9/t0XQoJSo
KBfNiR5PmRrFoaQsNCpxAtJBb9R9vJP1xxzyE98zFHTgtwhKY9Q/Wn74t9GH+Oxp
DtXk7RD5Ww4K265oEbBjlGefo7kAVY/6Rq5vRM9i62MCi6+0bKKslNitKKeN5nQd
VyZ0uaxF21CQdZBmSuF8wvcROKrx6JuAa1PFivDY/1rc/25nkzx39hTs4+4tb6KQ
0DKQa8hPrC0Z4GHPgmS1TrCILH5xjZom/WarfoVc2GVFxrdb98cgdmNFWdialXr3
yS4WEYME8TNC2hS2UkPxoN82CChRmFsBeMaleU9kH9NyAWQSdq8G3XsPnqZY+14a
Lx8DS1djEyZt/abgTTJVfjhx4XWTgPqNYAvUIXQ5OQytU+cchbdyrGcyyyPGAl8Q
TRGbo1EWSKH6/rBfcxVd7LV4eQ9ha5wy7GSxG0ul5zgvbuXOLoupfB5rYfmkYnDU
H2Jut+kgFxHJx+X94LFcgvUI+qqRhfCvUV8nzkxQ6FG7QhmgQUnVC1RHfVQpqZ0r
raQiaknhchtnZRh6zedvgX4ptFmDzaxmo6MmmrCkacQiksPnaQr5i6er8eCe5Vaa
S8sVh6ivfFUay8m1WG1WdjdudwYuHJc/e3vQR67mTpA6XF+R7yY+qM/IenqviYCo
RrlMfWdpe2ewbP+Zm17V8+xQPsDf42sWPViJhQvG7WHayhSW4CgbaKDb3yGMBpBF
hFazNuANz0CewQFibKc4fvdXhmH6tqzLVTnNV3wnCHrRjoE9IH4AwKs/Imo5m/fw
tJWovUc9yUCtFut8WCb9M8ueaES0GYq7IeMMSKOdt9ZRzcM9RxvbEf915TXCA+RO
3VO4GApar/gZAVh1xgbAtSToGHcMk82Q+6GSBz5xzS9wqem+Up9ABtCoPRZGGqSv
Q0HXPCkzeufnFeTwu9LW3XU8N1wicecz+2w6RmIHyFmXwzRe+2Faqevi0vMqZSqX
yRl7/TfbJUqjCwV58/xyUfecajdUmb2DVlo4VWWQNGUa86cVDNFcNQDIwfXzRCDy
mEYTsE9/lgNfEbyeINlUfNc7hkactjPaXESoEAGXkOCsshZqTfU/quy4HIyh7ZvM
PTAgHkffSfCs0OgNABDHCpGxnUoVb0VkcepzZ4aGDQ6MfeFCqwVWnyRQXkMtl0Zn
lFcPfG1t5LC/CHRnzbchOeYldcZIkzKF40wwJnwIQmbC4oGYYdzIRi7gsyy4M41V
EL39IRKQsb7/UCaIMOAfSWEwv/ALWbbOIsVfBmjzMOKJv14e22IDtvXvtYk9960L
7gcXQ74Vwa9XxbTT/td76FaJyCApKJeSWcQIJtySEyaLR4h8+UKrjzxZAKgeK8+v
/mwFGT98Qi4D6sfnjy754rjKuZUDelmRMA79yLYBnxXiPI+1RD97fhjKrX5+WPpS
9ZVBL52XKz/dMd1Jt2pYdgoFq0IWG1YzJXOUQ4aN3I/LE5VunFuRwg7v4/tfhV54
6vxOvMEqZVDnm0Npab/uyxGfGF+7qBO4Onif9liYyWOpgqUbunLPS9iGZPfLH1U/
bU1ByAW6zAKn55FF6WicVwfzCEQ8Np2irs3vWoVNZb6p0uPKrJ2ZdKp6NSNwiA35
m1mVaD/qnK27q7pvcmGqE6+fs/pSywxVy2nNKJUMxElwwG1W+RabVAG5/+0BNaCk
1k4sMkTWHKQIaJPKfYYxtjIrrSqVwPMLVHvftFJTRF1Ds5osybBKaaRYOI2m5ApV
9oZ1n8hZ7icqryfPcSSDHErWEu2f8Tmt29Qj3P9yNzidVFUZhnbzb9pfp13Pya2s
AYXJJv6i85eo2lHJQIXMqke63AxpRJ2nwjTS6WGIHgu98JK3LI/ShIadejOUdXCY
KT8iADvQKZBXP6uTSFI0hp1WcWeHbrW/loRobgIOhQVhVNL3WXe0PJ9rb1WdPjzp
xfF8HqMzUli/zoq2HNP5Q6ONoRn+2eBcKQzPdffZn/wXQeuRcOSQOqOcMZfo1sF5
uQw1Oy+4e6Fh7mNDEGkOuAjkhZISerkzTs0b3BtyPmHifbJ0j022ZtYDXTBQr9M7
cSrZvwwgNem1016l5HUwfdGIK4SiHHtBs8IWgYAWpfcMxtMgiBzT0of46FkXGtpB
7cIpmIbNxCP7AMAnXzrssbzx+dUAjL3MCU36FsjQq8ehRXXjhCF+oZ2Tg4devEv4
detq+KF0IL9/lubDArZzPFIfyXm+IrXagSn5N2qnkK4UPHrPmrIUbE5uv98FjdVj
JExE8EVJjrAQutR5hUpF3atPbeE7W/k/Tz+V7PoSEDLPiqPI21OEnftQtIWFNtZr
lk8C+0LYPM+Q0jLx18mmB+BA93fEa4o9Nh5rhF5ndWilPV01myM3AwjMX4zezA7V
21mzVWxx+R8xIcyu2KSTssk/FTRw643CapDr8s2HJMwyw72aVpFjAAKzZ4KMl+nq
TfWHZVmLPAZlSErP0vWrSAhUeE2wFIDN14CdMoPnjL3v8FEvow7imAsSWr4plo/6
L+BNaeL1Trf5/k5h0MPNcn8nwx0mJAxgg11omubvwEgFcUFGkBmECm5SHXkBmGCv
Bjf6ooMbR9+qFYhR4D/0EG2ptWJEsVbKNJPbelCScmRmx/p5RoshKsTWhojr3CyE
QneRr8rLcBRgjxnOVKdDJQ4w2jQYuuXmCKekyrJEJomYuuHRIXjdRXcJOL5kINv1
EAa8iAA7CkWpEgsrIBw5Mu5OQ+ib7aeUzweNxg80W6F6SlwXkXGfTxXC2aZshTjJ
1EfiGG3roAax3t+o5qdY5J+yin13HIU93cnXvHt+hyRGs7GkLJn/CHv8Vs9P/0BH
EQgIpNsoY8TRIPdPJMxJDjK/B9Tw0iK2+hexVjoSVIsm94+c7csrk34RR9XuYNx7
WGogsL2n+d4dgaI3ZaGVic2gvUamEeIm7yM0BzP6MaPuX+C1yGB6ohzEiuGEh0bk
hgBAl8OAqcceRrFJ54CDIpiak+C51w84VQCnuXadU0vYh5jFLpt+LpLKKVVupsl9
QIY5lQJrocaLIBLEHI0U4b6b+LSyqwPzIlp7aoJuCO7JO7rRDHTZNC4Rkm87G4t+
a4ZiPsp3ceKOA9xEXSjk1ei/k+Ne53Pwljk4SXypv10JytS1oC4Sqp0D8KfoSDQV
TE0YDBPWL/S6t8rsZXiuCsWZcejTV7fsJxBhoS1nk3J3fmhPpQ1hK0hTSbtyqLkp
IuQjJJLq7X9BP7cO9rDRgjbpiDEIBvfI4iWbNkY/r/yCilYoSaixEuHcCRJgnwWM
J7+QDVFtNvXf8mgSYsSErZmzIbOGPqIoRd8xMy6S2sRSUJjloxVa4iUSmJSBW2b5
yj5ujFrBeW25ThH8zZtv/MgDymkuoSx8N+egYr62e9Ds+6UolXoTeW7kGsN7GJQv
ov324gdUDGW7B5Ib/tUn65xhlQSt5mwRhL2dvDzz4GbDcEv0/uB5os8w7AqIEdSq
dHlcvE0qEEIN+MKPNinAzHvA28nHBd2x51pmKKqRqgNGBAMp9VDTC428C3nlUU57
seGv8xwEYpOGGY8cIoIL5Ajpdm906dIv+0Y+BnDWPrk8eDLWHQ2kLC0EJW8lP5G0
ytMwimgY85oevBxwYfZyCUNB1HPGptA3kgIR5HFVAg+1QvxdPh7pCvh488dNL34c
+sa0uOQpXl5pScZf1LV/NX98mn+Qh/x4oqOZW52sJ0PynN81SfrdAhLoFroFahF5
xwe43twcoMSAZhmPA4AJYcRR8AHHxcc7PxI472co6HpVGrsYtqkSMGxAZESEt+a0
k+sO0fODeqmkuZCA9+9JiGrTFQAgrn8iUAQbECLZUUZDZpiQi/GdQsf6/TP3kxAa
daaT9tislaJtcPxHMkcVluxX5USqQN6cTWhkHfcPQaMN77Uo92Th/On/GVWxFzDT
nNzdVxqujT2YK5nVy0pn9iUTgYJJa+AwgsuclkfU2y7GozS3DHyV8aEcd/bbNLUi
Kaj9YXbANVyo9i6dG9zCiyhu+Day6jE+0cdfZHdCNXtuIK4yiZ5dKcEZD7HraaSJ
MyuAOJDT6Dwcx9JdFFdne9rE639GEdDuAJcCEoxb6WbXLUgHoWZ6zXrtNtfi43a8
Kq5X+mOncZPI3HQSkXaY7MChZpiti5bpNHR/nT2mGX8hXHhfPYRkL0+rNWsbdcOW
3JZ8aBh1i9Y/CkDVNMnISZ2bYnGEcEb3WOy0R7halz9gqM8sRVrxqL50tuJLtZLY
3txpbXN2eV/HE1xQBkrqMVLhP0Yi3DffZsYO1HbMeodDZLSKoCPgBDKGCAIAUBWS
ZJsyJaEjIcC2ShmC10NkSJegNFz/rJLzjQWqgmoFlDMbMEz07UuZKP5PTHSMfG1s
r4T9Cvm/EkOq/OYR/rxXbOILDsJUymr+tyLQa4LWY/VUhQ/xhVHYuuin9mg+/aqW
oeRsDwLcQDesE0QHToBUuS+h8jPxgLTm0QhB4eAJqVzn7RT5yRnBx5n7HPVpxHYq
0LiCX30BhOSKkh4GP+9z63BULPzkS8xcPn68oHhTqI9eiNUIzxzoOS75oYIKJAqQ
gj4P2AZVwekWDHOLoE5r8KzSrX+2hjdErM+U+98OufEvM7+WwUJqLHTH47KjHgp2
s+iDBciSqgwdtSECj8aqW4LNRqv4Lk21oU0ECT0HJlePk6d7AZ7/rekDemIcMuo3
6bBWiZOl1UvK3//65ETXk5KDv03EXesnN0fIv3I4VPfzF1xRmNqlFDb2j5UHs9r3
kX6Yj2m4Eqdskg3716v83rBPhq1Ihxj/zLjptfOlhmi2ayiGEPgbPfPKflI26NTd
NIHnZbZhmy1VFx6aJTZ92GJ95Uv5CqznflhD8h/3r77h3M7zW4B2zV002Ekw++6Q
7QpYuxNfA3BuBtfr/k+ftUUcWMXUQrPI9M4xB3frVpt8i4Z9adkNX6R5/y/hfZIR
7Suk1PsiG2VaubzTvlqN30Z0KwQa41YHrq6vhfXRyaqfQGUWW+TfjDLDObsh+rgE
Cn/MejtllxZ8q9eL0pPI32u8xooKdtgBrg0Z8nbhGsVHQVdgIv2nFD9VuP4Fj15K
M/bj5WlpXXev/PPyCdXJ+ZWM6SVaxeye+cCs1WPOX24YnyKhDLlsvT1I6rtMEzuZ
p6LnrY6c+6X8mM86RttP9UIF/Al1SHzx0f+KceJ8x5ds0MSyyKcUstGyemqTmyWh
+NCpoL31TLo/Dgcpp36SjLi/awcF7BzqMDWDp0h6bpRBMhmFNEqcnlW3qWqu5kFr
HAkMvpM88EIV46sIVQdxbxQKWjGzlt3Z9wUoqzGw/9MgYHkIXyyOc1MyZQnsEg1i
lETiepeNII0spH56zWBJTdNkRbQHPd394OegfzFHipebzj6l2spCcWE2QbLG6YFy
nWxGuMI90y7D3NbiVqM36wYaiLeMBZKTXmmgQMXOpq1HTJY4o9q4OuJ1ZONMXhVE
/TyEjeAeRGzYDgtZ2YuJjKuvjXWzHoThRQ/RsYXm/2ZbLcBYS+Z/IjM8jAE9PjJT
MVVYvrEAy+KPoNQbRRFbyuVPxp0Xhx10avN6d0Ku/YIzLqiIRDMFv/0GbuCW+IxJ
X4EEU3OatY3JWsQNbEyDTo+QvUlUpSUKn1TYAhmU5lQS2G3g1GwAt3dKwBUgDze7
mR9CP4c9zOV+HoUEK6U6U1XZGe8DhMF6fNX7ZjSBdx1KsgSI22zxpePufBQ04ypz
T8eUTn0rb+ys8u7I1NWDCPK2hOZHyZ2kPCGWldpfq12wTO3F6y9fAi6Rol6FVFJx
LanxDTVG6UUZX5nU5YAhd8bIquww/pCTX23oU0HMVgKBatJnO/2NjOCvnDioRRHv
ddLNXY2XH7TMNDIA9fzVVBeNC75TZCVHq95iERhs1p1JUddnP/OQtfNf047tWZYH
irO19r+y1LxoevEHsqOck+CIyebfZVAe7WhvlMWddwQo4JSqp5qCeV7vgqSAHoMt
FGtUTgsEKvZAM56ZUlqa+gHGUVPoihBTVQNu49/n0IracfnIkcp8VchcIMKpYY6e
Znbp23FOLuj3IiAW3Ol9nF3mp785Q2MvkPaYuM7Q6OTudMaomD9ZJ3RE4XR+L/2z
ZEu+h7bFhS3A3HmjPsrm/M4Ecuz+KlNMlxZuyRHMBfnxmugyPfDH4sKu+B9hENAf
97YJuhHLSOBoAP7OnLv86Ns4JWptPEgh+EhPwjUYpO33PC6nFife5Q1rg9gIHi0x
1tVnMLbNUAv3vM4vvfFaOrcxYDR/cr0IZMxuOK7kHWFcEF1SNOkkV7Kt4Xy5qPsq
JG82ZxVogNQOMZ+xEbB7FhYOKl+b6b0YcT7aQ+3O455XdXzXoZg8/L+OcxxPOYlF
xmBrZ9/Kzj0ZnFF6Rr3TUEOD+Jbna/gRsc4MR8pPqocWgjtaJEUy3DJO8fSkad0a
toKr/QxFJl3dGH+kUi7qFxYC20bhVKkc4rZiXr4nujFoMpqrVF/gX1qlcn0K2G7V
nhkrBZwGK8JAYapnkWUH/y0JGBaGI5dUPhK7FSlUkNffAV8b2iSbEBLkgSABymZq
vd08hLBAXZPelCB3i16hgOPHy2JFq6ehHtP3GTOkXGCfdt7XBtbAAZ0rntdQE6l5
QkmL7IOP9ocqETmM48UMjdIfzcOgTxHNggRGf3G29lQ2Pj5TTNRtSyIiEtyD0mji
CThXOgum9uWPO+R0Tek8Dxa858I6avahjXvwxInMXnjcpgZWPJ7klNI4o7igJfE1
U3NcYv47oVQ/H4oro6p4FU+tEk537LQhyj57oMKZT6vlRPCWeSotsaSHgCvgqXpf
9pAdiNJLzy8ipUPpbribfTs0LUWVs0kZFPFZ8WYP6ZXjxx6orC3dOz80c0RTtVTc
m9anzwnNpKxyFoZgADujcvwCWqPJn3l/Ep6xY2y4qSv08PFPjqurccMhIuMAMJPS
KCam5KbiLmeGoxx9+0eAvY3OvAHAG+zY0xf/1okbshB8MGzWTFrgE6q1d6kxfCgA
Ny+txTw2NGKEBlKfp6Cbrk8AsNS6npdqIJ0hVXLYNHj4UwLlpO2dni+PdDQXt7jl
Dt1DPhxFs7gzWcRUfnUD+hmPLldrEITv5GijAMV16h2mlt1wLAtxyzxCl5A646Lx
Wg6CzwkB0HSA6HaMtpHZEFoXE6rITlafojxaoUYiIkXvSmWDAJdnoyt1eNEOGPQ3
ZTeVAVJSt3YRFn7lpOT85gdtkYVGeGoFIb02ufXrE9YNnkfd+nfsZlivq41EVvfF
UNjz6Jw9aJod27NOVmVJ1zryPu5YpUd0JTFDPROGruqNJTiZ5b1DzvaGNPYgd3+J
nyTY1WXYURLMxu7ZRvEsYhacbQ3cVL04zlREK2emX2qkFRGwvoKpsoIEO3LAfJic
ddhXQUPj1uPS1MYgsYAYKNHiGcHtwSFgIs4vRO9CjxrBvPJ3CDOgwPCo7zrRPWdx
C5ANG1kh4UDdyvE7gMso4vrjcnnT2ltrn4+H8zAvW0QUgapms/eKR5qkrsT9ZB/u
X1Xm6cckgJrPSUBKoGJMW9scrt+ykVmj1GXNeh5m8A/8sYxQ8ECUMoZlys2n6lpU
RbjEhFcCNsTK5uLt45QBUBiUZm3g3liRwsc7Tjp5r5VoGTjKnXow9rqNTfx2SbV2
VzP4rLuEh0PYOR5n4KkcxdStgL8xkQlOylxs9rGykM5Uqzpzqz3zw/OwsHZ3SJUe
pCA8oAdo0KFE0SWj1jX/1+Urdkj5BmlK5b8qXfS+quNNl7cdyCmdHUHCSHAUYxY4
iGS+l1GC3+1q1MbmINIut+lCi/AHBHjNQ/SPJmw11E8s2ibeeZmEnSl9kKm+r2eD
8f2umbHN83ZBri0OAGFwtofE/P8C5ExY09bpawi9EcHoWpfkKPn4M3iGF3Ez/HGA
HNAZgrhxLR9GVwbThU1MNa3rmGN9Ey8gmv9I2MxE37fX6HqFAStoRvnufWuPSr+u
9YuoDmFGax51eiphxZZHSLIVUUa1EN7dBzKezsDSQPtXuzkUYjdtk1PXcWMAdZH6
BhI7OKk7eDFKstWQsW5Vp7VlK62e7SQwIKu/IWRm0YZpx0xWotQxxius9w6wdeYg
7iGOuG8gg2DjKkRDBcfNKGphsdM3ABHWvlMZ3zGxifHm7jKXD9fGUlIVX6q+2jDX
4bIckHeq+iOSS85onq+3c0MS4CUBonOVclx60rp9Y7yDVUj0cWztRG+W8vMWbTA5
SIrTSot4YRs5UCfOnJrtXCefv2LhrcnMrrboB6a6mMjpwUmu7wQ1bk6g6C4Ukytp
CmIpY5+ryeM3zd8Q4LJa/CS0iZxxFLY6RSQn5BW8YrfvyL9IxK8kV0zsU6AdSsSa
zkTV2dSpc7ujc4u3QX7OYDBkrUmG6kWAsMM/2hrRsIGdYRgTs314hW0ZLuyPvvBs
Vbxih8kGRMaFjbCBwaSBg1195rUltJNjYKLhqP2fl0GOGt6AZGwUsH7Nm92UDVk4
wjY8acVi3nXJoVHTWfl3zuY/xO8kWand2zja668ibfchWFjFmnfpkrLY5bVPRf/i
oDqIzQz4JH0yQDC4/z9eyA26qwjjqAyT7ql3Q/T8eOEWUKAJnMotnnXeQkDhZrBb
w9MzESQQ/UrJI1Pc1RTCeN2LLMh5gSODSQuKj9P9TlwD5ZBWMr47kA1+KRF6Tpsv
tOCfu/qCnD77PE3eZGN6YS25KHj929y6eIrVYrR1si7aIO/1Nvr/H03wsApy0u5q
JrKt8hm8fESPE74a6j8rvvhSHujiPfMf192705uvGG3KrgU58FnYIJqEJHCcNZhC
bM1smcfksmLz1ZsQZl1SPjT03P719jEa1lHwI1Sp1q8s3R7RvgCEMMA18/6rAY5z
2QpoRHjHrO/icG/qXxCBKyaVvHgE2CrXwBjZ5/uM5V0SMM+CpaFyJ2AXAO94jUtH
ssWlPnNfo5RAUuWL4xmA0LASEhX7MfK40jkahyLiTsj9+31BuRBYYrFInH7l+lkl
i34IRbZdJmd+kgPhjKwcPdycFNj/Nvpm4GkZy9egknJEOGsMtyxXOsezVekj86Fp
v4lW70hnLA/d6quaVjq/pDRIp22rkZKjU/Lng9kTAwkWzSDO+r95o9wUYMkwzDqS
RLEM4CrkBOHmj3gORB3XMIE2opts03dZHPKlPAfeBGYxj8hwOKmrqky+ExvHCqrX
MquAz51Uz4mh6su0aVBn8oAWMQddFh6btkk8xuJp0nxaLKbTAA+3Oooveb+I0v07
vyBFtW31fmA2NP9zpa11UKDnRGrGmUBXPHBiDRwvvTzksFFjirID3fRgja89lnd0
zIsZkXrhDXoisuCQBbYz3hybWR+C4inZBN04Z/PeSp8ee1UQSURJrfp2u7k1JLhf
hx4gM8B2E0JTOLgaUXDQKtodsgcaVm0hgLQEu5gt3t3jSei2gNn/9TzbajbUYreC
E08ej4XwpFrT5WPIxN+2/JWRDjJ6EO48zLPa02G51QywwMcvwl6rGADh5UuWjtY+
+iuCvLRLQPPYZH4v4K4NcklaeHskxdMbHLJPkNn2I8RJADyQgFRQh/oPc8v0qnnv
1Hrlx2VPYb9z7N97GSwr8wHBiOd2o/ZZSGF3fHFWztW12rZr9TsnvbkMNpputnxx
v+fVxuhc9HDE0tibB7yd44GxbPAVqZsZkZHyuzR/pgJdQBlsnbWq/f2fZIQ7tbwH
LoJngV9nUoivxjyVJZxeT5da6toASTuz49QdTgJc/zDAnKP29oqBnwLqSFhUziRC
CLdvE4xt6LfRdx3siQlgOcJIlBrzM3pMJNdZyF1wIKyeaysRbyNVwPeacIIpa0Q4
VOiOd7CVVjNDf3Uvi6NceNqaKRAFA8rsiMo8GeC64m1xsLkgPC3vTgle+jXQvqNI
d4ZoAMEfPj41gQJRgYyLmCvisN0Z0RNbAY2B8HcSBik+CSHHAQxMXs1V34b09jKO
C+19ab29W7lCIfvBE5QtSxZixO7/vuqzB06NLpBI04UyG/RFFs/ekxPEovFs0lN+
Su0rzq1NijObFpg4UiTDyBY+6Sde8kGnqsIAupSj+x1slS8W3lmGVNsroNSxTLgP
X4J8h6pIPPQuYCScXUIu6sXesaHbU3VgZ3bXT5XEyBjQemKjg5H5RcTAkND9i46O
eoQkrNgOGcDt4b0MU8hchuko74wAY9zNwH07XMnsp3kEyU47sKzfyrNiB3suIfbm
I4tery3Qmox0McjnM6HeLRVwQIVKxg9oAlWPzWEBNf0wAJsLNLsVui6nADYQTSwu
4rH8Xt1G0K1cndoHl8VQ1+rbwCh3M8zNk7ftMMGeeb0ENZgqg3pCDO96SN0UNVjJ
JO4pPFtmwEMPHE2TKIb0E+eDDJn5lzPM+ByUteMFXPHXGOE5lFzWuJR2sHnG84T8
UAj1Mts3jW5SuKDrn9R1if/CPZ0wKXpVDooE7qPtK+Zmwz+euPhKSJDuV8Sdz6o1
m8Ay7Adtc9+rBgPfEyQ9cyj3i1z6nGaamZlWJVVhNJz0BVATVfa3E0bbkTgCiDBS
80oi0YJXJSzGb0rCkEw+nx3/QmEyA7M87e4G2VDWjjqMUUmeygB/cpYS+ejEQS2e
hq5aep2pAXXy6f1mwUoUZHHK0QxyS7B8U2xKVqoXmlfsnk5EzFsKxhd1AqcPXLcr
BNOtEkmaqgh1sxCibwWg4wawZetq0eR7OBa/8iaMSYXfI2SFe463nv0xqGAHrwUr
1xJzjGKBedFkGYDH5wemy71AL/bdiE/h7w0URLyFag7CdUY4jAZe4XdkJJv6Gnyz
SFQDgldcHuicy/Qvws9eaDCjRcJGzbrDzPUpX7mqkSWp6Uodj4+SlqdbIPQYXTJl
9r1YzaIRCGMLJkWdbYJ5pi2d9yS14uEJdK+p/uC5pWaRuea1sknS+o3HMJ9c524F
lJlEK/Y8Jg91/wNpBSZ5YqdyZkCcMsyGhE+ys7e3O+d+ItnhuGPUgmr0vroyZ6jQ
vosKcuJny+XoxxlFglbddXSOSSk2aqXwAFO1bVz3Tv/FY79s1/5O7C+XYC5gh20K
0KSFi4o00+n1wqolyb+D6x/6qndiio92DWh2tO6/LAWJomipmnTh/nQSfnKbnEl8
Hh8rLLl01gUiah4suFQVE0AS0ftX3gRUiRQyq/yTuomK9/Yf85eGbx0V6RnsX/3O
8G4EsELvtYrWhSoJaPaC8kGYRBNU7g8IzhJgkttef9TB5U8ynKBqJ3g+0r87nKPS
wB8joe6lPvjdkN1br/HKRjSDWT2hp/J7OvQR75lW22oe/RreaHFZ7YGlOwQIsUxg
iiLHmGHtrzISPWeZw/fbwFeWXZUi9Bokha/V/ppV1P3n31QuNxSYBUr8vG1cydGG
/SnkfM5V1yiSCMKBl/L8A9AHNJuS06mhWTs6VuwjP7J+BRwmisaPZVT4obcR831y
SBEQhOOV7kC5uLT4YLMYsAJX5k+nntwz1279qteWKI3PRJ5JUYQ2NbuDs0ddgb+/
SOBfc8neimdezI6pdijfd8oXPm62OIpnTiWLciraQA8qmLI8DAdbW6GLDNcVX3/J
h6Wl4BjaeKdl7VFwVLhnkzvimdsU0AWtxy5FjH4nXf7Bws6UU1O2zDjaR/VB3RFP
dGCXQc2RE5bFG3b9UjqUL7HJX9MVwz6o5ml5gIzqq4x/+0EVsIghdSfA3UfjTmp2
ZiaVUpodsHFNqnQcfEaqr5sk80Uuf5iXnK+s5ikjzsrqG+vtkykCDn97t17tLANE
aMnpNvPuh5HFsf/Teca0dzOk3Q0euY+PofsC7y2xiKwaJ0k6OlpaK8rQxiGZuiQK
iKtNRLgGawQkxA88xTp3O3FqBwDl4qtmXIilZS4z4+pZCKyx5oiwDN0Fd1ADHLQi
nblSA5sCjDTF8VzhGUC/1lyeTQJeJ18ENbBioUjgInmDJjVxk1CPqXwVI2VW/T41
5OuWJvZn4dTwyuM3UG0zHeoR3ryObBStgISGUODsR17uTocskySQOsBKghD0JCNG
pk1m4wBlCEmDGe9oJWupOCb7mAnm5p7SbYCi7FRiyjf2PnCwF6BMu6uazQZkGpp1
+Yyr0n7rLcxHlMQqwgYjnv86AxyOgdaDgwElwDaNhQNVRCEsswPaRqgsr6NHAmHi
eYxP1+ngfpXx2oGyO3JVXavEaLMrrV9Qxf3+cz4OenHvy6wq4C3sdbulq3/mTXpy
3lUYdpxKkO/Vw1fNtAGqAKUL0C81h0zQWmInCcazqtA+uwNDO+szgoWcRkYizgyB
RcdUguX9oD98bV8xT/tT1w2OjplDiZf88UHffIgEvtdrrdkkeXv+jV2Kt0W9f1K8
sLfZ1LGodCsCuAWMW8PTzMHp2MfziMavyscoaEcisyo2im/z/o5lnunS1uQKMKzQ
GboVF+p9ZbAuZRRrhcPv2u+mi81rBYnMdsoYwm1P8MBe6qjiLl9Nchl2opqbvRbO
zpN7bPUSP1QQwf8JLEBt32a+pdQT57RYCWL5PgIG4dCMAesf1TOfdn0yGMn8TanQ
4RYRFxF0LYkTpm+3NOUHYmO84l01w/delvOluwebhF4nVMqCu78extOBnve/VsFK
DlD/Catx5KrOrhksMqKYWIzvZFUShPPtvJilvZUzma50sCCi/zHaEUjAA8aYlZRv
LId+d3RHtriYu07H4s9j8n4vPZimlbgRBW5ydDyz+iCfsoelq8HCr6HXpYRvOhMb
ROr9WrnY9k2DY3nywoRY8re/rAhZRmsydsAxunk+e2EOfHGqzrypYmErk3Q8w3Q+
8wVClm5zjrsIESHo1VYaCvl+6t540VPUNn6SeQIuFGhzYyuzYbrgkvUhzWJDRQQr
6Lr5PyRf+uxe607ozZRaOpT/fbaHDWc5dSCBT4r8W9vcPijaTnbg+aip/KbIljf0
wJYFKgFm2ll6I3vGFwp+e3Zzk9+3KB1bIRL5x0mUCYEh/uE/pSzR6Siv9bx35kR1
rHK6BhhD/yADEVwD6vryhSp+oq4VxhRxzzLFX57TwSSKhl1vL2yGZY2hbclXFewz
RN/wy5CD7tQhl70w8oqi0DDmwRdMPQyTgavykmOWp7swo4ve/tK4Fol3K0nCys8W
TzFy3KvQFN8mhhx+z+uQNA9XhJt94zY9suzya084mpOtg7z4yAlTCyRQMx3crWh6
O2M3dkU9Jcj8CrHLP68QqyQqyycU4m0TxReDtCok8NyvGOiT6qDjkSMrznry6Eo3
V7mvxTqGWKxdJn/3Xz+0jcma9+3XX6lCbBJzVaoW50kF1JJyNLl5FVR6gs1zTr9A
dl/9ZG6z1Q2h6U4sDQRP2Al/TrkAP2PEZm+u9aCMN4nOYrXJLX2BHrYmUG4W0mPl
PpIF8SGdxqMsnnQtZMcgc1hJGRlu895mACyu7wbpR9HCIhSUvnq+5hZm1rJ+gTxj
Vu9ueBlY8sT5hVBfesKzGrKjUX385PaMhr9z0uRSsXxAIgArIR/wywaxZ6vJEa4N
gwUZ9UWtD8Vsm1qCTYPNTKYdegtGVrOtZXT0MlQjDsn8jkn5R198IMsGvkRvtYVb
01x+VSTbAop6jpbxPHy651mTH784G9ay4wutR2MWmg/fNfddLmL2lK8mzMQtqHL9
zfuCyWt7j4O+ni5KoH1AzWKeIN9krYjoDWrY4XDhK8f8as/tVHuALW13uJOj9OBK
rq8Dkp3zWz/3Gh6Af+G1+4ySKQPwA8IHkG1zPVIQHvp+NG/KhwP1rh9wceeI2xTA
mRtTd2SEgWkV5ur9j1QkVGHhGX0+xulQPlj+v6TUGaMOh8Ov/Sp8VZTZdw6HkX7M
3ZOyxgNbtF2shOZq7nsU87HR9uYRSg4BfqGjtHi+l+dCkD5GpvJLzxjSPB5r/ZGb
8cBK6bnHq2gsiMFef3EMYo+CUor+YWFR/eKNOO5kFvKSUZ0yRdoJ/78cteN93M62
Fc2DQ5r7SYLqmdVb88sx4I/AqIalCwgAz7zkGycV6N+CxkjHYI9Z69zq7BnNlaQt
W4ln1xhHppeleYOmIJQsgESfu3L7ndl1qg+oDqH89GKpURM4OAt6zniMk2nLckzG
fVzBNQgLPKWtWDmJM7Z+J325R+o3irQWrEBDEmu2K2L0IsZh0eedih+EuyKw+/OK
Jw4DMNHxT5D0qkOq9FyKH3rux1r0lk+vkohBLVHlg/wsEum0BYxWATTTqGP6Uzq6
PLkh4Epc/eZIDiwsyOHoqpW2Tpm5pP66UWbEGuyQ0+IChBJ/ONkScWRgh9uEGlYN
iptsqP+7w5I0CZTG/4p2sldKcMSvqGTECIN1Vjpf+zFUHQJuZkKQ8LRLDKfAqlOG
fOwHx0ELcs4tv/c0HymOvewIspD0FSz6V9bSnvWZV7GpL2MjuoIB0vPr8zcg0Vmn
SKjOOKNsjQvdIGf1ei/4sOM5JWWG2rB19Dv4GrCHe0M4qnuZDeLe2CGycMDlwrsW
QLNu33v0fyKynbe3aqHDq+QXxKiOBzR5Wrf89rc1zEovJd1+aSo4bWUKs2RUEBbQ
G42+KJvnJWEEivYlozn8ifPTkhWOhOaROpYpRCARqIGrBFlNR0HalS7PxP6gM1W3
yulWw5mjPw05dQiNJZlc47Q9WUbdJ0YlGZua9QRhmtsWPNHkQhJYXzUfSxa1BJug
c7FH93vwVrRksdTNbixWB0ELtVcXWZ/YIt1XnH9UkN5Q0S/4i+vYolc2nfsy8q5y
2vma7VL0S3zkd1P2psRCZMDc8ZdThi2XW289mQGMJQ6q/XryegJ65Dn6ZvMLSMRT
daaJrrGYXvhYwl5ghW41mDIYLMhsk+QaomSM3+Gz8CfFJMs8GcMxyGhUuIhPRg7E
CwEEbDX1PQxYfpihKOvRJ4ZJ+/bUPs7id5/fLezOxWjZg8lwQBr3AEOOrQkf8I1w
xBIggXIZVvKCza5kuuyN/ABYYM/E4tORQlOX2XhUj2JVOwkPh1zGEuP8vjSN4CV4
XwRDnfPBttT5h/pP+2B0B15Xz4SvvCILy5yMiGhRx7lIDTwF6tsMXVNu/grgrRVP
E9topShw2aE+doQXhPkkmHQ+nQMKf/EdULF6xUP2wgkph7CNqcQgzrX+1lHh2KwQ
/bnGl1LOmEr4xz7Z3XuEpnUsDy+ZlDtxFGXzVTbJw97Skn2+ZcSVR4kx07zwtCd3
uUJ78hH2gBVrzwdw3k9CSLbPnwXuwYZ1WGbfMfJ209dmkYBeIpSukyvD8Y+xgqO6
VQvTaIbIZJ+l4Qj+pVxj0sFpptfzjiJO23Icmoe+l6PUmNXG9hvouyrZpikEJekO
2yxRAqr5j7b9mkSPpJ46BD4e7klM1BIf5Pea+/9FhfICq/C1Rb5UcLSBVuXfqA4d
dYbwd6JvoZkU4buorgmZJKEINW9u5EJTWU7zr9TxFR8k4OwA4MkHV1jc77WIWcLN
kUlGUlblVDQ/Sug6TO2fgiFAcFTHo6KUlcJrujhTScvg1UqHqc36yh4oLiTAXzfp
Qp2S0Pb2Ox0jA2ni8aI3+FgU27A7r8snnOPaFgmAkHEpZ5/MZP+1iEKMmQ6e9EgI
cdLg2m8ydwJ3aK0nceV5Kwqbc6DSIYjIl+G5g7niVMoCJbchvQ9Cn1YZrVq/S5Lb
pjq7Ljsoo7YDoqBVEQYgCPowQAdwpKjke1kv2Ps7TxATX4i5fMpoMDxwdiRhPFIL
64ekC5t12EFa3SSx1FLj2Xjx2VoYIas7hujAB1PRR19AmYUmXptcS7bathe1HrU5
6GSeRDYdnqv1j8KHnRDwjKARGepEUIS7sbPiDQ9zt6knEEGmuzWFZ9DfzWr/O6NR
c8zcghP1xcr4ZYaPlRPI1n59Y9CnUAfK6M5cS/fZZimbTfQklawVW8JZ1YqE34tj
DL/EO6EhgHcY0RlmR++2TDu5fISCVoVEJHjZjRWL3aI3HYko+x8EGo7He0IRGAjm
jxBKS+p+O/Teqk94DYmb1s53PGJfJzHg1HkAx6cnWgEX1CKQD+xz7wc0K2LRRbI/
QhsjIg1gFvT1EbZHhxi5poUnHP1gmKHV9j4ORrfmrslM+A2y+LjBiZwWRVdeHclA
Et4AZsP3CMTkEtB1cXVq7UHlp87AdtvW8fdVTOVKgtLmckNHgzS3sICTko4FC0w7
hSs0s/yghXwU6XTuUWG5lvA5ak2gWi6/YWKF/VdPcPvTktxlSgHaQs/Wy+G5S7BK
lJAWOjVMUGltFEkmPSRNrs4amyqy3IAd/yukJZK1411RJJef+23Q9800LCKVDLDW
jqJOUyVCo2BnXqaNMS6O8QWkUe6w6KsQYJiEGq16YwusbKnrJQaaV169npBgnk+A
KQvKimc7JVQdlYaMVec5/sBwYIuPembTH8Ozi1B1mTrC1iHNiy6caUpLuyk+gMLM
CSMj4zmJ4bSoiJoeeRNlkh5L3xbFsq9E09VCRgF9UCuMFaqsLu/xBKePVL4RGXlS
g+m/5lySlwJ8CtBJNkMAUivQIV9JJq1cnjU6+LDm8Zi1mEqCNw3+N/WmLk9Dn6Zv
PaRYAT8W/F5dFKOsCjqFyNeKbi16dGol6vUGE1jn9at/YYt4MDbYYOl70w1Ef/m5
RnX5AHSQxZ1bxuXSdY2x/9UCYRPMPnz3oB91XDya0B91SALGW8lMWt1SiqXW/s/1
R1WaktsQx2cFUNdlqNQ09Icq3aZtqEWyNzZ7q9E01UfXzxhrWJMCXqrEdtqlElQ/
26ZoXQPDpXh8VbyWNs1pUL08lpRyL+YdN6z7ME/GkrBRcyiA56+LrVWIQoqeAyii
1rTc87xFnf4BGVYiAkd0qmKtsj0lEaiuviBodobeW6HuzA69EOiyQdJjFJKQJo7S
ibSQiWQdXZbkszpZi0Ni5GC6yzOvshjB7zq8XC4wuVs+H6oZau0okuhpTbAXhGYk
q4ROnijku589av5Nfopz9MbgVnZSGwAIhGY2OdRqyWMFzfOiW7DPexmUAI3VkZEo
6A+hF0XA99iI1hyqGisbUswUisfz88R6bYWGZpgw+n3wqg9afJNiRv4xnoJhVVGH
XAkJ+IVXK2Rd0afCXuzRiRIlpoQAfmHOdiWTCf7hXcCjbieo4WdAhGtU5y50HEDd
oU7CbZeCxwlf/7MVD1TIa6F6cTOHg5Ap6GdKryknp+MQdOzdxNQIQ2BGxCZERlCR
A1Yg6coB2vaDjdKUN3IQL2xEhZ4+tgn1ZB0LyFvkcuaxfBHd1zXcRV1EGSuVBir2
NWY6ePTPZMqkrIEshtk98yRN5szIuFS8YAtNBokYs3zjxyViEjj6USf5w3HX9YJd
BfyAoVa7x0ldvkI4IfMF1iCAh4/3D+SrqvG/d0xKx83bPOUItfjM1npWX9w6exuQ
TvO0zXiQpn3OEjTftK7IN3bXdmjZmMiqfp7Hq5NSG9bi95PRZPYDGmLM+AGekiuM
HllYivIgZOUQM+AYmPm89Fz+lMGVGiJNdkN1ot3P32EcSAFS6CoYxVWa84AhURJk
7f05Ng7DxmjrJfXSMVj1klJsJGgB6gc4HB7/kK5ZqEMboZpqdY2+13PgPv8pTsdM
BjrzBbr+qwdMhvOAtbAfHT3mR3E4f0YwaaDcm8CAnvwJs2qIeuP0cIlMq12aJ/KH
+YuAl7g6wteZpHvuzf41hrDs3APk86fUvo+tKZk2JbLX8/S6WH+ZKEhJ1Z5RCZCL
6n0mIdWxzWMIP/MVAHDvXJnohGb072bS6gRMd8M9BKDM2M10mF4+Sh8/pwu0tx3i
PWWwM290mveUjT8mAK+8/yZB537sg+UBXDHo2O0cLJry33W2SWQhNrIz5CQN5e1+
HlfGOGbVB31M/HLPmmHvxdibAPQGXd1hVw/Ovj0+3vNsaHcpg4SEthfzH5vR0VUx
P20YPsBDIgCwYZOvvhLrq4SEf7svFQGja3Ox7Gmv9wt9uP7i+8Bq2YV3ZzAC7YG/
kiPLPNQFCxjT7jy894jJ0aAUZK1faWK9q6Vw3eROmtReBawJo4frfew8JMtXPjwj
p2log97Qoxmpavi16DWiYO3ZXmPTHgL7H6Nh5wZoBqFZde3j+xYEDTK+JuLfECxU
OnA/6h1wHE9VCVOEu0umFoErSJZrMATSn+NzoFN4QEf6XwTMNyN/yqTiNky4E9Uq
lF/UozsED/CkL1Bcjgbu6CxawlIHrm3CH4vV+WdikkyRONXq/BEQJBUBH1JPwh6n
ESAzq2Ly3bk3ExGFcUeIatg6Nvy1pCCclfnP6UEDx/0W960oqchEQEYW/6BbcPld
BlixLg8P0lrJV7r2q9fw9ZhEPvABMQtJvU0haJSMPpZc4avPT1rIMqdxW5n/VdDd
FG2aIvsz7Y0vghVJaf4rcZ/v+0pDFPJuNOOYPBDC4KQA6dH6KSiN29Y7NQixBqtq
9A1ql0hSzjjT5EUe0Ys1JJ7v8OWdg5Qp7tptuKBLafGvBZwUCsQurNp2gZM7nLaP
3Ib9OrwW0IXYrN1GhXCNCZe+ZXwJIBjtaxXk0Z/lhQbVn4uvTwlsbUJ4XUA0+xup
04/PCgTaYlQ7Fy2cPwZf4ENCJu6BSiekPDzHDZcu45oTin2YBf6qTnG7Vke+Btop
yVL7HYSlZoLV8U/M18R3O7FdL8NGRzeH1NLVttiCzaV+h9ahZaOXOyU61EGR8CvV
eKPGGPKuGkYOsCIYaqKqHwOYsuTibf90HrIDaYw+QWTmvPrJB31EG28+1UwTBjEz
6I759HNO/p3LvmrrcVImZevW5TBjgftuGyKfcOb+1qtFe7M6lnnW6xZWOTbJub/q
60wykE7/SodngNeXtoOkgUYGOkx8ttEpm0XUMn6//shHvGgatkIIewfPT4ShIxk+
HZ6isOaueq+jN0seaUegm6Lo+3AqbsAebXcx0EXzXlMh8xShIFy/GVMte/Va5vxc
gB+WvE2HPzPM4ROErwDaSXnGd5OjArJGGxvedhsWNQ6U1WyjdqaQwLTI5LSVaPdk
BJhs3pNWb8j7Ve5grZDosbBRnsPawa5imbVbY+h6xjbujJ2RA+RkZiUJxuE1wCd+
xkXpqXgGTPddeLWApmmj7aWN1BMHGiAHAijjkhKgxftmJeRClCNvTFOFrVPOiDz+
67ucH4O0tp8OE5jkxJD9Yp1vKiMk7fNR/LH7QWTlXeJq/uGMEthiQixxTgNpE9OS
Ozl4UhHqcwtW0H5R97fIBxu7UmsNYpxB/o/pwjXWD8vaM4SECg7XRVNBi9HdxQzs
Nz7aR1aZl6zfHZCyn0GzmOCP3acVK5m/ekHDOsMngmw4gg9kKV99wqJo9rGYgLIW
syOPD28RFZL0KpGFTCW0+7zcvTEyGF9UBPYKTCmyCpWq04zFEoK0n86e7gZpqxwd
23JsOemdG3Iy/TGWT0V9HHhXZumZ+zCm3IuQunQbCupmtq5TeOINSPopgxvWq0j7
uAylusqTgP4l6pE1GJAaqfKskFr1+Az7V+56zMyqdkkRioyXJTnHHJpCfOr5dLHn
/yPzZaF9ynpwW35yya6yMhFurg/z8VXuNJzJ5nxw+34H6/mL5g8SEShNUL8Hjo0i
EID5kXlCTupQM6iJjlpgQwfv6exkba86M7hVqMRIqBPxP3JdCg9RdMXWwTaz1/ec
NLUBIzSGz+0krBm+5W5TzufSrG+N/kJjvUOMYxusK8vzqv6hRGW7tjkDGV6/BjlS
8hAYBnTtuJsrX2zjWD5X5BoyfZBM4Jfwcqng5WGiZQxiKmA5TqCG9V246/JfUEI5
WH/mYMSGMjsZQDB5d8ACO3Bp83zPNBNw1dGoEqv0YqYtvNI5R4VTHhjhUW3O0p0l
okhpQw0gzDkHV5iwfyg7/PKWWs7xrfQtHlrzE3PMn6lXK4s0+CdsZPR0sVkqaWl+
F0yiOVZG78VPNsQy/bujEKhfflwaOuXZyOksVBGjc7sYH1fKf+2YnhGxbTdIV47n
mDetOC6gWyMlFt0G/7M2UuTtfKoDoyxxQtcqufc8GMTbqH9RyvzYlo2FrVckphZR
mM+dAbqXoA8WD1urbLRS/7RA2UQqNBO4E5CbLo89oZFfruW5hXc65BVb+kZ5xVl4
gdq1IFHp0YLSBk3pNxkXitC1e3o1Xj8eMqCHLvCX1pGL9+P1MjBcqAjah0vQHqfh
SewLehNW3Bl1zMN29vcdTzHsud3FeWj8L3NP5avjnFVHmcfjdLSZjg0ouGvCSu6O
QfcGCEF+v3w3bCnLDQXnnD9AeCeAk1VCx7Df11+kIGQsvrvDC5gRmOFgVhtw1RzJ
rAZpzrV6GXDY4O6g6PcBVN4Snkm2Ao/9TScdpqOxpdpqNb5C8+wTUNUXjvAaM/l6
cLQg1Q0yfbovVKZ1BKJiKsaNLHnBFAThmFkyHNz46tJ0YXtuubj4ynNB9aA7GrrS
HnIJqiUzD2fPFlMIkY3G1/PtnZedKnoeuzDKy475fwhOd6NK1oH4cwaH0za72piD
DfYVg3XHj/oBZuh5DprhmmsHxasNWKrFVLrx8D6wSGJm+EUbdVa+lOaAVY9iSsfJ
bK0SpTfEzpX7qPq9yLPVq9tSbrfI5Q9GGYRQAzJyyZLwmgyZDZm+lrsXXjG8F1KX
W0e+FJc8tHBt2ecyT/6zssO8nq1WD9THWLcClrGfpyVQtM6BFgxrTTwx6FuIKDYS
nyWPtK57XjsapFWT3OeQX/7kLcG2Z5nz06pQryfmc7ac+9N5kBihVM0Rzrbq8K2H
X8zj1XF7izTDsketk7IdhZsydJsEXRYvQXrciwZbzEMLBPa7Cunp1hvtKi0nKwyW
vh03THQZG6dhoSSXY3uGri12sZdmxbayer3LL8KPEm30u5dDlmWVkeYJZ8Bj/AYF
I7ttJBz0LydGlBy2WKesOC2IN1U/B7ah8nej128PilXHsaPuWwWK0uerW/cOurQg
W5TSAxkOVgd6zzqkJKQ2E2WDuULQVu51yQ/R0rbwWQqvv21reADco5SCyI+rPmer
X9GzEAO7Easb/gL1bPCKLNp3DxuJBF4HLbvIWemSZPfYHbhJp7HhWi7ZRKw6bK/J
oPJ1zo9fzjfjZ4i5VgYXCrSoQe11vLyLkPVguSfa93yOOtovhl+9XZkJUALNiLz6
qQgTE9lHOB8JRqlLqWvHdC6HeZCQ/ExN0GVPfjF7zVwCvZ2GSKRdJGUVN/LKnNbY
QHJs2g8e0Au8zlUVhdjG8ruNy3m3iROk02Ai0IDAXIu35uGFEmml7Ltp43guoFcc
2hPRJ3Bq9EKQfNNsE4+GJUo69FfVV7ppQno9xeo/lp2wKHl2meRxNxjqBON1blWC
+IqHl/Be+XdtaIpGB6qWs2U90zSa4gSxo0zYdMaRee50uvcOPm0n3A/r/b46s2Pz
gQKf0yDxEdPzI1Ce/KCUCcrY5Ia463IaB+Zb9J2jMZBNC4fFCOWspkOuoCIkqSZK
BhqRlCi+sL2vbsMScotkO1lgPIZxDKNH1si02QZoq8GRtmyeqRGk41R7mdeT049q
h3Zn2kCOSwpdBZ46NNewUpeKBqUNzGd91Gmmcl0+pPOCWjx9dZUTuvWaYVNjdFBg
knwhd4mvIaNRWscSoBGXZFNq0o/5Zd3o9mNhfEaDOpqOB3TmDj/9cmm5ORtq9RcM
P70Rwgmzuxkdfn/ZPwSxwfxyvuMTk2uBRtpwbI+B9EOh6febUmfternwsGQEkM29
vl6JmanfyfaavBN7d5BEE+U+NLjYu09GFSKP9ywWBZ9LRcRXnYjl9PXK6DhheMfq
8CqKpJDlfYL6OuWNonhCLmwwCylwkHv/sxQodhQ9Sh5vxUFPa1Ufm5GbnEDwM4DP
N/igsA480C2+82v6Ilub61JT5sGccSmSf886Xng/roPLjUYs54JNgYPLuUNLIJAq
kC+6kowU3Q9CcfJXwfye8MdIcncHPcWt0TPsOTcsDTpm8kdrszHvIsPgqF+cTujc
a7SgH7wWrY3EQQjn2Wq9u9KAzcVo3aje68zwgsOUzJPmXCtx+HaMBWULMktJcBVM
qz+UtzYGs4RwY0Cz47J6R0Zy5ZCkeVu5DVY2xsvOfv0TBHGLc5oRJZ0mgkhotzni
wRd6j+/9WwwJHNIz6HvsHPA0DMpLNanm9FtZanKnTthmsvs6YsyRArmOF3sLF/9e
sWIVqf9qcG95Lu6mFTHkzNRpT9LrQHVZ86vdfl8Y3HNwiHV1T+TSPMTbpYRkVyGW
/bQgJ1PYagYuwCF45tRdYlgvBlu9xcaMrZGra90l8m7VS6TMsxST5OMeO4ze5O3l
m2w9APyasJXXG4TwNA1GCecJ9UKtfPxIFX75MdStJbEAL4DNYFQmhCQcWeUR8VC6
hWUl1lHjeJmOYtQzrdZ4szBua/bGBgr8qMhU0zG5xZA8FK77GXZ7qhubS/5L9pD5
Uy6DYDWjqke74HJ/I3eOgNsh2gtOsfgf7QYW8a0hp7BM9EBwxY4YK3vDem+o5Lr9
ZTmi9SuxaAXnMxriFcfIZfOqg+0nEjS8bgsdJqBpY0hZo8n7WbLe6ONZcYhLCyRD
YJAukETdHk/qLsQXCHu41JfVHjQ8RiW6IUA6nVFCk9ubIOfWnWlnCdsOcnrlKoHj
XarKIc0oia+hAplST1MDbPAKq6bzzFfYyrEKrIF0IwJI8+xK9uvicaLZa7D9AJUR
o+tKPDFrsyLvn40LNu5XUuNSGeKzPgQuvx5A7GjGoD9Lfgobtq1AGO7sSMpaFFVj
UKiTfSJZg327HQn/mHyS29HvPdJ4KZ7dXuxIH9yiQEjsdGY0U3PLLr+R7I+6vttb
3FvSiEabIrUzuUxoCmlg+hIDfKEnfKeZ4fGInSQxuASIQ403IagXH/9XKuJrb1pu
50Lc88o8F3+KdbY81st1quoFg7efh6Pryn4zbNscF8qdPRr4pXvn/PDS0lk+i35l
rNkRkxHNYphPAqEbmZr1Eo9Fcx3tlkDYkziIj50QUP5/UrieHRc8025ua53VIxvg
M1TXrxg2hg26kJbF06074h+LYjlvaiyxRKNxbRyUZdgPNMarlxb/0MvsD6G6tMXZ
KfzwdXeEE9DOfADOil8wzZ/JCPFJUqhExAnfTsY+myiBA46bDK9iGhdbfmb+BZy2
dhHTXilf3HNgw+g8BmAjfFsnWRf4OH2mCr7rCNt0LYbhfhRxIRZfH0YbqO1DT3ON
9JdnN9qS+x07qE7Jfex9U4P5OvxOpjROV2/qa6OtXfmaPi82ZdrwDe09GGNda43Q
zHcbvVzTHYS8YIh6zFizrUs00HXWJ6/PokUm4evApyuMHjqRoU0jJbH6c7IHrJF6
NMrIAfoZrVeZ5Wyo96ZdLldYimr9EkK5+BMdcGeBlTE6ahlzEIKHYH0mYyviNCUW
x8CrVvNeBMVMTz+xIU9pxi7yMTFecoSA6JKfmI+rK1cMjdlFIrDHOEAiHVSB+wkc
0fbInV7KYFCHlt0LBpazap0iTyCK43+n2gLKoFC7wO0Sq3dRyXmMMEJRhCFmPwSx
MqisGH3vV//pBXePUIDicYg98bAv0PFH72fp/rJhQFpb5okO8n/8kxKTMlNeqwBV
/gvu3FojU7W25ku3un76x+eQRWoxomAmqgNgUnY6TTLQTRjsddt6c18OugbIWETm
rXY+ZJdpuiuPVDNCoLJolJqOuocoIX2RmpjPID3FFkgREx6r2AEv82n16STCtHKy
3SoqLpJWLR8NzqSFgg7a8Tfk4cXWfFSZv+qPk1VTx8qEjr8qqv5oDzukdTMaBuO1
BX6ZA4HWvzkhJ+IfrK65T9hkYnqnMxjER5N4DQ2/iaXuRBIYQZdy2AwFO9+3DIBO
MP8qq1NzXGPs91Od0TTZuKDWmD0smDnM4HP1XA16egrqBpV1KuKp85pu6H86Xjt3
cnzB6Z8buCrg+i/TBzChl+UGc6JgCv3G/R9A9PUNLJ4PkhWWT5+omKjoMpoAysHS
VT4BkBq8yQE2E6DMNJGbLaYRkNH3UL5PtSVhmKCsP6PcjiILEKRTSaaL/o+YTMiE
lWAUHrAtt96X/imKf63JTz3QOOUYkKJm5fq89yX4zZD6ElkitfY0xV44v0sfh/RT
1o64mHsN4RAzUN6rCqjTxmG32IW07Zlfxi9Yk74+kCwrXnDm0fEGVdnUAoCjN18b
tbXD4sxcsStEoyTKelM691P8qHmiH2x0+6lyfpKEUBX7HbUDhks5gwF8vvXGHttj
uecsSWpCFBWiKYR3NCHHSgdMX6McX+FRAL7wbQCXH3PMVl5nezCl0KArF2ZH/THF
tnNpcJzIiw+ITXYuD4DJik9jYebJK36hbHwI2FwENcqJZHj8YN4EJNzL2eU4AuCL
lKWLVaULlOYzUQI9g6UCKRm5I0K6TnteRpBnwCBd1TeNw0NSVqlC1EM8PXVrAgm6
QtE0uMdpEB6+dcaJox8NeQU6VII4FDVhg2v0X4WMX2EIJ4W4oJHE7qXnjp/ZMNa0
O42zjAvtCHtxRr5bIk6A55wouj+4t8Q61PhmSY2biTBQT25SCtLOHi1iErahWH9n
40jTB63wpO2Y++r512xVn45qOWVJAWy9zQa8uRhUkaW+3yg6/0BA0OPmGV9BpSH6
/gAlP1vV59N7/BPMJB27WJSSXRlTMqQWocqCGaN2XiibJAjvcS/+2NJWbOAHUA8C
9Ud2EH3qgWorFydyfEitJaq56Fs6D/IgR89yRvrkcPVgyE4BzEAGOg6qd676G6At
PumJBh8vtHtmzGK/3846kE6g1x25rDyrY+7OqVbg/U6wfnz0VoI5lTgcJ2iitGVC
r/7G84GX6ebV0nSokgk6XE776CFSWZpUNLJzd0us4nlOOp3ipPiSJ4yhuksgcqAP
pBEZLMUbXZQWB98qsHuqJB18VzSFdJQyqEtbvKfG0w9ftbW2MukQaPp7lrvlDrnP
WHgernReQSyS3+CpnLVmk+A0qURPZvYF43sd9l+1ZaTQjVnMvJfA6cFa0uNbAko2
c7/l+cSwCyVenzRdIG840t5WdDxkSXmx89uUQMBEOY22kLb2EZQGJycXMnGWuQFu
dFQ96mhCW57hjspx9SCWw+z9qkDsUMPVyVyt9savtB7e+2N7Pspy7Oww+acj59WQ
0fbas9uHfi9XvuMbqufKE8LFhFV7p3Pzisq7orDTFggeJRBs5FgzyYyPw4cMtPCT
R6jvQFv/q0QyTnrmLcqJPL4Q6gkbGupolbgkPNmw3NLG7zXceAyYmw3BFCOESakz
bMO8fIZBXfD2qHnsU842WEp8nhVJen3cj7cjigOvaNgcUDykXt6Ut4r6Vx49H2wF
hSwS4oJlNL0OmLbE9Ynu4AjJ2dpNKHVerPwclBvkLADAsQKhYSwloSaN3txRVEDj
nGl3bBz9X40aPg0JOA79yKVETsFzsiXSuPR5F5DUUY9pVjOo76Q/ikHjaLSIk/lK
rXrZB2Lfry6nuGne4Nyzft8uiZzk5Beul0qB3OKxLSjYEQkz3pFQhbVK87sR6Qx+
3VO2ZRknbPqhDsjjeFtRqEzMZGbXGY6wXgZg/p/7pAytfKMZceOI2ys6yjL5mkhj
EoeC+q7JYPp3lyC2gcNa5FJvbV2rJh5gr7P3IJ5tHBb7uL520NqOkh9d1ll8pEpz
n7kdkCai9ZOEX1NE6yXdjQWO90epdHvWghO87il5CwjIYlhwdgJ1mF4VWi/L61Di
xkFwx0ptzxiFx46TY4aoq1M81ESJ2QrBSEf3UIiHXZ5TZAT7L+7SwYPGwJqKJ1T3
j9hmoazMjQE4O8pMFoIaQP+agXjDqw37XJAuQJbbcNipSiwiFw/Ur+dfTXL2b9LR
s7G983xTxWTMytWZfLQ9/WQ+0GPTIrfIz1BDA3U8PR3tUFZYMrGhs1cEndAtT9a3
q8I0xppgnkogegPw3381nyCw0gdd1i1E4IFBr+Fof0rAEV1WgPFr5HVyydc0AhlA
/1/ZZo0dd83LiV/Nc8c1TArCw1/8hMe1BrtM0NHCL4ISIY1JR75tSJ6hILthnwE0
whmuSh6SU17ydzBgC/kjNcI1mpKYvqfZoSYAaLxJi/B9/D44i18mUsxnQjcIDGTM
xNqk8O2DHrVgYXFg0c/b9u0q6a7iWSGWzAk7flUvAhLWoNt7CginSwmB2fwn866o
ccMwOJFe9pO2RNtk/2pPDl8jT2YpY7b2H4WVW8nMb/UO59GgqIY+ctFxGyzxxtan
G+SotrRF3xmu7YlIG4s/Ay9DQS/mC06cLYyMXj04/XCQl4/CiSQlh9/IFaM1tQqW
WWTXJ9cNh6ARghkzf1Cs2zmqeftfGlhtnquahKw3OUkmII3yzPEbQiyVvyHQQfLG
yij5BzM6vtcNUc6oUAitrg0V83gCZHbg5QAMkbPsan+kR1uhgXiQFobEMfSqJL3f
j4EVSrqWkiBAEcjCDTcIwRe1AGNsxLSD+XCf+zccEGEkjMceT2rQDgu2BkzFLtRo
C3h/1UdwD3Q9eNolRx1LgZmRESr3Az6yLFiXYUGVtSHbhnVr6rrVWqHGYVvvxoZx
E5Y/nH3tjYnu7ta0F0EZdQglhcV0UegQa4W3k9PI6Srz/rAmJTO0r7Zk7L/sqlpJ
XlwOD4qFa0CzFMU7CJjTvjn1GDSCpuLhWkcTU1zqoZvUi/KdvB2v4idf0Qkz8enA
hRtDUSRCOAANv7jhFDJpxqk3gXDnWXgNMT2KihCasL+I76LYYli11rQ6tilcjRF5
iC4RDnA/gAedas8adFkRgWS0uF3GaKUFPp92hXs/87xd/pQTTEW3OVBw5EfRgTDe
2wyXW7nJwndVcPyFxAWmbmWaCk1Notzxf/aMa4zwE3BHGr0X2w2z8A7aiyXxjARG
sB0kc30wCedD5KKCdLZD5ZoPbegvPUtfdr7C0PLKcHqrYVckqY7lp1VdN+3no3rE
8AATZrvyh39mo4XA+xUTQuRDlGT1X6ElplD7Ar2eu5ZPwIVzXF7QxrF+AHFwagFK
bi2Q/A3aCRBOLpJrq4n8RgMY4RQshhVOcdZzTFTh4ssqh+m2tX/LZ3xrJqMkeybE
ouSQ/IAzk1dk+1RV/0JdsmGV4UkoOdW9mCTL+PBqIzlCIkdFgA962LyUuoZt6+lW
rq42lbFPAnlk6U2NIb8yjjXT73leX4iKmr0rjS5Yv0F/kwFw7I9A6LA3q4fsEuPP
ziCXd6HepGB7WDSI06uXcHjy+tQrof8qHLeY4DFpTd0aeVQfhhYyezsLUfR/6233
bIoNvcMeR0+j2ly7V3I8w4ygUHd4EbPE/vGJkgzees1RMv4Ewe+/dxH1Es5agCHW
k9oUGUZGeYSCOnTeEVyrnaILUfkYDqetNvDN0ffHiAPnO0EPbj1wqGN+Y/bWzzp6
Y+uOiLMdgHBgyPRQwriq53Y+nGCOuiz4Mb8dTJCEy7J6vMhBRrgbVa7Q2DkUzh+Y
V/6zZQUfVbUMf1Mq8aC4gqmv1eXKGQ6HvGU4WD6PcUJynOww7+M1FUc6f7TEj+Dx
za3a4tLB3ErBRHTfu2kKTxEFvSzJ1G3G8oeX3T0PZVyqLppy8MLiWw8M0h2GHJDm
SMkemv7AOEIJPV7ibR+jflHulkA/0n9WrkFV5QBU1mBqgEoahZJ0UYtFSmGjvH1I
/q70HTsAONTnviS0iu7b7fdPqooMn/Za3CKuUSwatl307rExFT6zxKLP9lMa0dl1
lz1n8cQnouPFd3TtZqQGPq/fbui4+vUonzUP7BeNXoknahwtuHSzP/G+3a5cvZEK
mVJc1LXSz6feiQwfdWowjZnQVtwW7fpKTV1EZDUOaqCnasOqeIeSIFeeB6XKjF92
L844cyad8htsR0/bgqhi5Xd+5clruBPwnRx9mBQiCoiqJlVHaNngl1oWM73f7RQh
3CxXdQlAbGbmsu2PAGJONZK02Lp0JLDH2Zs7Oc4Mk5yECpJyMdkMMJoR7k9xhlqQ
EvTMv2D56TWMfJneda0dH93l+Nii1GIzYKa1v+ZiftPhTuY5Gg+UHLuPdc6uo8Tu
Vc0Tt6pCKDe4chSdOYu64f6r8BP0gYiImSe5rUHILDb8nGjRrkq39yQ09x/YlNkF
PRHEppBKdu7/Cl+nIwwifWdTpe2ofrjJAs2XqZGhHX5b3Z+B8zZU/Q1AMtcsg260
tX7l0Hebygdq+bsjx0fBpZ4UBiPKjChc3b8oaByQ9hqi0KNeOAlOjmoJbp/ozNLa
W3lV2NOdvt87p0LuGryC3NUcLciXlw0djqmyTRR1lSysOuEUejimiytJhIPoiHzx
PtKKSDluJjUemzviE8kd2CLg7Q4SfX3N/O4hWTcuKwFe/UoAvHZcSsYmFcEnewOb
JQjZOSFRJwAPELfzkLTTqT5DtCx28J4alrUU8feDWYhYhUwjAbleMID5PCSjv/fI
2FI4lbDX5f8a/4nIyQA76/AbZmika2GSdv3dFrJ5V53x2dJsNzNpPLIiKSdplIHk
YFXcDaR0ndd9Wd0GKphrty196HPVYtIFGBbFXWMsAFP2lFoMLOwxqODgNe3nDYSo
t+oN03DDaxeyVlPTSr5YYSj+8lh32WDgDvxo9L7UanxQW5Ey8x6D+En0lVfBCrTF
en9Bxcqlt1JslzJTnc+XDvMHhbilc9zng3Z8Ok/+hP2YrktQUgVLags8MT0cYBUX
Ek5Y0illfpv10X0w4A3y2kDbIQ5HGusOJ9Gr9QTDsTzSNX80ch+OaEvRe0rzYFWp
KjbLxvPcqvH6Y7h8XSo48tSdPVZk2xM53DRJfHb6yq1q+G/LfyyTxuo1Z0UEwjEr
WepXIGbCt0aeRmZjArudToBNAiWFyibHdZMCnbJvglWtsFukGLEa+BXsLX6DtUIu
BiS4GgSWeThrPClwfg43BUwWaS2XjIZGxTTBvCSFkuqpF3OTxfpwd/jaNOLsqxOP
rRs6sx/EXTmjeDDX42rWY+Y8qZe9ceJ1pNj/dknuk3UUR3jPSF5vuO+tHFGHxVfI
7qr4QXt3VaM9PVYBIsTJ2mP3Z1fE14K7DKRsNzMJ3EPbvlbS2jP9bSM6GvjFnQHS
rzhtBrGhfL6E3ptDjeiLUAzvBF7N9MsCjKNPw4F+EmtU789b+2aY2lmN1dmWJuay
/bYu4sXzMHEgmsSdfTYrCb+8wj+3ekE3WncIJastsyWvZunD0BFZEt8jyvcUMuOi
Syf4aghPicBB+LAHG9o2FZKcjmqwLU/fmI89mgnwSDw9YC1OQffGGC+KRJzYP729
C9sd4CBYOLE4P67+/tUF4YjRX175mFs2IOBfFsf18Nivs9kJa701fjKi9cJYbGti
IhtXxA96lDkeVD6vMwYEm3zQNW0UvIIpfwEgFLT350yu8ax7EHQtjxTLWvwuERFt
uS1a3vkUHuMgUpmnuneGUlBWA4haFRxk9Xi8H/QKhpzmObfAUU2YdmbZJ2QRO/JB
tKNq+xFkksuUITY2jfD/dDtybnRg2m+VZ4ZjZhqsPgzESbHdfkkfQtWXor5qbiIc
BLKzZA9yZkacMEKQ0pi+A1IIRO6+pQ5A8qkEzo1UVjxhWYjHxGjZOxPq/lFnSxO2
REGDi/aLdPhrH3ON7FkYndh35+RoQhKl2quoffjcrNZVwfzcfbJjCPKbF+NXddof
a6pPlZwSi6XvLwrbqmgw5smQYkchrrMlOL7806jC+iA+d0Sl/8nF2nrMpbi4McEK
ly3IPiQqwWFqMLtrDDzGzCiN3FZ6P62HRp5YwJC9uwj7Z6XmHq4q4Cw7pmZ+a5Hm
03DkBrXjEBC7LcR/A4Aa16T3+/vbgtd3C77p8pjp/JPNnO4i0I35BEuS2zMGG50P
94yjrewinVemCe1+XLxFfi3aAOhHjZPbiu8YrfQKI8WYvFauBzDZFnwMkPyl9TcS
4mI+BFnbJmLDXk7U0ZA5uwJUr4iwjaMQY5dXj8DwFbcxmtErTQvZ/wsXRsgPnx0N
IAtJCgpmJTElZXa8XICz+THzzRMi1Uw9zp0QlYiQi6JecAUVmKTj6YKEUcI/AP6K
QxUXpbesOUe3qmBi3a75E9MywxxFz9zJm/74UHV1xKKI6aO+9zNdwbRfh56bAk6W
EA4PafUVJrbImcqFjVqbUQK6WFLRKaCma0cwbQseZUsC4NeF92pCXOVsh5OcHMLf
sGBegGc9f7saoA0p81pcGz49h5ILsBq/ErjEg7qp20x2aNA5x3V4FYCwGueodRJK
54WiY/LXVuyy4CG/AG4sMqky7QVk5NIqQ0W0eNYf8Ltkyw9AHSLgLVcpO/sKh6Lj
+isMRSvZ9DCN8PtAQodUGKzGnRwov8eDBCDa64x/6aDvd88dtotRtyb0PCsjmpZA
N4t3/8WNptR0/HxkFjb9HEsAF6ROfA8pl7SDecOrtTadPmhzQuZacBthE80PxeSI
jIoJ63ndY/HCCk9UBj1EECCyGSskv5A1Jom6v2OIAB85nvCoJGCzf+SjbahVCCOK
Gpboe6oPtBsJZw1f2kDMdNWTJrHlSEY6bwTCmAvAfIet/tkkCUuJ0UdUyL6J9muc
qpYRl7Lyglh3vNlmf7x4Ah/U53XLD2PGTSQkNR9JlkktsIw8Worqhi106kF8gJsp
pQlGOEs6SRGBsaeQAqT4dmHI5sXgPljFOO4aR3M6IFioEdlUn1SUTXUeYq6NNiIj
p7FnfTVOusFXZhfsv7GYd+yqlbTifo4iVRB9zrWqdZnghYZmSEeoj40n74k4WJBV
pMiqx5uVGRJ452QCraD5FrTr52iQaB5QSg9tNzobxsxpU1pSvAyDPukiPi1rYQYa
GAGAPeMG+BFXxwyxrlV95KKsk0pcXTuG1fORJOsb5zycgXXaBaWtG24My1U3avtA
Bp/siR5tH3p+42fEfklUCVlvKWM6XvitGmBSwKD+s341Ct5C8sRrB76KFdo9K7MG
SBMxfyPa+jT//QQ8jwc+UcQdFHANKAp3+Riz8c2/ImPQEzXvdy7iC9iD8cnmc894
4Z7izDAPTDILGSgFPPZodSDESIikcaxW/FCajx5HpByLIghLi2uj6W9ZtOOt3DT7
XOmDlhsCyw927esbiJN0YlZ9s0jkSGK/zaqTtFCpN1soB/HrQveDQ3W3y0UlUuIo
w8SKe6N/4vfcs49ib+DbtP6UbqMIoB28NYPMTR0LcFAyjCWLwb5BMhqlxwdP1fTe
dUHAHasQQ+Ns+GGmyYHML1auURwbSnamTdUBAOANeEPEkFOPdR64bJeEDUgmUpZe
Kd8TLjPsNh0zf9Y+fXC+QKug6+WZ3F31ZywydssyhoMqInypMUWGYa1yrGj4n1u2
nANaufneafygVWitGB9n12QK1NBCJRWS0zPRlafxw4vPmeed6GIh4LFJTI9LZOC+
wZzHYwrsdye/zR+LFggMu6oPya2G93SiHImWWKOeb0gqGQlCAtvp+GwLWU/mE5De
X0ikdaWo9y/8giWrsQxhJllhSICtd+E8zT9pAPAdWUpCtXGW+270xvmoSGGxGRdE
CgH7s+G+nUFXJJg8G+QfVE85Ggxq1RyGI/Ca1171Cm7t9l5PMuub/NzdlIwoiN73
NZDxG8B9RHB5p3v8i26en2Q4vnbXLT0Ozbw2m12or1Dcz0uWW/vaNEzf1HciV/PP
okIqBN8MKHgKK2tsj1z+iFTKSaNPbFpGvhHQRdoEtmV8N0nyvhDdtuytfFoYpHVs
M5AK/dvB+OPkjxxuxyX1r8ACwgE+MSYo19LzR/gogBrrhvpJSS7QsrGioq0D8UsK
RI+Sva14kuIHWKSkGuOYgeqLYc35B5TuiyuO73gRCcCG+ur18cztRD9NFitkHNtc
fU0+G7L7ieUf2/6Q+CrUGdCgwCwCfENLuYo42xFXlBwU5vRgudkkc7B119TMKnut
MLzsfS2wpv+ZjZfGpkHjucGx1O7NRK7t57VIOH6gS9gyWc6Ok+Ht/RwPn9cU/AOY
iQ/DucPtwAIsvql+m/U8bSi2DJgi0zxFypnRzF7WrmKnOV600lMSsjmP8O147a0Q
CnMuCDGWTs97za/ZA+MIk6nYWKX9uBL4QC+NeW2qJkgoWAuJ4b/LD+io0PLRbFXt
JRarRNXZnxL/N2/Pw6FJomRiIdhOex17th3XU3Z2LcWyesI1FQ41+ZmSfcPVhQ1I
A6bnyb43K6TfVfnKrF0gXiKE1Bs7gAUQAp/NzrRMoTx1FUV8KLDPJfuzOStb/sY6
tF+ypKa5Bxmw8Srneuxq1uRVtxUEuY/uWrknw6pLtheKbyqXxw+93WnQ7K8RD71I
MmY6G9F6wVgtTvnuS6uqaz8G73NmL7ztquQFsvLZIfLk0k9QK7rSwkmD9YgYAKAI
JzwZX9CRKeG0FirQAV5oN06bCRlqU5ATUPn7KEVHOUSJ30BI7fP77mmxyrdF2blX
fXY+y2LAOYcR2oHO3empQ85neYnBWagy/5BGYxv5xpreBnQA86aMqBGWP9Bd51Eg
C/qm0Y8oPAteQFcT5dVmzc4Q3lEbr4DrtN26eLVmhmXrxYt/0UJTSmEtZ2mPWziR
r7FgZKXEAX76UIr944ibL7Hk1W57TRLmbWxHdvGfYCRiOYp47lA215MJzuSLAIAL
LGIum7mnJKgcUkI2KfLcUiJ4xbNt+ld1LwnVGv2DylGG1DaSITphQxD0kMXukKDK
g5j+nC5Jb8z8jvWXuyjTiivLMLV1M6MgkSFY/alcKZLhqZ7c+olJu3B98VYTo2R9
KYTUEGDh2CrbjvClCag9RRJPEi4AvodH9d+UCFWUF29+sBISNc23hcg1G4pmTbmj
TAAWXic5ykqAUb3O7gi8jHFyB6JoafHdejJakfFRLntY91f44ysjdFiYTuvrJqS2
WxDuso1BpgDyO7OE5loTCZHUUufKIAYL2pjYnu4rRDli25GJuwiooQgGalvvBTcr
sSrLOQJA9XawJQn4NPl/pd1Kc8JVQGj8/TmGpH/k7H1b+kc95fMsC32Z1LcGhCDr
lP9y0C6jizuu974KTSH/6nMyzq+UtiC+vzFBO2We8nFF+gK15BLL4Qt3ALT46fQY
K1/1+QyL/NVVFRoo+AuYm+XTsQQLJQoACXjP8+bzBjFv/GqUvLEX4D/27Fk+TK10
Vm9yvVercojVXgpaFbJMfVHJnmyiAcS5ui0R4KAXUduTWWJnTY6Sn5UpaOWAfY0J
kvpZW+S+HmOMOItnJrcJVePIwfHhic98+EYsXyucYG6teOFw7eRrl/sMSyoMtL7d
KGhzbqC4bDT4vHjAYL4LgNO4AanErlrW5RAvoXdSv2572gz2mfwb59F86eSWHc7g
hdG2TC95t1pvnhVJso+4c4K9m1m7aUSQ9T6J/RHT9in9e653AOS6O6SiNPdqEO51
WIMlHy04URazBbbZrfyg91EClx+RF2RAyXYhOLghFGjIpUhfIm2erkt69IFZq0/0
d6hrmksoTBMC0fZoIFcZElNSfD3nO2DvVHDQfXCuPYA/DNg6syx2iAXwE/y71XaY
Ne9oOkExdZT7n/nh9ZRn+RZMHl4hKi8zNz7RA5j4m+URPMES0Q88RZ9RkNf4slIT
/nr/NaD1DW+NAP98FnSdR0+S1LT6rg05fJOHqhLDUavqCrkP42DOX+PdWCUlE0Ua
7w4THYlvh7+XlHZ6ano8iIqib2KvNVVaau63qHCEj2Hz4BVgR2ojS85e9E6v+4si
+iTOmdH39pgXXUe7q0QLs6z7qLCZoe6gG5mo8xspJhzzEsDjRY1mjPz55zvSeUP2
B2+KNoazXN+F/hbafp45RLN5v3oyv2ss7FTgzkj7T/nx/xGmOHQZz5UCudMFiaix
loVgIMGQC9lI/bl9kr8rVaOTtIBx5Y9DxdYD9FutI3NATXox7OkdqvJwL/yQuN71
A1Ryj6I3qqxMqNfkyTSPiKQJbc7SIisNxgLOLZe2pqVj581j7h9QPqCQoveNQYZV
QnPg8SMkOu8tO5s0w3Au2UrfaODRIYUZozwi4plfCfthLMqHQo3v2df0jtRgp180
OxHan0e1inKvYCUj4uPmmjVqw/0Pbj8rMdeay1G0IlPgdRQp9Grxc/siw5YyEDlt
8TUA8f2gKv7BTUfa3oVa5gyKbbf+Xdpzm/w8D8qv5lekyrIT3SRSZb4nrYiirXyJ
09xD9k8ZY/DGOzYMeefwwdC42Y3tW1bc7A5Dps/pgbUks6Fsz4C7DGDPzGdPNaUB
yEcq72H76SK7BJ7Azs08yRvF4+tETQ3dpdyT3bjSkYDoASY2AIFVhpxFb2Uxd5vw
QQxxmTnSV/Xbsk43NhddYU8kwzH8epn/Ks9CYdzdsVlavCn+ZWYpJKcTeE50tbw8
Tzmh2yfhCGqfTPX+xa5dLmEqycQ+6cKprqGalgHERKdIbc1RVTnS9U0dDPHiHp4L
VJ+8VxPy6/0l2pNSaa2hqEZc8pAI3QPo5CdXTZov7gt0wEYVyoMZHtzYEaHgK5U9
TqbkYo/tSNkv1eyap5ivdKgvqsvwvOeWc2UNVn5xzbn9wrWttaUGuioKFnk5jLfs
/JdPwCVlbVwo3ZvnNmKwQ2DjwlZXjaP6CIB7jPqMYcFAZJBmRs4mD1YC3v1H2qpw
J/WzRrlaIVykZOKNAt9/x1UDWDLA8jNOUb7I1S4cDp9RR9i5ZM4/DChiJ/4ylZUt
m+yUc9GGF+1ofVoEEU6QK2yW1JaPXm5bzQRlq27iBrmYZbEs84j29LSghweYxZ74
uT0OTqRWBq5r0NvXwxxBSviqhpP9DxSTv6aKZZaDiQTXbovXJ+mGLY7NtLw5KcsD
o2D07w5X/XrAyLC0Mu8Ba+BBYHrMgYeXqnwD1WuFNLMY7c4boSt0EAIoATzOVm/l
YYd75EL2nDg1oTFhkCdtVvHxLOh5DYZShnqr3+TkX3hUZ+cMGDr8GDzx8KJmGvEh
IhBGS6XW5tfJrAmGfnwsMYMGUHgxXhpVYuv+RQWPi//I5jJoS8eY8qYi25/1QM23
VM//axNFxtKaXhwADvT0ejfqVx1za9di9jnyyt7KuCJdkf3LPZkjYDR93/wIBgGN
2ep0hF0g26MMPa8dy9C97xRsoEpQCnJuX/OKOVExODk+NfYDQIC5bVP7iItJQeK2
/5BGdehr1+b6xMFdND/I698gqcOPqhTKA8N6cOXVocTKYA5USuyrAQXAeydcoMgD
lxPIIW4EtQKCeIR/cUiyx1pr/IkwXYRKwDtw3DDCEmyfuG4o9rYA/rP6FEXXaUVp
c5u0o3+jHlivKeV21w4EzKo87L3j01Gf5SpvLVxT6R7P2hcMWUIXAoea8+8IpG+k
A4+lSBwolZQgp7hJTywRCoL0k1fCLBhZ9428uCUcYDfi7rjZutGXuqfyq+HkjE9t
40rB3SQ6K0HKTeNNS1i7ybVveEDrKjCnoGkeIXWpiPJdbwIEKDYagNMbTuHtIqaF
b1RqkGoWYJNXiz3szvRdT4EePC5Ki252/m7icwpdEK4eYTZqEKdWj4oEr8Q+OqVF
2qywhJCg0MaHCMJGGvVqoZYItBZKMFGRtOHTjrlY5JGuItWxyGR/0rxkAVLbKMc+
7MgPoWIkXhlSHyuEYXhzI0RPV6YlRaS3Sm8JBppSmLmhYEj7yMnKaaozCShOroHo
0RIiYsjQmAnJCCoIRU+ZPnJBAx8mvHn3cpGOh4hhCVUqyOfHQGhWMsP/yDI4u4Ut
Y9C/OK5Y5WdMl6hV7tttZlaFHnq0WW2wxojn0Y94zAU3oBliEQ8INgavVu67d3sG
vdlqIHX+KW3xOfztl6QbsXLrofUZ/NBXWWgmmIsFX09zYoMfVW6Wt8jyJb01kKRy
fUm9Z4awBZmZpiLcTvl8SaMqklu5v557MBpswIAaS0JPXfznarq/+6FnDflWfJTI
A7C0A4yKcD39mwv8+Ff9O3qT0wDiPNCfEobusMC2JVFK3GTt4j/ZA7vPBEaH7GnO
rOBhyjKNAcjvgBFW82rlKRREKeFpL1fOe4k2Z6k85N0+CF3RLNNWjaqdXJpoANE1
RvMBY+mZsaSw1ur5Tf+253E5hmQh5AQ3UZAjgau33D5fuNjGfPNj4zxkr0NBrP6Y
IZLJf/vHylULmyXI5jlfqcnIE8XyoAVIxUVlGex6kbTTRBb/hwrwLrQv9xxe5nrh
pGSIKEpSpE568wuf2avegvh1AG2eWDFe0DpFCtPcakGc2nHvGowp8l+kz6n+eFSR
Ccum5FHHaEN3+vL8S3kHmmNjia2oT3PhMNcXefbGJC12uk5A9xNp7Pqsqa2VK9CG
ZAGAtD+QUCa7NQ4gwBJodYmiCR2Uh/qITRgnTVmfgjdbHG1hPJxfD0otkjIXXOBI
/wMQbaGpHnObEtGKCqLCNmDBTLD7vXX0C6FWf4ZbZO1f4Jt5nweoEAwBOkM/YFs0
J499UHFIgb6wEy0Pv+Bq55ORqhwItNuRZ4IQFRCP6wS3sMrLdUf2Kr7bZcLEzu2A
cFWhu4q1VyzXXsalRNU1kgII5qJAI7rpg4cF6VxZ/276Mc28cR7+47t+jHtVPjv+
fe80e1OoMmsjX0Q9ZLMxTaot1AVxr6/jEIcM1U90Elrjx5PccN9XfS1NgCHzUxtD
WQQNQIKr1XkBzA8pLFlEDgeISmnxAJBzlY3iGI1jCDfgpdVqnjj9pqt3ToSoQnRQ
2GGczVOkMuv/Wt/o3PsPjxC2fkWBozxJ1vbMlapXlqQN1WyVuUH7GNQ2947w0I+h
zRRGbtwe2ejGnp60/+zXGhNQkGo7qIDowbZibjtYsdY7P1y9Gw0B3hsqIq20a8wU
qmi9JD3V72C/oOcjyz1jblcsCBzcGL9P0Sg+ioeUO2u636hdf8UI6/+2AphtMUlX
DjJW8kvAvCTmfWvSAp37YSUq22/kLk7OW6QgYaBZnGEKZxjDqU7SFdAoRxhxJTvG
b7jm+/SHiMI1NSnkijHrqViUT5VvA8hy26zIhVAM+IPRivzKMiJYaPYyGqfXdPEo
WP3GdWP/Se1DWOgaN4PxKfmsTZO4CUz0Q2oM4g52BZ92trjdKvUdReYngC6yP5XM
w68UahSuwUKyqaXyToTLeeRn52nh/q/qzDpbI2t9LrwO2pmOXFENCRIAIFO9TMAt
F64i0p+ZyBXF0dIFlvP2btpWgPJaTp6jZxPG1YryCDgycWX+1EoK37Fx7Vqh+2/P
RfvgIxDzgck19c981Gc3FOZUn8kR9EcZJwHVfLcDgM2rKQ3MOkQjJKtV+R93g/y4
e4ORKj3OJ+8Zo/fGJHZKLQENiYxw1pob/N/Hbp104gI1Zd7wNPuAwjG6X31DGRJM
xZq9Awmcq5poqxKBvnCt01yLe0gMdf+8gKcxUHe7tCBq/sDC0zA4eS08F8+4p8a2
1Gbds3cS3oqF6pC7XvkfKn47pQYDKVRQs/hq+qchU4WpJOUWHsz4Chgc8rLIRmeG
hgAUDe3tTQuWeBP3siNLW14FVo0EKs2ZF8A0tr+TLWlEKcK/pk9+DJuSEF4y5ClL
/YL1zZptO2Ljr4aLOdYfSz7AdSe+lsrh8Wp0hKD/EY3kbega4ktpy6vczIPxPk+t
XrYAe/aUM3SZFGrKFhfmjr83uNhhq00wtMe9wjZmm/w8E+M61x4jvN/C9zxGFw8G
fa5JNElOjd1lOXj0RcXBH68y9fbGM2ipDKwVlW4wzChY1F8ux1yjMhY7lvMZlhwQ
yC0RRzWZGBVXTeMN5r4FYW2GIsftPae1pAAKisKFOgEfdj5QUxHHdhjC/e8Ph3bD
bd+KKdff7uHd9knVrIeJYSO5+pctzjXeGs1UZVPwa04poRurFIAUzZP3yC6tRbys
NL15ChpKtkL4KqbnRgI9NlThIS0WvrDodJc+0jmeSh6ZoOymJvRkavOTPtq4GFIg
0y1SIavaOSE3JJcPPx9fYOl8gPGCPY+26bGLBrAa6ufUEc5u9A5C2amHj8m3k0nL
6Apb9quKlEdx5Qjn0Cnwxcoa00FC1LVArvtAwqJXkJ+VEMhqrPQHtlBWfjG3xoDk
JG7q3Zf/9UrWuu3azvHvXc8Prk4Us6CNmT0YoiatT3i+HsmMfl9Qari7B/a1qT+d
8zw4FvKd9iZff4hZ6HIMYfK+FO+uanO1YYSLmVQEklv8NtrIMNmLholu5qd117qs
J9mOi9N4vlp9AnAhNC9l/4wCFFxBnhEI+J/oTo5uI1s8bUKjd0jRMwXBFkfKUn1l
eG7i0dxrvmWTwSvNTmTuN3YDr8EL+mqKA4LiPlgwqfreFlRtfclEjNxZ3gAYIupz
pNhPwfD0QXdtZkbeSoz1njaMY7LrUqUMqXV0p76MCrs+Zvda4uumGsJM5SnVyu3R
/Nku3WRG+9PwcR79Aihk6v4K4Lfxy96lV9OnfIM/mIc8quMBBryge2WDNyAIvQ+C
Rdp4PBQ4tyMDETXKNCCLR7jX4SaaxU95LuPWaFFEtYbXrLz/yiRIaPXzA2aF4LkW
B2iMTNoRKt4/2WcBv6M5B0QNjVyuxuFA1j0FSXFnYElxCsOH6SMNoUtrSeeaI0Ky
3q4GxthonbbQJ/YaSfUwG7RuVLOxgQoH4mkAcs8G4jiVZwwSasvEPz9RbKUCL50W
clQGoLvN/qSCQkC2X74KIoNzllIEx6sCaj0uLmSQacEOLToC1kQBGhbBclmu/qTX
S7ltVZzVCSO4ZnsgZV5uDqjtt5BYWnkfApyk39ZBvCsV/TasPGzPD1j7WlrJktG6
pqaX46B5WxyBB3PK1jAHO+nRPabPUr+TALLc7sYLvrilh7AYr/viUnSdaVOygug9
TQBDbEGlnZWHJiJJUPjIf1ktFFApDJ+wLeAEdKZ47FcvZBJrNF33iSTSsJc08xfN
Vk2k/kzEMhJgRjAJ1w6tfn/n3+OTTamlF/RBe0LaLLgFjz4eWGRnOxg83eIfKe8T
meQe7YQnxRCUbSCVZ2gXIqGJUzuBKWP8U4d+q9fjnBt6sriibgDz87l7blzyQi3S
TRLoFe1NB5ifyjyxDpFxmEY2BWKC1FK0NGQY1ma1a+KQPKuwwvmKzhrd3dxkR77L
J8aod39cifaefdcM5IQ+G5j/delKTThEAXo6IKJaCTw6CAwQ6QCV7LMFK1UHAPev
U2TNtwp8I9o7xKkRI9XAEzuGOIAFL3b18hSBuEhzRAhgITqw6D/LT3KXgmIAuWqH
D7ZA4LZ+ZgwI9h624BtpQCRqbNmAx0LVkbwH/DMYnGAnXI8ra1XhtXcmxeqAqOLL
c9w74euQSeBQS0zem3X7Dffp4UsLb4A5WmvKKPeugEAXNjBuW2dCk1huVyqYaoY2
XsgxBL3s2hg0oEoAQwg6xKFdwjL2Q1ZNcRRgn6EAT/YhujH919meMzgg51qgOV25
xoyp3LJc+XWn68WaFjfTD40xRdYzglO69zl/PoLH2Pp6gW/GPz/ri2NgbWgcIaIz
23WyZ3Q3eU7zd6ka1lOEXzZpGt4TdyibJ/uOp0ka4xQkjYqY6oJAL1dbazjRmBlB
cLZ6+1h9IuYqJ/wIRZo3lnIUDogyolcz5/Gh+393JYcgh0kYPnLomjJwyjn9mq70
9UhxtZJR41yfL/ww8UtlblXzMYHX2rSG2JIB9bPTuVn3ID4t66hJJC8LVUtOF1+7
TuAY/8wrK6Qs8M47WqTW1EJ0di9NEfDYUxm+ONZMdXVE32eQz2NxDc/IRjZNQPO4
oKxd3B0hfNjXvt+NAuem6RGDwynJQVBc0oiH9gITe92tZoTkwrFC223sIjSelbZQ
uGQDY4reYWqcyKhmgxi3mRpkkjhgdnD/kDdDccIlNZBwgwkDfjZnXn/SKveArSNQ
r/DJjQODOVujjt7TCvHlokRtLk1jAO5+vV2qvHAmUQsCwsn0gCvn3+dCtyxbKMUX
nODaZSHZ2iVLLBM+VSM0AtRZzSNTFKXtmkdUPrZb25JTYZepuIgn7ahHwsI5CYP9
cA5bY5n/o8nU6FMkzM9HBbUDzrPqyaP4/nJu1GJGiLeP2gv0Zk43a6LvrzC9Ffgu
XzttAMpRQYqP/L1Q2F86r9pjhoLK4lnuSph16roUjMehM8KigMkIZ/bYMYfpqvHB
Rxgppri+MHHcxhRYcoO9Zrmy5baeZH6Nfh3CPR0Yk+BlkeiPIOjr5YT2iH2bgaIB
N9O937sjTAmzInoF0P4cuNkB1yG+8Thbh8LzME2FJ1WmDNXT37MS+7pKYp8hLX5s
tAkojjxGVwbNS7rq0TU8j2GXOzvbJGm2Tr9nsqHblriKh2vmOnNS/3+4m7+UvTkf
c5WyNiOCdPfecmLZgV7b4bGtnUtN0kgLm+xXddJRa+jzJxSqzb8IHPMLyf8NGuT1
gk0ny+z2XS8yry5M6X5384h524oH8jOzxelIFMSfzPbul5Dof+rGRl8Boyf1Myji
pnK2tXGlylPgvlFg71FT2UKlEMSCPems3lKRc52+B95lybIVWNzWAVtbyCwbc2cE
iLE3gHvSX4+ULA2XPg0zNVRdCwm67f6N4SIvz/9eVu7+3V7GSC8NTXJ6VRytqQ0J
ej6NA4YyVdvIG0XaM4V/1RjEruxsXYGOB1cb1rBDXj0lfJ9cY/VZkrevncDqr0an
uV3kNvtLvxQGA9GmE64QEOCNcLsjVfm2vbv8FARlXYMb3t1zp2z22DRMg2z/pqKF
d/GpabFWNWDiZNtkh3V5xvlN9t6DsfKJB5I9VXSONMFg3rhd30y+5rUUPgZFwkif
KgoQvUnf7SU41zf3vgRwYVqgJJNYDvwcReI/2cO2kNI8bXwxWwCHU8eiZMllLasn
gKEecKEPw+f7LXvnb2AjyBMoDXU1FGQnhAwAKc8HhFkRW+4b0QEW9NYTVgrWVZVQ
kH7YBXs+72Xs7PG7rbB+bfGzCk7ELvJzvVCIE1Xbggm56Tx3Gt40eLuxdv63sSYn
2FvXhCoPOH40rhRIwGEwQXgE7WyyPxilC5kY9+1DZ00t5ZgIBdfuQGeDzL8vHYU5
orOkL/6YrHCVotlsYyb7njRGBz0U1DnBSF1y8AI3A1RLqo5RF8KIa+xPEHSW5vW3
/neFGz5ILaL844zvSaa87Iu0v2i8sxORPI5OKZnOtqLCGrLVPCeVeL7ZrKxUfrIi
XJhN3/vqFjcYDpYO1cU3bxf2jS5SXoE0RzC1UrR5WoB+6H78nDYphl4xSFXFuaw+
zGXv8F16zj8iS8qrLF7eKsL/zDRZNOl5y+7Si18x47Vuuck/0hO7XJgrDbobUk8Y
TqLXOs8O+t/kDmTBPiQZZRughryEFHh7Y3BX114MEMcumUYdzzzQ2KlfI9FY5x5T
NUfpsVi/pVo8kfc52p4/7z4iHDL6fl8MQm5wd+8kUxu/WYHz1k2oSdxIXjI1WczK
+chzN/jBXpRqg91rc522QN1akqrb/dYQxFHziedOtHYA+5MvhtTx8ZuLewYuP5Yd
cN2z/YiZSuyyWSXbOaxXkvEWCA0tim5qCB2dYSl02oD2yFMMYNLUAzI9qjcktlkL
qvnVZ7f4W2OvsdQjM0yOgtRlktS3k77oS+JbA0UuutUeD6BxDT6M78dStjPPAGv8
wuPO+VImMQXd0pVRQiaz5vsRPZ9t5Dsr8p2pRhfLvDUIOb5AWjHWYE+vIud0dx9M
Av7zX7drfX6+OznN6aHcEskuoAAuvnAPmxgMtHIYQe7YTnpdZ1LGNFEnLtbvW8xE
UeefI/0aQPS0pvOTcO0+Sg2P+zJWKwJHSHwSWIKtT6Uq+mpcM0zFAr2CyjHAhMXm
i9atZ36m74DfnVP93URU70qjiX/mXuC30Bd64rfJbdBUC7BOhuWOu5hHiMkk2rSD
KRmfyaGOQ35mDl31JWWDBR3DSqaC3mbUReX/naMRIGdZRcD+gJDFRJ0oXJnuD+mq
bjYRP0g2+8cmEY5CsnTIoyDIL/qr60RmF+EWTW0ACY0sk51t19/vrtnXX1S6xV5L
Hc+Mplh9ERLQOwV1ti8pAw4GP2dC6iJZibWD3+3/sbSC3cNU0jOX7ICUr0OdF3Sh
2+MIX3EiP9x8fCldC07Hcv0qnnTTat3FMwX1XBfkAxpWIKaglkNdr750vIq3f+f0
ctyxX7ublaguY4tvAK1e+jqA3iBKuSNBI4y3ZutSPX9ikRupK7IUvniYGktHH8t5
H++w53BS81SCmCfazOncikmubxXg2ZbTahZXcn3cyaNbXxurO8sVrgmoOM6RbW99
Z5GfX3ujqdBW9ClRZGUEHR34wyupUcChzq+BWTu8KzRQwzUo82/N2E/PbpqUj6uG
b5FE/VhoV9WHRfs8rvrEmH9rNQz/XH55clkuTvgnRm3TFvF2Dq/0oEPslBrMbccF
CNn4Px75bhngoGFoKSCHjQmqjWAkwLpPDC/q6LZBCUnjHN4oMELCJ35IH3Op6nvE
VLBe3Jx9SLsM4hbZkGCi/v803M882hlIXUE7eMBsLJjJWWC3yl1B5Jg8Jus8FoyT
y4kzCtwNPiIXSEWnQMNOBfMbXwxv7cHu/3y0C55AWQdvgG5SwCkPAYGGQGWDCwdW
46U4okLtOvZ2yJRXrtL7v1rTULcY7Hti6ZDduk3A1fNkmTjOspMK8hkcWej+Po9T
rVj73DUPrU+HRBBPwr7oayGq/CIOBPQ10vnFnusToBThKWBBFjL4kuZB5dP98WoF
KkjzS0FUG0Fx+glMCbvI+Paux2KqVRPJjCou56XPN90LZHKqvidyfwcU/aYLjG30
9zashlBcey3cIWI1EhDwlO0RHL4KzC78ZRaV2yjVJ9v2nN6xhb7vr1yos9oDXiec
x3uRF5LPz6+sKeY53bnfFZoJTP8ZtqlM6u54NB37u9+Pt31Ay2d2AhBBi0tDeDP6
apMvWdQilEW13oLolU4RvR0AnfZtD5vMVQZLrWAHLvI9Ikt+mX3QuyeX9XTExgJM
qv6Sf+F5GDVI6iX7kkubw3IUD3JqB0Eg1Lx3OEg4A66rH4I7HymXKrbw4UBl8bPq
U09mhaFMufoeXlUcw2WdX7J9Gwe6RYG4Kxq/WDZ5eDftPpbSSrw/9SCz4b8aF9zY
uNjSopXaMBPg9FM5T8hCUvnIGTjfu+N1uIUCSXrrW15qrqdexWjclJdsijmxcOPU
L+tVjwUJp6Iu7yQ18Qg+xXKOz2ZmBreuNPB33FQSRMxiswYqJhHIhGCnjsIpfsNG
o3Uej1ZnBAY6OoDFPLgVxUh8S8LlG2Dq1wrs4eE/lwE4SVxLeno82cqbA9xDC/yT
rb6Muy0zvrfagkgR8CfS1zNzGFrEBhRrRrbsDRJerwRpa7ouRZpxLvacjdePdobL
j62k8/G+7KbUFGxbiDsdILzayfMrueGRujFA2scQUB3hrsRxrCeARxh07dzGlPzX
CdaygQzwmY5U6x9QP82moMjMBnXcU3bSHrUuMVk+PyPtQM2hUVPYZl3lSp4zfjw7
MSrAbz9hB0IlWz7UcfEsZm44ZJYszuGyHya1GrWGy13P9MQona/76gAVyBokVjo4
EZj57+G1dq6433ntYPncEu4vinHK11kQ2eEcCUAMviFmJr1hpdJKgbMKEVb+Lchm
OtSVi7sxUMc0zoh03QUYvxNIBSY+nffsNaRDrleCXO5vrXXqMIDa90NMwDYQp161
WVRmJsw2NqG8206wIaRZm5NzXK09xRCWg2idLn6BGQ23kCGJvNlMQkIlK1GPCAwz
q7zS2XOKm+ziolSEAhEZb8gagwEHM133L40d/6cN11pa70ABQ/GBax0ZH6fBQ41d
T1ZIlAU0Js8VskqLwiOMTrAyCEs9bpnp43nGgiYTYQ+VU3JAKsNruWmmrzYlBc02
ZFbgZYItfia5416hSI+TDd66iaNBoJwjyMpHOGBzSVIoPERP4nW5ZOciliaQAbCe
j2P8LmEJu5IFHT+vSlOIjGnyyekvigX45rgkrnNlI3g8rxMGqa14fi4PnsyXg0R+
5Bm+gpGqpnGzvDjkC74BfybOePlRKjExtMk0ybubBzQPLaGNS+0Pvnq9Gr470OVj
2DIJ4PZU65OWIN/8xHCipHvBP95bED/dmaEfL0QZbmcFq/SgudBayweYVjaumUms
VYYo8gxQdkoplat9UJnZxFG+ykjuYpsOtcUo87TkR98tm3G6OdmEZoQKvP+4WslZ
CtF6Bc4ywok93G+ZNJPC8nR8mt20b/M9nahC+7ncCkmn78ajL1LynGa5WuXmzj+R
9kWIpvzHAGlZNaQwKHcWYbAZh3auDMjuo2OY92sacPfuLpzrebkUih+EZU51RrHE
9mBMazuE7m3RBdFG0lnYq1UC8CZ2BSPTHoAtguIf8MENHJSCh2FrVkAkpMSzLFAo
ujFIDRlE8UEgofwmMw8c+h1iSctaZaRZNFw9BcG3+iMcbOa3liNpWmu88sXoSf5w
Pl6VXS8gitcxQe2fGM77p2jlw/stIMZEX0+ga930H1cW6ZrwpFUXjKyddNmKmmeb
08Y84BWkTQYrPvVBgZfovxBLRFIoAJmOe3DZ7lHs/TiWxdONsnoh2xuy2D4DItgp
QsCjDgk547TYL/75v3c8aKxWQ5ThGoITLQGWhpp/ZJk7DjjtGWq6l96LDywCnUyN
9G8ykVoJvIKseqszG2lpLzjr56qF3WqI7qxwRWL3UTAm8ZA6LzkK3F2Xvje+i3Mk
WfVQs9EySauyEu4xqDVYRihlLww3GH1BDR3f9c7dQRf8L6rr11qgfmWvXTTBBDjQ
gaQVBD0+eYE12L3qix55R4POqHHSWw3QAt3TJ3fmG6pnSR+outCmc6ADXtPtXxlQ
KDLPGS/i2mHa8v81zGoGd58i6ZF4wy63cBuq2ceNH1J/4DyvCqJxW0nO1Usip21x
+qGlJlL1/IU12WLM1CnilM4FcDfov6m93XMoab6HHWwvnleVYpqnm4T5eIkYWYbK
ARnoStLjMmWc0o7Rwv6LAadA0s9ZYbcvbmvUNrRuZJfiTg4jrFn6ji3EvSKMlomM
G7dycc/EtWsk7ODjRaW0hqEb4Jo7IQYBDMBwwAB+Tbg1bENENHtButMORqENO4c4
+nsZIvNK78pDADoHmnC3eOfAix60U75Q72BgHvDgNPJzHW1yhYitcHGxYjRbpzSF
4rxmGdcXz6VCAJ5WsBZJJhhua9XBnSpVHQW0AMRAY9A9fe0Wmye2tm3GNpBjfpuR
5aJ7YlkxhHYg76oJB1GxFMUUVkg/8fUL4jEkv3XkvPQmCkld8JL0Re9aOSPbGAF9
8SdbfI5kiWHaV24aafIi2Tk4M87V8M87ofSLktG9cjVIBeFootnL9iY+JgsfoAah
yYXpr5fXcCmucrtE4DuawB5cVzvAnSmFJv/ZPWKnwJuPH3pfZtl3w5yG2UG6QPMP
+OQ3+mH5l5qIPCKSoM3DCuMosDW9KSnXIW7WPLr9pwI53yl+ckMV/gL6gjb6EFiD
zsPxHPqLFjJAYTJQ3oCcBt6yCZEwH4SNx64i57pcEpszC7qPk6nFha1EhxbQnvG0
XmW85W3O/zpAMpf19qUrEFJTRkj25bYh2F88b8QysBtN98pmb5ri87ZMEu/ueCOE
6rRo6Wt6E0ga9NokicsE9l2RiFdnflGgGTBObtweiJ+20sSpP4FFiBgbw0tLubW/
M2S42vfZNPN2AvFxD+9b92vn6CvBIhQk3A6OeatzkgoaU+K+VMXJIaF4U7tyxcp4
Rn9Gtavldi1yKCCPlW5XBePxWaqdnPxAdEpPRfRPg10ufcwOsH67Do26xAZa4CKY
7T4AUYJBc+iUYTjOx4WOX4F5+UxgZI1S/KLzbvkgjLRrN2CUGLgAQ3aSIG6MsQ8h
ZWgq0q8WHLuE3+QvP+IzJ9zoHEYnEJU8mWYJRMJqgjXCq50jVEug2JOwGi2+GR+1
KYKDOhGUOMSUZAKfvNWy2dagatSgVMvfRao7uULPNfz9JYMIdXw3iGFjJBLjKjOg
NBvinwGOW2qhi9NhEYT6jrRJNmzUU/hL8ksoRNYrHF3hIjL6SyCyIlnciRxGDdHC
XCvuUaRAX83Xl1IXlGxDqEFphxLFEeFI1+yt89vaMaz5p40sdidAz9f/HN+Bxux+
GE80LyTE/jIWKpbfOAC8V1nSKuI3UzwW0wRdX5ykEEmXcj3j/uNYIoDW5aCSd4qw
504tGdY6MQXWAgZ8+P7WBGbPbfrtUUMhd3V5Uy/ygtBaa8AgFAbWcgF8RUR0MQC4
cW4qAu61dy78olMzKjmPp0YTnY4tsyx6DgV4FJfXEZkpgrSzu3hXTtoAMDaCpF8l
75dCbvBTnV5fnsXEjeKjLif0Xk1eWm21kbIJkpMtGg7y5hX7uNihYTzoMetmqCGC
2A9zTpInBGMqfvzhRpfW+44QOW5Z87z+37ET3H9LHQLcS1soIZNCQo1jtGKTZw2Y
mgPrC70UApwmXrQzb4+j0NwbpWrZB4jrGz6/idSjnASZAxiV+OVX+WCtC19RSNrx
eyLPmV+YkFOkCaumZUY51B5HR4Be7frni7EOojczeLTbIU8tWncEHu7/xWh52R+o
ZPf/wn2cXQ8/yXvplimzBDnYJYqpBxWQOx3bvc6UtGWVtdXpOdchbne8Sdai2Jas
GFKSLdX1/YAnsCBV1N93XqZTbGdiVy3ccNU5mFCRL/AN9O0PWoS9AIeYMlhfkukn
+XbUZQh3ZnBUOei7rLN/SovmRQfEdI5ojahhcuQvQDbxqpF91ZXNiCl1u4Y/PPbF
nYkKho1QQn5TfFICg7m4iCK5bLZu1YoFCgbfJVlvSpIamDnKaK0cwnY7mfEwqpI4
6qtXzGmTXGf2noryC4G/umDWcOGkKp9PtCgoZpjYZmRGelBlm0CWIVenDdsul/PX
L25ZqXAlhXOr65jx/vxGKcB7Lh4ThHVjYoDG0UpElQpCWRyHT48P8fzfKdb5v7CZ
XdxV9YG+Qub7IPclpuIHbPniWMvWNswpd3EKMuobh/8VrutHfmQ/vjA8+Y+0q1oA
weEmJk7yz1zq5vh2qlAZM7oKsbfrWsVLbtD//RUkO8a/MLcdTWQHKu6ntQHd+X13
cXAABhZ8cQxp8DiiDYQSi+qmppAsmTJv4Ks8YxxXoRMphQamxTjU05tzb6sfjVrp
hi5DDM19bZIOu3o1wjQsVxCBr73iErKxvbYe6BJm2xDqOmUKZwnev/lxrQbbzzAJ
hQIRUUot3oRpCyQkCygbDX0/DL/XLlQJdCurh6O56BnNJJ8JAMFCzbo+MgIBNhan
8Hw/gsowTv5Yn+LbJGCUY1sw8I9aZU1jTVSAB+cwgn96jDdRI4J2OFAG3aAAnlLt
YnWZJppKDplHKKmBTJhNJ2+YE9p3DZ80gVYJju45vVhE8w7M3yh7V32Lmm++fW4f
rICVQEvBGkVv3kjU8Hc3HT5+jIkVPra79NaPyqA1ZTW5SrswsK6UUUZnzPWMXE7k
GtAnV1cTBwtTRhJhzRZE/INicAiLdH5GwQctc3i3io1SPyrEFGsIx9kPNKZugdtF
caAYzbOEL1hH6gaRZB8aEEk4N5RiDU/YvxVBspoOSfG/ukQZ1MzQzXL+wub1cm4J
1mvYYYVu8uAq/eEo3dbpUv+bpFRBoZikjG6FTwvJMZLsh4ZM+infc2ttPwKnbNoL
K4wETVj7qMHuicjaRq2epslYTGJbHq7gkpmaXAtR9mySR2DH3xh83UmjE+M6J3VW
gTJBUGMd/6aBgmI+kRF6R4eoZEToPnxaBdQqxZ2hEJ8LOY5jetYIv9g0tqbqSJPK
3IlRr553geC/J89OLbCboqnszJak33o/VGB0F5fWhF6MvxBdXeWlz9iXy8H9EeB6
XrQb82cjDrbJUXgJlUYOcITDED5TLaGv06Y34zFPKj3y6WijxqiC4j65XnPUV62G
U9SNs4T9cRVBhgm350VJ5oSM1cFYG3INm8n0lQ+CG9m41Smjl3LBwFxgSxZMfgNj
5QNiHXqxZxqaaiCSYApUqFvFpRsVYyysL1Fuwx6bWqC1Lp8HY+1eywcmH+0dtz07
Moe7K8lZqyTFoaxL8I3Pbcr3evpqjDBbBTeDPQPunWFnE1AC2rz51EABg6UDQqhv
+i1AiGrLn+FNCHm+/d1L9bJmrK1DeeTf7hxE0vmXLIqdLY8QA48edtXkbZx6OEe8
rHav3Sld04jdKgYJ0k191WrUHL5Si+SPQhA67zhL1Q3PsE3fH5wiAcHZtG2Xsdoa
u84OnyqYaWS1ZAHurkwurreKKDCXd6oy6eVIlNHkl5/0ZY3eEM34b3ZAwzLyT7su
395MyWmQMJXNpJhjjN/tmY8/waEPBjrH+TusNVPkoQOsI6+KHqNU/E5m6+EHWiLW
d3Ld7dgBc+IMxg+b6Utfl72IcHxH/IFS5iKsEsY+pDPMxikgLJ6x8RKyIRVmuXs7
TxVReWCKsoWbtOQunMn+BcO2MIRMW3ZjqnJf5FtT/1SmJOdbM1eTe/GZ0txjhOBx
CW0LT4Unuz4rbFr33muLvKIgDFGDErfnkFMtO12/5zy4H0q70XoNvAtoN8qoZ+Dl
RHLCdvhzRqY6UmJ7L/NG76pfTEyHjGqfjlRdgkDpIUKxqfh0CgQOcMhdXRNVd8wp
swVvfdf4ROLpxtsczLG+/7rCbyPySM4Xj4Yqp+Kd34gatL0Ddw6wULSjQKobh1mV
br/XaEZ9aIJYs/bg8cELEURMs9MnB4XDx4LjRYxy8UizHzi3D1KJCu7vQmTt+G5h
Ld7BXv5u+VE4YIuX2ao2aDMe60EeCrln0rAmZUcud9dIdaxbHp6b55grQBRAZsdv
3AYGxnp44TuV3ydaIs+Dgh2ot2vZEj/qlDZwUvcPVI08yOaEZ6Di60lmvGL6VQJW
+gKE7YvViBU59FjUE8IVcMiXEJw8k+AIzmdRzjyTHIyZmW+KM0GUFgpsnEjxDGAq
lN+Tarf759MkDiVsEYYFEeu257rI7ZThfALu3shCVEvRc3a+nyTu6iRkr+z+jCrb
9dNrKuTOIOE4IT7zZEJN3EEVi5PXgEt6KI9nvA2XMlje677+8oN1koHMhxveg9KH
jYAsTzLnUqfLxcPreiqTbh0QFQf5vVCwrbaF6Ax2i0asGsCg9bOPmRM8XMXiEBt/
3DU74i03oPKIyFBF8kw5FKQdZzPK+k+2+HSCpcfWyIpt04KdnXO/j4GB1kg5MCFE
h6JnYlN9hhPImeGZ2EyQg3A5cr9hrlK3U2FVlpOcqIxtcoQcvVwxGanZdyLeaOBU
w7GINoL1f7Ob+Wszh0UNuVeuoFn3fn9kLg2ZBPWc4dAr2W61p61DUFJU+8dGdMWd
Fxz6m7vJlMmTwqo+P+yfsQveD3VVtcbPbvL0uPRODhs4G4EE/87INCDu0F/fn4/e
HB+tV1CMjBPyXe7VSJPwD7rrkJ19ygF97noTkGDRPeYedj/lKjYnovYDQfsUPr34
6671DdpnMxk+blE/KuZLwIy4DNwjooE++GQ4gJrOu4gaoSvcVDKgsuvTofyqtosJ
QR9TkhO9CDoPJvmXDYTactZ08OvXuCG9qj1YogqfWqHyETMKo8YmqW1DFJIMemXj
UgH8e8uPxc6I2g4g9p651qjtxfjppehJuJJQlg0AopWZche9KDxpC8aiYWkFQbP/
BeMFr3pve/YTJRf/+CCVyknQkdb0EwB6mzyA9PvjhhGJBiyOhYSk3cXWDNdKC0Ik
dJb+7wwu91odbY7InI2pPX8X7Cwdu0yLVRbR63O4DoFtQfGQYAKTdxqs1eHElh93
hG6VHTT6RNBd9EECBIbqaugbMenH9e1PtKKl6A8kLE4iOzI9IRwylSs+AufPippY
BFNOelfy+oXEWP6UGGEMgxipJ/kVPphaNKiz0fzyG+fhPI7TH7SeVQwLfOX/hHxp
XFzf8ug1Fyo8Yh6t0H1t26tbFl6nGGBNgeW4tGK+x5DJYWVmCTRktRqn7Ophe8lh
viDhrMDxqZZCosoE5cvWjVcHGdcLBFOmvhAOfoSHxG3usNKrz2gUuLxvIZJhSCDT
nIocnX9+cMXHzhMfy2Gs/UbWX7xQP75iMS51EbV6z9gUwxVj9S9UKqzl0M8NLfM6
QPTZosXPKjoV8IQ4vyjuWQ9tvwjr9eiqssXjXmSRxx93zUNIlG+CQCO7XduMOK2V
BGAU0+CHA137X/Rx2Rqp+5bDxXYNeswwuyrCm9G8ZcBUQ8M2R7BTjm+nskjptNpY
7i4J8aodlVBVRiwxZ7wY2NAU4fDRcsAEsC9ugdkFmxvt6ilIcr/C1Xj+rAfuTNga
Pgv6IKNq9eInPDkHtCDztDwRUgEUbL/xfVeZJ3e5WDB/SuZ3bi5+8eG1RjCOZM0c
bGTSqCPUxeTVlqk7w+gXJm+zBp5gkg8yEte2GXGOIN+ge76lm7P1nCBR5UnnimiM
6Eh42Y3naLc/3QkzTGeeQeCBXKxwWFd63eoVvU8QERziI5UE2reUL5+5HQDMJloW
lRfgcEFCf4k6WOPQx1RFNjzhpJ+ttaFhSzbXOFPpDnNZ2b2JOkljzge3xSE4Je1J
ljkqOY8xd0FC76heaYD27727F+8q1w1QPVArNmWavkZZQk5tTaH5PXP/C8t0vFU+
BoadwvdWZPL5iZIUATwTyOQcAqYMGTtz+U3t8f0MDHjkXXNUrjLrGx2u7FeAaRpK
73pBnp0vuSV8j5d4K2X7aYCgMa3IublzwJY6YL0o1X6kuDtt/YjqFnYjwLD6+rBt
YarM6SEnYh0J3BoRoh/ueYrRvzkzeUSuQMYVPUJzdoyFGy9sSsPdze6CWPZL4R8q
eETPWI/9fYh27+V3J2b11xUrgiZcuzlu6xuMyCGgYyIUYdN4/rPbx/hpUB7XAl0m
Ld7PIkS3vAO3lNileeR77JmNKeJ4urcRjQHdTGg9oMUhdhC94bvxLhzM/J320XyA
ElK46hxAOLQ726F52bAZOe+RV6CzusQGm4aysQYZjPcw3AcvAe9wObLGbPm/1hRm
rQuIaUvcTr5Zl5sio2xQqsN009x1J/r8N87ECJCW5UGmJaLweVes6EF9C0M8ellm
5NZKI+Zm9PDnS1YM9MxsWF9ncBSLHqu+4sQaqBos+aZmOjW3Gnpj2pSeFgPkNDFm
q1GbDScmzVz/+ZYzpfKjKIj35OpE9wkyvWDSvCcv7a/TSAdhDeizinYg2gR+wZsA
+rrh6KGK8mxuZjhpCXmOKcY55610Tszwlam+kyBKwNJGpw2PmC3qALmxJsnaKiRD
Si+VZFaFeHHlWWBURwtVWu4dfgAEE3PGPVQIOeKMM8aSzAvvrXWUUBx9gM7kV/VI
liAB9yYHY0KIpTVdIwLRGxQnY6f/C5aFD3FuvtvGQCZsQbD9EJsbSz/LRvgc/0JT
ZhAkUBt2DChN/uSyjlStQ/40oQgsyKaDf6b/rx/BoHng2sYOCQyqptQixZAKXJFM
rSbVuoEq+Ga8N2ZU1KX2b/InvSTbES55cnmrm2PDKu1VhAjoBcu58Zj+STDiuFva
EyalD+PsfANRRYs8bY+jicAEHZNSNCPX6WHczBZ5tvQESHqKgL1brKDRA9OCq03c
A+G0eTbfdeqYq2csFu9K+KQq4UtBNJH6d1f99ITyJ/ULabZ6rF1IWucfq7grhMEf
eMldlW46fDE2NABX87Fnu/vtfd4Yrxb5QAxkMIRtxE9YvwrSqjHW19lVxMt8HSA9
PfKpLmferKbOmaKwP9YjZa4Q6d3JUTeG/QLU3a41lBe7l6mPnOB11DdziDBVTOA4
4n2nD8P6IaJFKqhDUVNJlegiJ8hSzQ7AIcWuuujPtdpk6SZCJbyf/DhithK4AYUw
cdEKthwdUTCEAeT5mOFgTNmu6/9TxokhFkJolrWF0uYFj9yY4sLlVUtUkX81+R8s
zA5jNxfWHhEjpM9/zv3Beg/i4z9pRxLQLyVdVF3yIfpBP8sP/tcfIBu5oGyBIpVp
jAQQ3Tg6jlNWOR9SQe3hjmJx6gG7IdbmrVQh7lQVbPy/zcKD9LAYf86V+KMVs7nb
MqeNERbQcDZb3/M4qo3LR2n1jMDPfa1ePHPSEaTpPYnP/oZ9to1AhMgevdZNGVUB
RHp/UgM57T2XC6bJVan4lqsWEEG7eX5lCRioe1zKXSiNdEGwDAx6LBgODsh0kRHx
VVgTA3L/qOJm1tG0w5jUYwIQCaC+e66Ew+WMa08s71k+w2EbIq7p5+QMruths13m
c+8DBFmyvHQwW/IuCBPdV2E8WHPfPcMd8m/iD0A4o6goP0q7x7Bo+JCChutjDd36
PgVEyzyxRymBWmMDQKq6AaQMAk5wCn4qvXidiVZkeytWxEN+wH89BBpkgcmwT8LV
HmWOjehp8t8dvu04KpVwCgE7JWEJj1g0nBFE2LvwyqmlOTDiem2zFgZ7ZigtxrQt
oBb/XYkEd0YQMBAru9TjfDOs/mzDptWbmzO2LD/xDOKPz4jpy+AhRweOienrma/a
vZuVmQgsGKisH+CGtERI8VEmgDfCevokrcSh4if9n82NJC/cdU8CKwXBLgy3l/ON
AzVr6qANSaplxg28eIFXOuAiozeh0eW3Pn7JqQ2lVtrT7n0qINq0dMzFUHvE886O
lCGocgOTY5AfqAu48YWTjNF8F1vyIqw8yIPghalo2F8uUwojF0OZrUWKILVwyP+I
1yoFiRXnu00ZQlsi7QJ6zTR6HCQ05sovdIF3qppuo1dZCXQj9YKl+X/WF7Fw9F+8
u2okuuaqA1Fs3uVCRfbuhRndXLdjMv/1oZryOJD3VydIUBu9kBVBYXYeJafqj7Hc
gYU8qXdeacPWeZMv/M6NGd3rzXoiX4s4KwRFzgPemAuiVS8v7O2JKmQX9/mcGrhO
qXIIV+snnzuq4zx1448sxwTqrlzLUwNjnJSfmASf0F0t8M5403OTCFMkz6wJiB6V
gQLh1RXe3nXQTFsiMyDP5vFH/fCQUHFw/+sY8/07uwOh93L+4Lmu0HVa5nNgFWQH
AT5f/U5RD4F8l2JhV19eIi0/BoeACbU31Xzf4vM3YtHH7vqK/uGzCcq1ruBt2qXk
ScbuCmkkBs/wyXOqPtAVj+IIgKKjklYE2a0GqkdiU1zmCABP+lIP6o6eXSRM8ONr
t2pf1eVVZymXkOi3MwrFNEyxWSR+LGSyW6GTUOIsmgCddZkpXKTA0mW7dB83nN/e
kF+V97hwT57Z0+MHhimoUHkFGqQB2aqXq3Hcf87QpygBgoM1gTZ6o/265JDU+IQk
uz1ab6Q/DKNSECcSDzWFABAHqS8+VJjsa9EVYvFQCU9oYEGDUiVH56w07XwLQy4d
BAPPdI2+PpQsAlc9Y1zh0Ker41rp+EzJ9IZuLvMTBQUdVWFtS54XI9k7tLkubAvd
qn/ajw/C44DcUSBHC+Xef+psWExHO83UnMbzjQnHjZJw4r8/yZGJDpMDlWIZK736
bIsqLHQRRq0sOnjH+9SpA/IxilIgmTMCcy6LpInsmBtrZwP4g92bYFNZo33vJ+TE
H7azbpv1xNFclPbD4Go0jPkNvt3Y5CGVv2PoAosbFMWrIfOkTa5uUjxl7CXuK9Zp
JAWGC3Io7hnKnxcAq6tTB07rF0AHWYJnUQyN7gceRO3smmKqeCK0gaFEP1gGxZI3
zKFsRwGIPDXOP661T+0fCF8tBTDpy2oKSMnRHO0bMpr0G/cFhl9kWrv8EAJUSikv
uINDMcIvH8n8sGHWXvT2k6i4wFHTAfYDgerd/1F+1xrfidRgIYoP2pWdC3L2JZ3S
yds/Xe6pGT5q54BbhO4px8UJloxVE3rS0+abgdkhA0giuet0sN4Q3gtxU/CVSfqv
I7BreMhWKXlXIHRBtzJrGlmJw1Im0+OIDm4yk/KGu32RQie9b4p8+MQImc8y9xIN
clGWDfOt5ycGa7stx+XMzB+0BaOPVUO6ZMxRuafduRnNBFal2vKIOdYA+ihi+vnA
cx/MArnymG2hFil+aMGAeyDw66GvXx2Aq6QxDQC6yM08MSbYQi/SVWefPZ0iFB4B
ZgwlBtUDkXIFQJU0h24+FLQ7y5czuZpfLAtVrlDslis04yn3MwuweN1JJWR/SDBK
gQcFP1x45JiehH+9xpZ3GsGvj2Gq4TgwSlnhX1m5IfzVeU4xMMf8lHoQRajQL+bp
ErOQSIMBk4R00qJ4PDbBRautEjNSxpCq/4MSMSZexfQloXAk64dMlZFqpdFLwW0U
iDSllkuZiBxKHOez/ViDbAnWbhRi+fGjXFRlwpZbmW9egzods1SakSHJtubwmOK6
KggwAHggz2pyevkJQx7RRL5B+g+uZOCEIxM6dvZoa9jJXaonRHKGQsa7Hq469YoC
NCf+kBWtGJERE3Ey0NhEQ7Gm4dki8aPAviyvDhARTg7VLqN9RH5xN6TegMxkAwsI
1u+FgBPlkTFZ3seUum8lpmmpByT1Qu4gb5DpxXEa4FKzXxM+B1t+wjnmLV1rUJ1f
vOE72bLjzyizwFSLSWpD8fGyI//3nIRpwqCLJ8eLLMsBj7RvuzfJq2WDrzB8A5Yn
Lu7/rzWKVVK4vkOH1r3MpXgZwnoRvDZ1dJUEpenSZg+DhDlybfw99mDhiLsJR/Ym
JfUvEvt/vbMCARlncQrN4DNMuLbKH8pHfrSkXf7Qp7e9oTms0QKsCdoM+AbHsXTe
0RptdX85dV7qoUxoZw7gteTJcCPEEoKofYWlnsWZdK6dluNahidU+Pj2eOxwbRxJ
B102QUZv/DjqIRpy2U9HyeInhkOjL8CFQeYpRy5eMVfWPBSOBkHDlAzWFvTKlW1b
A0EKfpkyEd8Vtlu85GiWXCEP45/KsH1b6Ju5YFalVs7lpR2n1Idt+LPnUDoyKHPr
UoKtrJ+DIaGxasbAvAgw8Q163rfsh99NG6rrUCE1b11fROJgD7je7NLfOVI91Y6l
jI4cg6mNsW6B9OH7uibqA0PGTZ4sliky+N+MbOfp9uV9eF85R5LoXDhgWf32K985
9o7UMUrdthmxYvZlDHFtLp9JTtBfyHQMCQWZnnm2D4dIDeDCXPLbME4Zpkq9fw2r
UCoN1GItU9o/aA6sH9VgnTxFK3YrmNWQ1yg2eZfo7F8pqhztvPBhWYDBMcT37Bby
affdLKLH2FLzOYdN7unTvbQGvq/7++A0snGm8AGR8Vc+e/F1gLc+ZysmS3av8fBc
sWkjP92UunYCzOsoOIG4dR9uOZTaD9bI98yb+RsRcQxib7byDRR/q7Mug7QoAK+0
3S7/UuJLs+KxRq0RjVgB2DImu73wLbJuUT24WVJoTaFbCT34O42rHzrFgzGu2aQ6
rFI3qiKjqfn1MAWc6hDoi09PyGz9QSepVKDJ8fQ1sox+ZDZ6WrD6kMl8kJxijA2R
t0GaGUBn5sVMFvivehK2kNR/Mdx5cqGTydY77HhH5G6u1ePg7aZXZymjbTiwyhLn
E1TzICJ7h1timi6SgsSLuObPPJUQJiufG8B3U8NgJGE41M0IDvhoFr0YmcGi9PQq
8OKoC8eNv1QiU65BLviHBsVKkrBTi9e/+PqHD6d09c0g8iai41PKUixnTagNTauQ
5+XGDuRgopgD4k1bNFd5wNE1zk4NRyyLn3XXWV2yN32f55fZU2RdZqv4EaCOYt/F
IgJCzdO5h07mVE8uBxHz2k35+1PgEw2SpNv0aleClvsJLTT6AbOuYKMp430M6ab6
3bdBwf98R+aztkEy/H77XSICvG7CaStS4DbasCLZnTYYO6c5Ax8MB0XUYK3nPhN4
oTAatNgrJOBNQLR0kVksw6RglLzlxVaxgbYIQ8m+NSRstc+rolNDUodXKqvvACat
eMZHt1qO8EqPKprCj7MCgOZgE3qEpsnVFahKKcok3OqBeFNF6jE7PRp6ZQugZnXu
Cag0MfY581Qp1KdnyvshRVxkE1GtRKiScE5J9OsT+lfExwKeyNjGB6X997FlYPIJ
/ZrIYKf6VFbQRT0q/uIT69HUQ2iETC0oGGZrEG0L3QOztY2N6p5ZhOJJqaaygf8a
5FvB3AYl3JluO/1ur3vIBFMJf3+oEcXxXdC9zapUoFN69gn/LH5lJBjd0Z0BBL5l
BnM3QZuzdSmHHRAUskI9QD1swP+2aM7mkeIEhknMuVF0G8TvJsZYQy3Va8hDuBls
+FVBS2o29ikUA3aRLIQzywLQCCFIE+6TLxKNOwOnknP/GmhhlL9q0xgGP4UHxrxi
n/1vFoxXUxXYA9ERVoZy7AS2VBNlUxVFf3GqGAIHjczI9UUNliXKk950Dz67a3Jr
FOFiZkCuR3b1YjJb5+4lZj+B+Ippyd+OoiMuD3Vfg+W1noKe7HFBK/cCfsds6Sha
zSBKR6XN8QAnPm0Y3ZYwUvmffUQ53h/bY0d/lU9rYAVUCHJDxBr4++EFOIg0kAFy
kVfM7/56Q1ubbEXzS2ZiKHdSXGRJARSXxx4yDb95C9QyVCRXokuwaKJVnXTERFne
59ABTB3aGtTYFjW3MuaGQmLTnITebZYXc4oOdlSHVz5VYeIoUyWl5Ltn6BeLtZRw
/MNydwTJ9tAheP7vBt4z3w/6g6Bg72+4I1/9k8ojyAWC83cxqmV0SbRWSfkV9aoV
FsH1rZ6IHpNnV1J+xCovWC8ZIODBIUDmXtsPg5VV7osxs8W7zx4ANo5VthOi8DDM
Pm7+DfQ2+Or/rGKBYQZOW/5ls30+KNhfFCUzv5+ZnQ6e9sokfpkydNK6KevTQ6mA
hdBhE8z8eaLmvR67mcGVF1gobPInutGly4z8oZezbjTqP8h6kGfA6gcHaGV/CHB/
twArqryVw4M9KrPJIaKl2gulVhUgdlnpwqhKA3JVCRLO5SfD9VcTZQvFUGdVfUoO
lFHevxOSDdc/IIGnBxEopMA8QslmkVLxT47z8V9vIfIGwsDIIGEc94ZnhyeeXCM0
f0rE2X5XdLB3qTSZvcm7UBGXt+/FdNZUZFNxGnf9+ZtKQ5SWyShjXcXJh8YEhLEZ
vWZvHIlPhOL8FntV5ASGi2rzdP69UaX+bWc1cKg/oix2pXdObe0PWlUalXwQciEJ
kmHhuumq4PZTGAQD4LG3sF+EkenFBxlqtTR6dkqt4rWiJ40J/tk17eGU1nrDcxQ9
UVFYeR4wKrgSqugvwHRPMpNrOFTZSW50Ipx87cZdRNe6YB5f1/C14Uob2ML/kqo0
3r7TW1A0eRthJ0SKdqVxovzulyizki9KMe4IeRZDyx5XjKEEnA/SnNNw8p8cnVQN
CtaoD3a1FgjImoHEBayHv0lt+H4dl6Rlo0EadqtM5xP3JNiIhBoDwXHUlOR5um69
QU2sQuDe10w0g1IW425RTSkU88v1A8ilQoFBuUjaQtPgX6y2RRU1tj2y866M4M40
E3VaDlxkqUWxu4NZkc78x4NMwA2Xbt4cxDIxpwdeIdvXd04VJrhMdxJZafZTaRvo
4Ta63Bda2hO4H12jouvmyeR5t1vgmAJ0xOaxSLmmLT1xvRIMVn2GhoVBvI38zooo
oHlxEmGNVZwFb/rI2o+L9VIedW/v714nRx5pLyi0GjwgWv5ZOG2W5siiEM6qlLo8
urQ2V7KBPJs9+LprKafMiTXN7g4YiLfKf2+4CPS8+0K+3+YXHyniwxK0htqZs9KB
axNW9LKvXrMz3KWjgKWkA6njv8wtxxo/gAfSPBvtM0lZT+WveqH+9eafwg92bvHk
smo7/d0e84QH/GiRI/pcbeH0GyW6XtSUR1ggkmRPdRVFOsXR0TrhEwspdZUbMD1o
rv8pSBGj7iSW2XW0dV/qQnVB+NkF+JfXFZkwmEFP9sAIr6qn310u9ncjMtFq3KFZ
m/IQvmUhk4/kivPh5KmneA5vvtYQYjpjZgK9cscx3kc/HUtBpWa28ZJZz1jpeyIW
STXfmpFclpNotSm9Rgy3tc29LnOBA0LPeatXN+gYCIgvApQ7uTbuyR8v8YJNJ56c
XH1kKHt73ikLVXm13FP0C90KcTZzo6fXmLnp3xmHjtd3XLWljsAHPUQMf5M3OLrW
cT1gVZfAW2wqxSvZn0VakiC4+0nWjOY4luZVxYzOtqQqJoC5vYxef5iki1RPPcF5
9g/eQtYGuzAo3551V+09yM4L/vu5T0GaFRyGcLaEYKIlchieAS/BKU0AVMBpmQQN
wWiJcjP7tfPTOa01i1AbxDOoqOJny7sT87073LGsch0n7R1Ts0z85riF0mSXlKnq
c+BN8xRI/EzIkpxp08n6IsTnCdIPKspd6UYdoX4WEHxIOBs8+Lxo3k/I3GdtoM9L
agPTwTNqblyEdzck9tn18QRH37qrmPrvNB6fyaVS8j3c7mVrTIZObliH1pjHLgqV
bmQ3+lPX0qlIukXYooG28eBg7bhVGK+KXacDxHIwLzmse7+670YJCVYmLNTIvSh4
2rsPGqxHR/rzya9/HKQi8IBOgZ3J6AigWpExRcwkwPGdlghR8L3dJeJ9R55THwb2
Canfe+XaTMpmlovhkKqlRLxV8yVTG8/Rtx5Oki8mqQkT9i7KfgNLNavrD311HqcX
wOQPZQagtKONABhFblTpDItOuXj0sICJpUnyz7Twfr0PsPf8u7xDwkMPGNCSVUwx
6IU0USM14snsyp1OX9aY/Em7KtzJIP8neTQOmnMPL+smVjv+ScN9zadfmA1hVqAE
nogImxFOkPu//98/pwBZp5AS9I6fPY8y/J3WbiqigpwyzXNiRiohBZa4HEFgBeGi
MCzCOIdayBePL91dfFv2nrVgf4N19MCLpyN8lxtDFNBinWrrukTandj5Yb/7ipbt
AF/02uQyC8ulOokiTEAoNp4ku9yG5uaNyNo1xp8lUph98tEDqkmXTs/FH9LYOw6A
DNOLXwUjbABdQeJ8g4iZOHDUTMnUb9b4ueejn7pVJufofSmQ8QzhQMsZFaSFjrvf
o546ODpPIcKtaxz4XrxkD3bB5zpJQA+BcdwTwzq5zJD5Dp+VFv/XkmASKkr8QtLx
VsC9CxaNIzX5zXoFRMlCtYFCUhwqUtxN0HjVCPjP8jR2v2d6+zkB8RXAvIotI7rz
qhaJsXuKa/QsdEbmZlwAjAxoasIrHc8G8R/6UuYIJvbRHPKOCmaqikykoK+945hZ
hKoCkEaANZQxrhblhgpQxSvXHeWIeM8T39Gs92hD5QXKkBxbtp9IrYbmBYprYbCA
vV1QHty9J6lsl09iWP/iU8Gk50Pr5k9W9MwcduSwPoGrGkMz6q9+KP0CwDzVG1VB
qTJFL3MfwHjIiJA8WVSV0uhFVKpRgI1Y1stHtvBhVPBC79WYHrStnSCser5T7khX
XRjKjl5jhvi8U6457sjS+Tl54JMMMyEVOLTv9Pa8BdNTqsH4tLDcyM3DDYqEc6Oa
Yx4YXmkFk2MOn/PawS4Y4H85K70Ob+Hy9G7lTBBVldPb40W/CZdWNzQWtRVzqtXF
VI5b1KO7uMGdiZ2289wzrbzu93S2ILrbb7HPkS2NnljlOttfqykrqQTb/Q2kiR0t
zA33/xLkTLLybi5wI3aKSiW6IUBQXOSZXPaxu7Y8Uegb44LjIoIfUbG/4ItEpA7I
LaI9wPzBkevG0B0Bu7x/l5ZAVhuXqmjJvZ1gl/pMlwXHXxnoKI7V3dm/RC1IZ5QC
m2MJZEt16p+p9We60JuXPlARVihZ7WGlXw4gM6Yl+upT8E2HUGR1QIUU7XPHxDr9
LZaZnMzicR6NcXultBX1DyM2+MmCAby7yooFetdcvntjGT+krTn5mrvooQW7lgQ7
lFNrebgH9DGTri4UFL9WJrC34f8Yypb7xdZ62h6H1lmHKQvRgpdKduPyRpn9hAph
dYuxEJaOOlEsNkJJBg4h2t00YySiJxWO7xwIR0sA1Vdh+qCTqqF9D/V13h5dasv8
3ymRjRpqZLgmmLzQe3/AvygDN9fWkP1I/FNVli2/+GIVXfAlxifYNnB1GajL/m/M
w6dLANg/sbwFaO0VGH/j67W6Lz4tkw30DYP4EGSI6f9x9Hq7phmTG112jazl5oaJ
Gp3TktunaK9rh8OFT8noZ7z0csJ4w4LOl0hVf7HL7y9HhAOphj3iBgLhjvKlOc17
HuG3itmYMebh68/ek51y/EiiF28n8sSn6Zm1CzMlm4lidV9BegJ2hLF6aaGKIdNY
uISRUf1P8aBXMVw695Qz1U0MFNq98saCnML6pi7VFSvLoQ1IoRLRVCRv4vpHw8W3
Uan0I506mt+NWnQ3TomKRdBWhmbso4mabKxDsUQbKnRmykCNv98N6/a+l8LahzN6
ayh540hiALO/HPbjp+XURQERKXzBoqSYmiBHuzASxKf5dviJUBNpmmAJ6tWLjYEB
X4ZgcCOHids8+Gsj8uqnCm56oToKVtrUJoMjqbmUyXQCTyNi9ZDYMgAo9x1M2jEY
8CeiGMgRV0ZTvpFmERYnkDwA/Fr7CT6BirqwvnVK6IABXdlvwT727AvFVPtm82G7
jMnLWxQWA20N4ZHpMBBtmWBupWHTqBW9KYzvqscs/50DQLZNn3WHvI47JaGf5o1v
iffDan/h3YMhn6R5sbVzpykirPzgtp5/nuplzHtI/lP+CyGypefqmDUOKUnD25MP
5RsaNzuCQHvIKztKzh0oJwgBnXbkYQte3iVWikqq6G9U2wN/EwFxyLr4Z9KhC13I
HBOB4CJh1zSWebLobJcV49M+KTkFAMeL9WRAPxslPADW8G+NqNS0GbZHKHGZ3ZM5
jVIl3m/w0GJ3yad3DIWEUJEOmgcxhO9yazmrVuNPmLRdPZUzSetC8ostRp0vVFKQ
7VgP4dYYFZsmOeTWikPex/SA40uOAzd/nv6LPNzPk1e+HMAZh+89w0+vnOyfE/cU
87vTIe1+C6/3RCjPF7Xb9rTgDrQ80SdD7IBoE7xcTOHiYd4uNqqaaL4o2y+uxta7
kCBFP5hvHACxfI+1pJJMspri2pmEZKs1f4zM4LUQnhzdU/Du1fP+SzPY5/ss8JOn
S9OHBo8hhgdhmSciXPFpiFMgcIlQ+ScZfEM+sp4NiYoafPo6YRbs5AfjQATfWWjc
vlqMjgG5/MeOyVa9kYJvtNwo/cJq9Omu+K5VTcqd4AXpXdQoESQaNNASUD9SkVpj
6DxVYVnf8Bos1YDlnZ9G/nDBiORZ63SpSjUMKGVelMCp51DLKqeJI6aH6ZadS+aX
Lkb3wE/vxNVpB7FNN1gv091FosD2clDC5x9sRtaP6EqBZFXawrbxGE8PSebfKdK2
eGgQOHTT1oNAkVsOzRaeCk7eYdiN8ExOjy//XeaefizrD9dMUOq0PalBkFK0WY74
xZ19sHwr4h88H2TsmSE9PMUWfhEQxzjeLnTFyQU+FkHMoFRjJP8C76hKigk0FrOg
8CGf7g2vxk/ZDjiF2oE88fnyMckWp60Wj7E8t7VsTmUwb2kOnuODxXprtqF6W02f
PLc+A2Qv6pWYfLvY52FUFMUvwVobZIg45eKFg29zL4FnMJfzKnKwCrXl19PVuOS0
pjgOfpD4Y+Nss1HQhCp+4hd/usrzCkPG1NZ3IJVy1zysNpWx3CxnMlTVdi8EHyPy
A3dAPUB9QeASrH9xC2gdrZLlSdf3we3Qy1MZAoiaOI31QmppErHt1/mpDL/ySAf0
ELViutcMOQXVVmZjgs69tRZ3TB4g+T3RfvQ89usjgPrwYiRKcpzyhhVszzgbWG+W
XFbiiO6OykkcKRVk4tSUsXeZT486mXYwosQqzn0gayuAIc58coFvh0SKA7rDqrgV
cEy3BVsnyMwI/6hTlFeEC0Vy4qnFjDSnV/XgzcqfcnTrkmQSyTxnALl97T7kfy0T
LMWSf9rnyNgYzETpYyvu1tPAsoocWs8vpUEBmRFoc2dhzwD/vgimydv+32YstFns
vd4Ff0omTWM1qwfZOajgmN1z/M8qqmI/EN0sBdb7RRSkDgpPuR0cIO30JqfgA/Eb
5tOTQ7u0OGjtd7rdSY8mE5zwFCPl1cpmTrToiXHF4SSTPuKXPo82g+fNmvAwvnZg
Z7IsMD7F97V6PsWS8QHjBmcuBl3Q6n8xnv6zEZJiWFsrT1vTosicsttOkjJp7jxy
Pmd8nTroYTIgSbe6imSq4OvsFezjY3oFIx34lsiLaV0EfN+44nBN6TkFnoqfAz7M
jAbQCj1Aid0y/3xgCf0lXoVBFTHnc1MNark/tx11w58=
--pragma protect end_data_block
--pragma protect digest_block
JomIbKCSx+7veWI2UW1LBVe3i1U=
--pragma protect end_digest_block
--pragma protect end_protected
