-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
POBs7UbpOzLjfkSPb7Q/VyUk+X3ttcEMFVPK2zCGYgi//prdTYI49QnciTg6Kx25
bGfRItJtf328mT287riMNf+fUvGUYrg3ReQqdzpluprEHLhHArLMzBi6Mi0hvSUp
UvfhCqALvlVH71HLEeBUvYVRI8cdSCukoqJJKfjr5oVp4x1cUlowaQ==
--pragma protect end_key_block
--pragma protect digest_block
qVSyvCf9MeAl0mUmqc4rUHefloI=
--pragma protect end_digest_block
--pragma protect data_block
5xjDSGEb3Bgs9UkKm3wq1DaDrQVeuFw2nttHUtEe4IDxp5t7b8NDrMgpZ4i9cHsd
2LuSLO1V2QLVVRjB5/j+0wRKQoq/be3n54Ehds2+TAi7HRbK7ITPsq869z6/gz95
gCrOdjJQHf0yfSnazut0N5eGYpFJuJ5R08oQ4YcQWwXHfoizcXa/1H/zGbON5Kuw
YUEMd55qA2fu8nK9Wula3zLfofEO7B107g4wM14gquEKRG2W2HJyQ0OVW4gdnlm2
4UH/WtfJ1LVpYuzvQ/xVs3Z6fm2xSykila+ihE+nRkRcXP9k1D9bglEewlX61iru
Baxs5XXG+uS8h3FUJdHash9KMe9v7Cw+zJ9OVLZxKg5sI//Z2RPadZ7L810GJe4p
zgVH+/SugC9YQbYaaqWN9VtmqoMV7oNPIB7kKlyazGLOWeNS3l+r0ghcDuhNOEVH
w42QmMdFj9leTTzJOXoShZlNT7UyhmEpTYt1KCnV+zFC+R7gsfL9YBjCV8t95T7p
HjnzkumHMYr2fnMWGy19I+XyisVahjC+fnO52y9Xstgu8Sa8E6EWwYuDd4EAiym0
ABXrn/lLxxTQcT44C6m0H+C88HoZ55DX133BdBtzugRqLOjpnA4dI5b3gIUGU7Zt
vbbxcNgVRNRlTjpj3regX8S8U6/b3LP5R1Jl0UexQ3Rso91crFLolSFLzaENmm9z
RdH8zC0uqUa/P/hhbJU+xSDjnT+ktQx1TxaCEoA2tzDP/JmcCaLTJh38tuqtoQz4
KQxDTPANfxt+LKSEKFpgx1JtJ3anmFnQrPV0ShFKf5VpbpUU90g03Eghoxa2ejXw
ixkX0rym7LDphIhAn1N/730MGDH8JC9xpBzYcEaXqg7WgirXU6X8YIiXZaFGDPVa
BG8u/WILRWQ0tnGyuX0L9BMvvxQJO4LuaBErNWa+Gv6dlYhYhP0NOtPRQI39Ieik
ZGMQ0WnYXUz3Hc1f0iJQTTsuwEYnDX1NulYSnO6Bqta6uB1GhYPhhfwP5GIpsveE
jmeGoAXfnkjiUvTJ3dO0jfByQ6tfJk54Y+Zzxe94luyP4GIXew0FtbWfeHx2JV/Z
lPisgndhFM86SWtU/T8/wdkQfO9kkYLbdPpq4YKZhwCfG54BGog+Pk8gbn/Xav5P
G+XoBSGbVdqc0hhegcl0IJ3ZFstDFv9WhXyojqYsMARAW7UmZMApYpACvDN7IFxH
W/93Oi7ws7ekhMFybw5G6dUsClsaeo21MZpiWcpl0xhGixBJrlFPd/gOArYpF3v3
BZoKn5dUZ/U/DGQy6FTyIQkwVtHPq+tLDyX/3CYTnYtgA5RCac15cJV8XRFgrykf
8BqZJihVgOXbaT4PyGbfYXT3VNP8Kx7qDkuA1rCsw4Mq01kB6gtUDrdSkLe62mny
rCBff2piS1128EUhIVjHzTo2cdQK789B8XPCBIMGtMIW1xVYSvZsVY/8xsFmbzu1
1xtZy9/KZq8Xs0Js7KJOx0eumO7rHpo6JLWVt8SOAq7t5gi7tbEn2lbaoDcTNoZn
1FC2CwzCDv0fUIzMDu+cJ9HrJyrczdArXqlHlnqu0NS43+3DzwcrYZyxu1oscRNG
6nQ/surlmirPa2JDHE4WzEIzPsp4LZkUY1QZWBQya82r10QhTgWCqdPRbb1EWPVN
/hoyDaH9MezHeqvEDaSAbIXDh39kBZ93J5txb6UsXbIZKq5B4Pi0xGsBJoncWWa1
5G/02rXgjWJMNaKjjhohdGLxfVMza74auvwPB1M/CQ9ulphzSpMF2So3L9pisDWm
AUIh2iU2uneSaFw0OJquNcqv1bWyg88HptAuGh0XHV3LG8teSed+TFzqSpQlCdDy
XgT+89xpMsPV8CuaA00expBvGIUpyLE9p6jix3HbsDeOAQw2AkFYMu6kFck2DcBf
9jQlaxeb0IXKc5ICKMX/8jZBI2+8W+U2K5OKMSXvflmsX7CUcYIscOKlcemb+8k2
/dQbos7+CUV8yN7EuqUvLdsFU1WcErNFfl3mwRCecACd2SiBkthl5lJf+9cyfjl/
tPIxdYN2mzV6hor6uVxDJ8Y5gQToLoleCI9/lGeBACBdIncx1TbPyEG1Xy8N3IX8
VBSunwTs5gr7j4hRtRpOF1Cl9oQTUpONkiv5N3dJX5eMxFw8JRDwyixVKjbSmfBN
hQeowEVHTt1PSis3CHyJzQvCZ67nVJ16H2QQtEy7VOWZ1RcY0wY6aHh7r51EPEcK
Big34oQV2/NjcFOSSFtApPno73EfeD9UxH/PtPuusCuIl3r9jUQZOJuuNZUD+KJJ
U0k+VbADyo4noG0i4x/ALE3cNoxhdsuD4GOioj370ihUI9V2RMkl2xcUToLvls86
1gUhs79T+PaWneBs4NTfP8e6HqXwXV35G3NL0bppGnz92NmIt5Y4rV1BVS+0brlx
C0QS/SnXVCmrYYQTavgxqisK/StF+BeI0C1lHodZiJe8IvcVNjf5qbLOD/R18FdH
jNBhfkjdioiQ7RoPLx+QFm6XNe2ydFqmvYStqU7s96+LsUpelghiRffC2BA93GrC
92TCye0i6PQYPzbAxnakmdTxAbv6i1pRNi/HHguWowAjzxYxhA/E8OYTqUkdyYwY
j+z1kEkAKm1j+9/6KA67pFBQ8t+DygzqrAZ9BAMPBaUgZABJbMrxPswac6hQllIf
iADJB2RosxysYNYf1AxzKRS9Cn0f+Kluyo1T4xeK8TDBgiHTVs/sgUybDmxliYZb
RZXKuoRzYEigBKIxboe/+wepPPnHiYwJASVqQOS2oulNglFD1wRvwxjZbzt2jiLX
pGvWB2qffmBTweAKf8vRqeuMGCa0sSZetUAu39Ut89sL/XxUtwotJqUvjSDbDv73
ZDnNSYPacwUQK44Gx5DMm1GMAGdbKvuX3at06Xm9VTDsthN58Y4/in1p4XSLrJ4B
VwYq3OZn+sDKB/GMZSgnMqqQUJ9VtjmHR2zMftTBDcTLkc9D+apRKqV3p8mmcJmW
ZTsj9X1Wcugm2ZcAknfU9xNnHgY88Sxmjd408enbqxpn+3Jzakfrakb6JoEg+bRK
jHWFil5/JZCFho48jMk1sQQRxCBDJAR38nBbvyPqLpVO1C2JkTqxRSLeI4urzTXY
M30TC9pe2IKgepwfTK9BZ8GUkbPL0IjKSRlLrNcgaEBG1ujk4rmrpHUxAYucfRBO
4XwvTVBFW/TF9RJdx6f9Mcz639fOjdHG1g2JOf/bFEsspHxZgaA9ZcDGrcowprtc
OIoiaeHE/5lG06XpOK1eVMu1ZJjK6zYZ/IyCHjCnwzZArW/chwwPC90JBVmV9lnO
F8fXnnXrhQ+2xBW8/+bOcWB7NgLnNd/OX5KB4pUZuqz7WzeemmFWGcCWl4TFL253
9/h2nW03Cl+BD7XhpdHnIbsLWOcr86BcsYVNJ7y4rS98JPsolYMJDxFTm5T/wvhb
IXqsrDKs+WH8P5LfUgjgHmTrLv3H17UnB/saxJEOMGk0VHkhBXU8RLrLPCUYS5Yb
wGXpojxguMNY7NdjWRyPsLZfyRRNa4/xocQ3nul9aS50UqGiiuSurs+kxv6+YVXn
/ZuPHdxpOJ+R0R6W5ep3yxHlAOmpCrSobf05O8WDWRHbOgCZpoWBFuxN9SdfgRDB
SXJtZgQLjpB7HDyzRc/evjwZRIdGvWWbkP/RM9ka8OZZX/dU4wrJ1goolneuxcRa
PNPT8V5TZfxas+t4gSrY5CybXgpPIG3lyNFgAltsM0tkwxMoeCBOVrwkukYTp+2J
7OhIdKjQD+TzxjTIcxgGzN5wO6Q2SZswJUplWqkmFOWJsjsVTRtSrOeloMGr3Qy3
yqRDs+B1SZpDzq9oD8kXHo2v4bu3PyfOKcGDxzZBjxjdtn2VM8yOhONkVubgtvTl
JdvDeBZ4weyDMtEm5tysEStaj6fVy4v7LQJNn4J7hJMDv7FXcDOY7q/5FjUO4E34
mtkTw+xoM2BvfN5sTgheG4xljLlIwwx/kuRXTwEC3Cj5JgFN4i/Ogl9CvIkTk8Et
edwn2TTRxp4GO+KRT6FWDR0L1mYH6FyesS2SZyidtnqLRJ+PnxCAklhvSCaKo+hl
8t/soNQTdthsiM11uIrzRDkc9q24905YSD5SQWREHyNBtip5+NgnHEVyGsffglD/
zRB331RgkAu8Ds7iP4+SP5sKtrQ2Nxz02PQ62X87n1gEOGihEXd1RTFZm55wr5Qk
ebl8gPXO1O6zRTMcmj70NFJIej4XadObHtxBFmhsiUp8NuProBT4xpFYo9znsSCb
8WDaIWQ8JSyf9YEzbiOdbOcWR9BGf09SC+2QBOygyd7YwNfPMCoChNh9xy51ecaE
Xu87aSfF2MHTHj3fxipMlFrnIV1F7I7WZWiJmzd4obi5aih1ITGb8rByxsTPzp0/
eNh9J8aoEXMVT57K559MVh2YTLZ+rkPuB8jmZ0gOnrbQT2T3xWjLEigstc4qZh1y
x9Ug3pitgywKGmLC+/RWTUNoo8xEATyM8UZzY0Ec+5GpDn40BzPM0+F5wEkUla3X
X62pMIHJsxr/fdDLhpe8Ec5tUHs8xh7o6mb1j4MSi3llYw6bCLf4g/vgxfGKlykY
s9EDWkHTtGc0gaBn2YGfnG9R6TXrrFj8DcGkzlsJWukLagna7krwHDj6jNe01dXd
XnukWbSnxsXlWUex4kYvtUrtyXW6rGQWZQSgR6GlnULhyXyW8nB7t3qG1BzW98FO
GeGp/QloiNZwa3P/c/eRaM0H3VpVVheHhogWTQG606dWXnAjdWCiBoc3qb9eU87F
If8+sfc7FL+X2uqlAfvc589HJOU3rNOsz31HbX8VsHBc+ea3iQtBXynPVIFFkijq
g+O2uIFgfCsXNdSSc5JukJAcAjZlxOsy4RHBOuhyf/QqqNqX5ylmB7CDa+jJn6Y3
Ujp6RLqnwPGIU5J05IBxHGUoU133l2ZIxQP0HuHlz66Qeq8r4dHQe26RwR9YExnI
Xiasgy1FA9M9S5Jv9GUcEvWwhuNxqT7pl1X2Z3SehPs6eU++dP+wwZ4fUTSd5eV4
33sc6Il7+dT6Y2HE0nD+29bM3AJ6woo1CsY0ToqEVvKsKJMZfCB9XQETwdCfKOrv
MjdvnEPfbwJtm336GC43UZ1rbRkwiZsfmCRW0FAukNWbYnPSNgbfiHBMl/t7DvL4
s+l8Md54J7o+kxczwQrmmYySM9XGtnXZeoDTP+RrE7ijKD+uThZzC2h2r4BWO9Hz
6TXIP1mc5wAMa+FGoHY1Kw5vky27DqhhQxFLV96mtT7dEWSCZYJdmC3VaPnM3GBt
bYdBEB0MYv3v9yLjXsTbRNWFZY16ai+aM8Lo7p2O6OjXkqZ4qo8+z2nnrjX58NSw
HU2p1phsPj+yzQ/SRJ0z2nYZGY3Khm5RoZe3YFWPZX2Ag12Ubl5gwqWxJyp7izl1
ccO+9k/MEb0+csUgE1jBjwGyFGTIAOeXOq1rUVRYlbj9/nVQZ0bfTGbby66lc13p
NXAMsnl36U41r1Dny2AbRY3BiLA3L6GhptPLsCNPMbD/tu1QIdDnYZeIqtXQ6nHJ
5cEpBu9o61B4DIdSBoUbZ/ci0aoop4zlv0nvTZFeXL48kN82yd1QOYaBfBXuesKO
FvpNllgJjgjSkHTCDHCnktIAY1la0Vn6EiQUY1zYdLYINa0wO/qKpJ5cjM44Dvze
PxVHtVpi1XUUryS+853E1hgNVVXaYC5IXLtLE7mUlkeQ6OVuVmcgCju6NVhfU2sZ
xnzyj74JJK3oCg+NC5QoNfc4ytr8pjEdAFQrTtGM8N3GKNSj3HCd5f9m0vn7op6I
PmxHNFRizyhJbDzJYpONMBH7gaw9+pssocsnhmkSmJkbCKE6dRJw68tE1WBYYBSs
Fo6fUprb6DPtcQDR8u8Hu9VrZFYq8NFx8ihpcK8OwlZFuP+MALdXbEASmxijyXm6
1giGffSsOqogC3JS2q6ULHCaU8AWda+u+NEEBrpJvhHBV3RXUtymZyNIaXfG5tCb
IWZPT/ozc8RL2EBb2VJmZ9SJ3Q55eBe5a7Ec6w8/AJU984SXfayxdvjvlyhvAB3t
XxX48mlln36WM88ki56F5uSW32ZrhBkFu7nLehrWzrs8/zLUtVZ1kHxe2/uyDlPI
0VsfdR/1wZIvUh9g16bPpuGKqtesLWWnDdRzK3ideo8FwVEvrW1IFo9+Io4o1olp
YiMeXQzEIsb23BtA2n6EnM30XRJsxBcmXUCj7ULRsyIwf+Q6juS4psWESzeML1Ai
bYxEi6AEL2IOlVxO1EaxX6rBMfJ1zfdSRftHAc/odUI5vSgh3Vmxnj15d2nvFK66
m6MEvifQtOg+rOIMoV/En81ELExiS8sEeC0XsCfwZhjoSs6tp5GmojXvOnwtg5yQ
VhkAjxyC7QipK5/Gq+suKaW9HZJveaqBS2grazpuzZN3lvaHe86fDayo2LT2H32N
Vu4LhI36KmDdHH9VjlgS00gD4XlaaE12JLeu/fi4J5poFLoiNcfklt9WYtr/gFP9
uei0ky2qg+AYH9XYEXTRnA+u6gW7GkX7ekpADlrUnVqu5xfGHda53I9p7Pqx4toA
trl7+Cmny0gbCiWySDKgxsOu+dglazwk/MJyAXRafjVd/k6vxXmncvJa+fsp7dNS
Iedb/5YBLc+8abUdWBBO5OPsadw5buJ9guqT4nq34PpA23h+a1Sw32FgCm3PHawx
KjK2Sl/1Ii2+SZjdKeC+8ImkChzhs93AsdG1/T3ie++iRhvHcPtKCdHyH57GwrtQ
IixvhdKFrs2YJ0/x5NVYs8Bgm2J5QlpAkc68pSe5EJHL24jXj9/42lWPjyeWfi0D
nMO4AGkmimfVl1Q9JWcr8aRoEeIQjC6p4fzX3VjSjDbL/MuYc7ymUrki1f+8826T
0Q+dN1G9oppDbOL6IqP/ngHtXgBh0ZIbjSb9N7ADKxvnH7BFi/8egN0pBYnmWjhB
4gXE24dnl8Ds0bIB9fmd5h1uxzmSvLDKp7xUGKZqwhooCKaK/nG8clnJju3lHHqx
v7oG7bCvKgRSFfWxF5Oy+64QFHeLHglBoL+f2a+O1nSf3iq5HXxqT4x1NikQFLuv
oUoxYjBiFGAoJA814MwGA6T0OgToadHxrVU9doobSok7bmmzE85h1+99d/LzahPh
8SHzxOHy9DjtQkd/jW8iZKqXF3fJ+VMl+9DPpvU8gS8TxwRDJAlKdSHXRR/245Zj
3p5m/VfQyao7E4d7+J6AWDKTyrD0GRQajuv8tE9zu0GAhfuEf1iALf2jC/xcLpN3
7IFyMDsYJEYpNdm4zvF2wnuYo+GqdOpaWE0u+WqiMPnGv7s7CA5MkX7KFMmK4WUl
hN82WjuR0nXEmIw3wEh2IGctCbfn+j2aXrLHICV0zSGE6g/lX6RkINvDIg52eIxU
fGKviFTeQ+lgrPpplaDw4K0oZgUooD4JW4qp2VbuYMtQlwqrde3fYTdcyPLOqNn1
4G3gk5Ru2eA90tFgwE4SHBj2hjvLa9ecPXc8rzSDGrqhd8XjRGyc3kOKlkv3WlqT
anhMxHRhYrG1RfdbTw2mfyHe1tuDrpCsUu9J11mFXOJmnFmuKJY0hHnNHyKbq0EJ
aoVmvajvk/FsFF2ry/n8N4H23tMAp/jGN8dSmmK44/VaJkvXqCXiNLmT3uoH5dnL
hZd9enTNPd8mP0Dg/MgSkhfn/XNsGLil2gg5eVZe40XWo+oz7v4DbABJfdxKxUw6
43ZApQo3YpDVHLJT7/thXMT+xDDAwM8YL9ILKvnmWkvxuFAssFoKDrqHa5S6B5LV
gefmFv7Hwvy4+j9BzxkGIcpnyv8NyiU2+dXiMF0PsUTZiLj/fyJzex05tvTR+1uT
SZe3C3DpF0JxD/HLKGPixWI1P6y2OQ49VZGDyYro7PuNJr4FCxb10uGek9EocSJZ
xBYD3VNpugxg5ZC9/IYWJU+gJQh0rqOBiySdIs5/3U5ZFPM8CZv0laJnKMNA0/xG
fuLrJSAkP5xS9Sse7lNkY5FE3wZhjglKZBPKFpm/cdWph39Rs6kwV3nm7JP9xhJJ
rmeb++T4FFFZyaHOXm7WP+wjBgJ0LzzMYgGhxjUme5ygZ+HGaUMLsM6Qp7FmIbIa
x6wTDryMIwSQrkcwtn+sodUpSjuyDiTW4aq0m0WmxLwxAyC9VzMyoH9QMGsHP7/6
CPsuRfQRLfjnuErjnN3cvrC0SntDR+xOSzhW4HARdUr2W1VET2ZBoRaeVqk603/r
V3G4V8lteOtgWeIvaf9dXEIBkZFrWe9rSFf6LtX2IJvivn3l511U+J1wStQXwBC7
IWe3Z+4qXZg4gmJQYGi5UeY8EaFqhArb+nKQB18cLeXeEUj9Niqv6cwE0BrmjcEn
fqRhuLGBl0OnPKOcBTDqUINtgQo3hETBe+00iSs7gzw/ilfrOgnjuAJRS6YvP9f5
TC7xlMPCJiQi/2WGj8kTZAtaCatGuiQL0lrpPPfC/uRB4Hss5WBIpiQXTKFqwLj7
rRNxrdqAoB8Xy2tUuEZGqJ4GUQI93SY9DaFPlyYU34jRy9p1ZiWJ7m+U0WTAYFxR
G0i6TweQHh7SvbrmY7HXPDTNGLlTfIlPXps+vGodirF5HxLY0F5l/Sex1Hn13nsm
aL0+7+1gqIN06iszSeIfgNrZsHmaYZTCAhoSi2TX2ubZu7eDbfi36yF0w+55R9Zu
YzHXncYv2Y9Dip4ABNkglF7NZQ25W5JHtn/HrKf3KEyrMxwv7ZmyRNZJWSxCuRpU
0bAup7uSrL14YO08pJu4n4t4/REtSOVW7OvoQLQkrRQqJL6tiGb0HoLUZC8C45Qa
/VUzhF4+KyiXom4/lDIHdUyVfzd9o2LDmgM5GKTRwX1hXmikGvIU4+S2gY3+2y0/
KScoF1IdtQcSUtAVnXJui/PQD9IgWB6GUZACmR7hoT7SIt1U/1EkBxFaqVGJsaVq
giHDnZpntdWmc2g9YWqqUNd8yLxBDRVz6criHz8KNmL3zS9ymNUlZFCv189Hykm+
EytQKqi++He7QnKYRSgGId+fNA+fxcTkqITT+wnEJWq6t5XYmMBLD91Ds+WypFHc
tJQmeOoVtOgJCXpQ/e3+0KoAg4TSfQad6uiYPljiXtpNDgsGLN02T1t7AtnXO/Ca
z7xOLnFcMTcpOxrzjbNJuiOGKfeGKJ6doi52VxXTNz8yil5GHPYNZlr2rDkcoZEw
2MbHOIvcu2WyEVQTevQYVur8J8IS1BoTEMnALk8z67VcQKvfwuD0TyzxjNiMhIA6
n8K9yxYBsAHPOCt7toHdxRvfyqk0U6gydpOZ//wC/gy/GHSHTFE58cT6UjRhklJE
1zjhxrFvehPNY6AzrnDrqjrBSBp84/HxsUIqMWuEvb11uNh+tzHi2albGkt47ZHw
gDuub/v31rET2DSMBXicdqSvSZBkWNwWtpbiWaQIbrT2V0hUGiv1KIdiHUndm4f0
oYgMu+M3+ctba33PfAc/dr/ugMpBdhYcxSNPHl91r1wzbVpJlVvh4pKKeCoQZfu8
k3zW8S5z3/E22fiFdkJQp4FphGFJLdF49ueahjvvR85XpS1K/sZLF0uCzwP9BelB
NF1AN1y7Ebl5WDYvHcC7HY2cwne7rMuDOsdRbDyjXtNAQRi29KROgv4q+XCzXdP0
Vr47+gf1A6YkyqMD92YHCbamtgL5eKG72MCVj+Q3yqtw2FbU0iW88wopopeDfOPw
1o8HJNu/8+L3Fnhf0KKnogpp3AlBs1GTDK8TMogqxvxYC8xGAqXxXbQkOsV6qzoE
GRlmAFCS/VNV51UEBGdBVhmow2oGnWXdWO1pjhQ/sv9BwHekKU1KkoG09rnFyksE
mBpgdGxC3ZcH1Th19qJo1UFhcW7W1iuwiE6VDCwfn20JdrdWlhCwzgjgiA3O+JfA
+OWm9Cmjq5kqxpOteq3rZXJ7ihx5R+SHWi6ndtF7o633+JENF2ezBPqBZ+nFG81P
4vt7Yg8fwyOXoRXsEFAbturJ03+TN15HQziWCqLQFZKBRf3Dc6oshk93gCOCLBZz
j9Ln5h370K3NNeOYznxi8Pujq36LwkHkC2sgWX0yXGLGdPQ8g0yK/402GSU7s0kr
Ff+l0uhy4yPwloiK6m3KyZQnTRNVKDb78qJpwKMUH9v2k/UiBNy9UtXOfvCrQAnA
Lnvp7xvA+Rw3ofeRcsrABmQNadf37djnIIUNEJv3CC9kjF55WGsdSiMiCh8waNTe
E+tntYBU6QoQXFMz4g9MvtiPStdryZ6LcJbVOVPs3KpQt/+/ASeN1e2+dPy4blpl
Dv0eqz4E/IiN5/8i5+c7vfFxsQ+Zsd9Y1PBRSZws/hNrvidJ3E2QZNb2ZFRL2Isn
WSdUxeB5VToa0WTxgLLFC7Wxw79jgn3gGKMZlFvnXR1hg+Y24G9DBtZ4E0hkQoBz
Z4hGyZ22kZ8ddYD+kg6KE4nuKlyPDRdepHUyi7j3HKMeOXLaq/sCE+ckgUNkNWyp
CXztNkAIC7DO9MZEGkObkdQ5H7nGIL3ElaoJMGpeqoiTFgjYx8DRX4fMRK3d/zAQ
jzA/oPY4C9B4MUrgBZGUrqeUWM0cADCBTrcTPQjUNIPCJvsMGAmyGTpwXfxos2G7
1K3YdARtu8BVkLcF8N0cVn8E0iemkyaCltsacwSL9D4Y0VERdmkMi7U/9oaX184G
MU44VzeljevH8ar5ayez1XpE8BYUWN1g7qKGLCRyToRa3PnLPpxeMwP8fBywpYP/
A3krkVm9MvxqCThxOrd8mIDo3tywlhlz3Gk5of9z9X0XM6CuRVk/8UzMb1CUPVck
bO8B1aHc8sfQhhAGfuE2oPpsjArEgI5AEHHHAtHcWKfr9AI5Lm3rglxf7ZtZSdka
InyuYKCKf5IrkW1O2D1SSKwWL5BSE8acCnfz88sz0DfMkZiwGv9FD8rfJwmARklf
hW4ufbgFtRZ9vgTgLOTFvSwgk19bEg9CcgOGfay0abfR82cQlLaO3uH7mWWo8uGm
osiJDqLWeubOL4KuAJhSnVQ2goRTMEMepWT9Z8WKn9TzP554AMAwOv8ahwctp/jn
BeiZb8p4AZQI86nO1D4AxTqqK+6bbk5bCjY0KZpuxZnIwVnL2CQ32mj8qa2foApT
hqNJF1nKEI6Y6d112dfroRzpRuC7tpd56fmkSr6Ym37N1WPEcJCGcU/6JwWBrL01
WShAQzoKZ1vLMG2pqX+rWf4z4/jjYRUL7Z3bRaq6morFCqEWWegV58hOA6opjm/O
MqZMOXlSDCPwsBvfWzgbqQFUMGH1oNG5xotBa+FOjZkNpYlNvjp+gZQW6tWwMNpj
bzafoULSU/iDxDjPBnc8lGfI7kdeMD7KK4mKFfq/J3s/cppyxcMggeYtxguLree5
1xJNYTdZpJgwsOSvT0p77xIhOV7yMgUltES7/gQRMKZZrLx6oPR2z1mOTF7AnZ6e
ryiW+VriAZ7qXWA5sccBuEDWg6lvKSPq8iPT8WEp+bWZUzs64Y4jmO3GKIXv3P1D
JgwZ680JgEgjkVI/By401iZVF4ia0N6I6Uo8B8gCyrBnlxLwiV05gfi5Qs+PsYK5
aKozgT8vYPRCcLRgjecKCwBE60gXdleFzUwwsckVIBPlOA5A+rGq3opx/BEpG5Lq
GmmofaGr5FBlaQJxSleEHzeHk9dZrpfwrpsVvVr1kG94J5dhO7fLG1IqTXhsnArq
mvu/KbvohHtT/PPLick5E6RlKgdYYytIzCp2JgZDFsHIrqUZ/4iHtPRea3JBoUJn
VSwx9GtrY8HEJsaT38thx1H6L46xzklKsj+ijZmxduxSk/hYjAFFCp+IFS03k/Fq
LRDyeS+d7HQwoq7lQwuyMMAHcOrHjOm6aOH/5uqJno2E8Qx6gFfL4zQhXKE5ERDK
vfxOqsERQleo8BLCWgossiMCUEb9bC5ZpTshqkTue64Z+jckHHVSzntNOGk2wE7n
fn9BU0I4/hdN5RUsuu/MVC1jVNyuZY5X7T85hV+tky3xR8hDhGpHo+K/mZ3n+e2i
OiuUSRfkTEVCf06qqSSwja4DCu93VPZPMqAJLVulysmE6xbzY1YGBmTlGxNU3Brj
ylIhKTtgxrW98xOnZlwBQK6b38KphF86n1WY91H8EVhOZ1uP4mGDzzksLb0M9El6
7OzaZp9B2S3zrIfKMGZ356FR7I3AEtU51YBKm5mIjwUzhCEg3nVQ2G05AirQfcez
Il8otObj0SukDvXrqT5T+dKbWNzzTYIKDu5nGTyJyddlE9lX5iEKqWhsIgND0a8r
ZBEpD7JwD/3x33HYOg3POun82yi0z0MPRgy27+dEaROuqZmTRNWmcDrkKwhr18Qq
k8bTMWMjrHwowQz2MifieTjOQiNu2ZuXP99GM9MDJa4BOvi6xaOP6gVdk0Q5+/cl
C6yY+uWlsEuu12VeT5jg3853DI/EPJ4mcJlX5pBvVzcIa77/77hmEVc25hrN/d8t
3dQxjSWSgozQ8tS+yt5/S1CnPvEBufIRLgFLAVulrjEP/OvIdlR9FQCs0uoWWRq4
VNGXIY7t5qh0qh/J4Vlwr2HyrwBNyWwjD5eO+m3YgLSjr7ljm95hlEEGC6bj3bVF
y0dlkqUtly+4G7Xg4pJvT5iRtnJ960rtv2yHriCi9rnkEfkW+3VeuUMMqrVSOjc1
jv7jRJFmrbDDeEu6kwXp9aWazHH7nEpg8Yxsle2kSUv0Np/ehVm01thhuzwtq5JT
0ENOr8iGIBYE/s6Ibw6u1ozG08MKkRAl+59YopMtfMgMnb4fSJgHAl0oCp/42ILE
PFC57w3CDVS717wXSAYap5awRhw0ZoDVtlZPGBrp+wDiya5F0Pa8DPFb/qIdONWe
HgG3mLcWkBNQVBmZ4CtpboE/+GstT43/77tCrLzdoTr/j1CeLgz4OwVJLDfavuBq
OnP20Pw8Goqe+NbCRzINHisq8n81PZAia0Zq3xdSs+uYTodJzhPf+NGEVpKMV+Ky
ullsjJmAXf0SnAfyoO1KK6hWWyOxxFMdlhuzXVgnyvkHVxXRmfSaAoQ0LFSdHfya
dJ1VORz88KzZagxdXu5VNouash8zigLaZjqEVsMN4EVygXLA3NQD7RJxjfOkECCg
pPh5jGhnPTwFQHBGzpJZ9wa1H0N6BGRL/vtIGJgqUiKVYvhMgW/A+GFnsn345rMd
3pN/aupPpJ4XNbDVZpDySCwbClzoKxLwzydOefZ+oCoehYlDuoP8vAaE+evP42LK
9MSABt8Kuqu8FKDDx82jjvxRGC1pDLE2WYefkkjiJq2UDWH2rD56fVMZzSflK1m7
DjheYGEbcb0UFryV9wLxeb9o1dKztp9I77ifKQQuZtgU8UE/FPnaNFjed1gOwFPt
QDD1TmnUXVdY+3tpBYy9mbE80P/3htsYeoe45ZVc7cXzS1mdVr8sN2Bso/vL3LWA
VhP09AkPv2LbmdhHTTnXN6pswino1kbBkr4xf9Y3M1ZTtlQUEoGZwOYr9jSFVUfu
rwPK1QSD5vHQchHUceOJz0VEgP2XH7+OcJ0zpVB2+ZSsY6HNss9kz9zP0Zc2BT/I
c0cASgVYoxnptue2JI6vzpyS28oj+Ct8MGYMvR1j1pAQD4TNd0m0jfBYBGezMG+9
dK7xoyinrcLmcodDaMZIBJUipZDOHWH3uDxY1iTtrsARLSyFH5SY9P+InvYgp+GJ
SU6M8fwrgWBRUxvKc3F3l1FhLgPR959LlF6vlKITCMZMuO9qaJq7NvHZVUnJDPr+
B0X53VCCmKVQc/6HX2MJHcVPQ0MpmkX5nH5KGuIl5GcG0Vz+zDDNL1eoe9k6tUa9
BGs2HXr8HDpgqY57HI5wwxkvKaWdX1BxOXxoXJqfvojAwewRC8LHdwR3RAHn/P1Q
6nCG4qTabvylg0L3cYh1Z4zIaHb2nG2jDdEFKO38uw/Y77dOeM3S/VjoHkmVrdXY
YcbAfHmnzdx69BeFmTJdOa8mONu1ZRl2BBMvXmORepGDRa1w3GsneQiDx2YzEscg
ggNGtNsPg9cfsQTtBECtsf9QjI/kwutVlQBYULrnIxNlOzCCtOq648OAHg4tnOw9
WDPcja6ZtClNYTztTkE2D+Y++sVOUrZsVjIzzwUBNxUHiya0ggXH4dW+zmauX3Jr
Mu/fBevEPI+bwOMWzV1BWKlRlPaL4ngTZJP9v6dmRxbuLIpvvU7TPS0A/RTj1yE+
sPOwHf+rQACapzHAs2xPTtDChr7d5MVi0zeVED1/rczLrtN9pSgsBwlT2RrHogWj
OG9mZquqwQvLwpNUzcDbE62I+341LAvH8mlLrSq2rHfjNpQIYhnaT/sTnm60XVkZ
YCT2k69Wv7dn2KHSYNBM3QfNksFimHkPciT3/NlSkjtEhBZjHefRYkfV+jgMtc5v
xKY4vNmQTxGLL2FbS4kJek6CJUUKpsyPS5p/j7SDSMpPTUocCAE/2ZKldrCcjFRf
cj2qx53gKupawbR/RUln/XLq93suaXLfvIEc82pY9VO2lfgcTGNiFALLHYnLnora
HDgGGSz1ceLDnNvBL6b7MQWpMSlo1M8C9doRCIB4AoxFbQej+BpNAqTMdqZnGBwQ
v6OqLWbz0nKMUldA2uqQviZjtFrZKVWzraZ+oFTaB3aVO5i4u8AR1pq4QnXoBeVC
3rJycSDH+RDFuFZu1WC2gbJh4auji1n8oIYhCHwSaMSS3Y+WQfrSDCTAH4iFbIvn
x/wD5F3tu5yv01mdeXcctFDh7qGu7vFVxBh/Eo6YlCsbg3ORVCqAzaR2DSILAVwO
N+UO+3XkAFquzswUqoJuNnBPC4gcl9dcy/ctP0tz/IgsrpAFLfm51Uh5BMC4nMi9
KMD2WWJ7F0yF7RRPEwK4srGmUxu0vBy7xIM6LUbUzP9KIyznPI8DbzhZotBQLxg2
5xLIb+bpgSV46aw/gtC7dZ/gFRwanyfl+jw/qfDHlaRmqKo7vUHjKxVcisIS5p0j
TILyzRaPSp1N0lALW3oiZTRy/R8GAp3ic6Ue4QF6QLfrEQvzk6FGPLd28puahCEJ
HmSuVrUhi8bZMsnSevGG5hg8WokF+utldBHGhHqwuQac03y+dqum15C4ipsEOzkN
p9TRp1LARlcF42sLY7PTJO/1IjtRAiM4aFwGxhkUw+d9xLziifBjDnSNxt1Qa0Cj
C6VPHtAjROQ+Z9CY/ErFuF7bMmVqmEU4o+JXgo5bUJfkRMGWbEm9KSxZDJZlewvc
qct0kkMRWF6wTDYCZsXcjackuQFesocQE3D98dPOIuDeRzUobBAYMGBxQoTx7HM0
hANWunhAkNYuTdZTflNnvz9+57S6Uj2nUX27M+hrbGspYyr6BZeRnVFTH/jrOr2Q
T5K81cKcEFVzpV2hSdDtN+V03oQ2WXJBX4l4jhApncuk6oFblxzSgzlwmaWGmjhg
BZgoNaxt0rWA3eaIfLJWW6YjyAWLm75y1RcbMyUklN/XtbF5vgVRlXa7aU3HeHSQ
6yyFhhsrmvQ5VWngwBCSREtEBB/OhY9rqxU6y8qUworQOGR8b5mzooER5H06WXpv
75/NJaeL9xptwQK6G29rU+l8SiZ0fcuZqQtx3AaHosTH9s50gXSHs/K9uSxlbyl1
IcLhw0/EgOlku9JCh9sol0nIXOlEZqTY1khSiQCIv4p1vpdLSGfM6x+uor3+RCBw
b/ma8hMmA6MH/x8v1Slr4264YzpbnSC32uksPIfyYx0muw2AbIhyOwxU3E8S+aZv
jK1WOF+Cc5wBLwhgGEm+aWfO7xdGJSYT1qJWs5bHoJtTupz6W1HO9/w+/vIHn/se
lXIoWCaat5/qUOOD1cLssWdpWOWNn2+6I0vaSqLNtuai5gduuPzrjbNDdk1h5r/T
jJKm8wui0UqHZVwb3Y5boLsEelAyWni4+WJW7QderlY/nhURqFrx+hciCNhYa7+N
4AhTY6FBiSGvJHi48y/mF/j1Bkl4zXZoMd/L9TNlNMzQi6HwETPjQjusKtoTTU6G
bKgQ59s6oOFn2o4zePR86ErSiUXXDxLbB+8r1EJ4cCVydjYNZnAua1t+9fOyptsq
Z15cju9oU+Z7YZ/rXoM1VI4MtnVf2XxOVYgVcqupr4y6IiRK+BSdxKeFsYKh5hY2
f+eRmwK4G8bFTUed9lqUbC1zl0plDlouBy7Kd9fas6v1Ss1F8oFWjWVlf14QkwVs
nmk4xajdYfuMcCfuAXTOtlekZZngd8dUpjdt+lNLuHAkrI2nw/FixnyhxPJ/Jtnc
/fQrDb7mLFc0ua8SfGWUvGAovRZpgGNxtMIqR4lncxplaWPA7SUQQSGi472VplNr
fWNUYWKM4K996LWP3aE0yZRNuFBarOL3zI6+J5IRFLx/8Qq/kvXYuxHvn43d4kuY
Yy7XyUIrQX5O++uq80ji2T/BS2FbsgA7oG9AcxNuDvLHVFAXoZ+K2IeF5hdnGSg2
dON4P1fD1Nx50YBNU5427DcuIutwO1vy6R0sEa2Wm9LqEUBt1W6t6byuKKca74CA
4DoQX7C3RO4pSXBdFbJMbb0CXjoV4NikUB506+s/uvA7Mke38X5eIdLSXg3d4SUJ
kA6z6uU6luiLa0dKNBdV3HC/Lp0GabVA42ErcoGS/fMVgxkPP/WPp/OCo32KfZkF
pSSJdsFYFQ77bLtW+ZqUtKMrF0DytQhca+QreglEfmmocyaS1D4Nuo4YsnXLHfjg
wy4zjuAGHt8YFZ0B0Yii7lzgk98iY+RzfKJswCO+1mkfaO/dakIuQ55P3Pzs2T3E
2auhTq6RKRIM0hirY/9n3VyYi4ePcVx8wdF6ESdsz3zELhVCzeHLsALpmc8H4397
hX+6o/AeB0DsO76XpOW2ypAVA/38zq/DqbyoXm+vrY+TTBDdt5umhUynWv7AwkU5
Kzebq7P6g+LFyhrIGNs4cyuIgGoRnMrq9rv3dw0g4lCCivArmO2XAb9ZUzr/GiGE
9DrAn9B8CGeaW5vmOAXK6zE5GkZJ9psABfdMLxj+dgmc+nH0KxbqK4PUNF60yASY
UPdDEEKBM+fcs1GhCI2lICSsA4kFneBApT4Zw61jyPIuLAAiksUi/YEsb6Fffvsv
Xo+d55Y+8da21ir7sXdz81m6P6alf7siINYKlUewZVZW6e0a/YnESrIHj7ke98aC
PjqyRLO86OevWm04O6/mTwOKK9zib8Eg4+SB6ElSIRUHxoU6A/90+Fm6R6XflEIx
4gsUIidPW4U/b3Ju8WMqR5dX64YRAtGIHXqNpRp42JNvSgFmgceHOdSLX2NtXYqP
MSIAGz1LxAam9Ybg5+Yy0Lj1yPOC2cFT/FSc1B93ey1izUA956M9KApHpNAfyUM0
YY8f5Z6rgTMIcU2r1khxSSyHlm6T5a392UC/m67NNPTcUmI0aoGfI6eragrmZghX
LUFPvcZ9yOwzkmdcsmCK27sNV4dNDUfpClpn5kzYEVA+ygT4FhCRg/UW14WQEtE8
emC60w9adQ20nzECTdwqokJkovJFTHJbZlLhmDytGy2g7b9n7kEnFLsfZRV9opul
xUM+kstzymeBKof0du2KSvaR+iOA/VHF0ojNj72J+2ChxVxhtAAr9L6K6qJYZP5W
y6HCIgj7jvD7+yOs43I4iOUDW9gz/wZLnfhC/prGlWwmJ2XZBJOiraFQPwLNcP2s
/5bqoKBM87nFwkek9a8dZQ4557tGjxVZweXyk0o8GGtKnIG7H44r60mjD5SnIHtc
Ryldwp2bz/8FZMALDXaL6/y/6IAorGd6nQzlUZZLBSUWw+Du+8su3UuwbR1zWoZX
BII4JHNTHWORSkrXEkI5WXKvfeRRnt4Uugj04c8vWu5z+ThlvtSo5TLjpkJVrnbi
bpwD8WXoqj+QDJ3o79kHbnQguDLV4gHc6yvSQDq/tHBiBJSL8g9p0OdVD2ZEJ6yJ
zqqK5NVdbhTM7FRJK+ZeUV+9hUu6ksmSvJz10wk2B6LOEmmAWkKOG9X8seMQqiVM
KgIXDA2XLX7FvAAHfuLQlZuIHTH5YPVBDDhl6gZrlPAeb+0GpJ61P0xYL4ovtLKR
SrG8sPwTYxeSOe89WfZFOiaNRW9UeEhxjz+BEfQzLN067Ko5B2dmhofwwkPVz+hS
VllQvp0zVLaj0KQaQXk7v+pLBcOO8uydaCP5xkKd5atA3ZAm+pVlRaaphETA9UIC
6yiIDHY5Lf5sxJn7WLSua1NC+YSkEifsNX7/dtdEIEAf1WmAPXCZKG8Au200Qs3p
fvs2CHkAlYoz3kZCcXdidKwhjNwzHQupkGHXjrSs9iHaYfk0JsF1mQvIx9i+wpT/
g0R5tGOEk8m3ih+OOWHLTqtnDAtDTDSSlCFxITRYPhGV5Xr5OVd0bW72w/oF8KDZ
BHKoNzkn0evSnnSn3CiQQKTw7YzzfLy0gXrxi98CQK9bFryw1vT3TKvwslr5sm9+
5+rl7z+ctYUDnzWYfAj8psCSNzOcE/24q/d86ycSoBrAuruo6+qXcJN25YQBZGe4
Pn7m3nrpm1D01DIslrkR3zlZedBqdeQJxwq+T0SZaIimzUfmdZpn0S7BXjpC5DVv
ZX8uqhnkl8EGc/6naI5GNETEYNHvLeZLpHXUQUz34aI6lnjYW55v1NIFd5n7vVB4
ulCC8Vt3jRWiN/Nx39jx7AMykDnnIlCEBayjttLe2+HoTrwW4qAX3LLsyqelPixS
BBxxgUkgtjpHoS8YT8RdMeOYfSu4u6fiywpqprGFMTF4HI+kIQdlG44VWb5Tyk8p
/Grs/tzkzniiYHSI3GIwVz9uZINxyk/0e/K0eSLyXmI9zBRUmcOxSTHoBuxooXoV
yxwFN7nCcgzcLvLnnLRQiJ/3OLTR5HHK5SEOVJJAJW4SKSaeZiwHmWBsUeHnPBVk
wL/L34G9PtMoC2heFjZfqDeiqQK6AkrL1V56qqZF778RqwG7hQ0zBeXfWSkw/kGu
OJjh56DNsmzgMPgUs+fvUJzfNlaipT/twXMqrRZcstA3F8vJBrYZY9o9wasp96+B
UzgyShHTWV5zeg+8BZCbHSV1RPMOQsoxP56o0yOLyPpxdf9CG273ayd0Vb0x1SC+
Po4XxyEdhSh6S0y3bbtE0ymV8SrEW2bOD1aCNdyI1+ORgtr7p4AS0BO4SrJ13QeB
ZrUuWPswEbe11DV8weyxVEBERrBootDf7M7W9OVSpAPs2iPcXncSydiQMdczmVsp
gzgeVqTWGP21HVPrXVd2y0vq2sRdZ5SjNkp3ir28+Y8ejZIqMBK019UYgMUzJ0jr
MThpZFA3IDEpoUynsYMQ3E/lCyTRs9FgMn9jncpSe5I4AkopAYTqgCxeoqjAx37T
0z9+PfSsIX48gtjLb1TNc/pWGV9dZdkK8bjpL4Gp5ZGnysRCQMRp1Jgzq53jc6o7
SkG3Oy6piDZSF+JaIep8Yh4EHtWPNvrNBila8w6x6RDzd2w5zO7fzR5Pd1A4H0HN
3LOxokizsSSYDU2XwRHcSUCaUm6cOLxWjG4rMODXj5ewzDkpSclwids/p2FAnUPL
z398DAqMVUlrdvxuBZffLwyWyuRi8Ae7fULPx+fJYi5cfXpRn79ssFZPocuWUdwZ
lcP1dWkn/PwtAaKBXf8OqCN463BG7bvkvaiq4oV+tlI1RNyWEsCkzNfdNenY+UlW
h/UcpIzW4UmaykuHbM0Z6PWZe/h18q06a0BghKNgTAiu5ZESs8XvhpR89hz8fmPE
c9JzJQ5jXd2ZvN8BnZVeGH+s8cjfHRSiBW/NgigQGhLpmDL/+IImdqOR+zKXfS8/
A++U7jnQnefYRwg7YA+b9KqgflBAkZDYBJR8Y6CE0L78ZpB3OIxJC22+VYpuptNf
Wjt/AyGKyw2206+piEHG7wzgTIDQ8eMore9ZeTcWzD4di7WINI97GrQJsjyFdHYY
k1PMYD3sRa8RiNovj+U/kWIYrQJr7mlT9q7cmmgOQ+7JcpTOrV3LT4KC7XEBhp62
J/L6dS8fC4FJuXI38f9lNEtd26we+o75vbIVxjn84+Um/PCPEIuToTMNpNvYX3Z3
CDxGz81Osit5NgoiCXHX8pqP4Hb0ngYC47cRjxlST/lQkkUpQ43kTYmWgPrb3XbK
hyjHT4OlfC95CWnMpDEfkCdV2RYw3m37vuWqjpYQneh8ceRwBhl3sQGuCVd9gFuS
ubh4RwuLkhBdTH6dl6H53AVHrQWdtPmbZcp/jtU6PpdKcog62GW5vf0e+8vsPitI
e2F4H/jt2ruTnOXUId4N3rCv96vfZhTY/XT7qw3/Fx9Eth8j2Y/5ICSNawDBLIin
tWLkJJk8jiQSB0dgGIcS9hawWTi8TLHenFTQ6rdVulwcSscYtPpouXEJUk1qDggp
evWFde4aDr8LPWOJS9YValDdT6+j8LrB6TeR6t383SS1qG2WOt1W0HHaJogEn+ps
JcMp16Ue7eKVNPERzQAUNlCWdBi9aCRjqDNU5SSxsHj+tXfzYnX1gASybNG7PRlL
5f8h+OaYWnANfr2aAKHC2hTaAtE2aWXMnUat4ppvMgv92Uw08SmpeY7e9osJwhwP
LmAiUbvGjyc2WbCCM/VvHpu5oP/AsZXe0/ue03h7gTQYglYVSk/GoW96wqPQnPTG
ibIu3ZTfvIV6JCX8e6t/+rmuhZm/HwcscdjjA+9Zv7X2He6uiWtWrNSdkoUKc+0M
v0VGT+9mZ2qKWIR+sAoENGpM04xXFFUCduFkKJ+VH1BfjK0lR7XYYzauwVf77K6q
r1fwfklKNM8CeeI54AJXdBMQJPHBSf9Mzi2RrVdGahg8+oAaxR6wTVXUv4bl3LwP
6xYuR7IAyJCFWGwbfl7G1ZkY69MI2cogfiwae80UHrNvZ9DglymUAH2DgEr1BLfG
MHGbn5QQ8VEfxFYkg6gx3hfIfTHqKllYeZQdZn1x4zGubpE2xN9WhXKUQ8+EPYEa
p1lMvOf8LFhBSePj/CadRcC9s6e5BFu2UBZo+LbAj52cdDcT2LIgI5mWAw2j3mW9
bxEEyM+vRkIDpJvQybrAgEPj0cITx4PgBWfRZ0iYGkme03SXClbhge5iHanOwQpN
RTdcJFMZzIKhtgKgeFQr8a/ND1tULSiz6DcQdHRwwPvriinHfRPuln4JZksFLMQy
zZpeSlsiTgtTqe2EcwoilkKJOuuSkCigsKoTY6/iuErXEPY3OdMcyHwabFTFkD/X
mNL8q4iiwKfVI2q2cdXW7cmj0itViaCmJSG9OtYx4EtaTPHVB5QmtpQ0/CKPNDnG
uhgmOudoJY3jIzZN27KDwh5sjNGbYPzEEnUO09FabDXIcxyZU8/05hW+jbI1ahMi
sXlarKSvH9upkrEhitMVQvmu5vFNqOXLLDzTFauY7YlWs24p0tNwp9OSXaZtyK+6
wO6KmtajVpB+KseJytXmqghK3wXvX7Vj4MovB1yYmTyqkT8BwrsyE3fVdQ/NX/d2
aUpqbspyVUmEm6KOkWIp1LH74dc1Mh4i+2tpp3qcmu2gaitUzsN83jOR/a71sVU3
w8WtNqSWBwNbAHlA0Spd84nkJGS4iiExoP0VwuLrpp0grnYDs1Pi0gC33cxIiJQj
tmDRLq/PT1xQt3wCDOT17EAuINLEM9T1qwh8dr1p65rSxylWrZN6AvJJNCkrrXQU
s+tiEnwiZx45HT25kTOPxhhGIzPbf4LXYn/uJDKcZG96SAxSWR3O8dvMdAzQJVH2
K9mNO4yXj/ixDGZP3i1Z0Rye1Wg/Cr0ZhxzpNm2F1TFgDWOSQuysp+dkb8pebzOz
eHxcJTmu+4dQ4eWB1PnRhzzcouhnsMBWPlLZmQI10WltoBEK86GBnzbn3aZ0kcws
mGtNwzlW8X44D37p8N7f0vCuNZkeSY9iwFqBz7op4SaMJToXm+eVqQlnrAM9iLFL
VvPLnIVqdrJGpzgiJ5e9piHBWB3VoroKgN8BMQFhHlga3eIo24wYFSWjkZ4kFZ/K
pHcYByY7iEDm4g56kJ4rIUgdlx4Vt2l4QG7aAVCNITqiJdXtbJTKw3HiVLjuPrhs
5YaR1Ia8lDWQAlaIj91INh9sb0SIEqveytD7o50kufI1YZSFQ35NF0aR+CIt1LpY
iJe2s18HPeUQcrZkY9gzI/Ep6XJgmDBfkpYYeTijLlNmqY/xw7+fvmDux6JH9xRX
eHDcC6ZvV3UtvjcZSfw2Z4h3dU5nFusogyqljZsPrsAdk2xz5Nk1VIbh7sD7juhv
tkrR1SGZ/TNN4mijCr8iLrpPlvcjIb6B3qYKnXPG8pkwUeIJDBI8knKCzZ0cizNp
VcYpS6pJwRebnY1BxJD7WY9KFftXWHLxMt712HEiLDLtVYoeqroI3pt0iC4EoH/k
Rj6lXnhtce3g4JeJIbTqORDVf43a3J4m8w7dilGYvaPshA9hxabYhVwuj4R5ARru
ZVCHhQ+cez9VmSSjK1xrAKlqeHz5MPZwFKcke+vbF6cP5DJ9TlBDF3iKNRx0WHOU
j8A0uG+DUf9gWnKflpgOv9Z8bPcN63bDZBSJDWfkEMNgwwn+9kvFp2p4hoK3pzKL
ZiRCvbEYVq0NWfpVltO2UbjKceTsIMeA2jKxsPPx+5eBaS7MqI0O5jOdS9M7Z+mY
UyV51THa1K+EYxXSlAUb0nQnRQA5Phd2CIjqYtj4qOwdCrVJigvMzd0C+leZw8h2
c6/VRQRm3QW3dXzCTSc+ig9RdzZG2yzY1CDClWHq9LEuZa0Yn0A22Uyhla8m1oU5
LxHwqntjMjxWXHZM/HIYltbkppDr5bWUcFdFyESyU8PWImwc5ksSfqAiCfEPeFWp
4uJF0EuHFSzvz/2mK1fCMx+20QEOBUkGPf7zvJ+LkkWnHlc4YkwTDEpE3YTFAbDS
3yb11UVR9gKnQ6seuhqywD+SM9UoT8akPxG80gM/27WVQOdaiEIar+OkCUWH9EUz
3xZk1h7OPqqSGR3jckelX/U+t3TLgPmuVfokVFPAjTUWhvg1SEAZ5ydL4dk+qN4I
XTbSeoVWSEt+JSC9/e1Gq6jeJQTKxtHdhkh+YBOro0gl/t1GERJHisRgWHKCtlDc
PcouseI3AOnw+6krP3Ph5wFVHi89c9RQ6BJ7xA1/NqIK+23Xor1nBHrgdLTfzyc6
znrVFcNuVbHYu9+gfwnBpVg7YVrmNc78zuGVY1ZsqZrGCuIXgRdCjnhPc1oAjVw9
/PMpX/aNJ2jLi7HLkFBs3V4KCpnYHBZu7SDKMh8GdwoRmxP/71bfBeRM+YcZUpi9
T3yMr0Yb86kxg5VgI3WuAfB1VAqrAt/biFr+wZBPw5TsNpdbxZzERHRJirRllgYZ
/jd94ev42xK2YoA+Y/m7grZ5DS4Cebl8u4NU8U8xbLyfa/FW0f/yWYo8/mU5NvPC
ysO72VIx3cxVCcH2H4WkhZbooNuLc8AeIg5j2fc5fFqzErpy7tfA+tbJQU3FQCtb
/oqalrGfPNc7bFgm8sFC9600PdlFfmwWDswdvfEy/Bpmk6K0oTnk00wtTzR7vGZ8
by3WViAGeDzh5JEe0nyl9QtVuWYdOSkO7qklDYP30LAbatX1jSWcytiZzlXxAGd7
3wrrTZjO+tXWEG58vn05wPNfbZYRUTzI5sS6QLVj/I3mZVKiEk0X6oIxSAeqtPOV
uREZN1TpTGTvKTuVpCd97GtLpthK12zMQfiE+ZfK8b8nzoel/wXlGlNGa8irZnHm
AqWRknYTwoHjtEJvmBsepdRqUJV7hNHE6k/6X3wyofgXCUoHZqHCKrKT4teoBZvJ
rqLv2142UOIGVvLHzdqpfzeMM/B7eUx4n4zsi8tz8jEw7udENoUchRURLF7XIQKy
aSWqTX4LKHqE+zLODDD+35d+dZ9cl9phcWd32KTj6d8uS4TpTa5LcW7VvJrUOjty
qxZd9pV+hwH2ZywcQoPs8FcKKaq0FSD++YrrXTDnmEaoP0MAircxTdZ09o/4VEZI
bF4zKSGllcHWL2bze1kiTTW8qBF4GZMx9BRfljDIAAKY6Tp+b8R5LSMy17G1YL+e
gwGYBhmx+LMv2Ed7KVNikje77ChQWZqYPzH2GmcfeJzqz4JP0i+ypdwDb0w9ATwt
4X5q6slCW6YbHnALMHkPaM0rs0tTk+bEaMiavgikz08wfwBZNnFQ7Jggrr43Q5EP
QIa9FmwSvRzFYiRxjNthqm1BUcnK9JCE9FhJSq/tULqVbX/XY9yDAP1SLMHAuRS9
iWQaAspRaIXXRkp6EyCDIgQuhjSNdkDkUWyeTHRQjVylDYYzdN9CdWWywp0ZmMs6
2tpSvsi/A7K1zjM8xCO8RpHJUiogkT38J7iANhMBGA5xJFBQT+QrQO6Jt+dyOEA/
Dw3PSO30EiV6kHOKjJ4nrHp2BDCM7Z72bUptgKTP8PuIgO2E457h62aIjALcSl+W
jmq4rgBOxt6XbYOytjArNSykMwY8ElhVWclVo7XLHlaeYY9Yh4iQGY2Y628voQxV
mlkbUE5lcUC1kwIGbIkDbug5nIR8StNlVDEDzHyS1YA4Wi7R/n5SS8xQJF9nu7NZ
+i0QZEn6uOyngifXfjh8NFEVy5ohLFNCv+Luuhtsttv1LoIZIVlyMROvRou3woXI
FBF0pL+jK55JN7C6ziq3Txe5xag3D8c6Ag8ChiHdffEXOv4kqb/2SSAof4IY9FSa
/9pTfmMWJk08rBDVV/BXnX01pmgt+8SJizwSOsbTacWKNlJ8taRUyf/XV4v8Z8rR
7aSZhxPkDepN49LteJWpVwbiv6Dl7G0YwLbW69NmafenxXfqiZq5iwjmmfHYG/qG
ojZ+jnRDMH5eB+25JC/NI73KtB9Yw27MODuSJhTeHgFZj5lA1KmiLOIx1IEcRIz6
OX+hzfkl0sfD5BuxNJ3FKTSfkJ4nixwpKPYX4tskaY6NK5X0SonT8QDdFWFXARPK
xDVCY8ysNTfFlBi7GtT638pJuBpxTTiKBS55btdNHlXPd6Ejju4Q08JCedjJhyBU
FRDh7SAf69h707Ym0nZwnoEKuSYpVKFc/7qM/bUI5+o80wSco3UBv15nMeSyXO1K
TCAPGdE1J8bjFhA+OE7bDGI+Yz2m01pJqywXR3IW9uFjIGZG/cI/a2AthjrKC33q
ob/v//NCXfrdLvMXfQU3+jcP2zofm8rg5e31ThjMfdT9vVhNdYO3FMRT0M7e+j+6
eRjCcfCyFhtkO/u+pqGDl1P9x1a+KmV681DytkZwbn/8IJVikF4CQzPFdMVBl8MB
ET9qWAF2gaRw+mkf4GhlofoyqR3vcPOlnr9H991y6DRIdhQJqyqKo005Zd4QvFQx
qVhicgvO8SbA8vKz2UpM5hhsuXHJ1Y6kaqdQoxls41ZnSGGHcTz2jde5gkzCN+1l
x+ZE/nnPbLLUh938OMp07elWmpk2DUaFAWW+7zSdNyTTl7vWPfdVepIxP9gTefvR
zbrlh69BDv/VdLdsgbwpfV5+44RJ39j16mmjIjlyBxLpQfdez42BOebINJeXG7Gh
a2E7IbmQRP9CH/ARfY+BuVPwIsJoXl2DaOBahlvczHwwvbzdInd6qXEq64/YK3Gg
AvGrgUEQ3zIrf3eNU2ykloVJ3VUYCmwyZSpJSYdqESPMgAmEOnJiOBynWLeLzC+4
7zzFnaFylnTIq9Jvs58v/V7I2/LQlvmcpbGWVL5VepZsT+0cWBUAtQYkzU5uLVBB
0kfrFTSXRbpAt8kEDZw7IEuCwYJC3tQhWahxYmvC8LPYyhgvecLxGc1qn//0M7RF
QYF8kxoWgdx/sy73/4vynQ5pW04qBhXab6vVK2PwZ/WjjliMoko1iFg1Zgd/rWg7
PYomwOvCSfDz285S8m4eO6bXpy22Pdwd7AaSi5ZW+gnIucAOANnZJQmFhCWt0cNH
KXxUx7G/nf1AisieCkWMKoLWYqnXfB8Py8JNgo+6nii0tdKZAnL5HoeMmXExMV6o
ESTG6ODlru+iLL8+mxhvoe3+rQ7LVthrPR9O14CCyJydeZUDblPL2xavf7CPkMsQ
sM8KUudqmQtaYwU1EgzPNbZP4jw0rXp1K/W4ZiGxOaMvJxMbOs9vKZXCYHx+1qob
T7WJJ8DzXg6eo/m9hNw4Gc2+e+hqp0QGO1EG7wO6FK4wCVHhAqLMflYdlPJja4mz
aSP4yrHkNwWvL3j5Wo9/neShObb057JsMOLN9OnPMjsK6RKl/AOVONlIYbpn/gs8
K5u91vzFIPytq65c105oiPkzF6vUktWA4BxaXkOj8G5L3LaFoY8nENODxTZ2X1zB
tkpIIDioy+S7FnIj8S3I4+DIX/zrAHWvR30ZR4M7UE11teGtBn92/Re2VWYRAhUY
lwoErhI4LLD6aNzI8h24gCAZojxxU5SCI+qgIMIjnQ/FoNGWy9nc+por30NGAnO2
KBGSonFw3c5+7V/rJCPH2ZMg8x2XH6hCrPB9aUffXhfNPuUYES7wr92FRaMNa795
mAcqnlhbZFaeL+7IgH8+4CzvHBRDZMD+Cb4qjOYS1TjTJ4B9Je8JM6zc1XPiGaKh
2A8oPuq5GgGRBNnf5VRP4PVo+CGKa3nqLOgLwZOUGMp8MJO7TlQeaNRn0QkInnKD
U+obKLuBfkk5D1Ekx1T0hCOrCVkbMTtJeC4nTeW5ywc6z+3hm3uzqVdfmWbxtbqO
kbtrpl/VRGkC23rnA1hgRU+WjLu3qkp3apT/CCfiZbC5hB7TfoRAEpsVv20HWtFK
B8nC9VZzQP6L+HFt4fkMEnS7EJt023NSjfJ6cT+dxrGTLrFoVUmllx0AhD4049tm
CdzwZmu+1LPUU5Q6DNkhLDLsUN4cM75+MteZXPnqeSe54F9/jgu5Kb/mbJ6Y6YTK
vSjJCmw9bS8tch3wra5ZFPG5FrmCUBj4C/Bcd9w0LM4tkyTwFoCb9eHorojmzR9+
aOvfof6Smhp5bmPAlaiGl2+ooSDpNddrsEbvBr6+H02LtiZgxlLYLcRgfodtgmrQ
gl2oQpVtNw2PAWAvKau6qYYc+u4GFJ8xLqyQgZDpsaMBKJ1ogZFL7rdigdlRkc+/
4WVdcmYqDe+6Cs1KrNWBwSTjn6jqRWgnYoSFCfHf/RWbg/99Lrpg9/ayLYDMBc6Y
GnGEEv3Gyh+3AKJ/G7uHtb+pA/aOGbhkfZsiXsKcbHPxMU5IyUzm3QYdLqRBxM2e
bUiT+69L37wDfSmoKICr1jRTO+q1jTQXnNsQT4VRAyy5NA/WiwFGnC6RB9cJteEo
0BxcCDZbp3+QoZmEaY0h01dBv+DsDzuCQVp4U2tdFmG39f5pWLPzBTrJjGcrPMAV
Ymb1QlIsZGkoO4pfwQadgtnKjvhj4nauABNG6X9NL+ffiC9tgkCREeXgwWG0Em+D
jp10TlU+ETue4OZZtVm7w+ouMVKfzU8wMaY6xOuv3v8DGUXur9QbxUQeBpp3pgrY
XlG4X4IA7yX3hlLOAglMI7+/lGa4mucnDoA2Z/WLSv2gLds6f9LL0eHe4gAAWbtk
WsKYC/C5dc2Us1Q2aMjiNb/CD4v4fX5VWTbXks2wkpQ/8BLlHJqOGnub1/yf/gzV
nokSR0lYmKvF/+y5vBNuSUIYn8mRh5wEBcly6RHK1oI8XKxR36BY82fYFQKKj2rZ
KiEvEn0C261znzLpWtP90V+aKvwkXl6U9S7EMMOUD8lxdhXGG6rQzjwAkWlYgLAs
g8g9gNhPvwLihnmVHMylHpv1Tbc+AIxoffsdRYjSe60rfKEczClCnDg8bF2sHDIt
qktcCz9CDQ3hj09M65wk1DiAtUr0CfLhk6EUntT/oy75uKRl/a9jBcayd8CPyylQ
Qk7quS11xgggfKk+BaUAJKVJDNUHIRriAMGFs5pAJKgdVWC1XKcvuYlU6QpRdE8D
SCWHyFxQ1rG0/vgujEKmyS01uvh2DLVqbH5Vp9x6mehBKQTaxlZFEDo/YVo7iJZA
NLuILAQB85bjnMNMy5U4/8bDPLmznkG3HXNbq65JZsaZVYm/TRho+99duRqbwrTs
yo/vC2wQTbDm8iQ7TcU/kFYCVYQLiWgAR+hvdlKr+cR8ifHO78hSgy+h7bSexB/k
1Axj4poQ/ZEWZEhubdMpkqMOQuqPtto7vtJOWdwPPXXtCeHU0CvcM95n9+PYYEmw
JO1NO7ixxYzYekTfy4xytsqsBH8B027uGpZhgpessVm0WwmGVP66ehJXQ//AjE0U
Q77OmSPdt2RN0WeDHxU+hsP0JRyEBym0fYt5x9kOS2buklbCZ77MrG7FVTlrSDir
9UcjIYUAd00DuP7ZpFOTnhYymEJ7EYEhIivNa9ppdAHdgh7HPhwQtnRFgYEsa+pd
DyDpKi2e8UjPp45iR7x5zcA+sfb/6I1uFspJvWcfNcD2E0/eYlIBUOw0Qr/apmBl
LlbU1RyrN4IbHr17Pw2hQhg8q+mDM8LrxTdULI3EGel265Dp4Sk6eJoLGUO4+Xq6
zSjruBMNwXaINVt5q9gujXBugqny+9G13fKOXmC6qedgZc0hszo7iWwEmXjdzoo7
AasWkXj2BCotf2WyD0SsV9ruyiJNMGE4bDhghF6KDFZjiCQC0ysXS20Wt4NG8HBb
12olqW2gr+DkhW8CozJBJlAIkXKGMtDPK8S8jZgxBgbZ+r7o+5t9pwnvGyJUv/zC
Fla28ryVuXnpaE/7YbubXjKwC88/F2NQHQaCi0+yfT5fcMA1o5qkkR2EttPF+T2v
hcxRjlcJzr+YsE/WGokcGbhIySRSVWBFgvGr00SmKvYwt0o0pj1rBRO0be8nSQSL
LJYTt5Jiv6lPkbUfbYo9iYGasjpoaoxmTZR2f1CH8b0fk/jPzaEdwyOGMcNesEoL
Vbe093FlqoDQQqsqSQvlqzUDpBzMR2Vwc3lYkuUW+YMbQX376znoyQNhzIR4W8bD
a8llhi8QO8RY6WAjMG1ODgRr7AUNphVf1jmFWcbpUyeFYbn8J6JLSXA79Gjh7i9O
3iJBsewNMrlJpen9hNLTphdqfuMIsjrlgXeDt/DpsdRz0a8K8QVhl1BWkkYpTz0e
2pPqbgMKt1iWng84CiB4suwerGI2cw+8u5jr0gKT6SWhJOqM/tlinH1xue+GRaIB
dXPgEbA6FaCIxxoXtU5HCEp5Ji7HvHzOOfWwYCSp7PsDN/X80diurRUVoKoX7l/W
HwBoeJn8R1+WfTdbdZz/BUEpJ2CdM2VWK/HtpF74W8E713Nhvio3trXUZqHxqvJG
B2klhRxkB5KNfhLEQrLOwB7mJf7wtOlP9O+HELiE582wLEcLWuDSBxZSiH5FQV94
9MqksjJ+KFgk+cQJwpeALLjnA44rMjOrRzqA40irKc2OQB8hH368o2JOBAELnSHD
KK0sjdhld8Wl3GDazvgj++/XWkHIIe9yt30rAu5ziigl3yJNttAvsIPTjISlXje2
SxiNCfpqEXNVY6do5UZ9eJWYyX3fRl3Yse12ZiotfZiBRGj1pQ6UDVS53iEM0TyS
dfvS+dSh4ct/KgnWZHiZAhZvgc1xkNXulLC5tW0cReKCOJ6DfdUoQI490xi1uZ6o
KGDALP5Y0BnmGSaSQdg343ooFaD6ToQgII+Ts4erBHo0sTlC7MecwxFQBUASk3gW
aErVkKNowTfZ55r57Go1nfY7Gsv/PKktCENism+cQqCqslHxv5EF5NtYiXpALEiI
qYOYxiQv7gBM6nshjzK/deUf8slcveM88vBFYV+QIfUUbpF4FiiMjwMPu+wkgCvX
JQHTq8DBPU91PQB2t7Ep2kMtmE5hQv4CRSi6WOD50XoU6b4jUrsrX7InaPyDftba
1pv4/pVRWby+/U0qTBuiP4pGqqTxj8U9rYBCN4HLCmXt+2zGSfBmhDseoeIP2jZl
v3fEz7wfjajVVL2n2pb9Qa7A4Z1PvdfqgsD3MysvunYYprVBB4UTZGpBBaVvQZah
xLMY9JAqzsenH4uW99te3CgApo3Xwd8NTbBGW5GJxfrwbX4hyG6wy5XcIH8TKwNt
8XDL1SjhiezdAUyX4oHL4XdQ95jnqciHsDwXeEHnGMtz679ticYMZ1Qum4gAG/V2
ZVyaGR7igOG19CCx9VoeAz1IfI6CbBkh4EmQ/YQf/vmZLdSUGWNk0UqGK5iYOahA
LQMGEvRKTUz9ECLWi95hu7PQZGAaiqy6jDPvaKgldThQAq6vGKg5iHWCpXTeL6oQ
GjhEeYGVFKTKJIR4PCSVQ4S6u13tFNqNok90tVqmkepPWeeCdurZLTxN175ab8C9
0vue2M+Lzu5AYsab597iytGjEggn8mtnOToWjkumFjRw+j9Yudac0JTHVtq1ovK+
zBcRpsPUq6jpbu2ialiK5GIY3tkYLMfXqYXhw394qthKzbYEsZE9B8iv/78Z9Ngb
UC9qoPRHX8X3fablFy/gGxuwup16tajMf9EVg6qAUSygoTHf6yX6f97FNlaQmpSz
yTkbYD8aOkdiMAiWJcbtxS/QXzWRdlSBPevFvlWHLCsLK0t6wSIYuA+mhxGTrvdH
JzwuwjtzoNSBg68o3AKKmzjmByWUtUuudMPCLCfHwLmBBSDIdbVKzwpoUSE5kxXt
waN4aDWX2Etc3Gjy4hAUU6juOdbJC/4yUmrjV0QrruUv2NqUuTaTUq8EVKF+jR6j
5REJLlwI4OFiJ2i6mVTTsyCZplCk9CgsBjpbe4xBddDyfGISpMFGNDudcr+iHOSr
ft2Dkk/1/k7IJfGE3iXlbgsWIfdBDMSyoLqXoDndBcJMgoCAb+LolR+Seo72LQ3g
WT3SJDWmdb92Bxqb9OzI0uEHzC9LyZgCoANayx4z4Ef7/BeTDQGW2vgdDSti4dbW
ERrdZbWfC+4Hc+KqgYQhyX7vAOgVfv8DQwrRN23O35dPYZgTVn8d1vVbuOWej8zM
x6iZDtnL11BvCemdcLFj1nHr2ydAt9SIKDtQr7BqiAsvVm/IXsd9opp+0wBBSujd
tc6rEcsUwTOs6sSrGsxjI+dtSfy525eIKc/FwhNQZ8hG2uzlDH17yYP3ZktYl0X7
7tOtuTSl7QuYLnZC9WJDRPrUx/Al5oVvgF2Uy5oVI+0QGIMmwIrPqHhcX0s0qpXk
m0DrvWY6gcc8ADETpOqVWjZvXHVL/WGIdiIeq+EqWbjqrkSErupiWYRF7Udj6dsC
Ce4jjwcxevzwnumeClqhcJMIxKD6Tm+pgG2D2+68bzqvTgsBhEGxzGAuXdvd8LaL
A0feErKOBGFyWM0sBn5l84363T8wzArd6iOQzUX/19J378tzQFICQhOtkmqQkCe2
t8uk/hTAb/InKLFYAnOzNQnuvmxOj1aGUYkwTc3OLxJvjawKOZ7FjudWWgErJLbn
gl5yah/8rSFUYGh5dKBOEHXjRpDHm9IUmJSm+5SXSbIX8Cu3njEdvsxl73n8/qM8
aiY9Fgez1hEY9jh7RS4F6DCVLJIT2PI8z4H/r1LuvDPGR4+KbuwBFquSla3Akih8
nmMq/VJhU56tZpE8aImtYUFJuzjkhyx3mHyYtfdz5GOb+hx/ezvB/svfB9SccXUJ
MALh0By5w2O1pa5z9P6YmBs2CWpPorQrg7Fo69RtpUGICC7AuU8udxyL15XBDXtK
FO0OFRp+DI6FvmW74S1oSIbp+zHnqfnTMeAsKq4+A96KSNPj7U68J7n5sEAkwZQL
a7Geh2NvzLGbAqaf7D3UollQUNFqm0QFy3UZmLeDwOHdqMUUUP4PIvnw5G+P1nZo
/aKAsQy/CdA8P7KTb1FM+wQRHm2+KqLIp8t3c1kM+XA6VTCsD0cqq3YySKRNYaVc
x87Migt2C51sxY2eMyczkhPEPKlkX61kpQs8jqSSsF0zsCU2Au3opJlPLsXc5E4n
b+eWy8bP6cTYPKCsHQdKF/RBTdRFwu2zPGMmj8B561TogHFZYSNHxOmbSKkqc/tZ
TyW+gU0MSIAqKrQiTw5IYIPjnqgenB1MEJSNeKzNnjU+uyZ3w0mT0JrCVr3/ozex
uUSlUkdl4Bb2kNxIYtEiR3SR05+tW5ZdR8gWcu6NSvxugnMwwVEKJJMjNTamlzlZ
qjDXQadTuZNfK/4yl7gZBXVY6U99SegDYcuydzDco3Q8cUB5Y4k1LOb70BXdkDLr
UHT/DE8yaVuoKtlfM3KmkzOTfSNMBTKrEgIpRkLMJMMn5HH+ykBEmtKeWoobLqoe
JPuX+gZZDMSaqRqrAS3ZG7D0H7UgcvoNoD++8BxGlOaC1/sGPawr9qvUGRMkESQU
QCk2EFFlMYMUJY0CxZFAGIwz4PVobUzcf4ilcXXDYqXzW7qGGyEjxUY8fpIt4rIj
UWcRJBqpLdMcAa2VcSQN5+2SZ8FNJSXlb7wkdWZoie98dhygzVn8iV5Nj4sbDemr
bToDsmgVrhPhX0FVcM/60zuQxVyF1RjQLbwkOGYlRnhkxOCDodH0/ot/aHd0qi3I
5Mde85W0YuKJfK0K+lCkRozKzx0C7H8+V0FzT9otIoRAepbhP+TukS+ylon8zYKK
T5DTB40cqa4PyudS4HsUEvxv4+bif9RfGVpSayc2MtfB9SuRr4cZ7u5yu6FJv61B
niT2h2yQwtGNb55si5ilXiWqm3Zw1X07IdAa41Pt/mpbSUwtfq8kLiL5hriLAOiE
HtowAwA9uyF1hvjVOrTt5MdYOMBOnCC6y7gqcukST2ZmgQRzU6babIemufOxO5b5
dRaazuws42KrUyr8kPTEUuqdLRAUabPhdIwHBqUFTY7EvcdzeXB7IP3mpGiE+KwR
sqtQUFUouIURXptlfVERc6IPKqa7uZz8I21J+wS/TnrA3cz6U5Ic+YPntAtkFIYL
+R3kQ2VBfPdrsIm1k8fFRt7OgKC097qnSpGYark3DvtNxbJ8hkT5AalCtT1+5REI
80hyvvp3QSugtPTRjgtNQIsy++74Taa9ju+1UW5fTBnYVjk5MxNhl1+hTU9k/kEO
Rr0Vd4A68nik78YL1qS2GG3RCVb9AXseNHGGUZhqOtkKsobReO6guNW8ugpIz8+E
6zhERdtrSIXcpFUr/Hy1c14Uvlz8S4TR8/aKmEmZK4oXpSOBfPcgfcdC2uaibw2+
0TYeaMdnTfpfIo9t42bVC4LXj7epiVOS9NwZwSZlX0F6iJZDZXE/ITwgJho8PJBH
XQznsDaIk9y5Fh4xlP5sEJx7mGAsJ8QX/3Ibg9swfTlVAnv1/hcxQf8OU/zCGEBb
WYaE+3l8Ym9vaO7DzbF6yiFIC0/uPaXUQecNdlVN7mqk0Qp8UI6NC/AzzWtWTyog
XoJ5lmAMcMHZZUcvcddsXl/DzIvecvbie/y4xv21WD6tzzuv8BhL31ivbenQZxr6
6ve5fTJv9hOyeNJvI/QemJwcUPeAjbWrXz39BUVpFH/dupO5L3NWIlsjXn/hUoJP
MTJffnVQn6RplFEtRnvW8ey4nlqKgo7j7sy1EL6u8FvUpp1uSLTV35iV2zrT/HwS
l+kT4KpzZYNiWgSYuQc9fSFbVJte6jzgL/LtJYfQwnGmcCFhsdwoHMoVbx8ZsoGg
WqX7DAp4p7I/s32tzmThPUguV2stbGDyRwKgzMDB2w3kFMRqJ4lE/hZxtIZm4XhX
4EE9lrRQe/116vk4YyDMEsg/Xv5c/+lxclxDqwRjPKf1DcdHZa5Qit8pEjbNTijH
ryrGXnAGvzbH+neB73KFV8/wst/Oj9AnsHLGMjtOLTI9M6zEWTd8lRuyOXYOTyer
1DzZ6SpE/3/rnT7jOQBMn1e3tzCMakHwAOhrryE/W+cfNSehYrU9AvFnXXXo4sQ5
UP2lKnNZI2U44EhY2eGitPtmh9O3gX25PjjBXjNxsO59wMj1LNZ105sJJbNfRAcL
ei//xdsECCJ17jsJimRAOefsHuLG0aJhFz3kg0y+L+aknAC0RmJp457GrqUkQh5/
PakB0zaM/aW8qg51nOHQJBe8Zv7WBMs7QfoiaiZvMy0dcxnXAs48DLaCwrk1rARu
vw9sWj80oOS6yljOiI1UN6wCXa0StKzWSlige11FQZkN36zJZnbmy7haCVLh3NNs
WPldLT03MJ2BOC6pk0WLM9Po/c+4zFhqSDcrgAcIQW+XM1R9roKOgeIH1Q2ZcosF
ChH5q0PK5kOLfjrgm/8JXiCJcqgwVd1w0FSaM2w9FGAmTUmzF4Y4tOOKp7icOxMF
c6QOMjc/Q5o1zuoKVmvmdbCgWJFn0FS1f79E48DCiCv90I3S/XdVF6DE6NYyn0ro
kO4EscPT7WmxjLafxEN1MhJQRDjNN/u8DA+ybwLbupZtOn4gLqcjKEaJr7sLVkVU
t7zHdjB+0o3vO5YbugJA7V7ixWk8EkBrD/Qzy7/R+IPVzq8keiOfduWp9I5I/3de
oPP2uv8/oDanUwDIBy8luosp68Cmzq4+wRktw3hH+wPuRqQFv2CAw0bS6JrIvOX9
iC/nxx9qKZHLGUl53tzmuWH5OT4mBszZjXZIkMoydnZ92oXYAlo+HJEtaCR7D7en
a7aKAOIn/MEivmXKDvRAG38z3qHVHIxJ+4n7z4UNDA55FXxjjU+hlU7bHgG4rNCT
rAyICKA9tQKOKzvnk0wU8OIFgcpn45ZDltWVtZj42M15z6IpAJHwk7qqzA3Jh6g/
UtRke7WisYfw5B5YrV9lnnb1Hiss7f2HbtW5Hw0IyulETSkBojpEQWw2Q0IGsPq5
+sUtlMil1Wr6gCfpvfHpvHm+G34WbA5dSCn8OA+cxqiJgdt3ET5MMEvTO2uTmKqP
vu9eygAruNytt+AnpX23V8Yu3h2dNMylaG9qDtuqFhFE/ORFOIH4vEV03UmBaj2Y
vziGF1wwwZrXCoSMIO+S1MvfSGirOGdwi/zzAThJuX/zMtN6zLyQNmpNxup1bST2
OzIqeUU5JHWoiAK1cV5bLe8WynTK5s0TBnC897O4mVWVHrD5AiU+TdJYigJLK+k1
bOZI4KawmCVlIU5AgvqTMsHgFIb6d9rAOkAFi+jHPDwdrO42m7H4HAvZULG3UB+o
ah8WXhLuYvo3vnuLYuax7hlVqFBZByLMgyFM2WdN0C24cvrKg1g6qGqMwtqiiJr/
PGKVecPi6hVbE9yRJPdI1x0G6lyTc9pYaKbtn/OP766YjqhZ6H66ifbL+t6S0VUo
qw27MFwnXHtXBc018cIJGSZzts5yFds2wMYUHr6/uxdETf04MnITFd0qAaQDrVg4
GjTfRkmIEq0Ises6RLNUM159r3MCtFuMwELGdzTWHHNAleWzlHu97Z33mZdxm/kM
E1zh0XBeyAELaXsDJyzGXFIeUQbSHqbXB0EVciRLQvwE1qiiUadZ+fVRFOARLOd0
U4YLAofw1EpoxRBUQHFVJnwzKJdsa/gwwqrMl3ys5JFY5N9nRQdeuLL2PxhKolYI
AzSVTE6q9OKlIMPucPcRjN6lPdUirz3VOXB6cIGplYBGIfEHapCX6ruaxpBz6Rf9
x7lLf9AgLtGnRchUdkzSfnNB+ZrwsD+0d9Rg6w6WkxNmsmfOsMhJV1FQIE9Oui7K
sGRfkSeMuyoOHakp68Ki25H79G+oJkIBbow376O85oiUmoF845NGhDcN5Ea5NtTY
auP8DlWFUGv0Phi7h0OSidA5ZEZZJ2bQKOQOAURWVb7j/mNA8/nP9+7q9uvW5l+M
xYFCcWDD+Srjcqbz4W93fH08XnabNdyCqcS9UyMfnTeYSbmQy4CQnBHJq41oIKpE
4bBIBCVWsd/Lc6E+f27cO3KmHs41iGg02KyfQqWD7exhsNS2HR5IOQu6cgx6dZYt
fB7GXDLQTFsT4t84Z4OaL6krr+KcZ2w1yGFiRCUoD3ze2PbQAlO+5vEhYDk178wf
sCsu6DzQj6+Bo2C4DktTCSzhxlFsZKsEgIpjDJ7xNt8L9XCMgQZhJwXYzU1KjSEG
b5Se9sjeau1UzTNFZyMRvY5mVbSXlZAym+BCBzb/QtCLybutcTUbTYgowQUzQ9g9
RbULm14/ejabbWfVdcQfTfRAMr5kRjWbgjCqsJtIoo7xDY47oPsVk46+fAHRmYIR
YP5ZPgap3pLD0855rXB1Oz8Uomr3/dp1/AzcSNv5zC4aB7SHZIvMKAAXaUOY2H4H
aejVl5/ToziyRSeo5YYT8RFED1lyOd6iklrAme4eXLL35YbOq0aq4Rilo7XotUCM
eSyk0djjELD8onMzIe+q33ZPGENJCazAauLhA3g0JoUM7ZUkj4tBl4JIZHBx6hie
KG5tlCWbWczeAB81B9ABbbv0LnhDHdomJ9HU21LNYD0fPOKONov3i6HXzxHT84Qt
oXbSgkD3p3M77r1/t8iim3KSwV0cLpzvRDrsjxsfENB2ncFzonz8LUhDbhgSOzmX
DN0nZxmWP34cmp7Dkjh8gnuFwBgjNYw7Dg71BWj7hD8wy4I/9Lp+vbVSL0QoXhRp
bnt4YgFNbZ66DuTN5M1c+sVEmqED73g+HvFqF173KOBP11F/HvRt0QB+DYiLZJAq
PUi0+EiiqOahxrzdp0t9TL0ORDAywbnW6HyHoxgnArEPu2OY+CiaiTQ06GebnzsJ
dZ0CHKlBMG30heyouRslN7FBf8CX9ZI5YgATV2lpXfLA/EoU0M/utU3ZH+B4C5sx
2GcozDFiax0A1Vsrn4kwb8B0sKQgcY3wSVcQ8kLTfv6+Vjqcx8rD9TGb9BVC1nMK
+5VfLKlRDRSSRwb4X/uk+d0Og110w50Hk6DW8+tjx5T5NpSmLIebdsnRhrXqh5ij
ie/vFQX1G3kXfRvgTkqcEbuzKG6h9vtfUZat3FwJtxo8iZtlgENqp8difbZASoNy
OBpP+VYkBygRn9PLHmXYiimtqCXQdWfYiWfLDeuBASgvkFyy2bVROAFldodsYgu7
JjXmbJ/e4/r3CoZmtI4/aszWOVqycjurUIEM0ZHbuam6q/moJR8ryzpRzmbh1Wye
sb7ZG6dRSlQb0bFD0orXp2b5wZAKdiWw1lDYc6Mdj508pvFtmDSlro7jl4UFDzr1
3KRh+wH8KOZAx7ieaMU0u1W1JrEh1/jgW9K9BvOx9eJ9xwpafiFTG0qtno5VOQXA
UtsDtwe5XGwjfPU2R8b4SRIXFXRGRkpmYP7hZEsAt+5fpBY71jQdSZnW6u8gfdeR
/wLtq4gUaeheDzWB37uQcvcLMem+G6iKm7qhdndmVZziy+YrmymE2N1jbcJT0z3p
YiKCcdo+hQWwcIjNe0rk9AHGsJPbP3f/pPWgn/F9W0DN6a21NCl+9sst0ae50QXT
qWjtdLbfhbkTmFMAVsc98BUtNYyjViOFA30bnX+OlyvQ/WXT94gXKZ1r1788Xh7R
qPQdCkMwhZCVt916CrtV0hKn1RP+52EMhwvBg81G0ox4Pd2ftsZUMe+KIPUeX2/z
f1YYPbbETH3UxbO//e3ePnEGCKtzuqAf3mrTAXtY7056UMk0MiPd7HgJ/QSo3Zdq
/FnSeZB6UdGuQIJWvXV1aFQ6s+FOpUOdU9+hhdkbwbQ/Qcb8L4mtOBCwbMsqHZ7u
QPFzVqZaxvDmzphWxj49hBINOANUdtOMl/992HrZLR4tW6+35XCCzAZZVFkKQnmx
fIGhERhxZFVhFcJNpPqzJXANiuYpJCASr+yQxPD6q7icrG3ADfIoWGH/YP8b6X3f
WM8u25X0gHZkMKS8Dm2sKAzUl465pJM6SYT9G9VeftH0otJ0H9kk0Av4WXJRfxDm
VNmpBjVhTdQxh+q7CxIk0rv86bwAWVko4lh/u05jRKYIqDRRtpcfapj/hhM8cb3C
7Z53ilP6OOg3CiuB3rmCVS3oFgAbxnwGOXGcdfp7TCOrtPGK2gTlg+G7iZ5W4jny
irlsXBkoomR+dNa2htm12dkgLKD0W5cG4MCuKhln1KLGVJ2nxsFXgNoAKWGMKUEo
TfyzTKOhKmofXakJUlXdUbuNnSjzayTD2Z18iYNv4Vh194JBGJJeC8aL3PGU1fl4
HUJJ9IC8eSjvtw9LEzI5i20aOXEqHVRwWATD9Jbd5hYrdCqGutcc+jAFfq6mAExF
9guiptplxMQhHbY15Xch7w7kMReMKERHNtLQHlUUPMMQuDy2k2IJ/1TVUPiM4bEq
Z5CnaQwXUM0wARmsVqDWGTP2n7uwOhDGGPHskx6NO9HuL5vDF4VH2ozvYyi9rLnN
ccbsoepC7SyOBEQGfbQR+iGRF9iXAcIohNudSeH7GGHte19Ews17YDXl58HkHYaV
MI2USUZMWekpJs/NYWjgV0xFeICanrZyoStLLfLFFJF1Vk9SeNl/TE5b/RwJYvDM
tM3LOwYCLdYwuhrcrfkgG5LNON8xOe/BVTbpNP3oclxsiqg+eaEWuP41KJAY+AM0
KYNxR4v5G7nOWoi6fhyZ/KjPv9TeIqU4pEXgRDej0MBkY7A2dosPRN94I/JlRNpZ
M/TgtBo2C+b0TuQVxiBmZDv25ZlAjPNG7WPieLS0gfpLJA9JzHP3FL2N1AGx+kLf
2NJK4lWPtztMKYYx6Ce1HcyvHtQrhd77NOhqbWJoIZyp1G7kgaM1gDkKX2ulLh6G
BquFa3gcJEeLDBJHjjukspdTDnuahsjL3sezD8rqoOlHa3aoMLHHLrG4FbFVwqXH
d7751nAwmNOvCpjxpknzeJKqAnbGqJnK5zkXzCzXfPigJWxWUOGGd61EmIUGFDwB
2pD579L5nA6mXI/JSCZLUJD60Hjixg//NcMitgrrEuvAt8PK+sdlosmNC4znM/ZE
fE6fpFRfvI69/0gjzHYvef1JnPOFntG43X5bQpM7hcPfhyzKB53t3+V/b1L9q1ZG
2Hc8iJYvoE38RFtQFy9IO0eSOtU8Lclqu2ZodOnkJHmZRDmlgZbXHA2Pepzyby8o
GOAcP9w4Aur1GqWMENkyP1PmHfsKq2zvw8WKdPlXRKQpDjbgDwZi2/1JG/FepVYW
aaxFpVr5NLo2vrFZOHB6UmJYsGrg19C4r13sUo6rydtWOwa0T4gEvXCGwavJHXO2
NWpnU+mKYA64OXC/HboRMeAdxKfD8wRRGUFXk8Fmv1xgL9DHw9xwUG9DGWeOb8+x
cLTYQEe7Q/90KXB/tbI4I9/3PqQHXWzuvqPigKstVaqYd+sKz+qRZeNJgQrRZCPa
XnpdpzGeXVj+i/pTlqapTyDK4eAKxrdoDZ/nNKJMcjY+WsscmC2glpb4AKSXwzO4
CnjU8kO0wix8ZB2CW6Cqak9n4D9wRjDdr5Xs5LFVOlawAVFR1CQA9kdQFwBnN0cR
ZiHdeqGTiDShU8BwNCGMWakwe7mKHr8OjDDShb3vTpGerKFMWCftftcbeZDA67Fc
WfUK+z2vvaaAHMYhY5Y+3riPXnBwyWS55vBFHmTMTE2WBncD1rlvXg0nVtjJiFAC
7ZWwZwcJjh8eLw59SznfyPqLBkgaX2xeNxfF0xwpoJiqC0Z/5iXyEe/ZHFIKX1BW
UAGIikcE0AJ1QkkysBeN8jCgurafXfPbT/xcDlCglFFy2Gf/mmRiu7KrMdlXRMLf
/ad/VwlFQ7J9J/Xd+rM+rQFsKQyrGPc3T8MTCiT8Q9oqY1AIqWxNI7mfxMvettk8
aGLr9f1n5SqtGQ0zfzFPkEp0GdLoK1BiDKiFKjJpcrhBNSyc3eSn+fbJJcX2np5x
U8QRTwJOCYIoYUB6CiiYWR+5QHSPRb9AN65pwZx1nfYO/L8Bl3jnYV2km3AY30ET
AxKAMCoDhDxTKPur34n3wZfJdILYmWE22AOSJehi5KhwhMaNi0umxhwJBsnzjzC9
TMZrTNG3E6suNIFaEYI1R6J9SMD2kiaEEZF8WPwaON/+26h+47oKH/LC7W2oihXU
a22V5uj8ouSNJugQy7AwrvuhKm9/AsmDgREO8/7tvaqomgxXytBIExwFMkVv3yNh
W3YDlPSlf0ed9GJuy9lz7Qf//dCug6RCMS18acLELBwstiSGEclr8YCZB/YvffLr
N0FSSX4agZN7IRQ28hxiU6+f1VNC1SBEQItAj1lcGZepdUiCT5DfmgjICsYncbqi
XNdg6ijS36cazG1tGark+R5QXBupaz7If7zD75zIj1uv4NzY33oHAlziNQOsHbIF
K6iwwbV7CZ9cOOWNgT7uR2aKrJdv4IfsUhzx3GbHeCByzbc00rf8HsJ0ZtGo+31y
GRbuK0XJrBYSNPzdngj9ZGBvwvBiUT4z3HLASo2oZJt95t6PVlAxWhHBjXFGc8O0
50tLv0LfA5ll6v6PEFX4ztXp7hnTbQC2u0m+J0p8nIcdY6xRZ5vlPb/tsTC5rxho
e2o1HtdIwPxy2ZXXco2bAfSd9oyFCB7OMPUKBxNRKkcSLs0y7n8aaO1NDddBcBGT
V9KR95dvmsbo+Jl4pAcjYR3qOBl+GG7THD4Pb1ofxqfRBeH32Ks3BJS4A+zYy8yV

--pragma protect end_data_block
--pragma protect digest_block
nxEVpzdgJBV97nJqmhcGSLUqg8M=
--pragma protect end_digest_block
--pragma protect end_protected
