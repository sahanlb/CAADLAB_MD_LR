-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EJkbKNH2QNAA0sf01NnklseD8u0Iz4JrbY5BkcAy2A/FqgcKnU2tUcrimK5w7xvuBGUMJmRBQm+I
Z5jxv/DkVfPWQmhcUPemlz7O/znRl/bqBdHmfMxzu6MqG40TsnpKTyqPF6akNY3cF4aYliKZDGCL
MHH0Dpg3vIbaAV5QI2ZFhjeQoMdAPyEBkcFfImMYOIuvV/EEI4aYlNl+5keSXqsCWBx0aU6a6YWJ
g4JfisYBMM39Fm4l4H4PU9I27S90fxWDGm/1quLkiRz4rqttcfkjFKAtZsqWqrDdaWRtPQT8yk3M
Rao34P5Ex2Iyy1jVu9hw5ujFqmsYJzbtAifXpA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5200)
`protect data_block
dPp9iJNBk8k5OvxqEYhgRMcvPBqHx0jfWxtCF4Xv5aYsP4QovZivd8HJt/9LHMxwv4+P0gK4EnCa
veyG2jYhhY3IQ9hSdRnJJfnolDoztlOTpv4yWsygDRTV2Xqq3GUAeuxpY64yoNdekbpK6qdeQFwg
0lNRb6KjBeQ5MWlP54k73eq1kcS0h6aNFf3/4eUivxzIIERFjZM1KGiyzcQMMOWKrYBKsru6q1iG
DVAxTP5MWFfPTTm03XKpOuIPDx6PIFBMjHsw5CsmBCJgOfDoBrCo/fRZDNpFMMVzyce1ZwSuYEoB
Ce+TMJBy4vicvZBrnMmdE6QkmYAUqEgcD9bkDJ6eJiKwvtMF7KvoiDZc8olL9Xdnu8W30r4p6z5F
+0YsbtqiP6sus9KkIL4Q9DA+Jny8dyu2n2Z3GxzUzkZQJT+hVm1Q895Cvk3tkKJ36MY/uL+YEndE
skrAe7j8jJhrrnMhqkvR7eDf8AMCF6OC5Uit44XFaSv4W/ZQ8krfMOtS/gr6j6AKlr87DB2F9YP7
/ti7qqlG8Bi4Ma745bdHWkv8JsE6WSS3n8dzenX2td/kmL0H91Ha8EpmqjfQPwPcCfydtNuW9m7r
lA6Pwg1Yb0Bi6/6pLMgB2Ai50bqunQvsXleUlFYWIAQWuqrScnpWVM3gangWPyQuroMYYJOaGvHU
gcnllKLL387ns/JBChcZP5fTQUIYkW2dNrzqkOxyfvW2pJ7TrgfvmoZTOtk6JXIKuhGx3SwLAQhX
NQ9T/2NTP063wlIhq80Qy6tGDIFYOhL0EvBwQdNsgEcWnUwBc+GqkTSHl0yP5JcI0XWh/kyYY66e
9tNQk4TLU8EbZT9S1PaslfI3g47vLahb+aYCqsplKJNV0fx3dSHxUp2Er62/tv8lDPAqhyYCYCk5
KdPhmm0Tw2kufT4k2VVGidItJ2eulXhU8UuRbdY0Jw6PA7U1u7lrN538XYDQKd9UIyeNFPZwHr9g
AMvRFvH0R/cADSmWa6aAYRYi4JjdrUMFQXXzuf6FUpas/4sd0v5QeHN1CecKF6I98AIu68HV/pfC
8ah6zgYRyhCBh+txeYqz/0UgM+IrIk5M84xqEqsshLyfrhoAOFYwAhko2af95bs46GK0TV/gBaZh
Ei948ISxsbu2O5Mpm+3mLH/YRqZszUUGxPtBVqrEuylzWrQSz48txTqjk2V7eJM+HuAktn0lhqHV
twoY8+tREr3xxGY8skfQ8xt7+/AieWbXerzl8B8eSNx0Pf4ezJ/AaKyz9RWukEW4uvfsWzLp1shX
snRysIiUKQeIoLJ6of1MV/MlfBpl2/U1eyw2oAOmmv6WNfzzM8VoPlpBqcFzjnHy4hXBjExZVjG2
g7WE/mrzsASrv51p/t/Ng7b4HZMcweDejKotPdI6SzTK62Jjo8EIP7VKxHyumgNIKnyHWUGHl9ci
JEslGDdog+ySRbKAlPxz0B0uvNZbK+XiSHqImMZk4oubZgvTcLipUWJEg5Yx7/yKydDsWhFeBZvw
xjKlkGtKITWKiZsXB2SZUVSuya27+9eiOTQzGq6tprO32Z+7hbc4F+vru5gZxNa2ikF3vNoSOxW0
+95eLGaQDaGA9K/3c9tvBtJOkcPeaZGcxoJr8FtEUz4/0hLzGZufxQ2cE4Bk8l+J0vfAsbb0t38/
iem87Gz4974bhnTa1Y91KcGqel3kwkzq21wMt8yTQotfduVXQi9d10wTcrgqpReE7ZookWwUgFOQ
IOv64SFoWMjTriFGW7x4xGQXgfpwFCA5MDD87+7dTzVuV19MEbpNK2kBjJpAu9mByrQ08OdACR+8
MQev4rsiH818mmj55Hwf2wWj3P+EJT2Trj5hgQIsDiwoo6raZMlLupSgmDWRSQVAQ1qNHr1HIrpi
ImMh+dBB6d32CYoKqoq15EW1kAILFoXWTxGZdYj5SFmqR6qOx44Rtn72+b9/5lKDFVdR0nv3CBOg
DJjliwKxdRgDYJJvBTz8uiS1JXvHYnmWaw271EKYyxiYTnHHbd8/srelzCpZ1NCUJwy5WUfaB5ax
9n53DvLeUhYq00IR82U2yPJM9JSjmFdVaKp1mVUgrIOaI9+Vs57oHsRumQexYjLPld2nQf4FEY9n
UXWfZw/uIdj95K8fvl35eMQTzNfnjWcnfIbBeq8vbfE6TS4eiVE3UtCgGnUGzguH+JeBwdKiz0rA
HP0Z1hzL+327bFqWDAUdSxNOkqk1U7q2qI4bTcZqWAyltIVpSaj7fKHSTLReKM0CfPeDWWLygsDm
fLH3Z1VHrIXOUQ7QoQsL5HPS6LpaK/38heNJhj/1BmTB8UzRg7BlhUCl7ooBmzp1PUVQ+f7kqS5O
U3cTXZqE0uNHpOFNzngnYUbJowm0p25HaUohteXr4KLUZR1uqX70OFN/QNn4t9K+BT1m85PFR4a9
oNJgMlXR5ojTjlmzGEdTQTAVhC7roUfQOVHqm4gz0bYJkbAfL+L+s+UIzFS42lyRSyRTM9MGQKgT
I7b23eBeM8gFBOjYcYzkl7jEK6gkmZZ7XmqNyWKwgitVlMuSHamlFu0vDCTcmPfL7Y4cMldCmzQi
/mR4WEtRalaObCn3UfUFMjeKCHMUtYzpFCRUj77tGjA3VFQqte0et89Y+YHM9RedEf7JPV+dpUxW
4HNckRU9ob1Q3j/+fOlQCen4YxFkdFpD3Xk/ZCwQSXO5g4U7wUrSWXGGqPO3eJ/8hNT11tHk9n47
9jJtb8j9oDPEM6XtjbNtwFGmTK8WLs+zrUh7KavV52SO77cNxc4PEAsSPSr5w/Pm5gzgURfWO1Zp
i+S//Dyd1n2WtJJgxGBSP3daV1UcSED+bzbSS9Bqb6Uns65Mo/BuQL1Xn8JbKft2jaPj9H/ZMbD5
pXmbGHOEF+J4iAO6R5Si0vaq2p7pypaFlEpv2ZoqDyoLMZtihnrUpZSzDCUpJvArumIHpweqOX0d
hbU6o02Fkw2Bz5FG1/DrTfEBiQpK6ycmxUyvexK0UURmLoT9G0fJf7+OB+eGJ/7DW3fxeXPdrw9y
F8MHpGoTfFyOWTvz6g0AUCLIr+0i3hjhrjDx2tQpKDret89VVuj1raPyOpzmCn0k0K8wyuDfLHXi
TrpY0L4pC6/4unB7KbdQx5zIsO0IBeHTIFfDo/WalSpPZ6wno/c6SwHJZnkNyzaQuKAamnlaNSxZ
grWJl0pKrsoLys+6rHFDJPQioTTGVQak6Cg/CCwiPyz9CwwiHE3icRxOlRAqAJJRJOM097w5M+Xp
fmoF3NL1uZwwV2kfO3ctmfHtim0wabPW4tNU9eMXY/aERcuaj+0jeiv8PHJricXd04afYsmzrEmt
5bmKdvC7ToA8cUfD2hHv9wACJ9q+bx6CioJQWJryQx5nSyLvjwKtmbK8WAsBvee8y8hfZPDNtX9y
jvebV5kr41ro/XjgnlEt9zPYdza7HPRE9SqgH+pjJC8QEa4Qyv5b0hnfCDxI7/BDKVUmG//R/PCG
1qVmxEYqSNacMOwKKeAZ8+4jZBZDKj/9pGZISE7uEtpd6MywQ14KG/l1bNacuHq32tmAXHyJ2MJV
BrcH+d4hvD3Hqa0bgxkBRGEjhiCYiefRWgtpAS6J60H6t33711FeeExEycaE/iD4GiVKLO0ROEfa
wOVIJkYqfDqhKiybdO0YMt/p37rObqK2jLLViTIqoxEPlQSvKpuyRpfRJor1JS7yMVQJl4OtBm5S
niAW+BtdC7nw4xPtwW5PlCJ3Eel8Ik4Obm0hbwkgJmUacY/RLqIzIuFu4Z7dNXzkB/0690R1TZjr
cbxo0lHg20sn0yhUapzXAXWmPY92KBdsArj/MU/tPgyjxRNRQOd0GhEPd5za667GvnDJlkzVcWDJ
jI0rvePXZOrVCCLts57YyGcSF8iAsT+Wqd22A8HjfT46/tkQZ5u8KRrz0L3exH26V5mKsk3w+ZJb
yLBpRH7ZUe1lSiuhqgUaxCxPYEIyL3C/nUTWz3DVjKyq5cXVfg1n3G2LAfVUNQM3+YJJr1rC4X9b
lUKo5pHChAPrOCrpJPNI2rqaI9RogR14FTt84Y/VnoUvNoonvYmQQsTAw84a1rLzTAcZURDAvsR8
SwZkucrLqhtsFyp30+lzKxW+udlLwYUrkOOphcOn5xCFU7rI4hs41uglVV9ORVEJPkHThayz4Kk8
3pWj5sqZC06IV+ymDSTG3Q3zsQRe4d6JKgpqfv3Wcefgql9EzddjVy+e5yYAX0qDBBiaLCBCul1q
L3c6/wQ5YLpQjYaBYyku8+lyErrfeN5xOb8gIn4UsPPYZCA7aEXmUP5swgTp/PFE/nqenK62Sq71
BqxFgzW++PXXsX8j56FF8Wom1rSxUSpAr7SEcL4L0WHsJXi91s0rKUic4QfIArRGUr4puAw66sHZ
rpQkcBxLqekRp+V8IztynVQuB36rl+cPisCFgQGP8ZexzeRq15tVIyCeFOjA40TD7JzcOgjBlsGj
hxrfGljc7sAP+8KBtkIid3JxABquaZGuf3CEuFDLgCQiAL07aNVdhny41GNUW5p79xVfQeHEM/bV
5JCgKeujLnOGx1bjfvfgkFAZRh0AQAJMlqxOvQ9fowX34aQDt842memwT9E5bPXBo7nPeS+K5pkt
ivdOt1S1OBXS46uWqLVWF6DoJ4rVmz8JAbnlRoBpB8/qe+61FXbDOlYzMet4ssHEL3WItxTSQYKP
W+Biy+TN++vhyM7UptStd6GJucP0feuccBP1mzen2OmBMSe/aaLW28qOJjqwQwZXx9fv9ItszghK
vGlyPcxt1CFcQ1VGk8uZqLL5lD1JCTq3yQiLU0W4phJn5Mqx6x0NDma+0XNyeoUhFlF2dLQvspJN
dCZNOt3uHeMPdJ8CMFlxf4aSv7JkNQmfYVWwnuts6BZ0U75ivWrjlQ9x/zi6fhkjZLQnJH59HK9X
jfcepxBiZIp5bIm44waIIDU3r+ovldoKGIcTW3n9YL7bNAQUdm/3f4tLxNm+7kbyKHt6GjFX2akO
fQocIlC0eLl1dkG7DW+7rONQfQffkN5t8iJsbwg2rNwmxtG2FwOMI6RI9wixxU/nDgBMvz9ZvClT
Gja+ylG12EcvLh+KmNY1ML1j1YTdLsIfhiRejyucCtVP3hryzDM3yWeHk+y2hblSmZNTa5oh0Vw5
Y1MvFFLKAQsmv3mYSVN9RILkhgcxy2YjKC4aq+f0laXf7NxDWI8jSGg8lKUQ6Vv5Gv62HRquNQ6F
Uhbdc9Hn0bBD8eEuL2EjFtQsOPQbyNwL7W3Yh1rLO/JwU9UcNenIxMTc2YIn66/Nhf7J720VSK4H
uE1ax/bqJo/6N7NrvKDH7l6Y1bCtyorEBUqMQZ+6BeZ+2Lp59VFCzSnhghYowJYYllFWc4DsxJ0l
W9k3v6kSehg7635lCJa9uyH/YRrK98b/8A7pQ84JXKUspYLnEYfLUwJVYrlIaC+AqtCUIaulrMs1
pIM616cDlKHdLHnR4r//Q1nrYekf3I1khqdIeVPoL3Z034fN4OMx3ZN5d6sBCc652J6WnHRBy/U/
jBAhIaDkgkCHZCcKy6XYAlMtt6krqGmWCyikqeF6FCXscv2/UCi1VbguwvftpJbeeMPkLrsm3fZN
J7BnFkyTD3486evTuuOAVJ9weTAVvuh2OY8GprZrlnsEU+UZskY1AtVhr3jFUHA03K+KvUPGxoa9
3r/yTLX4obmPMuCTY2gN/TQUJDBwxwI6I3RTaoG0y3026j+Hm3HvtVH1s9xLzLey1UBPPEGxLCSE
LuDQPQQV/WPT/DPNYeOcQVSw4142Oc76RtC81YQeKPOCEr8WsLElXXbkreK3QfxQeMmi4ci65ppY
nQ1SiCSfFFjhgsjozkNHRag5L2p3L+e+/SbkxTsJwwzO59gGXNtJ8jkdj1Nxu8/nvfFVl0WK+lIR
uZrkTs+c9KHDeN7l8pT/iUQNAYqVU1cXFdSXeO+pK5LZXmkOX6/Owg2C6UgMvR1Qb4bRPV7r70wm
DVPU+3foIxrLMt9p1Ar8HoWzNamgu2UyXHFYmLzVcRTOKkgG9Hm/3w1/CSItYBwj3PrVZEjMrpOc
cLLF+kkEX7KfppEAP2bab5ugvEp1sq4WbVf7/M31vTIBpCGS0FHAPabZdS2YZq6n8hNe9Mnv/3WH
/O2EGl3YEty3Au86giKpv8b4XQn/jG4kdRv1NMs2TzCo9/lcQgJimkwWqgg6YbuvTKjbFS/9l+Ec
IJ2Aqryw4KTcekYc13O/17srW+dFhGIm7w+Nsf2IQOw37iMDUVb3z1bjCfiVnrlPsdkjT7QwhCzF
8icYCHVpd/J916kkIIDp7frj7GwTk9pmQOeKhexODIhufa3rIgsjNdA5tm74IErqInugScWEP3jT
3rerFvfWodf8bORJcA2IOG02j2xBTbYtEDZor89XlHbLJxfPWSGhc7oSpL4TQN6ZuDRN8e4RBaNY
Q5r4HNTFUUHyt1iOTjz8fb6Vm+9dXlohazro1xBTqZK7FhziFi9PeR7BJEBh0jwaDx1qaDCvGbhU
EJqicUX2zQTzNjbpopttk22fNQekKKScohIsnFaHllZZi1cJMjpUgrz8raBAETPkHvt23NBJzK7J
p2H8dm0Z+RZsXzvRyzC/XIqnI8PiuHnHI2WsgMgDJpahAr4N3frZEyRvTPGQ0H4AGPdJ7PcTxS/Y
9m5tGot6vEPjbXN9MTSeAjACB/tXi1kFPn6fZk0Eg50a0P7ZZXMmgaWmftU3Jb2HQp+hLnQMar7Q
jOSl9brncW2pgMsuXxukDPduD80UiaMtcJPLN3cAZ8x2cOhFxmZdXkntGPocSgbSESgLi1mBFTqa
X6F3ZLvnLw9USliXZoiyBma6lxQDnfuiKWAJ1mEp0cF0FLT2OVKLg5vP4MSBlcrR/ZnY23k4FeGH
ZDNL57Ary0W81OrvZw==
`protect end_protected
