-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hT8uGhGLb3mcCC/dQpPcKnWbB0745UzNM6X9+6bNDn7ARKZDvNuKOy8EX58lKkcnGJIbONDaNBxq
66zhrmOcfO8i1wgMsBc5f9mmITCA07YkZHmF7oPeX8ehBB0JYID7QtVi3wdCaq2IC2gjd+jD6xqT
USnpYbAKE9NjtquL1fQYxZWK5pql4Z1FW7Ne+ip37vVBcEZwwa4OfFF3S8IRpGvqNFL+Ulipj0qB
QOTJgkQOl01ocE4Es7nSk7UkjvHZvMgmfmXlzBGOGNWnSLMgE+pfkzkwppLSg0DzvgRd+keah+cM
aI5//vgDAPw5bNoYNBNVEeuktDOGzl4Kxr9QmQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7600)
`protect data_block
qpgw5cMiqJwLb56ig0EwxAJb/Ju6xlOt7GYRX6oPC8Ya1VY6pMFqGxRX5Skvk5bGiFJJzKfaSJSb
d6n7dY5OwJwtX4gD1qaF4vtLr6Y2fMPXQV+/qLe6l6YA8am94PjmgZvnLeTX8Q86DTAAv/BeAJfX
4T+eYgRUgNSR4Xa6Gr1VLrgQxWDfenFzo52+evlxScAcGidwr61K/HI4mMaJHEDUuvKFCVCuRtXG
5L6vKHT73vMQcEDOgnw5rUDPrMk2M7FI7C56USpH6L7cVOOxmbKzHTxjCzbs1ICvUThyl7PTFPlO
zTABp8/QfvMWIzOTtyQ0JwYE3V2xE4wwDKE7X0EyTVstt8dS4wRwjXgQ7LEzyXc4ANETVuSW8Zl6
fw2+LA/IQdm3BuVD9EfccrobQrtqE2xQsfiWTfoTq20CzRnNJt0gOUE/Msl7hFPBmStTnh8Ue8Z9
BPZ4uuVcLmD0EuWJphKPxBKLPApfPECFdxAzJTDQUZgG9WryYwzYZY4KlS3V6jobSwup+kfE4j1J
5cS5VILGCDgF3LbtLtSUbELgtjroYxYwF7w/QybruBZYxpLvGpi7YAitf3WFay8joGx89p4fgWiK
7A2mEZSc1c38WsK8ipTshGE7crausckE3qeef7bSDDta0O6+XoPP2vkB2SowT8H+4sfhDbqFt5Rg
hxjvaBuyib/Qbj8AJSmkLu/xaV8swsFRsZ6QJ3OdFTDG/LqShyb2Tcy+wuJ8fzrhrxN1GqzJ91t7
grkKZGV/8w0bkgU0V15XNszznkSxM6HBIeDjkzLl0nOn9b/FZ20Q5L83QyJDEKVovtZPlenkxcCY
KRc1rvlNPHk+gtCv3o5iD5f8lJ72R5O6Migm+o0g2+EJFNO1c5KqPj3hpddKsLdmkXJAJH0TwdJv
fCMQIm3M2TnUQqihtCFmbMupM/Y+ZxDLA6qQIWfLbBrG1e7vwXVOAhQxA3N/cbjh5iVeCx/CzW/D
T98kWv4JOnpNUG9D7O9QQN2MARloedznoozv0MEDjopeo416O+zfzLDPeL7yfYu1cvdQeVLDSSVM
PQ0J/kniJH29E90YX9Y0hCMO4YoXuIcZQzjysfuiGWutptUR1Nzni8OvfPeBQQlCYPqvp5P3Vluz
xdUs0Lano6/HSt6Y+l7dNZdV3YFkFM78G0KIMde+UKikYrzjREBknJS/Z64JwxoAbSyzg8YWoD1T
FDjlEq3or/P5iH/LEbawNf3dF7Yyg7f9Zx5RfIfW5qIK7PD6V9U59d6/xzPrlxe/7CYPK0NCLrX2
qppUBwLfZX4ng2n9qzIKR3BUnAPkg7jzAjOPzS+eRs30OxftNNyphNCr7zKvYxWJOQ9Q9YhW6uLU
bSjXCEL29aJytwIrqqNjj+oVayCN7RFr4eTckbMs7la7oY9WeekDGigs1qgTlRXljNvkPghIRJlh
UoU3TIk5kQuRZ6FV99r3QBZ5R6H1cGvBDfLNpPbjkE3ex/ilZeRpgNMAgp7PsFw4pOrXq874ksad
69yixHsz6JopL6cAeq38uuWHRVTNbzBGAGFjx171bI0yWMx6J+O5b/ox5Iz+0RrxxBEbvP1gLM74
DnBDD3fKW2XqE/GVcyrFTLiKQKh1Jme6IoNI+TkNHlUziWm1SpNisBa4zC85Oa4F9IVYRGELoczc
0BfOKKGq2QxLUQUEbqs436l14+mJbk2S7qPSVmoN2oTruO5s+Z/ogFOcOflJzP/9V/uyaaYBE5yS
cmPllgF0czEBwZeMCkkThfGFmdnuaujDidSAW93n1a7wLtgFpQCBMEMXOyu/5h3Av1bhoJWuQJC7
RZd5NOna2Pefam24MsDNecx4Tt+mzjV9hCoEtC06NCAXgIOHIAJP3Jvv/djJqwV/iyYpU4scJCtR
+HHpNW6sxjTsVo9+ryCE/+nTpjw7APz7iSuGGrGgeNarFagPCdxtsE0wUYjteRYjLACeRB8CR4xd
J0iolpVNO3vptcxcKmFDthr2hKwmOecmECFX7DqGfDJf6Iuj2W5BUWagAo0PQrPXeUt4KsPEJ4ux
uIO6jAqlz6OQEm/9TCcC+QOMjJKJNa8FK0gPoM4xVHufjG58DxpIHQ8RsWtWi3KvaGc2kJB/jAJC
u7+9VDm2cNrIZH+miHo+o6iLqDNVQCNvrBv+ybimERAtKjFCyc8/oLZqRPKiKC6hBoKrfFMkkRLW
LcIhpSUNbFxO6vmEkA6IQpyq0QgE3JTY8H2eoF6iljTd2AYnaiHuG0Oy7NdqdXdLApaMzM1RL3Lr
MZMxVAG39YPUhqJxbiZw1CISB+bzZpn39IQYJ8IWo/aTzNsrhXlj/tOOLSaQ0Sf095I+LVqyja/D
6kfkgeMZTF9Y7e0NDzIBgV7W46sCB7G0fKQk/OOf6yOejlEI1mb631ZsWC+3en8zNiP4fBzhUNpu
ZTjAOT39p+g6iZNbD0HOhdJyvmaS7FKCcqZek/QDfBHS71ZhLpwHQ5fQRQS9CSCYWYE0GN1PVjUR
ai4LoKTgBrOTEKn5YJsQvkVHQTepFjN/bNMi2RpwAph0ARHKdt+By+9Y8QOxrKRQxGRD3s44/0NI
it1KswB7+W8CDGEPp3LPzXwAH9pz1Ua36CdJWoatjpzFmJr2OzmkibRWNtpSdt9elVlzvndWp3EF
3rmgdzKDePXBbcsPvWItQmc9BClbkOPo9mFEBtV57xD6ay3R5wCPo830+pwdDBMTCfy2wSlU+Fil
qgakTSj/RoAcrqwLiZK+a5WkTmPYfx0TAlfOK3M27fQgkJdiZz1WmSQYdaHC1QXedMqbZiiq6b0X
1/s0jQFkGZmgXt55TP6SHv09iKpVwmlymKoU2YLCbHzkDIWF9orHJjinY1VmTeXXOvSRwgokDkTX
sana7R+SksHxnASLlCQR8dqqlNN9JQJ4Ux1izRJ9n0lztYEY8D2SeyZPt7+sbqkAn9YP08JvCEXd
cGm+kPwdvuSEuo7En7y/EMw+YtFk1KCXKIH1GWRqFVTkBBlFELq9jZp9Edm0wu6uSRAD1s3qRX2u
FK2tp5eyKtpffKe0TgPi34y16M/Ekp6tiM3dd1+E+6TytoGFFNMae3oCT/+ALI4jjs4xnwbZquAc
f734N2QKQXMcVd2EXo80TuqzmruB2BD5nNwnvTM6tkf+vMYLtVG9LlaB2aXJt1sDw4T0ME4QQI/3
rJIxlUzHw3WJJ7Rlx3b/MBrqvsDbW0xXyrrDx8ajXycUpqGhegReD0P7k3IydgVFY3AewLibfNfe
NhKVSXXHKt4+BOIuQ7Y/6TJrNHfOq0jdX+udSjsUcyQx+Yfb5fj+wRkePYwDJdrHzo11Jss9mAmq
zhLdx2yTxh7XucOBQACaunqIqRzQzbG1uB9NYNX+gGKs5j4/OVKNv0iPIsgKg6ObDSmOjBn/E3dA
d7GSvGBpKR3BGDUf2GwK5SrL+SQOsw//kBEy+MDrLLq+QKF8BQg7hXg4TqD3c1FwVKmP2OjPN/yB
/AJcwOJVK1rifDf91l/Ozql+VV6G90x4KJgJcgXf53Hbiykwcm9iXuaKoq2sZWFfxr9NeJg9MATx
YKRDmAh1X+feduIg7R3ItSfZep+d1MDbTPTMHq7CZeQiL/nr6o4tBLTiBHP6Hi3x7CvMq/PCmZrn
UmsMSQsJbgy7pWKCUzE64/6eSF4tE5Zk3IKubxF3Dn8GCKU3XuV/XhWS1lsMcTodRYr2l3Tp6OEP
YN72mI+q3IpH/vVytjJm5VwjYGqJ6sXvHsBVOHxo1PD9fww9qtiLpNCIe+ph08I5ahe5dQc4iYUx
OkKKzlaqbDjz9eVXJLmx25GVSff9MgDO0oNRhBXdI8eNTVW1JHmwJmMCRT71CiUrNJc1JgmYePRY
tCkhJAmZwtJIcgQ+hjLhmK/wBKZPZSE4XdCTasKZzWdbvUsW4ALzqBuebeBG/eLKsovp8kBG2xls
fETj3XJMtOnEtR58TEwjgJXkmLMZWYUbW/XkFdFpIdLv3+H/UbO9fKEr1c5jKFaV6HmAlPlXpbF4
niAHA1kdarbk6sDJYeeqPn6E30aED3kYata9i6/UIV9h0J0cS8o4Y7N28R9FK/fy6cmATkq5qHlx
KzUHhTObA8fP3eTMIR6OYsovEsu82dCB1ujwV+OpNp0vvqGtowNT7RwtsLjUv1ElgmficzifNJIu
FE7MDqAHbUsFTWnIc8aVaWru0HJ74j5LPKt82BSwrXr7kLI8P5mdkTkbSLqursPaqupwftjbJUOv
OqUcIfjZUN3tGJLk1K6DPUo3rX43MFDhs8zV7uaBYCUGWk5N6WFOxzb3sP7qpj5LuxM3fg/I2UbZ
630MzQ0R6KAb35q3gC7n4EvmnoYgoTql4nrc50hemg0bg6QZmMKueF0BfvzPC4fk4StU9/PF2wcc
Qri9bXA5lmD9wPj/Ip6mzwcO/1oGc1WGps/MfAvWhBh6OHiOV2gBIlQJfQ96wveeN1jO5lsLh/nK
Ty+we7YnemK4Po3h17GiTuaV4f8dlB2FZ/DUQ7oZU6yn1f73MlFC8q+rWTEVpxq8Y2N9NqpYUXot
MZYOgQb3/2R3WnzoGdiL7cbE7XFsBcoi5crUr1gV9+OJubPjxM0rKrPTaMphRLlPM0ad53CCotAA
sjiAqn0jIz4BkFRri/trMw4uaPEo8LdoO4uZC97sfYxvS8SCp+TwLwyDdvGnje62B61taj8zvKir
qtNwRW9IxtTwxDMmWyEV8QRvRY/mVgKF7CqDMly+Qv0guDynRSVzE7c/jEiBpZLbesc9BxDll4QC
mZtxq04bT4eWBUe75uhf/MiqwKDqPlepro6Y8ElW+SRLZgNVjFemNYNFtAGQH3NVAA2v+XKVoRDH
vu3dQJXccrgvfhlghIZJipvdZHV0tpbkzJ70wEN2FJPW8Msy2L+BCEvnXWQomTGUMzZDcGgyIayh
JXlUH4OoqbAVog1NEjOo/cmxQrDBVtCRf5EPPpAryPI+SkCs3q07VkTgC0lH9Z7rY0wom2t6t0pM
yK56yxbuDL8QdvOaFJ5wHwW9mkTriR4BFqnentsn40YNRzPzzAQrFcIpFWxhZDfW11tpZT12Orb1
S5PHsGaOmLxB8ogxLwyORnjgtGh0z/NgslkYUF4TTYSyMVrZNvbdOfh+GN2n+zTbekBLmCT4Zp6f
4jYVoE/i9FbTXxLKeuUOPHZf/Yi1Ow69JD+90F67JrRBU/eWJMFc0ikeNSrk9mUzRyg8Uu4KgDxD
TOYcOr943f+lErVunQbo6j5f/3XGF5mPUzhSzS1RXcLf8L5HpmQGHdiHvOZFTrauhCNa6D+qa5DA
uyIamTeE4KiSlWp3ekRbhSYvshC3C0fyid6fd6zyfIhnhTcVyC4msvdxFofCmEaEFbC66HpUIr5H
3zKDconp+TjIcuh41vKoFlhuMl7PrPTK26vKN735XHDQNW5A7CGngiCQiOdCh4wiVKzlf1t0fISX
L/bVX9kAA9QlqCIFGPzYSZ0pt2eKPs6J6d4ziYTq+Sv0UnaRaKsjk3wKlpi6mdHnkGLHW+OzetJb
GVpItYuLhGvoq/hLm8QJ+gnFBCYPjbNI2qfSGAcXDvQ6u0ppqai8Z8iH1UY8GtmEIa5Q91iMP9Jb
8QIKRe/y6JMjBMMqGDYduVsvaePghMFvQhegulpe3bpMkOh60Go7uRkN3xdyBAjKLvkjFpMNDPUT
rUCyjARiIViK2AAm9eAcnyAu02haG9nAow5zkq5u01e4So3AFPBBapXVW1yavRGPHx+ReuUVK2bM
hEBjwFGuVDAzELAlg8NwaHpwlwr/+Y3YYxBp6e661PlujYjglo1zfdee32w8dQIIvTnZVJBYi//v
vWcVZVrZuEUSk1bSbNkOL1CnAvCzYtL+jGkHSG7RkxUyI9+F2/2gHHYxKjscTnNxRpppQkn510zL
0CVwj3nqhnNkVyo7alg3W+TXljvTAZFwTAg4QiqFyZYMrYRhfJglcmzEWQiCvO3KEKVpauTiLdZK
jVBuwbFZ7BTxn4ROWNH5lxUqHws1FgxiaxwV8aDcy5qF4E7Mwmb76MtslmHT3t0nVJxMFUJfesWe
/hhANkcTsTCkpu5Rc6jU0Tgo8OP7Z53ZHGPTY8J898blHcln4AXRFf0yFnGPR9eFl91fR6xOUJTF
BBpSabivDnmB7SOb1j4StNs29T0bbices+mZi+5yAuTSs3oo9p4wz7+tcxHkbDECl+kS+niJc+iH
jKvAxqw2yB2hTDocn/PJ7eKndPwxRIV3D0vuVLvLXGCP62XmM1XoQ6VHqygNWrihVhASDA/HrkYb
orKFTGJHtiJ21Bv9Du8JQDv1ejBRFeUG2wwfBrUA47fxYanmMEj5t+AKDN8lkihLIe/OC4CEMzM7
xULUSww1A9to92nrptyNQO/WKfqK0IibQ3QaFbKT7H1TQnSRicA9dKdZTJBiY/Bs4tbz4lLET1Su
OVxyiG6pyIcW4cBsmwcvx/aWMTNbRNVmvMJtkhHa7oOcAoy6rO2REsaSR7AM8Zqv5m/V05waWpwG
Nc64fmDqUi5RFiEfCBCcWRboZ4dNqiCJo1z5N4c/x9PwokZyW47+APW0vnC9k1EdTA08QfdRSmNp
yvK1w0tGd3D8CF3CW+cKXxTxBpVYucwaV13sbW9sCTRqlw6mRdQGeW3rfWXndlN3ykoRg5ofsxlI
k+O0MRXCs6vmnhIBNAkZhvNOKQxn561O0P15bRm76Nxf0Z5ZIuCfMxB3sSerMcB7BBktMg34mFSd
Sv/ABVl0kU0TzVp1f+ZcH9B8YHgBQbIRVut11911oTyNIgmEwu0MQXdvG6MPGDxXaQKakZcDLp/e
uUgDKdVeEqwztoPhnw1G05eSvVwHCCmJn/rKXHJJE3rUnWLglvAXd8++4nS71f7p5fHKozHBSKNh
UiMb9T0j9rCgSpvfxZx3BYeFHLs1COsb2ZyY85jsxjKxmIk6FOvmK2hKvwmZmnZJlRpr83KUUaFm
CnPXzfkdGCWIpndZ90aYrW8SBCjJS+F1imjJ2QxT4qkCD9UbIzaB0KRS4OriqwJhjYd9ybipU8Wa
YwakklFqogOLsNg//vOBmxc0hKqVhOAYGAKa3QxPY+1Ckk5LiTQFIlg9I95m6IcXJOj944nwrrHZ
1vyBfrw8qe3rCQyTbTod9vHiQViT+yDzDDc37ptMGakUHdLghZz122dHjwFwTo976J7oNkL4EN7z
H2AXwSZ1Zx0bHw1gUXqw3et57+n0I8ULffvdC3UUl9Nxe8XtZdwevVznKsvtRHsSlcMzeuZSMenT
1pFPOLv8KZ/3kVg0TSglhFG8zXb9eGatG0H0VAfn5nctx98Fue9hGGMgFgmO9m+GLtftOW3AEz9Z
A8RXaf6Yjg/OFoLmpGBZ2uFjTdGgsg4NY0JDl7+93rsuAlwukOlPN+F91DElYetV9VlMzal+zvTU
1yUUX4eauJ9fJhPS7Z5IcRJNEQ8+2ETeQj2cljkHw8ZyHJap1prftlP8UeIUDJ24gGzUVSGi7erI
rvFQ/9NbXt9N9Bgq9GKv+Y3cMhYALtPLuovTcaDXqrthMETIs6iJTazPEPR62M5IPZTJw3bAYReB
RafQriwoOc2PKD6qaFQ7hoEV/1Hi6uXBZ0Us5nqHe8hkhRCI+A9yO24SjTv3SFRpGr6vBw8EWOXM
d4mKpe/G0uW4NtXPAuWbdqqbM9vqhb0WUkVFmCGq6IcXunfpeFiRss2k9QEdmXyRsqvNlv4/K2wJ
cU/XzK7pCGvLp998pb4mXg8INa7fG7AdQLNI2YFp1hQ8mYM0JnkkNnuILM2kAz+8rm0IysvyMKDS
aHk3/JO6uMqClTgvobX3LYOmyT3o10uTwJ5yDnkB1bJYz2LYMBAVTIpwwlXKuwxOI2j0GT0HXcc5
SInom0YEJBX9Zn0/BOsXwjuGaq0ZNkA/agYV4gvvyKa9+migg0B2Madl4G2s1qL0idQKhYxTNa+0
tK0mHjURYaDyMwr/ytDwOG6DE496e+z8OIsI2CQAZ18YahS296zTXmJITkGWyOWCZOgTM/EGA6Ij
cGdiohXICrhHEnb0iM9kGqJX1J4hyo/+2AzRJUuZoP5Io2Nl4Whzm+KhL64M0e+k5Gfks19Msu+H
OX1lF2niy6Neq2uEZhkIQRaCNOxLEOwY6feyssNfFjMNqw5UQfLSxo1GoO4Ufz2fxvJjexwGqKJg
31X6IoqKsNAjQlYgURynT6Qf4IZF/Zp7HPZ9WxB5NzslE15ds8OPgZXh9aJmZCNMajFJokyvdESh
hKDNmmlHTtSRL2pGk4DigmEPLwHoS9MYd9zHXIOhqCTHhNDoIcEOG6v/LduY4qnthiKM9ICei3wN
MlySlMjyeruYGcEbbiycU9s8sBvHoV78PDgxDRRm3SOx7JBmDPzPmi9kMQdDz3m3DSzJTvnfTTQe
uQszs6MR2x8CwAF6N6bTZe0LS5hmwlpqGbXly/r/JMlV3TRrcrmgqYtpj3/Zecn5CitDl1wO80vf
etaMxEE2mBiJDePPsHVFhEcpMANz18P1tX2s5MusHOqvh/HR2B9lPrmW2+VUHKEWzJst03Z4tfRR
xFbjTHeP99lv4n0KrCCeNg/+35Jx6FVhMapJpuLlruP87oAZXiCt3ESPsTECVyRYKpMrTutRgOqi
7u41nCEYgETc4jLGV9JFwqNn5LJSZmx8VP+N4+89GNaxOu0PArJwD5s8ArwovwoZAXYZdDghcEBs
x76BjwBDaAwbZO/bPHkamHFmV+T118wmSbSRzdloLd08A2FMw2A/gCY8XJH/d8+kjMScNhIlxlHw
LfQNlik/Z4Y6AWEvjzmjgC4eSuuGutMX+vrcEm0D5qq9py+hkqaaskLj3pFzzQUlpsgPaK54v2UD
CM9SZWbZgbzy2aV8CrwwWZF9HMbbKusdeO7ARPGdlIbGVmQ3MZua8VWvJCIp4zVnsvzoZzJuh/2R
LQuEce/5R19vcSatbeMP6QzaqIdBoBpZkLtDN57ACjRjn7uUdeLhfJSZeUDydGYiAP51gBWTnedB
9OpTHjLsEZjTiLDXlqGtx0MTutWQNWW3ikhz/Y33+Unzx0RevV8rNahDo29wx9pfv4BNIVMK8ZO+
W5xBYsuvp2PepybJ7Oh43zM9XTh7bNAe/y0W4/KzWhM6ewbCxclwZ8JLhw4CwrA8R+6CRy6KxkLc
FAnKbHfHf0SSE3uzAFo4I0wy/t1mvym8eJBLfrcgmvweUNbrw7/aukf4NmtoFLgBpSenZrOcpatP
h0sWsgh4I5qpVHOwcuLaXk+Iuz3faWvit4kdLq69+02txPw1cAu0QCKijz5xOx7Nqtk6RyK4q8BM
K06at19PxO0qrW55ptICBlFsGXCj2YMIRrYprrH72FLGkMljmTwg4Dk7fOupRfKLQiVcyAj0x6ml
2Xox4eKJERdYKo/FdhwMuEjR+Oo5SVp7RGAg3cywEHlCs8gIvILz/IwP6JbYiFIMUCJqLJJ1hV8V
VI+0NIJ7yIjrdyfO6nvHQta05w87AyKZw+n3mk+vD9zftp4q1ytQr7lpXuxHnNHzblEEtfE61OzT
dh6Qob5bRA2cM/CJeNVrLoYJAv8KfIRJ72Pperhjxxc5Jqpx9DRvC5H9/O/kY0rmebJXaX8OgTnG
aLnQgJG0fKpZIsCnRCNh7G+qD/TsZAvpY3DmUxsAC1Je+uRu57AUvei3aj8x5+mYPRvqCmnNIsDt
K6ShE+5NYrGKoqh6/wLr9//AWAZLYo5N0BbTnxTp9AlpqYRGr7QHdioj5ncaQ3qEUWSL7w638Rgt
fCMLrAnue7/CaMxNtJ+koDC5pAEugwn8Cnyyx8QzC8na35KSnBu1nIweM2J63o/6jAV6QqEESXTD
3aHhVK9Tsl1sHrsK0p8rR/J5qu3Jq/WJxKPbeo7/6+53+KN/8fIBRxAQvl6VZtbUqqaqPM+dl4+H
RdSLrtLgSBfaZI5iLUj4R4nRg8fBSrN9H8W19zLN2waraZ8a1sK6VMmM/ORk2+vzOheXja/CQZD9
yALLuYhsJXbJukRYwa/9kdSbMHmqGtdkI4gUky3H2BTYT9jEINllnLrZhN1bd0E9ZkPAXOvOGEBa
8fN4DuGxb3kSQD/UR4es3ZPZ0A==
`protect end_protected
