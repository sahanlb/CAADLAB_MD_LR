-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2IVD0kNnpAZdBXcE2kgi77jZ3BWPgAbdqZgQBiaryVm/F7L3EB/rDtTy0DZVEvEP
h/FnxDf3B9sr6qz15vXgjmTh2bvRXDts/H2qGkTCluzT9evxVkIicAQcz6It2QLq
Y58ga2YrS1Edt9g3CyzIeA+nrRfVABSZcsVBFOypKEI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 11536)
`protect data_block
q+UbtOiOit3bA1YZFlnxRmXmNHO23xRAsl+j+q+1J+EG/qC0vqa3ZAoInkaRaB2S
L43kfm3iZJ9EnuE/Z/UWfeJ1Drj/i8OHZKO7X3FKU4HFNYFGOzsFHFMM2m4Ihc3m
tQZk/5K4AjrM+UnLZq6Ay+zZrXwTkqjMhrYnQVfIucYbApfmc6feFQNQU3T69+43
FCHupT09LmgM6Ox1IxIsen2zlE5RHNYtqjqAqYUK66giThh7bJB6k2+YV5b2zbV/
jneTENQ132LwmXrGS+JTfeleUFeA9YQ2vDZToLG5YXo0uKaktjB5sh4KZzcnpo2a
EvHqVOSPCtqR2Hzu3WWDeVV5Kf1Q6zA23qtHoZFJUYNf1P8uKOtXKfkX0Sddy0qt
MnXZHarDAfFVpD7BQl0bdWI4J6YHl4jvC/m7QQmnQPNDCSrEh+7khghcOQe4/Vxa
Ac0um0lz/AkVAwUFLApegdJB6lvPpGkAHPmnfZZzDip9yJWI2TbBD6d7Okp1Uc9u
TP/8xijhbYibvMmDJyjtyU6jmTOqX3tS5jWISfcVOPCq68ObZ8IE8RPCx5SRhCAB
/QmK8lTTlcb+U9i3xfsrxjKbJYb98ijXoRvNAtXC5IX1m2sBaCXuVknioCcZ43VU
2pWv7Orjv+nZiqdNXUnh+PMkL5cVWBnQHKapeDEZaEUiNofjuAKpyni5HV2hm4An
87BZArefA9bqXnSu7XQpExkRNBJC6N+kqV7lbJKWdxF8gUxktVBxyXitdhRoSoxM
Ctop39KYPV/iNdBnw9aBaT4TOi/9UkUwgr2xC0no9s/sFLU22y4F3QsbZrVzI1vP
xhqJ/UVgW95UZK1CFSs5gGuRo4cXiwOwplectFuGRs37HNRIkCObTVb6DCo+mY2c
ZOueZq0T21/An1nMoxF9jPDomzdZM0W0OEyYURiIw8+c/pHiUzlyw3/yOXriFsic
CQvIMDnDDN3b2TMMu9CrzwbY1cHU3ENmoglpqPkvjrZ/AEKR/j/3MM3FMeECJOT8
mBANSqLoWHIk49c0UEeE3zKGnFyR6qh53lSZTt3E9dOgLXpqnRj4RnTwhDvYKLPN
NmsOumaWDVJkdoKQ01IrbUiLoLLLI/1yUQ08AFyf2wy9UBuFiaQ3GjGNL2JGJ41h
KK+nfwmZfso4Xk3gLDiP11mSA7ryNGqC7FG5hna73X/ZAvFxzuMTttu6UiF86eNc
RKe388obOyUiAOs//W4OHBD9E1UzjTUik5cgzgzFWdgYcmDzqoZWnVMrJc+nKntl
TODgFyp90hdm259ZzNXlpQwRRB7F0GaOeIMmIDsXjn0UHTiImUYbAUUTJ6r8nkRn
yR0ntwDZiHyC9tCZNQlHiSS7E+Zo99rxGq6rB/gwshzzUNMmzuH89M6xA8x58r3Y
xXyFiX08y7HeEOYxId+5CIoniZb0Do5jadRCTf/fQBa+xYEC50FfcoShsyR39IMA
vkiOnzw0KwHKpmXQMPoe2QLmY1o1c7c/w4zQq6NDNczab1dO7EgXvJE+kpuE/88r
90wthc+iNdQsvxJnFcBHXD2KXLL1l7bM2klb2xC4au20xcGeq99u8G6kSixHRM86
uTYoPukWFatweOpK2MdUePwgVu2jIayC0QthmiWBJe19hrii5XaggeJQGRWJuzlS
QsPypjvpvOvKg3rl26eMJSo7mdvqi63BC6+5q45AIPI3qD1pWsdTHVi+/WJyIzsD
7dP1nqfR58X2RjUoDeOlQ75Mmcvwko3GaFNedpv3ewKtEa9kYRkp2/AgBi/dZrO/
2otwTgRIJQkcUwaSC1ZFV70lI2t3qNk9g2l2WzZ5G8Tuiv5ziASIBCXxAytLRuxb
wXTwdIFM89iAh2ghWks8mO0i73FkFd8w52Mo/4CA4rAW9Hpr1CenDquJxkuu+Djt
qU9VQ/mvuVgCmm/YXWKLmqyDsSgAZKnyXV3yBQ3huNsT0IwRUPjQOzGZH1R8MfoM
agnoz5mYPjEVBHNh9cnde7xbq12WUkIMu6uZP/CHM4t04XKSJ5mqfbeqDFNNygQd
sZ59ZWw1tja9Qn5Y5G7NbHh8AZ35Iqhy8idoXtT2sbWNnEjGMfqeq7w0fChuzwxV
7zReKi7qR+EijhE0ZIF47oCg+CBLk5MHUfijeFbA9CieR7jhonxY1Z0T4Jmc+opq
Ite19/9TQljMFnlkPHcZkO3+Z2+tVhZlJPrfihG0fAVm4Gzke9WmzDNyyVwIW6Ey
ieNDicTjvRH11PhB7vbQwtixwufP9RlV3MfLqqDMIrN1x/Osrsi1sI0aA6FKDm3y
W8ofEb9Qv7aNU1nzeeLLp5Er5Gc593XTh4es7J5iYUN23LUhaTodbBrKKOly+2hr
EzWu6c53koMlu4tZewz9F3nHquOA9OtfQbpxEYQ/O4vl8Z/ovV5jOMgKT9/PL3Ql
P9CCGwlgSXRZ/yZJKwtaT4F4dwkaE89EsL1s4GaSJcl+wpEpCB/gH5R2Lb9VMPo5
e0azB1euYP0qiAp82IUMMQFvFdpXsw2uLHILsINRejZmCX+1Sw5P6Sr158Klye3g
X/lC7yZzD01wfmFfUpOzrF4OOt8H7NIquHtfJVkfstARPInzL+UnzMdF6xbIVmz2
nQ7yttapJed2lgJYRK+vmwXDpTFO8JUYZK8IAI4S/5eyWU9q8aFbcOB2QR1npS/9
ZbRHiKt+51gjZ8iEC1wDLVPKOg0iiaLwhB1WgH2x2eivrCYY1fwuBN5uhrPIX+4n
M+8c0tauEDDpyfHTkG/RKLnFDAMTC3j20PS4zMRGbKGmhq8eg9E3d+vXgTW3Mwt8
bbm04g8P6waZbI0CETmdGvlwc69saaSrMPrU8sVWmqDgjrcrua282/N366DCFkuH
CU1sbPpsF5vBzevzRX+rjTSx+W52MlI30vy5mWAiekM4LbAvvyoRrhwRjSAHMurE
HZvwEICovitO4lgs00s6mgadZ79aAQChfqcPaFutM9+QdH9gA5o4SjSxbpsQhc2N
SOkxcZ3HerOH/DpY970Q5aJmlYu1bEq31omQiebJGv+vpXo2cchnp1fIoWqMi6QW
rnmFPI9KV0gqZktNaTSC1XRDm+osro40mJtPQiUdIcnqjmqp/3a35CNb+LIwhrjF
NDDU48ARjm6IWfNQWYD2Sst3QNJvPvJyioiBD4oVvrUHnqtGICnRQypi9jwGeyVO
28Fnyw0iIFx0sOwRDJEr+qDzeN/a9gtAlEKiSbxu8uZhOmfJFTMszrMTQ7DR78pm
ANBVYPrWGqkkfSnys3zzQ1u9yMNcZk30Y81rM6ZAB7kmpIpdYpnaxEuLaUOv09Ut
BqsFdcYDNtMoI4sDBfMY0uopePK3rvMGQsCSNu7aF/mUXokviiU+iEeBG7lhOCDq
KMy5aeMtdyJBGLntwUsmKwJkqWs0KOAc7V+vDZZMO+FtyADnwcH5flD5RHCzjIgB
PdIBtDIk/KnvTGH7l0dNQ5x1tJslzZJZKpc4mmn0bksRkQlv3SVh+cK+ywJV6PZE
aKEdI8i0u8TPLsvqztDlbjd9MA2cOvHLaW+Bq66O10PhrWyjJ+rDIEkskVN3XcS8
CKq2DUlAsFOCLysYdePQhDRC1JBNUezhvLHlotDDM+TkS7A5UriaMqx7YuwhleaI
oTJgEWEKsZcLpaqrmztWN20LIWyQ29y5UydVf1UyVFkwKRlNmlzSjpLZw1xxQrvQ
sA3Lw9b/cnA/0WtyyYO2xfI0ZE6JZguOYnwDK+ATaFsVTF7Rq3Lh9u0WwHB9IuE/
7X9EWC2Te290J9I//o7msnlsOmpWlMVIJ2Z7L+y6rwWmCngx6T9rh91pUsB+hdx/
mCVigH9iaH5sjtCxMwnUKh6kCi0im/fq8usDizUv7MrBhXukAm+aSk00/lAX10g/
X5hTuwxveE+xI/pVRDXok6kLTY4yOL+rExOw0hkfbBWWxpoDyv+/M3VCD/hak8Au
LcDIJZTk3Zokvd9KE3KYvdXpTVR4wdQ8XpNCPxecYfJbacWAkbWvY9lb7Y0uLHqx
c+zyxQ8fdkiP/XSd1R6ivEEg/PPdt/n8vavyRC5R9FLnP9/MhrAiEN6zg4Q5pezp
X3gGcjE/sNuCWLrhW3B5PvPRVQdzpSN1C6di8oLIEHw2iC0d5v63RwABxxFiRk5p
6ZZYe+XriAII7aiYCAAt+hwwVUnRzw+CeR/cu+bxWxOvYVZf1bZpAbsJSCcrFjcG
8DKnJEhQtYE08+/GMWMhZ+FfrwqXSnsL40vUNxPVOe8NcjGgwuaZ3VS1GwyjDa/u
Uw1BPxhOhRPkxAUwFwaMQlZghiYYibnynhEIhvFWe+NS+cCHjlS/tXRKQfyIDifY
48cgeeThaX5BzNOr4c0VIWFHoxlhpQEjPqg4jshqFDFovKRQsjYdlFKwDBlC/z3f
fn2mjeU1jfZ0kgTOGpRADzEPXESRMlP4p76Iknwh3LpuotXYvCHH/1JOJBbf/uUY
UYDwWcTPu2iUu+vDSUy/00DUOOMgpKa3X6G7UakNMdKFr21i/85JidWGJSPyeSRb
D4JAWHrWSppmnFiPRgZ/fvb1HIuan9WXT3hYQmgIF3aGtMiWHq+EpUOF8q7yEcZ6
lzbs6bnbTk9GE9ivr1KUEERoE+NYBbOwFT5H/bL2BXfONyYZLWiYWLR50SaPRY9u
cq9lK6jrrQ6D9SA+pI+Bq+KiyscCxXPhnEApjw27Oj4abv6rmfEZEBU2HPeYgbA6
G32YCIiIGwNuckiR0XP7olgYqXgZmoaZSJyLPSpJsYAoQ1lwFINRR5fvnya85W3i
plycXTY704+5jw+JNsUvIRzJPSyzDk49/kVMwScTQ1M5yM62CE7drcSKk79ndNhw
RXyDB4v1hf5denoyu4X1xleXpMc+xFamQGvLEnroh/HMaONND1tix6cAsoyw1M89
CPoM+14uteaR57CAySyliObO8Y8j2z78F3NU5AYW7tW6Bz0t2SQrztymVg/fies5
kpQsRDopCaHigVALI0Ie7QbFtEWdIbmgx8BFIDZWHjODXOPT4f3K/cCoPB67WjhZ
vRtMJ8paTZriYXgR/bXBncmZBYsd7Jb3RLo4NMJpru6LUjgF2OPvSIO9DEg69S4u
26WkUn9ROvMuyaDc5LxDvx45XPgVIXfXHOKEkyhl5ve/50HdMSk5A+bz7oLEPZ0T
HjXe2X94pC6QtvPvESNYRLZK/wmOgraykj7fFVovkcg108iR+vBCoeEE3HNPE0i5
zaDuvYS8PHov//UmTir8a7BBgfadk3u8UTDakTum+X01YHMHUSlsD4USoNf8P/89
eCDD9zscdu++65+abaXnh9JNZfPE4YZSeQ3LndTZMU5FIL/wYGN/jbkJ0sAdogVt
GETd7SdhddvpCBSTKtKgR73jpmhjwAs99418whtOgtL0bvh88EEoUUw8KbzOktCR
COclzZs1Mia4uwMbbw1EDpGLIfny2p0U/5voxMx07ugqJhAvZSW7UkK88G6q8YPE
7WkQQTX6FGUPomDONHxoiiEzN3LNtkTwP3BpnZQjMoqy9x4tHTHYA489fnFxUwhQ
qYG1rN+9alRVYsd/k2OuaQfM6rfgkZW0jbbfZj9aB2zPW4o4OhQ10u2LQxt2wWnB
T8Mngfnq5WB2kJIXnvJdAqYxnNP39JP2UxTIHVzNhi/NdaiSFNLXzYDq4vrl4qku
k9yC6q72TBbOMP0jwgb6/4hH5ut6FpkCXlMgiTNSQsDV6U8VJVPv3yQnKCV2TT4I
CTt+LWVdzde/3v7FilpEwBUbp41JJVsOzfgx3xSdadZUrbmCFlCd4mLhj9zryi/E
FvMtcVsUK7DUK8Y/RgTmfr9FHVltI4G4RaDSdUFcxm3pI5WxCH6FK3/f1KdXzJ3e
lC9nNHI1WUKvpHsqOQlyQtCUrJiYbZrWDFyohKU05yIGP6KmEEmyMy9bKXgmSKH0
LVFRJoV5neKXNT295qWoL/BUBrePDWWqgXZzUU+ZiHoB4trENaCsFKv+E0jWMRlW
NempqmCQt2B+uv+al6b0vPXn+gUgJL574IYFs6YzJu4s7KPmCxQb5lIbHVsJ+aEa
0shQt1YHReCXF3hKhWttcwo+p+GVx5nXW2qdHC4KE2ma0EtzIljS0DMDkk9t6oxx
X/v4gJyomW0bNkV9sqnjoTw9ftAJGRRGYcyleYtSyCuMpsuCny5QiTzblwt18JDl
4ycasHhflPIxrH3smSfs1LbTK/2FjrVNcfI96hU/66BxCK7eiuQRYf2jp9JiDyKi
RWvD1ITyXfMMoROfnLq+eTOh2UvayKteBkruTJyMc3rm2IXZjiSI3ec8+aHh16qB
KLrBV93qLstbVMRSqzTScDky/vCWS2Cy3HN/wKN52GkH38YgZw0Dqai20cnU1lwr
JQ9h7fE65qBwtmVOZto7TUZ/1GMHSaUXkoUwPhD7lefdqzXyFwYd2YqZcayOmJTZ
/CD+g0HZlYZHSQVcZRXnQum2/llTTI4+zyBHSPz5Y77wUIOAx58vtSO2t4isieUa
uRo29fCh+Sw1GuPtF39fnLN9kO9xKnRwGpepgVCgLKLgH2nGtlbT5fA56sTv6nNB
Hve48HclV03ibkcTzqUPWTwOihzt/tjD1uYSl8ObZuoRzuj7HwyS7C6tM7cZLQL+
/jld3BMXok7wq9bdE3oWTpOVlYqfH90Sp48tHobgafOk8gWhBw0s69ZOYPINYzTu
aDZor4eTwWWxrM3U4eKrIaU28x31yeT7AxMg6ezLetxcz0RUC7xZgi2GhW5aMqRt
eq6jM/azDR02RwPnYQgVidmbbw/yXp9yqrNxGTum3ebVqY7JPkl7rGemvOCtInP8
v/mh97Hott46GxEQSxR3sQT1TSGPHe1JmEtEvcI6/GcZEV5u+HBCev7RJ7n4nmxB
bC6cen38sL7Mg3TvtHs7WbITs64uGPuEdajdp0gnkOQf0b5vweAcr8VlLsuNb3KO
wFYog16Noh3gC72AKUB+lMVpQUG9J5e0zdnQ7YSZzPy3bdRpwp9CU3qOOJsjmgQU
rcRTnu3XzrzJ5eA7DxNANGtYYerl25kfqGZ6C8Ex82UC6oOfjh08Mx4FJO/hSJZK
tHFv3bAPyodpir/DPYgxGvTBPTdPejz2RP1WzAsE22WnqErLxtz+c1ORQ+k6GoWK
0Bvn85MDBgy63To8u13CuoAEXdAZI3rk9q9QyfY0MozeWZEQBssHKsuxR3SkFesJ
VTBTQsr5+iZgcQ9TpiXx8JbRpgyEX5Vf44jKe02Mjb6d152uyylcDFG2ZItf5qqe
FczRsHMcagxuAKUAQYNkuO4Ivw8+wAxFTfPvlhcle/iZWdsbIxxUhhywcE6pIRfT
SMLl4BKqbDvf4RD/TfHNPC3EoVlPh9KIyxWMeQgxvkjiGlzPUGvy/G2teaWQZ1yP
uRT9n+dH93gWE5inDLzgNDnm4WIlgEjOOvwTfs01NZEEQG22TVueMGeJv0UmkCa0
3f+HcJ4Aj8Ok81xW98IB7ub1DXXTudHmQsK26WiahEkkdzAYuIZDUIjnXmr8R7Yj
N7Pq7zhrW6N50C0FrWPGt7et9koQp7/R+1RdFQSFy4tJ4xYuYEQCD0GoR1zmWNn0
wIpeZbej/3TA34uq/oJUt9v+159jMlf2+naAGWsz2V3ljhom3u+kJDUAFfLdLy0x
PE5kl3g5v76rQjpP2ZDVMgZw9Ye6koxdC/S1aFnzsafHYdiUP/w0nvNaaeSo4uo0
jA2X6TjxY0PGVaHrONKmkjBcJKjWnFiHSBADx/GQF89YN2dyCQrgdCqbu/Mx28jA
viCzWeWs7tsS5OxbGXcyXToguGwgVY4zo01nrq/ml4LwQYQ/zmMDFobexDcS8IH7
IWztLDk+EyGjf8IDMBPLk0z0G9VAxBksnEFhXy8ViZDkQxZ3XaYCuL/iSjz2Wx8Z
v7VQ86uh7dCvLEZj+vf2q6I1XMpcsNkD3HWOxCG+hmpzEc1KMgxiJH267h7WvXIx
Iha9ZxDTtlZQ/qBqX3TG1UHm7yRo0hXa6RMeTDiUWMPoALO9YGlxkQQE7VMoTmHX
/yGnrwKsJN3u5goSI5PsgpmDuMdT+2QBQp5xk7janK1NlsFPirT5kn4tdmLj7yNu
ywZh7A20dhVCzdMJKOQ4cGBZv9JAO0v7955UmJuYsoKRcA7xaRw0zoxA60fGltAj
4O9slLu8XW7I8vxSk6GwL4Kr3pobifXLWJgC4ROCOh7XXBF63nuuMr3oipYvYwC2
zj31uejZUTv38s9YwzcyACIDsSKrYmrr71wSw16JPsO+GkKzCyMsGqUPz0u1L1LF
kNqW5eqa1fN4k02v6mQI7mxAizLb5cwC/4cgHt1WgoNFSQO13fOzQ/kl5lJ9se47
JpRuzJ8dm8RVmaq+fuY3R0oVcN+I0r12YDfxVwzdXZSQc03v18vv9euobsT8Umj6
ELoCI3UlBruax4T2BEBBJj4j05cBGR4TnfGWWTn8k271ZLJqHjhiNb6IYhsIQh0P
1+JZ8XmNnJjz4+FXU2njrcxmeZqQ8/2rGpC1zXyOuNvglRxYs2bi5MQtNv+U1wNM
L0rxh6YHljTvdjhzaSNMpr7gqEDqgt7HlYNV2c6ZkEtfNeUPvdtINKETANmF00gf
GQuBDWOAvlhjJ+z9belmK0EArAz4Nrzi+MuVuk2bYW+QY1NsemnwIayxwmJqQIJh
sMKSEsuzPrXX9ZsxcLGcRMp/KxmiD7EwVoARs+CoJ3O0+cW6S3UgHetJsqVC9a2I
oPcfX4BMCi70Iw6D8eGj2RUsvTjxSWfnD01jZg/hkIIITTl/za7+1/3C00RuhLAI
AOBz1nwUD4ldFe+kN3XjX7zwgkfeho1oSyv+qBkzOjrzEm8AiBa8wxzzUprSO/b8
9GjOclNGEiH2jA2+jD6vdoATUgGX6UFG//he609Ds/eAoO7YhFKpF/RnijMnWvCg
CJW7wmNIA7HUV0BkNg+RdimawmosxBwo3Cry3Lw78NN9fLU9UOKKNaMTUYj9CJIT
6IlZu+ouyg+TU+1KvqaEwI3hQTCUmc9w3jBImzUonI1MuRqomE9CUTjVZyntLBUg
+QYuMhYKZXSzjhwyxQbEPH2Nl2ZAYHnzLSpPPAcbqsqHKe23Q1c9YheM3oCjpGAg
M3Ej3V+9SMT3ZXKxVF37bY/Blx1Y4rD4kMlQv1WBEPSI+ZQQ+y+xVCmkQQkIJ/8z
RNWfRRI/+mfUreGlQ9TmHMRCQA/gPcQ2PkeYB6yo9hQNtpC1rL2LWBE6TgJfaQVg
2RLc9Syj33xjzaVllu1lbLZArDdFqA3UUBQ/Ob4luv9ehL1m5SYxRxxeoIBn9Zk/
2n6nJQ8wnG2GbuHkYAAtdpf80FS4CE9P28bOzHO+/piOVoMTbNMSfoR1AVq9wRj9
MLQoLjIN0eoWGCi5eTD08YT7FspXqpiNLIXNLgpbvMK0+q8lU9naYo/Nawx+7PNy
T3G/i/x+F69UyQqDW4ENRuk4cUlRTfZf9dF7IHC4idCil1CbF3I82aqbnWCEJuIz
4gztnMG+T8enjN4Si8bmt8n0RNDrr8lW/cIsYCvquX9u847+mOYkPTLTGUuxwB51
uGeDmpfZo2yx5EqHzYpDtfmBzOxvLGDmOMg1b5HIni0Mt+Omv9YfpEoO2q64dTzz
q3hCxXcyJK16zwu2KQC1Xlde1HZS8U1iqwR2QsDcDxaQs0POwus6ykNxNX9wM89i
3hBB2o/h9kRlfUapN3aixj0R+uwmaCn3tOte9JcEX0M712gH843+e5uYxxo0dnDP
JHrIBqA/fjFr2R/We93ZE0c2tDPXHM9kj1W1s1+qGxFNisphm+A4CbWV/zZorXl2
ZhSxUsdCpAKmxQE8OP+ixXjsOTLpe3WeGlqSfiFycEzFRYbFI9JWlUXqhdMjqp5+
vyHlq99zK5vT4Nr57Zj1GkOC4MDGaz0ThEONhynIjsOw4XPk+W+7Cwq0BuAldF+r
9R0jfRDNcjeMi4MrLBFJheGSeoiC0d/OU7JJivNrVEKvn6zs36VBWm12JzbCP771
sSQSaBgdlih1+ubd5K4s0++Sr6ks6X5rNpY8jlj1gQpB0mHByQfs+d/i2xfCUCw2
Vrzz2SsToZRApz/voO02d0JHgcI59bNCtYni9qp9tyxObvnBd0+AUoeh+f/4q5iA
ualvj5T14rLDmLLE/eHqkVkel0WRjE1svtYWNiBKTDvC4dSCed3xJHXOeU9G43ME
hcAu7CBZ5s0dKmTno8lPBHpXUMxJRqafodZBxxY0CMxSHIvGYPcABUolJwXs30cr
o9mpmrB0jRst84WtfCrGRfJUBo15vtqiiqRyTBXkJRaDk1NE+7SDWtm7Qy2paqDP
R+0O2Ic0jszePppToEHe9CoDpnTLmD/zlPSGcdqUveJICj2MtGrz5lLyXYAgblvh
DiALD+RuNdR1YBFN2M5KQPXzp6lkKfqujo5L97hiTdbXv9FKBza5hT9Ck4BAkThJ
8fquwQi3J+joBVFRyhvNtNzS3DbFNyXMHMrpqCf1+HXt98OkcQJY5PAdBQp1XLdH
QTFn2Qc8E5ne5nReYdhudZJSySLps0ihG+OP7NGcSSzINGrhNUQmClxdVlcqoRLD
ep/09gHiRYOOAdzhz2ImDb5fgSj2ZIDrcUhmFCQ20nM85y8c4JrtBIO+sZeZ8g5s
LRt09LqKvsAURt6oFZHO5yAMAqkZorwKbtKVxqkjJFFFzFgJdX2Q79UzTGwikSzD
TeUm25kfApcZSnscsJMMlJfeg3nW/tiQFpitDda0qBKYMWjBRwgvAkRZsAWnCqZL
goPoWUqfLU4C0VzYgX4S6bOr/P+DD3780loYzW483NsNTc/m5nvyHQ1z4XGcrduy
3YfXolsNgIVbk820i04yIMbh1/zO4OjCBoMSatKieqjgr/gega7mW3c4oiIcl8sR
N/Afk6pcaMgcTeSyI6JIukzf1M/OqeGufdEsq/Paces07cK0G1TNtkgZTTFLRRhc
wwqCB3wgTxIeG0Y4ZpgyYlE6fPR2NOsFCyk5ieOXOzqC8HLQM12CebicLvqixg6I
Izi0fuvoM5JD8MaoEk9NbiObk+Dd0wBUwfh/lqtVW82TxqgIM8Q1hlZa+f757a1+
grj/uMUxATXEc7xQ8sr/Pltfn+0rPAeh2y36lr5wNUjzEAtO0mM3r4J7ESmLDuJZ
rvnl7vMOeK/ndkSkD/rPZ84pG0sTEQiQYe+ZF4qOyGYbpknGLtkql3hjmYqFJ/dG
tx01VW/rIE8lHjwR/vWnf125ObyXP1eerxh9K2zJCvqMgLym97Z9e0QeyjaDize3
Kw8pS5iIXUKoYBURFDlu+VGGdJk96CWbhdfxzn8yV1uVreZO3lyvvS2RaXdHYQ4s
D2h+McBZVx2ayflWv35RfuZFDN8UFFkv+qqXlYdTAyY2X/mdJWcWogAt6IPhfxAQ
TC50h+CDJiOgC07sInqqIlXJzEBPhBQLALP7Z7wsRckNa0d7UqCwz0G3S/r+II8t
IKDKjHleMEzuO4449Q7yYitoZw33FcEqH+EbhB6d2/G6glIpqbeUdj+K3OXqzxiH
G1a+S1RDYNlTmeQ0k14xHmo1NfHjK0fZxxkQ9yTVDV69JEHa/NtuxGDbB/WsXQbF
WNJLq8hd4PB7L0f/qCEwzsJaYe9ufOs0PENxJ32bNUixEfjMHt8XAobnWBOMbiNO
EHz7NrkDTyoKA5pBSMmwMpW3ezonby7T3DTAOldSeC+tnxSJ+A7JuZrq8VwLGCAN
VoZaW9yJh1LUnTK6A4F817VfxY+GuBXte5OQFAijvU4T3/4fM0YKx1qMsYVq+F6i
+v4w4SOd+PuLx41rZkv3bNBFSAo4PTwSzzbrGCkCNeC1opy+s2qeBixlU+KGD/DE
9ruJdcEXZhZoplD1OCh1HYpTZydFVfJHCKgrk5WInAH5VbvdrUcQuTrAuTPKxgIn
fxb2f7/wq1Tk5LnWO4jU1IHB3ZJTjyN3si8XZC9WlIvLK7rp1NKUx2Na9CquWmP8
8N1e7+oZRwTCNmDDsMqAEOlLZZWOupwmYWaFpkv/M+fN5VBDi+UmMFAa1JN1hChN
jSh/pKB50dZmbVWkgtYxrD7t44pV1ZDmj1HbQZjlU+kOMmYokGp/LDqV0s1JlnkH
H5EIEZoDLAeN+BNFJDuKhOCKnW+b9QPes07YGnGLpBOLN4glWjze57b1zMgGOPqx
SZHe8wsdryr0M4rGU9scVzmXHI0qguwDKIkMXeTALk1/57YwzWhm0mTwNWcptmXF
MbVFCy22gb7F2Kh7+RAG2nJjAU7vP/H3XlwkEWHRqVNVwqSfHLq86hwHJMnHatJj
i2y051soTSixk57vxT3LEdlxU06MIWoPO76CYDF8uj7Ob0pNox4gVn3s8yeWeF0H
MfMhdZdW87m+OHgnVRgUgPA8Fko5HbJGt+NtiBXgY6yQqsXTEbSwaSlOHbyTEb4b
Idn0WMw2Diip3n94Anaz5ZZ5x8l+PAjA7T1HDHO8rfcc7bZQ11+RcHEngZqOxzis
jgTll9QeIpwrTmAXHD/ELLPAg/xHhrRDZJXTAsXzT3btWTLVDgyG8L6Gx1rqvc9V
fsHnyixv3fnfJBWrpaMfsLzUDFeJPQY61fajDvPhOlouvLXeN0lpw0Yrfia5qBTZ
KHBMlX3y/V9+5wf6CtOMyFnR00devMour4DGkP6LSlXLEti6ay2g044dIGVjN7+i
6mvyTxh7LOb0rc++uukvjzR6yXQ7kR4+HAE2pAlc4gX7N1qKL+kQDlYRNyUq5LgS
aUvSDYwbmptO/IlFBRPyJgGqTx8p7hd6ydxgDjMZjx61/lDqkuR5DCVrJCf8ok6v
ByvBCiFLGAZxHMN64Zu5G0OUJkjK0BYyMNih9v/Kewbo45hpwsJprUaWorSo77gs
47zAlJ8PcssFOWO5MQ29oTA5I6hS5SZwuioDcYeCJ6hQBDg9MJkWztfrzLMJTBR7
izQWyNPiC8GnqvfjUk7VHKdOewWbD3CyRWDACS6IFzp8KYov//1KVX6PWQPEw1N0
Wmhcxw5Mksm2iRr4zGmoq2n3FUOgThPH6Tq1HGdBajgsjTdqzd2woTB2tB3V1zRo
bSFN7Pjg112IVZD4ehM59MZdTKxSsOA5qen9mRXJI49/5Z3GNfl9/Zb8ws+2yIfY
btNZzIFZwZZ2mOznNlgXwh8IpwZG7AbsfXIqV0NgBb6dpEilSw15zx2OuNyR525L
xie9Md62iZ9hSsDmdETw7IKqAzrhGZqxfpSQN4Z260LT0TWciik/HwNL7kpsh26A
oJejQ8v8qdujmIYPWqhllkfxlx+sCjF3ECq+zugQJ34QdRT4UhZVjUws8DPyHWZD
bl0/N/SYuHt/pPMDKTb7mW5KfV1gEoWjf/na+4MZfS2yR5nytVHwhW456TwpPswW
TeqcH02QtNbtOXr/sSgUgWarHCL6KxucAQDjugrfg1bmLlL82EX3S4UIdd4UDczO
ESswoAaMy0r29UTOm2sGsWpKlAyVeBmr/crAytWNvPC7rWqtiS1iDhH/S+IXUzMw
BqnuGA51lVhsXnTvnKjCp8j0uvUdJACbKXE+ci90bMCsBdgqgArtf17+GJ8aAits
9XgsERX4cL39nVj0IEYdgUprv7WyJT/oDc8FvDCiZ0aX3t4i9qJUOSyzGuAuvrnU
CjXIzzSxCvVx6W21PBPJ72m3IlbBa2y2h3r/k9GSxfe5mkpEteIRKBHpr8TxbZk3
5T4ErurXHlRJHZjALZBScqpw7GFa2KQAL1Y7K2Ifto3DSMmlasL/MTd2e4IIUpIm
mgdGfXjuZLzNstfTZ+AF+IWah+hPCUR5gbEfU01C4AlTFRKuTEPdlhlnfMZu+nCA
ig/DfvJycMLdE7FLZXaBLDPzp+i5ltCksxixNqgIFpPMXTWmYrq4v+8Vpbi/56Co
j5rgpDgMx8yHPsIsV5npGATMIcg5lMIGa9o00kbwNcVZXHnHr7EL3heaTgOotl/o
7triOa8wM+f76x4HRfvjyeZTr1cpqK5j+GhtQqlvqiI58QGc1fqkQ5chx/AFujYG
Q0h5JYc3UKC2+nssNLR1TRZj7x5JbYpmNFigPRaZPbTXjt3OEYbTUl0xVeM0WUhB
/u7fPt1NX2KBe1fU+Xx0gvcQ6t+vpwixDvxoNUH1aYPcEPMvJ9FcbwfAEh7jt2EW
uA53F8WZxzusDcMEzWmCPGdkd698htu8THUurBJhdgCZgVN5fz67Bq/1VGqa+MKM
oqzP8o8QZuPafQQQzIrWlrs/FBPZehU7C8Ul9ezaaHpxe56vAHOS8ZQsILuwtU8V
RXZ4FGITKiT+nGFd/ckxjkslea4tHvHY/3DvyIBKsBGCIqcM64SSPFDq+rhPvb9Z
xCXgnEzo3g2qOS8qx5lP/8numRluXXQfVorf12LVF5NI7Nt+IXq3y/nhqPUlbkXh
8X5++bJPAa7DXeTqWJYfTIImiPnVWoDrDnN5/S3aSTHswrtayHAu4Qd7JzgqMgKa
SUIDJll54pJNOkgdFKw29iXpXQNGLdNb3ugJo+KZF6Hrr7VUu5rCt1XQGV5Wiyil
MDzOajoKmDhcSnZ/Q1aCcOfas+Ceat/HEm8YwOmsmj8kbOJl638935JTF/0hqXXM
5yA5imJdwSDhVQewHhcGIi/40spJ5zPXgfNEY7xVoJShyKAFS4gFU7aCCh9LbzTk
euVXPWrG3yI6fm9G1Da3ecv+c82PB82c2D1iDG4JpyUur72m1VMXEznT0tgPc7+D
I/CqczvYfOA/+VydWxSonq8NtKU7sLqfonyd/nMHWwC12kw4bO5tX18xLEi6uhUQ
lHqNAj2SgksXONSQwFtQH+XMi+45Rx2x9Iv04cYEBiLH3nqSH82huk2vHgk2e0t8
OzZmRX6dAmp2MwAGu4mIIds/7OoJOsrhHXYP98JDwU0nzWImgq0IES10SU39ZzSv
OejB/Io0BiGCgOy6QGY/AmLjrhEXmwtu/YTnsLpyCBuVDwuYIwSLSwAEGvOnshTA
2ZvH0gXZB3XG/ABpPBi7gxBZUDsu9M9VeFBoKlMHo1rMuumagoaLcEbjUVVgvTMu
E4chgDLyObmSubgcWTkppUNoTtkdySR+Kfu8D3iwvRFsW4WNxoYMahJBBtXmondY
bKz296yE4LFxDqZj+va1cH3WGSfLbmyEUNLvx+2WWECnNoOEVopFwxyQzlh9uZkf
cwg1vlaeXZMDjLqMrbJk1EB0aTscw71co/fKjaBfSY/okBljWen148wycQgTHe19
8GtccwECvI2zmptoLfkF36VnzA9wHaOkPmcYwPkSPX6LU+Z2J56pJ1RCEvC/aBGJ
h/HTEUzWYA9gTGWY4TIB4g==
`protect end_protected
