-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
PCI81sDXfqBJrc1tl4aX4im51eWvzekfkTJSFu8t5iPtrQZ+fbu+EkDjiHOZNlUS
Elkc9uRO7bLoIjYV0szaPcJAnnYQZD7Hz4gQrLZeQMh7pX75X8asPweaKaGTu/8p
iFtB00lrDOsz/2wHfpAxMcxFTHyPYa7egfHfuX2tAw4I8ftk770JcA==
--pragma protect end_key_block
--pragma protect digest_block
o+MAG9K+ozE6asVJ2tOp2qe+098=
--pragma protect end_digest_block
--pragma protect data_block
w9WNxt7WRDPkKBwKehgXf64Aur9ZI6S57fE4FyaHQlg4q8+kJQDKkoor9fCFOGpq
vDK5g5WhguJD6WQbdAxqxVyPtFASGtQMOyI3WLJEhHfylzxqfP45QnXlYrnUvuel
BYL1otxSCEWgcb663nKRclPR0+99KBI+UAc5HAynespOYqHYRbO5gBu4i8ypU6yZ
X8pcjrn82MPkuq+vuKZLZQFhkGrynxtfjZsS1i05soWErByPQ/0+FdSLDhTjo/VN
2AFB5hDxlypVuAVR3CLlH6bPtro1NFwEfvVg/7Ifz+LoMPJ/XM5/mLrnkQEB3KQO
Hxe5UAIDzXNaa7qKwjuJcD+uDD3Yvnw0fT9NnDN5C27PltMo+JT0SJ5TYS+gam3Q
IIceoh5qYB+yBoy8oU58zUrCQYCes88oG9QKIPiXWALy0dqqfX5AIYc9AuQghLEv
ytXs/RzMW9XwVGaX9FO4OhtAEJXVCf0y75U7A29JYMJKt4tsWXQ1njDdM/9g3vYb
17VBS845xB61R2vUoDDXSu9tYFifvUH4axPTkuu1mtFVQQpd1iNxi1tTejwlbgfN
oXhhRbbcSQhlhsmtfl5dFP5957/i5VsrjNIR3V5LN4tpBBCqFBDFXKSPDjP5yvA3
X+zZitGM+4+8tJH1e9JLFqqh66D4LKJznXl7+K7ZJ2aV2R3ZrPus3k5na/2mKqyO
6cBbvwkTmZhkhx6o+XOCgcVjDnXiw5iRYp4CxoPuMLN8d/fAiFCo1IP7aFThNzUM
Wd3ij9sXcjVZGu5WHPnmkuJe4zuLhEJvBtcRBoAe/3GiAAnIHMGGg0d21TLIRNqo
/N1eQISiJPq9B4eOpyLwrWkZKn37kM1JmCX/7zZCJE9ajoYd9uMqYMOQqjTGeqX5
/s/YEYjNzd+BTXeyDf9NXi7XkcNbXf4gWfJekLkO9yIWvRID2m/a22zXFpYfrGjD
0YdQyGi4sky32xnIERwdv4pe/l8t7PiTQWy7VimvfnSBLRQC6FgLICMpIyg/0Jlr
4tOTufIL53dr9GthsjIL5imwuJmUPD8ZOxo5QS45XOiywge+OqNf0/RoX4sIufDf
4E0dH20ZDYkrfZrujVB8hM41h0Uzh6ZBD4J59px7O1kwc4JcX6BThfrrbgaRelug
rztETIMquKdYbZC1xpuByw2d6qtQYdSTuy0yZuoVJI4BlviGREofmcchI7lVEuAy
J6yAhLS2IklU/7wjv3WJhLOh1tvPBEkE8BvysNmt36UJbZOR8SX91qumzJ0MYGrC
b4ZxIdlqMlH2IfJQRKKvdnaP/B7y2FN56HfFkj+gZ0x23ScKL/qq6pIdibLjk/3J
wTWqCgTq0DM5FBu5ro7RuYRfGFYO9hL/gErI2lUNik9Ie3leHbEmvsSGca0xEfPt
Jz/IWyXHF0lzHtcfQxh8YGptDHsv3iIPhZ9XABd96JuwSb9FhjqpDO+Tosi/gSYc
63nD3m9vNIKb7xkoAc8GHJd0a2EvXd3affwGnQgmdMI8WRSedUdvVwAql5dDHRtq
aTvVXfwLTzPve4bSTUmBfIgA4/VPNpGmWwFLZ3fUm+fMhd+9pwNpohyGRlmDyTNQ
TERieE/sSlLvzLs66moJvhPeQI+fxywmIV+AlUOspDnz8ClAZas7gDGbEcwrkOBy
J4vAlGx3BB/aLF35sC11g+Yd7J4Ci1Ftag3pp+9FkruczAWfzr75GHcdlvWceaQP
p1gJEIfv6hluF/hpCTymv+i2m5xIbPkUE81YQZ07aLxesQNOi1QAluIJ4Ou+6Pzb
P6jiywVUx8wW4E4qiqwjxN9H4m2Ub4ImYHEccxxXea7vex2wl+4D1SJnDjDYn/2f
xlVBv+CQ3nH5rbEt4RVA1KsQAOcLl8yhftSOWRPu4oa4nfFJxeqKJ6tbceOoFWDH
aEE5ZJAr6ZvmOkVIUGT2qFvJuxOMu4hoUKbqFPd/k13Z4vaJCP/H0mgo91FyyPPf
2ldP1a1z3C76gzMAO1BjvLSfYnNjP5MNvxMWXNZByPyFggT51cV4XzYDgVm1QgwH
ZsJL6WRlRJwOs6CJZ2edbClvpiUZYQPb++Gj/Pis2I9HQricq6gcdKa6H6M+03d4
C59y7FQsJBuec2xJLllL9rnP9q2nsJo8A3RsE85C4BqwH+MLj0yNiqvBxo/c36qY
fbbc0LsmlPeL9mWtEEWE7Tx7J6ieiZGt0KSZlrD5gi1VleIWn6mcFUcrF6eDgYg7
wSz/wQzwlWy+MN2HJQetvjfY5b1EzVteWKZIcshMLJ3fLVzPpx+PSo4+I2o5+NZD
ukIXbFomGvXGYgbNkKYeI3BlwH3kJjrRuLnmjdA5knfkkCBXUQ6nIhC3hlGxzoOT
zBpx3xVaH8kevUtcQyp7IU8Nlwgc1bQwckGxabkqgMkGKKkbbO2KhPK1xKtKyDp/
Bg2qlPhwiayEdJitz5jIsR/O8BTdzthuH2V2YpkPqc8cKRl3bnjtNPH16ziQeJNh
8BpE6OEZ8l9EYuhwxEgYpAOkIFQCisSrXpSKOBDEqZnoeA8THJfAt5yUw4102D04
v66jCZED05vlnTyoFVLkaHjLxoKm3b9iKL0hgb8m+52DZrkKmaiZ5Adn/w+QhScy
5xWVCHFNlcGz/kL7/GxipSbcqgHquD/WIwIovLxk3JBDHowrOBAHMc1+FE5PidUL
pX5/aeUZENz5E4m57ZiNYjqgOcmCml1/7HhMasxEAzATakaohkdmHM9qnKFLjkzj
dRWVxQ9n8n9wDZILgPT85AQqgfPNW4Y6gNnk7yA5Q/h2sVxpDTEnMbDnNNQsaA55
yIOgw5GVoxcS+QhkZmLWmFp2XBXOnaxMLplgZqyyXycm5uDXCjXNHsHi8uGAkN9L
Y2yZAViaOZTX3QtxRGurHWyM/EZD3C1WBHDwDiIE3ZgwI0YJ01WZaR8Z/XlggTkc
dAamoKG0cPI1TKmREWwy36ZJNzHrznIfkFt7+/VODh4CPeVIg/VFbk3jUMvVB2xU
9kDa0rfjOfhrEbPuxCZ6oHkU0bfSvJmWAOrmCzMSgGR4bBS6iZ5H3nNhbWuNJdhT
6IM0xhRU5gl6iuNlssmMY58gA6zgGeLjjZC218Oe+ByFnlcb1rXgXdm2Uo6AGW7P
6r2iOirQtxcI2OOPhuQohB5h0R0avWK4P93SDKFTEy0VOzR6dRd0Y+YeawratYcu
fP+fu0b71OdFduNtClGOR9MkDTzDUig84ekY8UePwyiiRfEjTBsTLYps971o+r/O
LmDk/1ynPcOSluspUZiuqUjRrn9ajoriGmugoCLv535PAft4daTguLFHwUmkcL0b
2ar4mW7SZI1eLd8UJeP69A3Ja2A0MGwP06J6yxOx5uVEidR3rPq3/DAROr/OiYAS
ZFU9IyGnub86naS5DPn9Q9AmsTuaoIhKkZn/2uNUhpuiifVVDlNtQ9yEU2wynuOl
frkHMa5eQtwq7R8zDRysBegbOV9rg/g/BnDSNLQVLsSjxJiAfiv/dWdPAAJtKJsz
OT+qifyUlOT5SbLyKr11PQtqWkd+679sjNQN8hXzB19XHAMUGpIqNgivqLKBxJfk
++ZBjZyYUdzHaeydy0hibLvR04+5eH8kI/tkiFSfCTaaw14xqihwEKh3mr4/29u5
cEUQ1KaVxE/g+rEijgi7Ghc33thm7rHchLlQKgK9kZGCuFkByup44addBAgQNUGL
wWoiwYzbl5pyaGg/laL8wWcRLDsoU+TjXYbxoH4GmKgy0SOsfGwxoxVIUa12HWmT
k8C3VpaOfZDU1VQk3qsKcNy18vLhk9kNGGT2Pfu/UnpH0QQ0UaXHvWuYnfEDy01k
A+n32qdeIEXhfYIujFQ7EvOgWWDuZrZGPJgfGl6PAZNkr8jLM0igKpKJ4djZSn0w
Uut0F5l5j6rtjPWxYwphkTsmDMSCfsL41Zmbyg3Z7LPy4F35PrHLXB2aZb/Cdv2w
NbHk9n+1cMn4Y1C90k4wE0qmIOwoewXRQauS+50GJznaXcd0B65vSQH2LpwrMzjH
yY12JbYw+GeUuxknPYjsNjAPIZ2RC2LykR1B9EA6OkuKB4M+kJdgoj75DDCaFWJB
qV1OSfWl9lvhQ5S/dmi8uisaNZnB6xVkRg4pUNrA1S0iIsJDX1NhmXt5mSpz3OXw
EZw3sXpBWqGU7M8S9ZnizCuj1VcNqgZ7zITvH7rtMJBDViT0Bp20VaBr7qoi1vzc
gmi5GHj2KKylrfONowlZRwbdTFbGoot8N4DtTQdV7A2Ao4RnAOUm8o+DEA1ujaMI
tPG6gzdd5pmIRCmT/zxY2Z9xe7v0KWWHmCQSXhHdCra1d6sdc4BkPCcN0kk4epDy
kQyw2UdVshdlLNmOtzJgT+FJ4cfuycK/2M3/LL90FsyrEs9UjtZYzEF9cgpFYTzg
t2yFVmvbxJE/OH/cOgaDvuIr2/3B3gId+1AKNKBN9TX6KWXAPp/tabJ+6VgM4RDR
8zR3STxgwpBk7J8Mr9dkVLn6adA3/H+ERVAUKZmfEgFznXRe/JIBDbb5T0T8kEEL
nG2wKySXou8ncppnw5hPoyxWIsQEEMiBygFO/qpyrENlLlcBUqzxNp9aNLJeAyVi
f4TVyNuisH0hOGNN0QpugcWGEaOv1vR/S7i31MSzxjSnckF+qJMfykesAA1YjxjP
ITOTDTMJ//xawFKOMZey44il1mlK3HsGiGIMlbZUlXo9RRwnRflC2qFdSqbVbWRE
05TMg2o8h+nhyeEWAt0QN8sbHSe+A/BdLNobN5GeaOfWp4avxNYZikLQPsHOetpU
xQujos/vRSiWqPFR0vUvfXfsVhdjwKk7G38kmNl1oFQ2Cng/mhOPr4TUOL997dub
0haL3Ya1OXZx8gsU+S1tefw7Km6odOLitAAnR5dzKm2M4H7W1pTR3ADfIqqvD8oT
+bqkcUEIUv8bVDxsZ7E6hzX/RtlC6uwtpXbx/hps+qG+djvPuf3ON+NByPQT8CE6
0kkcQYoxHDP4kfTQLHkgWo15w+yKkUTiGyHBbjcxmuok6fpNIp3w8UNv2uReRTqW
H02ACRQIU/3dAVW8dSmutVMtZzHR6eEhI+ucktV//hAwlKIpCXiayNnPERu95rF0
lNWrWpmN2F0feSACS+/3A/peE5KDHipfJInYzC+i570/h7kUcNt1OovMIQxNCbEw
9ll4ccNSgdNcd8MJOaUr8+xPz7gncC+MmCGzHxxqHCQ9sIfxwCMraWbkdmD/RwUD
1DhXlFnSvRuOf5v+Kvtg6aMI1cDlj15pYeGFYmF8l+JucI3I7poMkPqXX0loShw2
Qbe0B5u44ws85DC9dzhubOOUN7DAfGwyZyoQeIOh2YEiexIsVQjJTp3KGXMgY1Vl
ZTaxSuXN8mLr68IjGP7HZPjfbIdVoL2WBTZj4wQZBaI06m38i4FNW2monXo2zdQb
2xu5cJMDVLMq3xExZ+g8ccml5jwEYDU/dN2XKHqUWcMycRBqs5Nsf2VGi09jQxNk
f+21IRlgKUF9M9TJLBZu2/7KaIHMn6I5O3W1t4ZUJqjgweVSxlgsxGrPRmwiuRe4
oVYDF3Nrpk7dllbN+0RJtCwnW0sMCP9lU/LrN3IHXp+pC/TAuGs4LF/j/vPDK4FB
k6lkDJ4oUloG6F1xOfJOfNa3Y/MksP+jcAqtW12K2Bp1TULxBEXcmxnTamCe/xZY
U8CsXJkANEtCfnf7q61WdJ1iKyK8wOAnY4D8KnDLFh5DTBGDUBox9/gIZAlkSzZx
LiO1RbzBWhJoUWuRKC7skIy0v4qHXOpBYGyF+DTXlUHwr93XcpyzjTSytx1AN+Kr
yiDibeSOPL34Ts/lckzxxxwjseiJrtyTilQKeH1TJdDa0fcKjdUDAcss91Zbswlf
8yI5RkqjFaFmIU5/qKGKSbkB3qo/iqPx30jNbu6WpRuNJwhnYReTKmr/yEi7nPwG
R7PH66jdnf2eONxS6SE0Ob84/mWOF44WN1FPLetfbPXIA16U1Ra13pWVxPMGYum6
lKd7ZN18+p9bzQyqcZCRHk3cjaTGgUpz8T/RNGcXbN7kNyGcJtnERdo08vWs4kxb
CVut9wsLAovTSlQmoDTq7LhL57DD+ZmS7gOAuKZjDGX5P9zAOS4Yk34UyNHmkh+X
Na2yciQ+6JFONF3yyFOmKKGbHq3eS4vd5kEekzaxsCY7MVn6UBAbmqBbQZVUE7Q4
+lMokqJ+aDnlv1gTv128+zAbF8gN3+pQkDX546aYfSC6iOAqqbKGRfW7bwV9CphC
QthuAnNtd7hXkR51WmxvMd80gkTXPuq7dXCrAqoGbYGN4Cdlcm5VMS7ZSls1dMG8
Iydp76aMmofZ7tUroyiOkrsiUWXzSdXvGevsGt2eGvETwIV9kJy90Gy5RRGD/CLR
YLAKqhBq0B4Sn6lg75/EkLKafSfOfdQ3Fn90eDctEjK3diw+iBqo8orC/kasHj1D
EHiRg/mXyrW5Z8fnHiDgz+8VchmePiyPfzaMbqOz2THxJHk6+L39KNoRbsf00vBc
XntAuUMw+mepB7ptKCVxvPENrYug0Ab/wkkcSfI0hE6BxUui6Tnuv8ij1FD6Ab/D
OSlpqScfdGc4gF7YQpHTGZOcXFtZqkThnfl1l/+nqqGnok8Ob7CruDqBzBbCv6D4
4/mfEOav30JxwTIYSKjQKkYfG8SKWQPDR4YxJNCGNuODg9zLhnL78h2EsgyBJNJc
6WGEj+/YU/N+/5T39/1aMRG9WWpRfs/E2Jte2W2VNjf/6gHEwfLvwKQWOMRdo0Iy
QaKr3W//kLTXSG+swOGOdVdnJMorbB8W3hRaQRzQCEL/mmKrSETKmgZNG7S/CGTw
vWQVWg9H7f5AHOofYZLNDoAmMq0kOhYhgD152aUWN1t/n7m7ao1MXs6+a8XxUnWo
oAjyhQE179BxuNJjfe9FTDz7kARAFGAR9Db37TEEnjp9d854d+k6G9FRpxAH2nZt
SBJCOwa+Aw4fNS67TyoiFsxH8CKtUGymwk7TGfWGTZMBPp1oo5f+gG9KkwrXX3Xh

--pragma protect end_data_block
--pragma protect digest_block
oheQWHbGEwps7P7YWKR3aDIf5n4=
--pragma protect end_digest_block
--pragma protect end_protected
