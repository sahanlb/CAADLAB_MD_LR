-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tvM+qCq2xVJkGyQmv8ysGueyTLlVF3kphKmRkAi8UCYx/iEPhTsnkuWXBhlpRH4SgW81TNPdw5df
5sKGVeiRDxgv+NjMFzgmBBb6fy1A2X1+XMI92Nqg5Pzzk6TqNAM1VIBz1hIxKc2If39tSCCgPn2A
K5yaBeUGyjFPv4e5H6R/YqQHAz3yme5nmu/ztRAhKmOadGKOCXzv4vX5ro4eEatMSaEWpjifuClJ
tGQyiyX+EEtnUlTSZxzb5NDoZKAVglEau7BOoaeKgwLyposskFpe+fGRKIPrYJLjY36f7Luc9fD/
zIg9QfywMvoMGlwQV3ruI1Q2KhTQMDT86b8g7g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23312)
`protect data_block
DX73ZXaBY04EcM0DBasTe00gAS7/bMp9VjlGIwrFB3PvXEw3xivlEoyF6L35KgFpgMekEqvbIlUN
XyzEJPvnq1DdzxjXlYepDbA5BFx7/OIECAVZBLhHSv/eaJhuBh2amnJ0KdFqxb304RJP+euV+fJp
40F8XYa0B87f4yiQ3MEllNtR+g0sL6FlaUzFpSMe7nHBQZI5pk6WT3yL3XvECTeRlw/8TVg3VKbT
qpx04w+Dh8nTDZQ1DjtthuNXMnGnUudr5hvp2XRfngnU6jnRpOUtCJwaXghoKHaDIaqBvUjwZ9Ua
2ozV1lb0t73w3t//vsq5ApSoGH6w3AMkzb57lSEVraB7jLbIjD0GC6Rw80pJSMPbIhoIOARJil39
LW753LdAfejtLxOdMNndUjZRTXxa2ASzuZ0ghMQFZUpJ1nbqna8AJDX98aDnv+eFtLja5DIrhPNF
lWR6EfRkCZWcVWrmFDWU07LOvwIK10XcyApvAHwjLHr79Aqdy+vBEffoywie3IRIQXHFAIQOrLAl
0EV55gNDnYieH3o5sj4LMzBcII58a66APjHogi6Is717yc1HXTj7MEStze+T45QU7VYgXTF1ljrW
PnMrMlxKlSK271ka8hD/7DWQAhA5zZDKmQNYJboQ6yANM7P1K2yuMAlxltlC7WShgs93FpN6jwWD
2IVJV25Z9ihkKr14viJv2z84OVHsdKYMXhXE0NGFzqlIa6LKb0dYbOzKOEp58E8njzstYftj072C
/IU7FHFjDw0qnlhaG4T0bG2dqOtPAxGkRopdPdbEc9VzhpD8sH6NYZ9YRwWBt6o5cYKLkVPWVyI8
cja+coDGUxJUTU+NfpfJHxfZv4uWq9/s9dGrPQe+3yYhrYj72G8l4FJnoQVkN8YFJEmAEE2cSLQ+
J9XMsv3Wmy72wZI4IaDAnq8EPynDUysshYoncAZJuV3CABYwQwMoKWpIhstQrIHDzhO+2FOtxvOG
Ddr3u46ng0p6JE2M09h7IQvZ4fd8r8pStD5HYatZHRNFhEVRi8oF+q1McXqPzxfeGCefK7g522vx
tqzquv5Hns/I107fLmOCMT05KrszOBPIamGZ7QZ6IfOaCANrW2cbp9BZWOcbL9VsUGH0kjDimX7M
xukfqqqs/tf3SNFAX/w2AZotsiSemxKoS6JdAUv5cagyA43rKPrvzWNsJBkrhulPIEIP8pODDRqz
u4KYZx4199p6Vr5GPi7hDdrbYlqcfgncqRccfntPoCGaVC4vUR6B/xvx4YwwaCjQcixz944fI94U
dqyKXdM753Bx63tkwIC3ko1v7nvSyR1xmQNoyMaI15CGc0YOpOGT4ZGYfc8er1OCXpJjbt2Enh8c
MyEpUYZjep4vtpBf9mKcXn2D0FTW6gM6+vJaz4jC/aS76XHsBVrepdzAokg3aAZaj8zqpR2Ijikc
/M4OdR15jfdQSolxke31g/a3cu/RXzsJ15TjJbXosWl4l5XaJfzfZ7mNUJoDlomL3Ra+4+JT4ktX
CANCWn4c0J/s4DXxzIH2ZlsVE1p7SrS9jbcD3NBGOiMuYpOCRc2nXvodx43O01GdFtbZHT9Lkskq
pQdh2Wrk3AvmjmogKyGx2P8CZB1bvNCwIABHpiS1xrs8NCW1d77cNUk+aZstlQMEmUdltwVzTVNB
0a3IroMpFMRcGWeqKM2RXj3gVXjB0mk55xL04cUCQT/kJMP8UfZOUhW/Arm9EAvS8BPyOjomvxnm
/EhZMQlUNuSF6qW624pfotDR+u52MjAKgOnBvCbtys7nFB3U6eNfX1cKMV77FcC/JGwK+q+ZSJcx
1hjiMgBzMCPi95x6n0n4NuQsz+GmbtAZ6gIT0EXnf6XcHfGINjzm9o88nVSMw4NMAjwS5NqOCtIk
fGXfjo1nGyF3LotcI2jBlTknLin76Hn+SCquTr/7KnmTE0c8CQew0pX2mpBDGaQA8lcJoAOwITlP
SKrSiFoWURV32z8ecdPOLgeRnjTelgZBex9t84NxNi57s8zyTgc4wN65cuG3YirW2EACsGjqbxDi
WZ8eSqWXS5jcx/4J2E388FzwPdP1rFH2AomC8pnWavwYWp0gLGFRqifJAX4OStKsMjA37W0al/lu
NSN8Ppq55bjKPKmsn6afBoQD0yeSKgRumpfdNMPdSa03KZMv1hUckUSFr3YKVE2ilzLGPzWpm5wg
JSvIWCjeEzRjkfFWvu4oOmifFdHzDJUFYocoJ/iP/sjvOTao27z7aLRlK6wyUseOKejvEo+LbfaW
ePdev7nXYJqt7mL7e392ePk66g4jSVko1WF/ZY7osI7NNLiHW2lXgz7/8yrPXYx1WrkwcTwv23ZC
4ncS6HuGru529SX5aEfzQKzhrlFlHo49OGQCcG4HOBJJFx0CoGOstbr42l0fiG7fWRrRsYEP2GQt
9nqZ6hNbBys1Aq3u1AFCRCAjIv33zgcgARd8cEzCvdX59a+K/eEtCrYGvdioEEfI2oYaXvkYqJW2
23Ixc11zDDh+BBO/aHzIhHurbeBR1M2SKS0lk+ePlcdwX8hPUwcYajKD9GA68aE1166sJ4q1V6xY
viB9/1sHn8HHsgYYpc/GZ1xY8yCTPmrZpySLVsN4apDCAT74J7Is/fVikMtfxx9raxDmKPdiH9KX
7i8vUnX9rRfemByOjWWnMSBopCFxJyuJ70DA5rAYvztNye4PWCGUqSMwValJ8BuhxfpDy2oUhd1l
R+rmBsFr+kDPzipSRKk/WHvzOsQvW1w+1cK+ucnG36TAhxU5ir1Y1U4BnYeI1yPCy7wzQIudaWDq
LyV8pJx+kj77VL9DuQSDz2YbrsuL3Hn9QbUIJwFJEUlFwTwT0p3H8MLuQi+IdeldemJTh4V4DL+l
2N6JRPRS/tbm7IFveqAHB1rdDtGPFVeR/RH8JhxYJ6Vpxt6fmnqMUhT4XdnyaxslCvPDbENI9CBy
lyG9c6Uhutn3V0lN9Jc/x6R8uDlk/AVENRAU0BU9KaAnoalwUkqZ1IRV3pnjbgfiIBROPGQQS2vE
5QhvYAXjBQxqsCZbu4wEQ9yJ7PkXnSjksbxrttdQn8chX1ounNTI6Yi0voRENT+3J1pQWw6uVxtw
x3OEiFNfeczht59pXUCwrmE6nVoeE2e+bhxchXB5MFehB3t5T5hAKPXoxnHCLE0LrREOzn3wbEEr
Z7Z2uLAm1dp4E34AOgqqj924Av9J6l41/gaEzz6bDQSoGgGESuU9eZqrU/RPeFdPqwUi9dJwvzON
v82msNQUXm4M51n6wZ5ZJF4w8sRX6KnQ/9pjkcmcALOZFqr0k3G/vZOgv2ACtf22APjO2VQrcvP6
yf+saC/mFuR3g7Y54tffcs51nH19ouWDrnZ8DCtbtBDMBovjIU5BL5JrMAvshwbgBDw7RfVDRfr3
NG3d33J58/WkaOza+YBA0cNhB4fyyDxAUPROvuccOfIMpvNpNUlJaqW6xfB9OotL2/tVr0cUbXd8
WLe0+7+eGiJmGGjcu/9UHKPaUhJ/yU/KZCFsCT67X1mQ6sNudq2kGxEuceym8MpGTUh5wN9lo3aE
EU/Lao7QVz0cN8IFS/cki9iQyoACQ3hKrRIPdWvddCwddpL7LqCxZ80peoNQ6SZyD5uBLNTA8R4S
MkM4uNp9xeM9sOrO923P3trYgwiixZNzDyFTMu23/fmzRg9eN0e4F1v1DYJRbMKCoLnvgXLmCNyz
geBRess+G047Gh9b/oj45Z4MJHrzu7Ihv+nwYFVfOgK5p5JGeV9M2uV65nIX7M5Ej1CR2aYDg84Z
gS+d/JvDkAH6S38r0a73itri1ADHy+wn2JUUmrWHO13/nCJn4vvB/lNnc7WqmiueYwfRJ+o4SCRE
UScSOEdhPHenqc1EUT9f1G+T40v8aYbGiOYlT3HN2dScs+tcC7/QPqnbV56aDJVa5FVrL6kHf8Ev
z7Q+2zoNjFrkGLZZaQzL063/SJazZr3CttGbtaVS8NaAkW/GLQXFwBKp1Gp0ourhCkci0LA8sFhS
C2NujFmPdEoP84/lDZ559k1K58qqkRrE1ctEAxKc22X2bVvKRlKHcpsvYdugqXJbZuzn35Y+BAct
z7pfPktSGybXwh4bB0vbLWD5OEi8OzvROmXoZMmH+n1ZKdPM6yY65a8JG2s3f1uqIF4QbEIHA02s
zVlDBTEAKnKTS90AaWK8eWnzjEu5EfjCPh58WhmYLjerJbN67oKlL+Ie0r3zNywW0UTfvKdyf1jJ
G2jKD/TAKa23QOS+vvNjgSUjAx70U0mOBDJ5qzBaS0TxKoP1wRhdYxDmDzR61BmRJss7UJp+8gx7
EAesb+NDuzSx2TGXVd+70pRCtJHWVQw+TmYf6hXK1mTWfamuWx3vgk+TgwK8AfULpS0exKU2+aJW
qlWFG8DgBr4WfwWktScrEqPI6RyJaZaDfQmGQBUxJ09q/uNeH3YHpSW7ikGIQ+DU1S6bSWuSunZQ
IufJMJf45OkAmqhBjDS9G79Cfd+bp0bfv002ZDjW5J5e9qYQunsAoxS6Jy7Bumc6L5T/v4Io2AV6
CGPHLwm7rqM67PEEIXbUAUyp1HofE2ym/eNdhENHKUH4dADP6DleaPPs530t3OIbzdXLKeWN8iaz
5ZU/1Ar3z4BTZ4jjDG7Os4bUZ/xGiTKb4XEawKiUjAVtxiedJS1Og0i9C/F1zVt3SJ2AEsJ9w0fK
qn3cllTdIrLoyz9uzE9BwyYZWD8y3VuA6j7a6YboQhgCvn/eQbVJVAYHdPRtz/vjL9pFY8dvZ8TV
jLWyJmrcIApmoiREd/CQs2Y7hy7h0sbtroCtBNaUOiLRCoKz7pIqP7i9Ba/iYOaA5vuLmzAt6zo/
cf7dm5tz/EBVlB1xTWgRe3OogD467Z4LsbenaybmhHjIk0fRpC+GhDN4FGc8FrzKfUoQFAXXxtc6
APAqJZl6wigT413VAT7J89bXxLO/vYyrQ4VENY00/g6MG9ke+QYUdxa2xTVE0NCi/AjyKCyikMnb
9OUeb0vjcc34xrptXkDC5cTH4AdP3Qj2TSUDIwRjtc2jPtSCzt45CGKVprlorXT12fILg614/+Ae
Dqk0+ffVftQe/U4y8qHDzSiLy2avi23Hgxc6ygzExLL0w4K2nXsFcgtGav12X7ZIaacuSB+UET9g
2gyMCRanEVFtSQWCphvQyOWAgVzD8x3+jFuk0tvzTH1kQD+QWcUmjRqpv3+qdkIkylETHyEetani
sXswyVxpLEr0W3FJjaMzimcv6TfU03eKeIWePD5WfH+qcZKhV+Ga7/rCazA2BzuzmI9RN7l28sC7
Sc3NPSO+xj31yUEoIKpcG35XptE2buU4t/5+aiD6aIt9GJU0qHyW2YcHyiq1e2VgY2b+rYlWmExo
HC0fDpzdWjnuL6RJ6nqei8yvFpcIIsix1ZzxqueK8VuXenn4guovm8Cabd+vX3h6c/M0+sGvdFVV
Hn7N2A3USy0Z0q1ljZfgz4QFnLS3KexOLlkCpRm+aOahN4G3LRfZ3VXLO5be13w4mT6AGgPSx9Sb
Q3/Ulod/rekbzwdfaXeEPucdPqIg4S2aP+RDyLMplfEPOh7YNaSVmBuhaN6eGP4Ongus/2kBtZPm
Rw4ZmprPWAU5p+24wueSPdkc9Uanqnp32LpEeeTTNe7r3/kOy1rPf0Y7YL4Ng8hojrc8L3DsjOAs
JmpxewsK3SGQlbMSDHFmpQMQWJmyUeHoAQjqlkKDY7UrS03t47pJo5ac8gdGlEuU3Ll5rhRZ5gpo
kZqA5eHdzyybkokrTN1xrrXCx34ePUI56vcYiOd7oRivMf3RqjSPblTMaKRJRIONY+LmgE0Es0vf
Ky7nkkYdPPutwGp9coV09+x2x4M67Xqaxh04PZhnCo4BOq7hgO2jiEK4W2pxwvr13xcLvzQJW5WR
9G7SIALZyVyLT0deRxhZgD4vuWDzlfuM0v/Nj0ML9IG/Y1RW7UYMDelYhpwSI52TV6C9aEt0F0Aq
bNc0PPqYZ4xLNhBz+fbtcBAml1aX4jozRxuhVcxs9xbhmIOK0RS5/MuVYWy6dfRQN144cOn/QyWQ
nWOwMizMLDVJPOgzR6H6kgHEmR0sVaYpdW/jOggw6K5+K+pJjhgB6UjmmhZGtpa4IDsZO3zHHoxX
O6SaYRZbBpZaMl9PyqdqyBF4cLkAYJfQNj/+nJr0kaqGmmHZ7RcHHr6DQkqahpA2/XSvf/NcFFiJ
hmFJWs0BACLu2XBb9FJkApto5+fC1P1LyhtQwCOK69mAzxKUnDAgTlNRdnSJ04eBGhCre0RYEPTc
g15dh7cxZhSLO+efcUwe2gUFgOm6KMT6JagV02JLNYqrb2AFl4+zADRzW/nkNmIgOP7agtnwKiX4
m+8ONtKKMxC4jOudzvl12OGjp4QVHGAwgslm1V/0DX/XvheiaCbMKxgrlrXFRHeZpe1pGdfXJTGw
rPyF4/gphceQw2ZiRbDEH+FAs6RUBQYVpSIvcB6CdUqXSXH6o/Xz+MZPEWqxNzPR9DXd5HP3XxXA
UztFCfAj3vitXV9xzLv7QQoeJLg6oy11dXsJJlYiQjro0qmufY9IRE0a8UbhJpsC+//TX1yxfcqx
a8U0sxQguXzbR62Ga9SrsZlNCpaSfspOnehBxODQcEGjRFmXm8Cpck3vJpujYoNewzfkwlrhzUlA
p3bH7s456FElmnqGe4ZcM40XIX1xFY7KG7D063G9fH3bfdjWAMT8YmowD7tpXCngcto8q02lIDte
tXc2Vy/NN1ERYjjZnYG5jLndBv7z/hTzpJE1G4erF8YGSmRl2/IGE4e6qHSZn2yHm1sddYrWfaZ/
lbjLX27LH0LqtovbHA+JtpFRWJgVojURA0wBcMI/Uu6Rj5YbOdnezUF/TGXBj5Xuj3lu5gXkrHji
UB9pJIKuAQJnofs9cm48dzLIpt7YwjLcpNimCK5KIwesuDHsiF2uTa2VghFBpFweGaoUia6YPIqK
YOEHM2xSS7CMR+1A28cp3Nm+sAzntjttc8ecxRP0hJ+Q4jJE0sCYvf+n7Ho3qemkpqPT3ndo3FTL
43Z5RGEXBbRvBOC5iMuyPIAqQOl/7RC1BZB21i/zcUgIeB2ssr/uF6BIDLr/9m+dFsMUK2x0nAGK
lzpxMFk7n//Q5IyxDcREFPvOb7EMtPPvVxfyja5di7wcXpK4dVEt3clrRGtbbAezMEjvpoB4gh1w
CPJKmmMfx06mvwJ+RK8cvi3ji7pvh5lM6fPRf0a7RX+qC6jvqh0GD/2W0vmqML+CnnIUrOcfL2RH
N7kZMeL1CS9DZ2vOELwikWqaP9S9CkGr4+dYvjWVkz/y4NZrrTxKkS+EN8Vk6M/+iBLFYOzk9794
7RKfGfbNPCXXoJhsWAf47Bvwt/fiM2NWtv5RDDZbXEYQ2DKbnYnyq/dwnYjXrEiaIqqpMwBJXT8A
+Q078tJGJmiE1kaM1HwMmmNTtcCumt8EYuaXG3Lt/0JG6WhJ7f3y5RNMUCiZx8+yOEJZsaPKl/+/
2SDbcWieST8yDspZfwrj6OrRGG+pK4zC5cxbTf4NGSimHRq2igFmscDcqFr6KNkpSt7GjUOoQ0qb
N6IJxzyfdD4nNDr0a/YYgc48uBuqnlwxxY80KbsqjTZ4a4zXJvQrqdQY6j7NbrRg1fCBbnSVNvfZ
hJo/61f6vJtde/w+2uvLMsNxL0teTfq0/Wqtm0ofOdM04ILdbn/XU4i7Dmtjbj2U1tUp6cyosiTF
FFIlf2xfUvH6d6Y+8snujkLjsMqnOwXzt3jGgBCaDFNpnCApVEGcmGUiqCCF11mvXdC/qmpPTaCh
rFEbqQq8zlu8Jw42Jf3FKVlFBKJ39K+dTQvs1vZI/WdbTt4Kq73WdlL1dHeF+v9gfs9v3bPDPixW
3jKfM/ZSnF0jnveAH3HvYDFfYxexy4j9aerq9ipYen0mZTs2LUWfAlbZGoR06xjYTQ1kq4YlWbvZ
8jXYB8imHRjI+qc2awn3biBkd06BSTJJp4daokeNJ2DRUnBIptUaZfnV2AUkJGBkMOVCjjsyaAxw
Mh/sc6jL/0Au65VlxUE373cMkeQgQ3BsKLknDMQXVmu5Q2oatq6Leqgg2MTC/KXPbmzWOPW6HSbl
IOk0i24LoBAJiW7ifwm+e4glpFabTnGOEICbjfXe/Q8AiPyRM6jetwbK7Xf5rfo6MZY4FKOITBWu
fxXadVU9gzgq+uAZ24o9NCi8QPB0zX0mz2nvd6xdx8JXC+e4XbVKvOsv10uPZHU1udQrfFAwuXMA
DH22I9HJ9OYD5wqZXXgWGSoiFog86Min8RRbEMEl3NSp16PwNKC38UysxI/GK99q+li86CYJmB5X
lpr4gAQHx7hdNMM4rvN3rnQE6l2ohyGVk9fxyTXvOiFv5hAlt+AEVtfVMY4Bupu47N9FdRZo5uwC
oU06R60u3UD647FFl+ZuhrHu+eumjySNRhhgWZJ9oMmdIMc8SqltdDJHirbBBBly//JHfiBy7IsU
TbhyK9bOl5J/mK9b9g1f2EavUjeJKnbsSORfX7Erq17u+HF+LU59oYOIm5rXbY74j5YwZmR4OWTy
5WeE7eE9wLlTaCQFAYVriebuXV5yRMkBB3uei9PjhcPzpRxynUtHMgDRYtRlEUJ2R/ak76KJxD6/
WycLnooLid7j+kKtkR3EYYTSj+9UgTAcg5W2P4g0w9bDymf3CyD4O4i8o6jtlxczpV33WxW2k4Pa
VGYPqEuipteVb4ffNHQkZdg0aAYsCB1u0+A2mprOETR4yzTJtFaBycrfLJr2LhFpcabLOAG30m2C
P2va02jOWHo+tUJJiiUwySx0LUjV/ACYE2yLKZALUfGEKfljl//qzu70bPLSC5VzH728waeIVmAr
QHVaQL2dpHBv+Feolq0k5kqcYqU7PEHuVF60CI/mRYrrxD18oMbdhj2gl/6GwUWnsi4yruCNkL25
k7sL2GE2MxZ9hktCJLk5FfyEU+atkIKX3t9JgHfsOfgoX4k1PfRN/1RrkYQ5onXrpcLZJEgNIJP9
+yHtSf2ksLsM9WpevLOz2mDBVU4oZCbZeeLETFS84idGopKz25UfyxSSx7KaOh6iwOlPRvohIFBl
rQczNLk19JzkdM9IAf34DTsXxwqGAiHdiXrZg0ULE8tFpdU1UudNcFi0Q04UK5yuHNB74h1GPaGl
y4+A8tfxwvFdfltc0EFsK9qVJE/ITqveYlOczkwkLbiH8qDIhzd8w3vGfXvWRd+GXqOqRaCn2vHV
Hbd3/ySpUYUXROHFfQNgvsOZ0ztnKBjF5mk8Y+kcH9xj10RmCAVTTSIs4Ev+2U7QiVp1VovDooNe
N50JupCiI7liTXmbeBl8oIYaBjI5H2nvNEsulHRIRHIeA3EbjHXkxdWJ84SdBO/BhbeattT69+Bw
gEtLLwPZaOWwPGrgT/50DCL9+PeAGVqCoOfdXzqz6ibcgK8LGKarjIKL+NtM4rLnzsWsVvIewe5I
pwKzmBgz3vMtdpvp9M5dpjxFP29V7qPuZn0wVTD0FcxJNE2LWBm4jutyz6J4enWmgvs7H2Wwl3Vc
H+yXL5bd5zc6Ya5eHp53k2K+Ay+jYW7A4IHxKayO1TCfANqU7Ju783LGN+91sv37eMZ0tfGxZVxM
f03uJR8FoTpDlDQHerygLhpeQz1RFtw/+X/+OBjQPHOV4M3dVtsXNbFW+za36intb0EckA57P4wd
g09uveP5ZuCkGz09x51kcShZ5j/wPnrYfsCflE6LuC/wj4/+JV9DpW0kHyjc7f9E+Uqmj+h11t0p
ywB8YF9jCt2l75bA0LJkwZW0XGK5zYCjYVwDv/J2q5I1DG6zroCslRFmHEl0FzmMaxc2Z7Fbt4r8
Ar4SSyDuuDZnTAPhytJS2FeVuO6n+ltNn1KNzZkzeVGABi2S6pXLeBfRltp5FEjsOeafOlKdql8j
fjIMVLuIgrmK4NCiSZLfU7UZwIJS1r2tewuaGHkgGfgVHEiG18oG6rM15h85ZCBoVq+duDAI0x2s
e3dGeMHUSROe/L/Pv5PQUyDBeqbu0bzvJa+4G0O/bTfoO6AbNcssNWX6SP0umwBi1+jdAlTI4EYq
bAPA1mtKxM8PVfSwOpZ84tZvJs83aobuIx8AeTgl54OApkrbL6S34XDiuJtDTfjhhxwDNMny3yPn
9wDoDdRWSy59IVQ7ft2FmVsQYTNo1WJRRjF28TYyfbdylR3bQszS9DBl/7U/v6A9IDc73TuaaleC
1g+1HT0CbH7CBTwvkD62CQYBIqKNjGuUz95lO3tRgfMMjezxTkFMPS+klbRQhnyow4HxndmmFw8x
exP0Uz0x7gNrhtP/PMCmVjW4tI2ScyKA/ZSDQOef8sGtSQAY+u+3jy/7bbvUVL6pai+EZ14cb46g
3dSEXdcVtEFKJrQqwA0IK/AFnmPFTVz+QvJ4LBsS+Ztt+0+Et3JqHzQZWu1wG0a70W1uKCNwwPij
2grae2mlwzdA9tVPktvZeyqdBHXDNY/AkfPsH80QLDevkvox9FPLjxsvbLn60maGFIgap9d2Ut7c
2wGiAhff+NQxvLiHdzdbek7QZ+IROwVmrgbXk6Fu3YWi6Qis3VYprCoU9Ls1e1dKFnUy8W4xt15N
KiOs3ksHoAqq2h+fhociTM89wbcPiorkVWZSg44B0W2T/kSLqonF4cGkIZ06OFjp06SoTMYMi2PE
I3mFo69WHX/dAegA8b6sqfcGWQdVT2t2cJERe0+7vof6qJxVaFoz+UaLOxTenlneYCV+oDVscNqB
MXo/wCJsCblvP7W84bG06fL43ikvnUavlZMVxeHarXrxwCaVKUlCDWqMoMzhJ+tNtIeR2LQYWPO7
9+mx4XGEm8jIULlCSr6WushgLK/J7b+HXrbZFma4j2NvgibCbWoNFsxUajmhA7xerp/ai+uWOyLl
uwBGIQtRX7a8LqljOhk6m8K7xHzZ5bEq7GnEFz+3omLpKLJwtfRXEDffPTrNHlIUfKpK/T7NCGRS
HKvBHFp7PzgMQzr2NLe2M3peK5cmOQ821Ljz4PHH/CEPDaBL73+/gpU/de2Vm3ovqibnYegIDZj2
AWunsS9zSs1k86T1mZji7UmSL/U9fOHVsCh9JDcuPUM7fNftDzvegqTN1vuV/Lqzv+J+nkuQgUEt
fN9ho3ZV7yIIhjGeQmmHQvQBtxEm6CojS5BwDewqK9nigQ5BaoGAx7pnw/6oyrlVpirLdKsVSZ6h
cahZ1cMMvAX8bbs2/b7Z2mIY4iql3QmIVG0Ajjug9HLAgeI3TNQPfAzBoqcvymAsJlJl1GfYlsEa
A0xhaUcHG1rmg6F5uKOxDNGsj0cNByY8YP7I1XV3PhfWjgu/UU7fxTwaiVEpjqQz0+fdDQG2RVq6
Dfpl7xBCELqEc2unQi4ImrYiGQxUqJWRFWXGim+zGFXxA1b52T37r3+ZxwQiBAj9HU2BSVLOqIvM
/sXss+HS/gRxylGAciiDKShHHekrgCXTzpHFbLSVTE8WlEiOdx7DvweE7XDkOwGC68JXwIX4GupC
exqcn4U0Vt6NVDjIs3ZjsBIwagH7GYqL7lS/EScl4kxhvuP0K8k70P6Q1TCp1yVnVLsO3agu45Fb
akciNUcZ+rva/9UY/DgQ6wK2f1HlAyTG4CQrfhg/sK2GMkUDrQ0bC2OyLJ4ps7dDd6+z9MF1aN1j
O2+TJOZ9MjyFN3zFgFAG1NumTLGr/WENA3oLf6uM/rDRpEZ2w5FXBp+GPaLt8p6dLdj/RpxiDp6l
O34hfF7WBTcPdqVKWTHcQDjqLpqUExUge7g/jrv05cLAzzpkZh6Zgd/pgyAf479eA7wJ4J1qo0lO
GMsToreyBTeKSKY8/K4878an4owkx9LoFRgJ7JLWGp1sO07Dz/P41SAr6neVqL77LG+TwgpB/q5B
4RBqfry672zjs6S0o95ljRlMLL05byQX1oZ73riEbc0H0EDtU4ennsTezHWoj62vEOs2UCQqg5QJ
1NwwUTmvyMMG5s5SSxrVDilfR2jXieDH5lmiTtVqThZ8WhJwUvBjDoIXaWvNp4pPpcr3SkyIlg7t
Su4zCphsoDPyDeY/p3mPT+bDVhhwIfuCPdWsp8rB9tLK/lVrf+H+NMT+KemV7arPBKTBGtiTt5qt
Ih9vaFJQx9V1PEmO/j2TcuTmeemvZGreA83h4SVRlC7ocxdc37tgM11o/8UI1pFgR4SChOEec+Wd
WWzZYg/1xoebqIbTVyigQIY423RUlUf4Ns1VBYRJFnxUa8gJY8jjezpNzxdDujaweGV3/7kfUcMj
1lXWFZj3/VeHw33qathAbCX5mtWpZJMC0+QmfS9yzip6Nerk0TdBIhdv1d+3qTxzzHzmbFEgtTDj
lC4gkSWeakyhvx0Qx42hEucCUfZ9TV9db7E0ZiP2moI9hGDWinr7QQz7ZSsyk/yvXh2gD47vHWHZ
toPf7GZZwzOfD1MTuIEn5HA8FatvILeUlKxqXe8U4ov25p8qLlSqHRYxQImB45abpWf9wdFgNak8
yqBiH5VL1mqBE6/JI02V0B8yARbcUgjySJHx3bWT8/+xl1XV122YYqOypGkV0AL4yZET8xpSv4fr
lADeZjKBO0ljcz+oJRmXmjc8Sw+bLUZ6W+6LA3KE2mXLjXM1ctqqejrKIz4OJmyCs8HCu421RqBS
pQmKfA7BM9aFX2wj7miF/ZNXrHyr0J1h8Ultrnj2n3FYe+zuOlEoSBx1Ta1uw0PidZzTHqV/3pCS
JrwHrgxqC430K1mrmLIfVs8RUudBfE+X67Zk6oZzAsSTME+G9HbVrmXyOkRURM4mbtd9ftvywRH0
Y0uMfALuJpkiEthfbSZfRgPzgfab6e6anNrRSpaIUMlmhL2sACTBH91a4Bd3SIj9GowA3pNJQrk3
R7gYel8f1HjT9i5e/rTC8FOjirvGAKZ2TL69kjSi1r6ng8YbxA8NOyBNQpViOVBGFdxM01ZrXSf7
pV0gHtAt7PnMLWG2sYaDC4yJFOngrd7zTZJNI/H9Bo9QhK6H5l/3jNfKcHlRoMrje24GLAOdzltR
6+wb1orcLC4+95bau9gF43gJ98Vq1lBPi9HU/yKt6baOYjTP2hHzwpqz64IhtaB8Wzw6FMzDwy5R
wIw7Qm7ZMjemeqbwCuLnK3jDN2jtgYuVfj4jT/P5bx+5lCAat6QWSPzCI+FM/a+m8p40yQTI2Cuv
4XMztLbYkQTPEuPQPcMCNmbm+qocMf8nky1nZsFA7jg/U9lzhlNzyyoMG6lJeyrZ562eJO2Pr7S+
V/fLdOaoYKceKpKsz/u+8faJ6FgJ8GYzqvHGZAPGU9S2DP8sWVPiA0J7Hjim+ozjiPEuh9T1THyn
4Nc1eKFOYq5w1If9ddfkBuB6B6hJmV+g5mjcoclx5S7eF+sCqpdlA7gOWZ84batmQiz0KcAT8yWy
wHt3eW6BavIzaln/jOFcwKZ2TDhUFxMaFqBBjJYIQNVvSSEeBhNINi2rEZZvvMHdyoiLg2Qw16cH
5d2bzM8Iaqf28y6gEe0eTH9yTYbej9+ucBbcahpEcr8+c73eP4gV07x3Pm9JYJbqR1ddOeDGof9K
rqLc4ha+4lvQUY7SWFsW9Fpvq5hr0yVBQ+O/Z6jdhm6ovT/xIfmmuZivB/qgh8f9lZ47ALwq33q9
9yOyIH05+x2c1NUPVg/1qtWCKX4U+Wf7uIl1cCW7t/xjnZSKezHFVY99JOSri9WuR1Fn7tOa2xP8
SIwzwd/80D19aJH7h+qROxLvss1YIdE0HDr0Jl+iwL4wjZEIa3cj6xLbVPOHLxK62ipqRmBYD9m5
k+4Yki5RltDVzOYJaAdA1wVoRdu0n2+uBUnQP+YEqB7D6ykTPEFrUzdTjcTdpPVyeFfgF5HsIj1+
S2AUkOnXa/dqR2iQhI8QOZUPZ52PIYRPLjXeLbdZwkRz8dFZifJGRr5S8JPUDIm8Zs2qRWfIMEZB
KR/WAm4SBnKY7HHrT0uosIwn11SFFKfJX0FL9nQCm42FHTMG12Ntn3w/oguAb4pbidvo1ibWY8e5
yww2+eZ7SKHjZ4/SubBrIQmxdWC0sLNc28AcJz1k/9J1Iq9+4A6ohMbQZ+VcC2p6wb75yJmG//jq
BgIwLSFvzu+6rL1UnGXz6AtklgN9LmnrjC4BlQkyAPVd/N0VWu1VRJyYatsm+VWi6/mcrWoNA7rB
rWywFDULKx9Rz99En/C0aZ06WIiwZb0Ab1lnXTIGb0lcXnlg/FMKVpiAVlqI6UVdD9fNLlxpuKRf
wkkTrho3EAw7/clno8jtKHP1vXvtWsXrm/VBygph8F8xbhTYfZbkmRwyCOmriOs1gc/J+fG/iUjA
2UT9v/moTKdjqguMSyh1aBddWMmuqTl9oi/0fhm+D6gYNk9b+qjjegQVOMhLshtJ/c0JSW5wd5hZ
rfgCFoZNr9ei1HVQsQPllaaY6ggVQzEBR7CL6CTdj7NOIraVcymrvyhm+ywElinj3oy0AI9ago9F
MjNQZ5XAayk7YaOWKym/1uL1qxbLWCaINFU6SKJFzxnyKyuqcgpn4eul9WSHJ7h9P8sxhDF8T8qb
kc8HdSNmMiJyes8M1cJKdmSA9Cwa+axSqi2cfF6n/iB1TydUHHp1Zi2CBqOlkFrURupTTRc54UR+
Ip/RUWmUm9p0d/groXswzH3MkqZvzhCRibrlcbADBkiR9IhlsCPd8KbReWOuccdbvPDtjTfiNQTu
2djojD7IL96uBYaDAYl67KeW88ACgYuchZStoPInLgyN0T3CeeioJWCSvY0qzFywevXkLHxWjeFa
NRLKVqfXbNlD3Akmr9j8NCb0lmVN6lN0r4eS3o0BqQx6Sm0i8Hj4j3A3JYMBO+RgO8jEOFZIHhAa
i23+RivVfCXBmHoaVN33a/K00097HKlETUinzDDJUvAhlInzCu67Lm2EXyiIA6cjbEMggwe+FQ26
cfO2PNT0lxvnfE9ppSZZQoTyMTPUgLHBSxqvIDwvPMOHO3iN6N28gl3O/mqB3qPSoV+1uDQ4TDb8
WqYxonnFOnr1rjXGf0bPO/iU0ks8nF8hhbLCe7YQJGVI3x6JQgQ0HUw0OnhGVvzA2ICvrp8uWD+j
hdi4yHeHodGwY6dvXoo14Tc0RPCKuLpAw8dctC6pEp0jlh95NPXOL3jdb/syT3VNAFK7M9hJRtvw
AGsR1EuNNYdjiZ9Fnw3Px005tlQabplLTGqVRQhe3subnWMcthjrEvzerWIottTn5sR23iakpDNH
Gc+ezWmj1MLnMRHLKl1w4TPVQ54Qg676rk6PtOnQZeY4ZajRCPaNPDGY3PQywRY9UcxJkoUD42vM
k2XI5RDLOiDyOI39y/BCIHuQqbtwgZUTdM+OMJkP/UngyN0OVfFx0FpzXrZHGsTsYiQAEh9FIUi7
45DQcPnXD+7cwXVgmVQx/5CIqRUPe2xC+eQD1w3TzwcLjuRI2LFF0sP2/nuXKB4T5KemcUbtUFtx
IEY7sKs3kfuwOJWzMMpvcrHcDMA6f0li57ibYIDw0wN2tUxL89ehRULQrbnLh0WNI6tQ20+AmNRo
f1vbOJJYrL/of+eCAq72e9ItX6HfKAdqlj2j+qWezQ1x3xfqAGfm9UnUIzk20PzYd71YeG6DlTLr
wy+tAcfl07aHUG0R7m/jG7yqRRyIYn50XwdCnHAmPkv+N4Cdvyq4/gzkukh+a919/9Zs7zs7Flid
Y9XXr3PpOYfU0dplPl9WpVYpVRiqb7QFK/b+XEQZa35Eg5rgijNH0lYLLQcqhoimYO9v3k2A4oeD
a0f2nu0/Cmas9VavZU3/Y5ML08ALpup0/tO0eV1SzPXHuCZhWiCbD/iiD/XSP9Bwu518HjuSiikJ
xon2gUwBU3C2GpOXhtbcp4NaUD9lOYIQGhw/LtOrG+gXE+lZ76GGDIVMfSPSvOmMnS02R6ycssE3
L5WoZuIdsiHhIjaMW4XJGveBFZsEd2aFDHEWX76AZuoIX3VoAY5D7D7tXD+ot0n0F+nmdbMA/yEc
SAfWZkskadK6JsNDiOtf0oJUg7hhbarX/SMo/Yoa+dkrmrdoPBYF/xvfZz01CkEFbfDLVYhJXLtd
654Ku2ba9jdIlXx2CXSFZQYF/WnoobQbD6X6+nl3hM/XAWVuTVYxZ/Q/oFThKys6IoWnh83zYMFb
bq8pGHTyyoqCK/kvioWBNWsFOJ8daNZ/muYIqT0MyyTHUhA5JCSTITOA22DODyQrE0Uj7dYqkeai
vBUQ2c/V36WFirW0HCZyzRViCH1EkW3kVhaqgYvqiZGvyV5Ghm4xQBJe41C3gXLZejJa3JjxHzwC
Yb2qqmor85mVhveIeKdfXoBz1YoR/brOLNdszRI8CyypevX1tq7iqX7PPur1GiEgPCV30EwiOrdu
mlrVaNXbRRTSiDWshZSG0fETG6rmW/21yMBpFvyv+ecUHhImlNjjiyIGx3n33svBzYmE+RWeG4lb
+7LHYt4zGbmU21LZ6gNaSz5lUtKY+GyEUDrBoAnfx/CT8xp/HRiqTTzlIH9ld8g7gNG1hjrlB2Nh
2LD737PMYtaId2m1OsQTGAUd2n3yXGxfZPjhYx746Dd48V0imjCBWlS7h4csVjJvJhMP2kmXhV6y
B4rLfa8S1Uwtktk7UsJwGSCxfuS4BWkFUXlTSK+Iejt29c5fhnHCFHw2iM1r11WMtUKDKWH1FkXs
m5/kru7lgIL4rxLuUBxR/hVFHyMN46Ya1+KqUz4Pe/cvLs1f0xvv1+UGcaoo1XHapO0il562O/ei
aQpJu5qkao70Zc0CbE9JKx1mleWLe6U0VEiPO5SrRtO1dj6+bETp8UM6jBIOkJwk70gKT8WRkJ6g
39YwrPbEoG9LAxwHlbyodZM/pYxVLYawqfn/LaVl5mpoLDadSJc0yVlFtVnXW8LJFJ+zX7KWURsi
VMoze1Txx5mdlyG82ePSpnSvyldzJ1TSKjmGbIKYjl2WD+wZP5GCNObwl2RQtKC3gtBSpkVUZQDD
WiI8oG7CJ9l2h43waWwm+fm38NsMRm0+uEUGeqBcxMDRicybWoE8NehwmD5hHzpIjmys0IfL0HGR
/oJP1/dzFytCXfDaRPJI+LaMk0UZv1cClHyddImw521WEhwLJNkw0bJBgqqk2sS3X721eswRKpIo
yc3UoM0L1ox7ycRLLj9MMLfDPZwjuRwemYhuzOuAHnTG3180S1BsP1YXCjVh22qQnLgUTE+cIiGu
7O9AAgXXCXa+5TN1CFJOFhbheZTEhN7CWV1xGXTPgOF/WccnEEEpYh5L0XdZ9Xk3Jw6abg6OHaR6
F9N0zAnIBygoCzHDxOdJYXMO0TaC2R/Dd+lYY6yeoyfvZh8Ky++FgNv80hW20QL66todD3S11iBA
iR9kKPje3E3d4RwAGVaHyWgnPgn1wpK1I+8nN9Ek/BvMRm7XEDE0tHd1ruziPKwzLiOaWe7U16Xv
AxPHVSckK2alf5d0dOfgnMs+/ybusw7OaI3MQe6FkGM/ZnSNKvvTPM5+MvDqsP+fFToyhVKNgpmp
BiKOCqAtLp6XPlq2S7EDkXSpJh482pXMoCE/Sf6SBVdJNwJqP3XHO/fLkWZ4+OCBsZLiGQx1Dmml
m12wvfdDss6DEJRGo6XuMS1yF2HsiAtW4abTW/NsKjuf7ehiZ5JXtpe3TScIhlfEbknl/8xQsPvF
B5QjBWV2m8CcIIHsu70qR0yFNU/7xBqqBVq/BEUgf3bCAVUTQQIuprl6IvSoU7x/ZcejgRePxNbF
mzNyu2OSl5MT9Q2AoQKBuxqtF7C9qGOqVzsTd7DxpQ1a69IDEvwhP7wNHXfZoABg/pq8y8JXu+dQ
ihhiS+2NzU8Qzp1JxON2dn2HaM3PM/eXrTBw+fE0c3A8Dsy13HXTQsHhlLccRpu1wsHlL6X7BnhY
LSkSPn7GUuUhMQApJQiaUONaMowG7c6MulCV14n3wOK9q7+wmIi46sSW8vSsX5TQujCUFLJA9Q+M
P+rl4Iqjppb7aGcWYLqgav4MIC3ByCWw5b8pi93jcZ8alr9DtVGugr4Mbn0YLn1UTQ1o1g8BNigK
LtkfXqJ/KXlr4HskKwYj7lQ68WBI7MyohEMTZOvf8Cfup7hD4i+ZOiFYCEigR03FTqzO0kMRLEf8
cJ2iPDwzMypauQv4fZMCojnH2uE7fOpWdZZmiZEeI5/HwFIj205SqaQrCe4OQpyxmfNkNuyVcGKf
1YFBwkQOU3j0uK2+5yvWDhlTqlB1gyNGIR4r478b/RigoAl52pPMEITAnc8Ojul8o+V6SWKs+k7J
BBixsVnKcQtIgmyqDDfDDMcALczbhMkbNcWqLdOMdKQA0R3RhYA91R+Y2B4h3lLE/xeVsS1bmF4M
PS8teLRXZ+9ydEIgezb+9LikDd5AjIzWmU97Oux6IPHgStYAEYRYeh5Cc/efvEhvaqJnPxo04JBv
Lrs4vCQyOqyQP/VjYXV5MbR96JdjHxjOAdrNAS2MrKeCwJRjkOYhbTkEypfSgD4XiDq68+ZG8TOC
8m6XCKdqK7rsAgtijKwIaIMRYrUx+mkBKYIkq9dgbTl0mxXSJ4rTFz32OMEZuVyujKeWDk8RVtks
j0KDyA6gzEtExdmoR0Z9eomMlToqKBqmSeb+sHUuhzfGJzjP0Z6ECbG7hVG/Ka1u93MIZZL4gAMQ
lhfekwyEcIyWIMLXVyjbmTErKUzwK1VAp3cGq8pEJAlJw21rJGRLKlgDsCtHbyDGKjCNEpMndcb3
3frv/35A1twxwfI+zUHRMBjjj1gCiTIpbeB995MPRCD/jMNoRcyoEwKcccmiCUZlAqfaBYKD66Rr
SLflc+ByO3RA80STLkXUEbHFd4JVdXIRvqc4HJJJgfqEmG3hgbTA3blnE8jxhYmIGFIHl+t2l6oN
9yZVJE+tCOP/66LNlclUz05B1/GIXHcBlGUadwRROH3onAjUQ6yADPTBi4BrFnZVjOZ81qKZ6Taq
RvX6PbhyaIHOno+v+BhSWwd+OY8LV37ma6YiJnirroXXtBBP0IVKZEhD8sGFTfFKVFMh7wbXVsmN
jMNRKluF0vqKVNSHr3QX9IcfdZAwetPdJ7ZLmXP/U94Ay9QNukM3lcM7hK1ObdNL327Ws3TV7p/I
19Rsc3OBQtKle3u+rRTNUvGZ4tfsaLBOcD1bvi1d5SgiPqVJtHP5kFJyPdhECm9E6noPm9RcDJXv
Vxk7PtcnhJjgqDHQtzgJn642j0PcSMDplGabvV1Ox1EbzA5W57iwQG+Pt9lcl5WI3RloCRax0ZEd
TA+vJVfhvHR8YlZn+Bro5mpJVjH03oNIa3UlUwCC6PdJqQD9aaSkVr1dxxoeg3WuqHVcHdCo3wz0
kyJZjXwypP3pgxDiBjIlQr/9KEaGisruKemlZmXLjg9i/QHIH5oSAZvwGEMQFQ/triijNDZQTlD+
FovxpSHJSmuESmLsAW9bkt3ZpoVvFsC04YiCVULEU/spqVDDEX7UYwb7Whep5dpyZIJ9CQeMoB84
XQ7D6fK/YIC/ZGBXZ2p2/vQdtQz79iI3c5lPU2tBusmRJRXviED4A4UKQcjqu9SvCLNjCIEElxR6
KdJnVFIFgGmY0lu8OMf58MpCst8KQw+6W0knjaWpAXMyng1o0oEyL+ID0HhIjl2oDoyC0TgRym8T
FIvUE2k92FCIBBEeMyQlP434cwqKUgHn9Ht5PWALZht3TMhkRMojJqVvOHuTKX5wzZjNA3HnT+mC
4NHpP9yeE35n0zVSJyqBa5DQz3LK7aoSuknNAUss3HiZ3XWszepcYGTehS+c3ycOjtjHcf4FOHZj
O3JhB7mfWk6MtczRVN4cPLYiuqId+1dBaZERkoo9lcBuEnRU3iTO2U7dbAZsCmNWgYaiSbEUxBSh
QPzCrJaq6YKPam3KbdwHL5ChKrpKQEGI2D97fq2WpAHBso1ueXipHTHqfs1EFY/ngAhVEam9k8ps
9lBZl+2WzauI3MGvx/1ZoSH10OXNP0x3HjFgpkGoywvb8OWJA9Uwdj5FK1MVgGb2lUTd5RdtJjEO
IklKqfoZO+u33p/unWoxbdZMA0MkdWZn9ogESoWM+yb1MPlpuMEEXn4aQ5awNf6m7uAj+e6rYOxf
CqBD4+mr7LdoAKK2DnGTRxzE1iXA/pUelVqXvp8jFmioDczXpqdkkRfurIePa+R06ONW0TAv3NsI
a2oLbZ69ws8ckxutFl/YpQzFPTsss2Ueu2B9Z7U6KLWk4n1mI9hB8eRCupwIqVOIAIAM9jz6W91v
7NgigjuI11budJUBRxDqxAqj4cT0c3YyAp0Tb1Kgu87a2I9DYehukbaMG2IYJH9Kjg1Ej8fNPZjy
W+TPLB7/VK04SdftqSqJFMls7CU+RuI1t/Mvk1BS4pJu52loOHijTZXIR6Zqgy01eTpIB456AKfS
W+jJ3Hz4jJxMKVMf3iEzB6pnbxUwlScgkhVn5HNaCd5PhVAEF6cqXLFF6sVy/VsvQVVD8auWVoUI
1pnVHJwzok2L5Lp7Hkn0A+f3zJToDKnufp4lsW9x55lgY7iswlk59TW6f8iDhDCdiRANs/+UeWRw
sxgtfgxBiHN4qSZuQlnmK6/ojP2Ov+XfQCgMscxlK8ScBKcGG946pqQrN9IpiJOGvPF4RriIYC8z
mwDgXa5D2zDloMsaTFM1C88hYgFGWKYGECBAm9Ehk/TybabgUAH+AUGZ62G1+Jb6dtq5LhXIgnCt
kPjQ3PloW/eIUv69XAJKo3UqhR4BHtfFggtRCr1S2UyWoq3+sXYUVh/t4wXfAVB87GlYR8Lf5QJg
ZVyhMxp6o95D3WfMDpt9F0e+hF1hQy0hpM1BANJvT4Tskp9dtS7crk5bTROvNWi+jN2GnDLDl76G
HM1u+Xkfmyi1cvCbTCz8EX/FTEZOt8wQF70KI+5DQQXq21X3PXtAIHDB4KHKOEK+mFwKOtUrEbBY
pJMpXnAfPdvdFqLXCfWRfKykjONkVCoGUHZcYyeESojQ922rWE4irxC0xnIf1vrF0kL5PHBzAALe
I8+Fh8GmgyIcV0d45CnclwLD36Mazg+TUzCsC9v06YWP/mEbgzJAlmggaJ72ITmdZ5VQlLWE6JaZ
WI54lo7p8m8Dw+4fPQha48ZzWdwB1uSn7M1giI+KPFFtbiBVMHoTCRkcSbB4Wlg1up/uC2+AEOtk
kzjOG8F9qMUg5hCRgyiIsScBBPKWg5MzI2Fua7Sr+93p+zv6YAV3UHuVSpvHh3iXK+pzZzwtCYeu
/jI7u8KUsCdHI3tYuomhgkld1Xket3fjbOMFKqVbAQhOYDWfZx+IVRt1KV4KDRvt3S/1AOS1n6he
nlrNXmrqYFfBtCBs7fSJvNY+/YZeTK56PPQa9rvCBhOiZvazAHG70b1e7w+GEF0fx+FMyNuJbPuT
EjIgRkpTElApngwtpsX4ksvhdDETEVhIaNi7PGE5oViZ/elxiBuNZzcC5fudmHf8VqV8EBZnKcZV
+HQmGSpnNSebxMlbzj55tMrk8+HXiiQK5jA33hIELcdo8+VxRsBY9bGl1XiUyCP4ZG4uB58LvdsU
lAwci1OpXtFV2X79izZr17M+nrqLd8A7VG2bpkwvvGAyqe/zo5t3K/zeI2kQoN4XSsT/jQQrNC1K
O+8gP4igpvaWlay7JpTbzoFThlpZ6KYeOg0I75fRAR+rIpQijgKlMHI/lb46Dw7+YbMjRkBVXM4R
M5lZjkAv7W8rgz12yqyBRBWkNoeY3q7ew6A5wvAnbteKygE7yAajqCqyEkCdsWYN85bPLss7dAji
PxZndzmL69SkFLLSHufwvtNDpp/d2irGSTuTEOl81kDMuYTlxHWZDhMPG8Twmra4CvNegWX9D/zY
Qn9M8kVp5/VcKoliTw+ZpNPYZOg7SHLHc0Jl3NA0y+hFJCIZLLOgeEXWKAHILRmN+BlJ3h13eFgo
hDBoYEpoxVFYuUD0nigEnksgOZErJxCkDz9SmnFlQ/GZBihQNI4XkPMLNz5pB3d/XdM+42spzE6O
vF4pQGErOQ/Y/GLuru/yNy9FVrhgBrJ1pdxKbrZRaNaRBJxoqKG+BTXdbaGagAe8RlyKJdLryBV5
gw+6lfBEE9RoA6tWyrTNtHpY5FSJGeWBofhzeFw3McQaZNogXcXQBwMIfkG6P5NYAH2dGh2oJloF
/8Gwwr3Ho1iPhIT9iw2cSupFWTK8Bwiov10BDxM6n+X3KYVWBrBit8Z+DqOfOcPMj7fSftezvTMx
AXjHpdiu4hxDpTqmxv/KsZqOT6qBIZ52ncA9RwLFFYEIo5gUVbV0lQRo5y7kM2LSQAUA6HO2qhVv
+SgzrMS6kQNqw6nezFv+RTB6gC6nSIMXFIBnwiG/d9s2vRY0uPfX6Dou//q6SoOOA+o1HU54yJ9C
Egpwn5MLrEETTAmfc06KmTIV60N6QyTBDhjhRHPkjGk41ZhPXihQcqadh/ChApPlc/BHbfHpMmvG
H5Tex78GCigUivmhhhKLOZcJw4xPEf1noTdqJtBdHoo4vFZSZuJv615RqbxU628opDBV7IIngNjV
o4e/RRHOp3zIWdvN3rrhCFUJMMwqrIbPZvkENYshMLUNQLHJloqPuntjQ1QnvYDZnD1yi1zMypdq
7Lnl6fp7zJ2dqzZycVvWj+f02UpNv1S8BYE18HuUxiD6H41Eg7TGHsO7QJtCEK6cRZDA/wk6YI+N
X8KQISXj7UWTV/X1gdiGyGfuXc2BRXALTMLDSR2v/NOMBU1+HzQDCcMsZ9i6JiKNwPQKM5B13YMV
c0UtmSb7xa1RPv7RMTBi779mc0Ak1cxNvyupxYdVI5QCBXy84FRtFU4Fwv0LiauYdvu7wNXDlG3G
734mYC//QI8m3jm0N1Qb+q+tSq0e9vsN+ildnCd3gTW9xsZwDKaEMWAaQM6yMScgYqyxh6uqWrvK
ZuZ9KEvWrDCyMJqE+TwWyxwO37oO9Xjhhq64YhRtUxK61ddoCzuKA8oP868w/pc4j8QMTG7BQoJz
8ej87W2IQxiATPF/yVHARbRzAvWPR6qlmz3qwYTjn+CZWjU7kEVUXMIfwRrkUBeYsf2MVdq0M/35
GPAnYlE7Fh1pPkn82YvQgfhV0Wg5DykKQBm8hCFOCTWPwMZDdn/lAYN7IXnpZ7G/yAkN4rfUJ+ry
TXflfa/zglhVSaDxjV6fw77A4CAAtueAAvLaSopWjTx0z6M98zqTqptJRAI5bkwhsnX/mHfHXpVE
sFCn8RRSQpGpoWlLWQ0GNgU0JYiy0RohZCeCcOqkGRbfUOdRWgJeDEn8i5P5BMggu+OfzrH47rSr
JZR9oN0KHIad8YakWw5AV9MMiuvsQXhfSI8ojbvYyb/pWykPp7HmjPJgGpyOUuaOzXdPy5YgmQaF
ktQx32DyUKPZ9WwOX2VLCR31uTvbDGg4xm8bx69S1bUIAg/DM1C78U3w6+XxDBkFBstUg98/AyZm
TpBfXQNKL+K3cfSCeYlT3l4T/II4HDgUMACOXBGmnb9Xf3BVWTs00+cakVFHxVYcoKwqo+lDOQ4D
5+iNfBU3eKQLZyyOEuon2ZG7Y27eyP58Xkk6vPjI5EVkkVpratXUhETGanpEZdyZmG84PjiSza1R
jI9f5eWu6UtKVkx8ejUji3KlDtw3jjKehPEsh5ZcLl4eX6BAN7j3q8DFVrtxfUSdQxuB3jzqYXz8
x3rpSPm5xeM7p4bhfu4/wOfUIERZ/WsUu5CEio5KxXmt+LrJKLp0KGuO/cQpwq+QO/MavTgBVsCN
0GQEib4iISiDdUK+QscW+w6fpBw7NHNgcyL7V6u7F8aDJC79mdzvQ4+iL++X4H8EWWWm8AM9GBNT
9glilc/cwou+nrP4dut6Vn1XAucD8rlCepFeC8xI2WIZDLz5kO6+2dd1jKzW1q8k/xCxLSsi0uVq
GozQOc0q79ZTdjCr9Wtk0lEtUJzZX4hyOtXO8/+qZbjT9rWGUCXqtmJ2eHGYxEDFweMNHeGvHJE6
u3Ttp8h1XKWVBlNzLAYycK1MeIRyWvafcbNNvQWMP/HuKhcP3V8iKsLFDtFvKmuICxXVA+SP1KPk
rz/4Baq8npvJcUCBb8WnRUu6AOwUJYBy9HH7ybc0b1WpDxJPTYTi7uqgWE+YsfWGWoh2RC9xVRZo
yIf1piOEnDO77JUmqgBad9zUbv7XdAq1Vs8XnI+KSvIXFGs/9y2+WsuXdRl2XLIg91pjRyWLEycJ
2QEPaeYtoVh6HN+0CNT0U0zTKy0BthHUsKxgqgmbhyBZ307JWQIlzEaHd6itQRfrHFwIQaRpts47
WZhUPkhWRiAHiMVBSKp93c4Oa3UM6zpJ5u5O+WZqH9OisMa5JE0N1+wp+few8Zd3IrZYaOEa1IIa
/YVcNNnuP6X/sJFX6YafEq2Gt+INEktFst4KVIKWDHJpNbQMPMnwO54PPG3kJpsRfDJF4PzJ76vU
RGfozZkgKrqk2U6ML3SOqP+rfdLCNugE+9Qa2wnTtUNObiic5H32c+BjNQXNrr1JrIVEjX2yeYpD
Xmr3rQv+ic7LU/+P87wMH/DPwCcLC0IGsfPE1t0OSDj7Z3GrB3bZRZEFtA3xIVf8svKr8KIQyAcA
HiKUlXti8ajMFbmwob2sDTvde6ojKcr3p2Qy19vFrYvqYfMlR6vEXatbvIfZgsNdDLf+Q0dHvQel
n9MC8D1rE95/YdqYat9Z9O1twjR8O6uRkAvukiAVTZ1Dd5gX3eys6WHT9L0oEt2Tezj/VB7sc3Fs
cXoQOQocH/AKnfdCnT61G+ncTRE/fOSVmUnaGMFWKIKhm++Z5h6pA4tVPd0/g3T7kRfFdneCpdQs
1PeHJxpHaqNMxxlixz3TPIJ5qq1UDA9exvnT/HR1YjFPRxRQHqjZq87joxsj+l/HBYmxIOloYHsU
skVGLP9i9WOQUxbL8Fe4Tv9KKOkyPseyQX1QnQ+nppdtXzd8GAcYKZqh0OZWoaLXgeS5yRhDyePw
yXxh/xieAcPNoXA6jfQ/XTADApdCSaBsvJPXDwu1K6mXqnqj+0mqeRP6k75n2aM4F8lIap/WPvBE
Pd1iKzhp5P3NFKMIXzYsxqR6hs6DpzTzAysK6i6YQ//TrHaAzplTr3qsjqbkrHkiPwHDqS+Ev5r9
O2CeXE8lcILEAFqkwDc9peoYXPGCWn6z/JCMQCnUPrvSLK0wV6sPqtSYMXPuzUVMHYx6BE6kmO2+
cYuO99iEEi4E9P1DrLE2tjRrU+oETh2CKF+U7F9JxYxZ0TpBrcd42y9iMGyRwrgr2DtRsd+RW51l
P+FqfFB3v4SddMHVle8u3mM1lvvHID/WHZQbyOksIFiKlCmbMEFEafuCW8XHmieI56xx6fwEBlWZ
WgvpLCJCE0l2p+w0wfuWjSj+wA7vNImyXArrc6PbqoYCdH5A61vhAOp3ic04+sn0pS5nJm7siAKt
2ikVshzsawOmcdTnsWEVPLqT/WUx49NTB6TWeHppwarepB72019UC6183TszFXatXJzxBBVpPuWB
1vYxVnB6+jgWn+X4ErBSuH3ZAbbzkQ8gVk3kTGlues96UnLpTPzxMn+S1Qy3ml9spow9TJK+BfoX
RfFZ+gW6SSHB5sWgyaUil3+5IQtimlH4n0XtnGf6ZaC4ZKvKI+CNqT/thVsL4hTgQeJxGNznc6s5
b0YnEQ8jv1RlND2HWFh92C/3+qNd08sITBFAvG7/torgKFcvYKZCFCh7YZd3sQCbzPW1MQPk9zrm
wgWl/U5+xOqdTRbFWzM5sAlxLgDOlAwAHeacj8ZgFS60m2tVhzgyTVmGl6ffSykjI/fj7GegOpNW
DWL6IjjvZLQfh6MkjG5QJQuo/y65cyEbnzUAYHiZAcyAklynj5Qp1ydYs9Z9NoEVfBbEmrBBP9yC
bzNaqT9nA0II8FU2KSLaMlXKq8BjbFYh68nGRlo/Pd4xZ/gOZSFojs5Q7psGTrGG3xNrB90f7DC8
by7wArHNqB1tWgXc1HD83VMujpfhCHt98jaWPKj1d/owcm7tSN+2QXCIfL4F/3NsEuywcE5y0pA+
Z3pkbkvZcX0F51+mmqlfk7W0RdUCPPJmNarpXbBHGTD1u1zrR68z7AnN8KVxAPugygsLYVbQkVa4
lV7AsE4F/EhQT7wUMfNFjEwnKGzfGMcSW9YwuVG541ydBsPSn/v/MWhaARLTcZX+X5C+DYKp4S3R
iEwOof3lzlXcqYOyeKhn9aRLPtKymN6HAcui97KWkuZCNYR7y1pcaEPK53dQyLgyk0/Thdq5LoNE
1EhG0CBeB8h83yXN5QTaNLT9d3I/KGkL+rFM4voExSU9JXMQ96MORsBYlSENrYoDic7ZfEtHy8MQ
rHMElWz0nw4/uaC9sVUkMTyJ4s1fE6MSQiwPHKDTtFTtECgxUeAhM5yIoSXY8e7fXsGZsCV0DobT
dGN1191s4Qiw81jgjxjNhnmb/drM6BKUAYZfwl0eFvI/hPaq+c/IhbYSnnH+X+ZRksUvtl7UAxC2
sWkmnT/m9xaQwAoatpYIji9HYiN/8K+sasCklsdlkV9ncRSjCr8Ao+qdZD3nmDCW2iS0OkfOzV3t
NDTr1GPqaub/sxyYktBk8j8NgMaeqtYb08l8NQco2tWp7LEZdAkmMKX+f4s1YrlJyLgaMUCwC++R
AO02yOaDyQ4l2Kykuuc+nx5sZuWDi4HWLFtmzNdJ9RLJKI67i40jEdSeDewDn5CkHy6hZ7BKLGD0
so65XDeEM5QJPm2YiqtjAMoJpn2WBOEA6j78WzT0Az/XZMQj+gVqGbx+DazpQjdCMMV9GUc3Cgeh
cq5rQDQB5qTRvl6H7/pVlzQQhSV/ay+xsu13r323tH4RwUwOejvV+ubcOKAiBbJvRoyEDxRnaGhg
l2H/Xa6c5399dX9SHFfCayLklh2ix5kb65/5qhDQ76A9uafgITSTQMa4ltAIqvnla/sPLx8ary+T
WAsQQqZMOUHkfIcxXeXUmAWVRute2Q7wtTomAYcCPDdRl2Xe4i1dhZ02L2pQoQYUjzR9ikOtBCtt
CqQ7ie7P7tChikt1A/De5sxP1Fk0oZmwXRWAcS/mWG9j/JQNkaTVGLqb2mZTebjg+2P/NfrUzOjP
OLIug5Mvft5Tebm2vsOoGKrIy1H8kCvgPXTx/cUyKoUlEdT2Gb6PK9zZST7PuXJruHuvMZVdA9Oj
9o225wHOby7d1bVAHm68b6ij7LVFr0jtfdHIjOGuNhDkymH/LSKfnyknt0IkytD2Js8LyJQkYyK6
+k0jhLKPTxCHf8sEMuduwpvEX7BnNhX1t8M7C+Ic8GpE4Ja7dWhgeoNwFlA3uxk3Vah03wSWKkTc
pZIcpr9o33zbsRjAef1gWNqtvI/r8VT4jQzX13FEs6KsrloDdCXOG9gsABwmqn3YoBpemqh51rYL
q539OZT9/CHq4TGITmTdyFKqv7iLwoY8t5MMQATF4AOFKvosY+jjIurnj6i1OVUeFXUZotEBLdEe
Xxyaatinc1lpT3LhbMQS+IU4rhwI2GBxTxUCMdbRxpRF5NzcQJZf9DYRxZSCZzxbA4BckkWWxrFR
cJsxavhTTF42yDkrQ8FtZJL+BPxcvhx3jR7OH3636uuktXwzbPLhThgP0R2wsP96F2Q3pVLIacK0
icG+T6SU4coP4w1AO/GX9uvGE1CX/cYB5uywxLEj/I1T+CQwVpUuoLpVoBKfVriuLR+wshPpo0QN
+9Uih0x/6JmgIdgpymXhatalgFoR3mr79GHoPC1L/mTN5C71Qg/+EoJTNMzEB8UkrLz/8J4wR85g
JqgA8i6uB9Nxi1SjnKpfNnD9mxWB7gbIAYCZUSvwKaRx7YwDrkQOnjfzqC3HQ0Vm7do2gs74O1v2
EIi2zym5PmUszIe99FGHAhOrs7QvXTVl+1K/Lm2GVjZdrpAKfi0Y6AgnN6xRpy2axtNpRRmjktR3
YpN78L8Qp4G14wKIqrELAsVYrS05U3wFYSTvcialt3dtuSmaeAwtUABCcY7YXjhC0f8rKZO3GOmc
uPXSUWjGui/tk7n/nd4BxoRC4smRb+5Dwl1ugeJLZdMhgj4unZ1SUYNRmqZx0c9D5YaIV9lJPrGU
knvbQT6IoPPumlMBZtaTstMCXLUYZwUB1JdKHRKmszK1vt9uYN+vZ7bemmAgNjzR8re32gcQt0x5
XIPSFI3OBL1hecC0u3tyvMsZICFvnWgho40JBb0FsVEAyqgNgl+G73EwKmi6r1Tg/xZ52ivbjWRu
QMzV+M+OYq8LEIlaGStKZrIdxC+uYaRSDxsPI1WUz5HCDG0zKL0ALExzy+PESEK1FRHSRCtMcrUp
G6li+jhpBJ9zkU+0G1UHOmKh9oHqd641A8cy9oTbOMChX3Ev9iFk/jayOopkvGkKcNrpAPTEeyOO
4cVX8/UXv9pcDVtOdl40l9BFWMpIGqD6kj2uddh2SW4fa+4zH78e3H4hHdR9do4MIzWaxmBoqYUs
UBRjnZhn0X+76Do3rw7jObPbA3mNyU8BgvVhykA7DGD+o4cDmqIv6CG8liiLULSRBWTLcxxqDLKE
miywUVYdmJpgNqNYbK0qbszPiMSCFa8z5aty1Ufte+6JF5ggB/cARCpEBgezgRKikD5w1cs2ckTb
i+0UOCS89yKvbCZZZ7cf9M9uvgzEoLJd2O3uFHrKn6DKfpZmFTFsHfSfR9jHpfludzfiZJ1tHjxW
cZUQgo6SgN+wCwRL/sm51TT4+aI7Cy0UiosLDdi4RQL4xsGPVPOAQjXeSPppaWWvNnFT/5vtH1BJ
kInEOrnG/QN5u3LcvAgPut7G6hUtVS8iEcYV9E21RfS/kkZxUph8A0Nmw/oF5V6onbR4+s4dyAoG
uO9glfol/LsTkkJS0LX+8ZQtdUwCAqPRdy+sv08mJJnENd0uoPlwMIubVgua/zKbg1yOA0jgKS4T
lsKQZHvw0Z8QCVZDkHV7tyvAVTbOFhxIwn4913u3FQ5Qn7j/ktARzCg6ZWEHL1goh3nZbi6JNhCU
mwESaGFNgG4U9nwq6iWq2SkK64hWeFsi656UEBsrw07H41ximh2t2NMscY1hZL82CY2xI/F19tFD
9yQSOp4rtbsVeEJsI3Yq9ZtHOOvdmKcI6lbj1g4myDn9g4LvKY+VNk5WlhVKZXjUhHfJFFViVvnf
wfhSQuTNUTK6rTYIZxgdxkZj9X4QcPdCRqlWPsXUVomwjB6Sem+smPWqDSkSFzYuqNxYriUk7cwl
h27pB1cQmbYY9tuw9uM0/yF5wpC8daQHoZnXL906wV0QjZq5GFdBFeMeibJ6mnJa0MvuPn4B1qov
tiNMmhjjk2yLBa/AAlOcOp0UvYoW/ysPXK8zdMW7FzyBw0RxJS6hCaqwBjEK9FZ8NmHXDcup7t3J
KdP5HaN0i3osPtwKGzuTz4twO1vSL0p9qa/sfmH3ySIw9kc4eGtqXz6v6n3Gz5SdMOkTnGlvUm0w
5g0LASMJ6HlAnyBAsv1adfwTmDbBke1V/HKKJir0+f1hHlLj/pSRGbmazEZQVDlrLWs+4eg8OJq/
vdoJg1akVVk7tn2L9uqu/cYCPlCBCHGoSTASxbVFayUhbo8j6JG3ObiraVozii4eB6/Sn+/lseUq
iQMZ637SosirmQaz0uvzV1uSxFp90ne8VtFfw3PlRVrZXwfqtZAaql/nMoabiukjgd/cHF97+Aib
wivPXDNgsCSz0BuS49TpTqpm4lFUxkhLQ5rEIaQTL2UXNL3bUvgSPGsiOmwOC4kWIDrC+feH54KU
2QHRhMfqAsZAvmTDqSXZDWEhFL5rHzGFVw6Yl8oovOtLDZQ93CbQ6bQKXDehXaCWqPx6ffplYi1L
YJD4Ke/g0MD5wdKy6UK9JfVE1XrLB5u68t6pgFMBVOxWAaE5KnUfH4FbwD9aEEzu8HlGhxYNA0dB
3NGtsfPgBWfA1qOp/IcIuF1r1LmfKf/XcU2nwxgeXp9wPZtFYtiEv5RuavPhNrasOK3jVQlPlE1+
35xk+uYIXKlzFCk8A5m++X8BJkejHWmMjRx0owll9VQKsjL1D08YtythhGkhMcOvvDTnDLUPPT1x
7ke9RysWrnfa/R2vv9Q13MuIxFtw7htkJ46kw8zjjshrylrc7m1WpbDAdeCXcv9C7OMVuLMCjHLF
WNU1mAd8pZu1HE4oxOjKO8B4sRgvQERnXZ4iuXKqVayUi3/yFePiqecoYT6CGh2oeKGtSDuvCIC2
zoHTohBtXr/RSu9stbdYNh1hm1O1SobCEHIwn8gFKw6BcG5FeKOhn0OVgykENclyPvTTL6S776Oc
OPUw1/5AOzV6Ikvw8ct/kyu9roCyhxOPQ4VHBEFlaklvkMhjiKzcGA0sli7zxi76R+zle1i8WJdW
cT0XvDG6tSSD5yqp9AyxU8Z9M0uKzs157ksdU6XQKQ3Yyf8dnREoIk1LEDN9cBhLoBluISPR1y9U
v2A2dwIn9KIO6K27mQUEoPC8ME5g08OEpRm/T1MUAObbgh/aki8p6SJU6Wn3xic61v0qrXsIp18U
ppxJNYFyJQKsP7Lj9wkM4zveV/4hDebqqMpQkHIcPccuufofZwffLzN2RWVXN/tch/4LDen9GEu2
5uCKVf6t93EgHqhWG3+PyhBebuB44NYOqmn5FVmKH+BT2t+sI8ohg1o079NnjqlQJzKfvE+rTO3Z
XdS7/3cDA/N0WcGzj+aaNS1Gomkgd57/CK9hgtRAXPj7SDxIUnfEslL0S5YJF9SeDNevSXjqKdpq
6WEmpfcW46qneCsshgFVYSMS0PibumnmpZsDueGvnIfKM5/a0xPWi2MMdXtdGQ5QVhyrlyD0G5XB
39PZy1PgwmJzfLRPZWuct2HUQ5zL2cHGO/i0BwMTzsX6rm9CbhEBAjPRid8GdfvFJpDJKR3+4CSK
tembqfGezMPJE3ZLkpZ+/MYkVkf9VrZGsUUiSjGFr9SBL/dkL4CANE73cZCNmIgxiDGw20ALvvnF
cWVg+yYpkbYGK0vEU49pfOgOwoZNVShSHbdD1z3COAWbiX2EfNTeKmHSifeG/QKHhaqzTvMUAfE=
`protect end_protected
